
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1090 ;
  wire [3:0] \oc8051_golden_model_1.n1092 ;
  wire [3:0] \oc8051_golden_model_1.n1094 ;
  wire [3:0] \oc8051_golden_model_1.n1095 ;
  wire [3:0] \oc8051_golden_model_1.n1096 ;
  wire [3:0] \oc8051_golden_model_1.n1097 ;
  wire [3:0] \oc8051_golden_model_1.n1098 ;
  wire [3:0] \oc8051_golden_model_1.n1099 ;
  wire [3:0] \oc8051_golden_model_1.n1100 ;
  wire \oc8051_golden_model_1.n1147 ;
  wire \oc8051_golden_model_1.n1175 ;
  wire [8:0] \oc8051_golden_model_1.n1176 ;
  wire [8:0] \oc8051_golden_model_1.n1177 ;
  wire [7:0] \oc8051_golden_model_1.n1178 ;
  wire \oc8051_golden_model_1.n1179 ;
  wire \oc8051_golden_model_1.n1180 ;
  wire [2:0] \oc8051_golden_model_1.n1181 ;
  wire \oc8051_golden_model_1.n1182 ;
  wire [1:0] \oc8051_golden_model_1.n1183 ;
  wire [7:0] \oc8051_golden_model_1.n1184 ;
  wire [15:0] \oc8051_golden_model_1.n1211 ;
  wire [7:0] \oc8051_golden_model_1.n1213 ;
  wire [8:0] \oc8051_golden_model_1.n1215 ;
  wire [8:0] \oc8051_golden_model_1.n1219 ;
  wire \oc8051_golden_model_1.n1220 ;
  wire [3:0] \oc8051_golden_model_1.n1221 ;
  wire [4:0] \oc8051_golden_model_1.n1222 ;
  wire [4:0] \oc8051_golden_model_1.n1226 ;
  wire \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1228 ;
  wire \oc8051_golden_model_1.n1236 ;
  wire [7:0] \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1241 ;
  wire \oc8051_golden_model_1.n1242 ;
  wire [4:0] \oc8051_golden_model_1.n1247 ;
  wire \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1256 ;
  wire [7:0] \oc8051_golden_model_1.n1257 ;
  wire [8:0] \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire \oc8051_golden_model_1.n1262 ;
  wire [3:0] \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [8:0] \oc8051_golden_model_1.n1279 ;
  wire \oc8051_golden_model_1.n1280 ;
  wire \oc8051_golden_model_1.n1287 ;
  wire [7:0] \oc8051_golden_model_1.n1288 ;
  wire [8:0] \oc8051_golden_model_1.n1290 ;
  wire [8:0] \oc8051_golden_model_1.n1292 ;
  wire \oc8051_golden_model_1.n1293 ;
  wire [4:0] \oc8051_golden_model_1.n1294 ;
  wire [4:0] \oc8051_golden_model_1.n1296 ;
  wire \oc8051_golden_model_1.n1297 ;
  wire [8:0] \oc8051_golden_model_1.n1298 ;
  wire \oc8051_golden_model_1.n1305 ;
  wire [7:0] \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1308 ;
  wire \oc8051_golden_model_1.n1309 ;
  wire [7:0] \oc8051_golden_model_1.n1310 ;
  wire [8:0] \oc8051_golden_model_1.n1312 ;
  wire \oc8051_golden_model_1.n1313 ;
  wire \oc8051_golden_model_1.n1320 ;
  wire [7:0] \oc8051_golden_model_1.n1321 ;
  wire [7:0] \oc8051_golden_model_1.n1322 ;
  wire [8:0] \oc8051_golden_model_1.n1325 ;
  wire [8:0] \oc8051_golden_model_1.n1326 ;
  wire [7:0] \oc8051_golden_model_1.n1327 ;
  wire \oc8051_golden_model_1.n1328 ;
  wire [7:0] \oc8051_golden_model_1.n1329 ;
  wire [7:0] \oc8051_golden_model_1.n1330 ;
  wire [8:0] \oc8051_golden_model_1.n1333 ;
  wire [8:0] \oc8051_golden_model_1.n1335 ;
  wire \oc8051_golden_model_1.n1336 ;
  wire [4:0] \oc8051_golden_model_1.n1337 ;
  wire [4:0] \oc8051_golden_model_1.n1339 ;
  wire \oc8051_golden_model_1.n1340 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire [7:0] \oc8051_golden_model_1.n1348 ;
  wire [8:0] \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire [4:0] \oc8051_golden_model_1.n1355 ;
  wire \oc8051_golden_model_1.n1356 ;
  wire \oc8051_golden_model_1.n1363 ;
  wire [7:0] \oc8051_golden_model_1.n1364 ;
  wire [8:0] \oc8051_golden_model_1.n1368 ;
  wire \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1371 ;
  wire \oc8051_golden_model_1.n1372 ;
  wire \oc8051_golden_model_1.n1379 ;
  wire [7:0] \oc8051_golden_model_1.n1380 ;
  wire [8:0] \oc8051_golden_model_1.n1384 ;
  wire \oc8051_golden_model_1.n1385 ;
  wire [4:0] \oc8051_golden_model_1.n1387 ;
  wire \oc8051_golden_model_1.n1388 ;
  wire \oc8051_golden_model_1.n1395 ;
  wire [7:0] \oc8051_golden_model_1.n1396 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire [6:0] \oc8051_golden_model_1.n1557 ;
  wire [7:0] \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1581 ;
  wire [7:0] \oc8051_golden_model_1.n1582 ;
  wire [3:0] \oc8051_golden_model_1.n1589 ;
  wire \oc8051_golden_model_1.n1590 ;
  wire [7:0] \oc8051_golden_model_1.n1591 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire \oc8051_golden_model_1.n1738 ;
  wire \oc8051_golden_model_1.n1740 ;
  wire \oc8051_golden_model_1.n1746 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire \oc8051_golden_model_1.n1751 ;
  wire \oc8051_golden_model_1.n1753 ;
  wire \oc8051_golden_model_1.n1759 ;
  wire [7:0] \oc8051_golden_model_1.n1760 ;
  wire \oc8051_golden_model_1.n1764 ;
  wire \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1772 ;
  wire [7:0] \oc8051_golden_model_1.n1773 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire \oc8051_golden_model_1.n1779 ;
  wire \oc8051_golden_model_1.n1785 ;
  wire [7:0] \oc8051_golden_model_1.n1786 ;
  wire \oc8051_golden_model_1.n1788 ;
  wire [7:0] \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [15:0] \oc8051_golden_model_1.n1794 ;
  wire \oc8051_golden_model_1.n1800 ;
  wire [7:0] \oc8051_golden_model_1.n1801 ;
  wire \oc8051_golden_model_1.n1804 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire \oc8051_golden_model_1.n1825 ;
  wire [7:0] \oc8051_golden_model_1.n1826 ;
  wire \oc8051_golden_model_1.n1831 ;
  wire [7:0] \oc8051_golden_model_1.n1832 ;
  wire \oc8051_golden_model_1.n1837 ;
  wire [7:0] \oc8051_golden_model_1.n1838 ;
  wire \oc8051_golden_model_1.n1843 ;
  wire [7:0] \oc8051_golden_model_1.n1844 ;
  wire \oc8051_golden_model_1.n1849 ;
  wire [7:0] \oc8051_golden_model_1.n1850 ;
  wire [7:0] \oc8051_golden_model_1.n1851 ;
  wire [3:0] \oc8051_golden_model_1.n1852 ;
  wire [7:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1889 ;
  wire \oc8051_golden_model_1.n1908 ;
  wire [7:0] \oc8051_golden_model_1.n1909 ;
  wire [7:0] \oc8051_golden_model_1.n1913 ;
  wire [3:0] \oc8051_golden_model_1.n1914 ;
  wire [7:0] \oc8051_golden_model_1.n1915 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff0 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff1 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff2 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff3 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not _44029_ (_43100_, rst);
  not _44030_ (_18190_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _44031_ (_18201_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _44032_ (_18212_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18201_);
  and _44033_ (_18223_, _18212_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _44034_ (_18234_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18201_);
  and _44035_ (_18245_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18201_);
  nor _44036_ (_18256_, _18245_, _18234_);
  and _44037_ (_18267_, _18256_, _18223_);
  nor _44038_ (_18278_, _18267_, _18190_);
  and _44039_ (_18289_, _18190_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _44040_ (_18300_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _44041_ (_18311_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18300_);
  nor _44042_ (_18322_, _18311_, _18289_);
  not _44043_ (_18333_, _18322_);
  and _44044_ (_18344_, _18333_, _18267_);
  or _44045_ (_18355_, _18344_, _18278_);
  and _44046_ (_22218_, _18355_, _43100_);
  nor _44047_ (_18376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _44048_ (_18387_, _18376_);
  and _44049_ (_18398_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and _44050_ (_18409_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _44051_ (_18420_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _44052_ (_18431_, _18420_);
  not _44053_ (_18442_, _18311_);
  nor _44054_ (_18453_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not _44055_ (_18464_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _44056_ (_18475_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _18464_);
  nor _44057_ (_18486_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not _44058_ (_18497_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor _44059_ (_18507_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _18497_);
  nor _44060_ (_18518_, _18507_, _18486_);
  nor _44061_ (_18529_, _18518_, _18475_);
  not _44062_ (_18540_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _44063_ (_18551_, _18475_, _18540_);
  nor _44064_ (_18562_, _18551_, _18529_);
  and _44065_ (_18573_, _18562_, _18453_);
  not _44066_ (_18584_, _18573_);
  and _44067_ (_18595_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44068_ (_18606_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _44069_ (_18617_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44070_ (_18628_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _18617_);
  and _44071_ (_18639_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _44072_ (_18650_, _18639_, _18606_);
  and _44073_ (_18671_, _18650_, _18584_);
  nor _44074_ (_18672_, _18671_, _18442_);
  not _44075_ (_18683_, _18289_);
  nor _44076_ (_18704_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor _44077_ (_18705_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _18497_);
  nor _44078_ (_18716_, _18705_, _18704_);
  nor _44079_ (_18737_, _18716_, _18475_);
  not _44080_ (_18738_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _44081_ (_18749_, _18475_, _18738_);
  nor _44082_ (_18770_, _18749_, _18737_);
  and _44083_ (_18771_, _18770_, _18453_);
  not _44084_ (_18782_, _18771_);
  and _44085_ (_18803_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _44086_ (_18804_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _44087_ (_18815_, _18804_, _18803_);
  and _44088_ (_18836_, _18815_, _18782_);
  nor _44089_ (_18837_, _18836_, _18683_);
  nor _44090_ (_18848_, _18837_, _18672_);
  nor _44091_ (_18868_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor _44092_ (_18869_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _18497_);
  nor _44093_ (_18880_, _18869_, _18868_);
  nor _44094_ (_18891_, _18880_, _18475_);
  not _44095_ (_18902_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _44096_ (_18913_, _18475_, _18902_);
  nor _44097_ (_18924_, _18913_, _18891_);
  and _44098_ (_18935_, _18924_, _18453_);
  not _44099_ (_18946_, _18935_);
  and _44100_ (_18957_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _44101_ (_18968_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _44102_ (_18979_, _18968_, _18957_);
  and _44103_ (_18990_, _18979_, _18946_);
  nor _44104_ (_19001_, _18990_, _18333_);
  nor _44105_ (_19012_, _19001_, _18376_);
  and _44106_ (_19023_, _19012_, _18848_);
  nor _44107_ (_19034_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor _44108_ (_19045_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _18497_);
  nor _44109_ (_19056_, _19045_, _19034_);
  nor _44110_ (_19067_, _19056_, _18475_);
  not _44111_ (_19078_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _44112_ (_19089_, _18475_, _19078_);
  nor _44113_ (_19100_, _19089_, _19067_);
  and _44114_ (_19111_, _19100_, _18453_);
  not _44115_ (_19122_, _19111_);
  and _44116_ (_19133_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _44117_ (_19144_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _44118_ (_19155_, _19144_, _19133_);
  and _44119_ (_19166_, _19155_, _19122_);
  and _44120_ (_19177_, _19166_, _18376_);
  nor _44121_ (_19188_, _19177_, _19023_);
  not _44122_ (_19199_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _44123_ (_19210_, _19199_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44124_ (_19220_, _19210_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44125_ (_19231_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _44126_ (_19242_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44127_ (_19253_, _19242_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44128_ (_19264_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _44129_ (_19275_, _19264_, _19231_);
  nor _44130_ (_19286_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44131_ (_19296_, _19286_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _44132_ (_19307_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not _44133_ (_19318_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44134_ (_19329_, _19210_, _19318_);
  and _44135_ (_19340_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _44136_ (_19351_, _19340_, _19307_);
  and _44137_ (_19362_, _19351_, _19275_);
  and _44138_ (_19373_, _19286_, _19199_);
  and _44139_ (_19383_, _19373_, _19100_);
  and _44140_ (_19394_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44141_ (_19405_, _19394_, _19318_);
  and _44142_ (_19416_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _44143_ (_19427_, _19394_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44144_ (_19438_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor _44145_ (_19449_, _19438_, _19416_);
  not _44146_ (_19460_, _19449_);
  nor _44147_ (_19470_, _19460_, _19383_);
  and _44148_ (_19481_, _19470_, _19362_);
  not _44149_ (_19492_, _19481_);
  and _44150_ (_19503_, _19492_, _19188_);
  not _44151_ (_19514_, _19503_);
  nor _44152_ (_19525_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor _44153_ (_19536_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _18497_);
  nor _44154_ (_19547_, _19536_, _19525_);
  nor _44155_ (_19557_, _19547_, _18475_);
  not _44156_ (_19568_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _44157_ (_19579_, _18475_, _19568_);
  nor _44158_ (_19590_, _19579_, _19557_);
  and _44159_ (_19601_, _19590_, _18453_);
  not _44160_ (_19612_, _19601_);
  and _44161_ (_19623_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _44162_ (_19634_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _44163_ (_19644_, _19634_, _19623_);
  and _44164_ (_19655_, _19644_, _19612_);
  nor _44165_ (_19666_, _19655_, _18442_);
  nor _44166_ (_19677_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor _44167_ (_19688_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _18497_);
  nor _44168_ (_19699_, _19688_, _19677_);
  nor _44169_ (_19710_, _19699_, _18475_);
  not _44170_ (_19720_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _44171_ (_19731_, _18475_, _19720_);
  nor _44172_ (_19742_, _19731_, _19710_);
  and _44173_ (_19753_, _19742_, _18453_);
  not _44174_ (_19764_, _19753_);
  and _44175_ (_19775_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _44176_ (_19786_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44177_ (_19797_, _19786_, _19775_);
  and _44178_ (_19807_, _19797_, _19764_);
  nor _44179_ (_19818_, _19807_, _18683_);
  nor _44180_ (_19829_, _19818_, _19666_);
  nor _44181_ (_19840_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor _44182_ (_19862_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _18497_);
  nor _44183_ (_19874_, _19862_, _19840_);
  nor _44184_ (_19885_, _19874_, _18475_);
  not _44185_ (_19897_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _44186_ (_19909_, _18475_, _19897_);
  nor _44187_ (_19921_, _19909_, _19885_);
  and _44188_ (_19933_, _19921_, _18453_);
  not _44189_ (_19934_, _19933_);
  and _44190_ (_19945_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _44191_ (_19956_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44192_ (_19967_, _19956_, _19945_);
  and _44193_ (_19977_, _19967_, _19934_);
  nor _44194_ (_19988_, _19977_, _18333_);
  nor _44195_ (_19999_, _19988_, _18376_);
  and _44196_ (_20010_, _19999_, _19829_);
  nor _44197_ (_20021_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor _44198_ (_20032_, _18497_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor _44199_ (_20043_, _20032_, _20021_);
  nor _44200_ (_20054_, _20043_, _18475_);
  not _44201_ (_20064_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _44202_ (_20075_, _18475_, _20064_);
  nor _44203_ (_20086_, _20075_, _20054_);
  and _44204_ (_20097_, _20086_, _18453_);
  not _44205_ (_20108_, _20097_);
  and _44206_ (_20119_, _18595_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _44207_ (_20130_, _18628_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _44208_ (_20141_, _20130_, _20119_);
  and _44209_ (_20151_, _20141_, _20108_);
  and _44210_ (_20162_, _20151_, _18376_);
  nor _44211_ (_20173_, _20162_, _20010_);
  and _44212_ (_20184_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _44213_ (_20195_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _44214_ (_20206_, _20195_, _20184_);
  and _44215_ (_20217_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _44216_ (_20227_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _44217_ (_20238_, _20227_, _20217_);
  and _44218_ (_20249_, _20238_, _20206_);
  and _44219_ (_20260_, _20086_, _19373_);
  and _44220_ (_20271_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _44221_ (_20282_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _44222_ (_20293_, _20282_, _20271_);
  not _44223_ (_20304_, _20293_);
  nor _44224_ (_20314_, _20304_, _20260_);
  and _44225_ (_20325_, _20314_, _20249_);
  not _44226_ (_20336_, _20325_);
  and _44227_ (_20347_, _20336_, _20173_);
  and _44228_ (_20358_, _20347_, _19514_);
  not _44229_ (_20369_, _20358_);
  and _44230_ (_20380_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _44231_ (_20391_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _44232_ (_20401_, _20391_, _20380_);
  and _44233_ (_20412_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _44234_ (_20423_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _44235_ (_20434_, _20423_, _20412_);
  and _44236_ (_20445_, _20434_, _20401_);
  and _44237_ (_20456_, _19742_, _19373_);
  and _44238_ (_20467_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _44239_ (_20478_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44240_ (_20488_, _20478_, _20467_);
  not _44241_ (_20499_, _20488_);
  nor _44242_ (_20510_, _20499_, _20456_);
  and _44243_ (_20521_, _20510_, _20445_);
  not _44244_ (_20532_, _20521_);
  and _44245_ (_20543_, _20532_, _20173_);
  and _44246_ (_20554_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _44247_ (_20565_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _44248_ (_20575_, _20565_, _20554_);
  and _44249_ (_20586_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _44250_ (_20597_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _44251_ (_20608_, _20597_, _20586_);
  and _44252_ (_20619_, _20608_, _20575_);
  and _44253_ (_20630_, _19373_, _18770_);
  and _44254_ (_20641_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _44255_ (_20652_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _44256_ (_20663_, _20652_, _20641_);
  not _44257_ (_20673_, _20663_);
  nor _44258_ (_20684_, _20673_, _20630_);
  and _44259_ (_20695_, _20684_, _20619_);
  not _44260_ (_20706_, _20695_);
  and _44261_ (_20717_, _20706_, _19188_);
  and _44262_ (_20728_, _20543_, _20717_);
  and _44263_ (_20739_, _19492_, _20728_);
  nor _44264_ (_20750_, _19503_, _20728_);
  nor _44265_ (_20770_, _20750_, _20739_);
  and _44266_ (_20781_, _20770_, _20543_);
  and _44267_ (_20782_, _20347_, _19503_);
  and _44268_ (_20793_, _19492_, _20173_);
  and _44269_ (_20814_, _20336_, _19188_);
  nor _44270_ (_20825_, _20814_, _20793_);
  nor _44271_ (_20826_, _20825_, _20782_);
  and _44272_ (_20847_, _20826_, _20781_);
  nor _44273_ (_20857_, _20826_, _20781_);
  nor _44274_ (_20858_, _20857_, _20847_);
  and _44275_ (_20869_, _20858_, _20739_);
  nor _44276_ (_20880_, _20869_, _20847_);
  nor _44277_ (_20891_, _20880_, _20369_);
  and _44278_ (_20912_, _20173_, _20706_);
  and _44279_ (_20913_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _44280_ (_20924_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _44281_ (_20935_, _20924_, _20913_);
  and _44282_ (_20945_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _44283_ (_20956_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _44284_ (_20967_, _20956_, _20945_);
  and _44285_ (_20978_, _20967_, _20935_);
  and _44286_ (_20989_, _19590_, _19373_);
  and _44287_ (_21000_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _44288_ (_21011_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor _44289_ (_21022_, _21011_, _21000_);
  not _44290_ (_21042_, _21022_);
  nor _44291_ (_21043_, _21042_, _20989_);
  and _44292_ (_21054_, _21043_, _20978_);
  not _44293_ (_21065_, _21054_);
  and _44294_ (_21076_, _21065_, _19188_);
  and _44295_ (_21087_, _21076_, _20912_);
  and _44296_ (_21098_, _20532_, _19188_);
  nor _44297_ (_21109_, _21098_, _20912_);
  nor _44298_ (_21120_, _21109_, _20728_);
  and _44299_ (_21130_, _21120_, _21087_);
  nor _44300_ (_21141_, _19503_, _20543_);
  nor _44301_ (_21152_, _21141_, _20781_);
  and _44302_ (_21163_, _21152_, _21130_);
  nor _44303_ (_21174_, _20858_, _20739_);
  nor _44304_ (_21185_, _21174_, _20869_);
  and _44305_ (_21196_, _21185_, _21163_);
  nor _44306_ (_21216_, _21185_, _21163_);
  nor _44307_ (_21217_, _21216_, _21196_);
  not _44308_ (_21228_, _21217_);
  and _44309_ (_21239_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _44310_ (_21250_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _44311_ (_21261_, _21250_, _21239_);
  and _44312_ (_21272_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and _44313_ (_21283_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor _44314_ (_21294_, _21283_, _21272_);
  and _44315_ (_21305_, _21294_, _21261_);
  and _44316_ (_21315_, _19921_, _19373_);
  and _44317_ (_21326_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _44318_ (_21337_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44319_ (_21348_, _21337_, _21326_);
  not _44320_ (_21359_, _21348_);
  nor _44321_ (_21370_, _21359_, _21315_);
  and _44322_ (_21381_, _21370_, _21305_);
  not _44323_ (_21392_, _21381_);
  and _44324_ (_21412_, _21392_, _20173_);
  and _44325_ (_21413_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _44326_ (_21424_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _44327_ (_21435_, _21424_, _21413_);
  and _44328_ (_21446_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _44329_ (_21457_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor _44330_ (_21468_, _21457_, _21446_);
  and _44331_ (_21479_, _21468_, _21435_);
  and _44332_ (_21490_, _19373_, _18562_);
  and _44333_ (_21500_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _44334_ (_21511_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor _44335_ (_21522_, _21511_, _21500_);
  not _44336_ (_21533_, _21522_);
  nor _44337_ (_21544_, _21533_, _21490_);
  and _44338_ (_21555_, _21544_, _21479_);
  not _44339_ (_21566_, _21555_);
  and _44340_ (_21577_, _21566_, _19188_);
  and _44341_ (_21588_, _21577_, _21412_);
  and _44342_ (_21598_, _21392_, _19188_);
  not _44343_ (_21609_, _21598_);
  and _44344_ (_21620_, _21566_, _20173_);
  and _44345_ (_21631_, _21620_, _21609_);
  and _44346_ (_21642_, _21631_, _21076_);
  nor _44347_ (_21653_, _21642_, _21588_);
  and _44348_ (_21664_, _21065_, _20173_);
  nor _44349_ (_21675_, _21664_, _20717_);
  nor _44350_ (_21685_, _21675_, _21087_);
  not _44351_ (_21696_, _21685_);
  nor _44352_ (_21707_, _21696_, _21653_);
  nor _44353_ (_21718_, _21120_, _21087_);
  nor _44354_ (_21729_, _21718_, _21130_);
  and _44355_ (_21740_, _21729_, _21707_);
  nor _44356_ (_21760_, _21152_, _21130_);
  nor _44357_ (_21761_, _21760_, _21163_);
  and _44358_ (_21772_, _21761_, _21740_);
  and _44359_ (_21783_, _19220_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _44360_ (_21794_, _19253_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _44361_ (_21805_, _21794_, _21783_);
  and _44362_ (_21816_, _19296_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _44363_ (_21827_, _19329_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _44364_ (_21838_, _21827_, _21816_);
  and _44365_ (_21848_, _21838_, _21805_);
  and _44366_ (_21869_, _19373_, _18924_);
  and _44367_ (_21870_, _19427_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and _44368_ (_21881_, _19405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _44369_ (_21892_, _21881_, _21870_);
  not _44370_ (_21903_, _21892_);
  nor _44371_ (_21914_, _21903_, _21869_);
  and _44372_ (_21925_, _21914_, _21848_);
  not _44373_ (_21935_, _21925_);
  and _44374_ (_21946_, _21935_, _20173_);
  and _44375_ (_21957_, _21946_, _21598_);
  nor _44376_ (_21968_, _21577_, _21412_);
  nor _44377_ (_21979_, _21968_, _21588_);
  and _44378_ (_21990_, _21979_, _21957_);
  nor _44379_ (_22001_, _21631_, _21076_);
  nor _44380_ (_22012_, _22001_, _21642_);
  and _44381_ (_22022_, _22012_, _21990_);
  and _44382_ (_22033_, _21696_, _21653_);
  nor _44383_ (_22044_, _22033_, _21707_);
  and _44384_ (_22055_, _22044_, _22022_);
  nor _44385_ (_22066_, _21729_, _21707_);
  nor _44386_ (_22077_, _22066_, _21740_);
  and _44387_ (_22088_, _22077_, _22055_);
  nor _44388_ (_22098_, _21761_, _21740_);
  nor _44389_ (_22109_, _22098_, _21772_);
  and _44390_ (_22120_, _22109_, _22088_);
  nor _44391_ (_22131_, _22120_, _21772_);
  nor _44392_ (_22142_, _22131_, _21228_);
  nor _44393_ (_22153_, _22142_, _21196_);
  and _44394_ (_22164_, _20880_, _20369_);
  nor _44395_ (_22175_, _22164_, _20891_);
  not _44396_ (_22185_, _22175_);
  nor _44397_ (_22196_, _22185_, _22153_);
  or _44398_ (_22207_, _22196_, _20782_);
  nor _44399_ (_22219_, _22207_, _20891_);
  nor _44400_ (_22230_, _22219_, _18431_);
  and _44401_ (_22241_, _22219_, _18431_);
  nor _44402_ (_22252_, _22241_, _22230_);
  not _44403_ (_22263_, _22252_);
  and _44404_ (_22273_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and _44405_ (_22284_, _22185_, _22153_);
  nor _44406_ (_22295_, _22284_, _22196_);
  and _44407_ (_22316_, _22295_, _22273_);
  and _44408_ (_22317_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and _44409_ (_22328_, _22131_, _21228_);
  nor _44410_ (_22339_, _22328_, _22142_);
  and _44411_ (_22349_, _22339_, _22317_);
  nor _44412_ (_22360_, _22339_, _22317_);
  nor _44413_ (_22371_, _22360_, _22349_);
  not _44414_ (_22382_, _22371_);
  and _44415_ (_22393_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor _44416_ (_22404_, _22109_, _22088_);
  nor _44417_ (_22415_, _22404_, _22120_);
  and _44418_ (_22426_, _22415_, _22393_);
  nor _44419_ (_22436_, _22415_, _22393_);
  nor _44420_ (_22447_, _22436_, _22426_);
  not _44421_ (_22458_, _22447_);
  and _44422_ (_22469_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor _44423_ (_22480_, _22077_, _22055_);
  nor _44424_ (_22491_, _22480_, _22088_);
  and _44425_ (_22502_, _22491_, _22469_);
  nor _44426_ (_22513_, _22491_, _22469_);
  nor _44427_ (_22523_, _22513_, _22502_);
  not _44428_ (_22534_, _22523_);
  and _44429_ (_22545_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor _44430_ (_22556_, _22044_, _22022_);
  nor _44431_ (_22567_, _22556_, _22055_);
  and _44432_ (_22578_, _22567_, _22545_);
  and _44433_ (_22589_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor _44434_ (_22609_, _22012_, _21990_);
  nor _44435_ (_22610_, _22609_, _22022_);
  and _44436_ (_22621_, _22610_, _22589_);
  and _44437_ (_22632_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor _44438_ (_22643_, _21979_, _21957_);
  nor _44439_ (_22654_, _22643_, _21990_);
  and _44440_ (_22665_, _22654_, _22632_);
  nor _44441_ (_22676_, _22610_, _22589_);
  nor _44442_ (_22686_, _22676_, _22621_);
  and _44443_ (_22697_, _22686_, _22665_);
  nor _44444_ (_22718_, _22697_, _22621_);
  not _44445_ (_22719_, _22718_);
  nor _44446_ (_22730_, _22567_, _22545_);
  nor _44447_ (_22741_, _22730_, _22578_);
  and _44448_ (_22752_, _22741_, _22719_);
  nor _44449_ (_22763_, _22752_, _22578_);
  nor _44450_ (_22773_, _22763_, _22534_);
  nor _44451_ (_22784_, _22773_, _22502_);
  nor _44452_ (_22795_, _22784_, _22458_);
  nor _44453_ (_22806_, _22795_, _22426_);
  nor _44454_ (_22817_, _22806_, _22382_);
  nor _44455_ (_22828_, _22817_, _22349_);
  nor _44456_ (_22839_, _22295_, _22273_);
  nor _44457_ (_22850_, _22839_, _22316_);
  not _44458_ (_22860_, _22850_);
  nor _44459_ (_22871_, _22860_, _22828_);
  nor _44460_ (_22882_, _22871_, _22316_);
  nor _44461_ (_22893_, _22882_, _22263_);
  nor _44462_ (_22904_, _22893_, _22230_);
  not _44463_ (_22915_, _22904_);
  and _44464_ (_22936_, _22915_, _18409_);
  and _44465_ (_22937_, _22936_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _44466_ (_22948_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _44467_ (_22958_, _22948_, _22937_);
  and _44468_ (_22969_, _22958_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _44469_ (_22980_, _22969_, _18398_);
  not _44470_ (_22991_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _44471_ (_23002_, _18376_, _22991_);
  or _44472_ (_23013_, _23002_, _22980_);
  nand _44473_ (_23024_, _22980_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and _44474_ (_23035_, _23024_, _23013_);
  and _44475_ (_24376_, _23035_, _43100_);
  nor _44476_ (_23056_, _18267_, _18300_);
  and _44477_ (_23066_, _18267_, _18300_);
  or _44478_ (_23077_, _23066_, _23056_);
  and _44479_ (_02359_, _23077_, _43100_);
  and _44480_ (_23098_, _21935_, _19188_);
  and _44481_ (_02546_, _23098_, _43100_);
  nor _44482_ (_23119_, _21946_, _21598_);
  nor _44483_ (_23130_, _23119_, _21957_);
  and _44484_ (_02703_, _23130_, _43100_);
  nor _44485_ (_23151_, _22654_, _22632_);
  nor _44486_ (_23162_, _23151_, _22665_);
  and _44487_ (_02884_, _23162_, _43100_);
  nor _44488_ (_23192_, _22686_, _22665_);
  nor _44489_ (_23193_, _23192_, _22697_);
  and _44490_ (_03126_, _23193_, _43100_);
  nor _44491_ (_23214_, _22741_, _22719_);
  nor _44492_ (_23225_, _23214_, _22752_);
  and _44493_ (_03363_, _23225_, _43100_);
  and _44494_ (_23246_, _22763_, _22534_);
  nor _44495_ (_23257_, _23246_, _22773_);
  and _44496_ (_03564_, _23257_, _43100_);
  and _44497_ (_23277_, _22784_, _22458_);
  nor _44498_ (_23288_, _23277_, _22795_);
  and _44499_ (_03763_, _23288_, _43100_);
  and _44500_ (_23309_, _22806_, _22382_);
  nor _44501_ (_23320_, _23309_, _22817_);
  and _44502_ (_03958_, _23320_, _43100_);
  and _44503_ (_23341_, _22860_, _22828_);
  nor _44504_ (_23352_, _23341_, _22871_);
  and _44505_ (_04057_, _23352_, _43100_);
  and _44506_ (_23373_, _22882_, _22263_);
  nor _44507_ (_23384_, _23373_, _22893_);
  and _44508_ (_04156_, _23384_, _43100_);
  nor _44509_ (_23404_, _22915_, _18409_);
  nor _44510_ (_23415_, _23404_, _22936_);
  and _44511_ (_04250_, _23415_, _43100_);
  and _44512_ (_23436_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor _44513_ (_23447_, _23436_, _22936_);
  nor _44514_ (_23468_, _23447_, _22937_);
  and _44515_ (_04349_, _23468_, _43100_);
  nor _44516_ (_23479_, _22948_, _22937_);
  nor _44517_ (_23490_, _23479_, _22958_);
  and _44518_ (_04447_, _23490_, _43100_);
  and _44519_ (_23510_, _18387_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor _44520_ (_23521_, _23510_, _22958_);
  nor _44521_ (_23532_, _23521_, _22969_);
  and _44522_ (_04546_, _23532_, _43100_);
  nor _44523_ (_23553_, _22969_, _18398_);
  nor _44524_ (_23564_, _23553_, _22980_);
  and _44525_ (_04645_, _23564_, _43100_);
  and _44526_ (_23585_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18201_);
  nor _44527_ (_23596_, _23585_, _18212_);
  not _44528_ (_23606_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _44529_ (_23617_, _18234_, _23606_);
  and _44530_ (_23628_, _23617_, _23596_);
  and _44531_ (_23639_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _44532_ (_23650_, _23639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44533_ (_23661_, _23639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44534_ (_23672_, _23661_, _23650_);
  and _44535_ (_00927_, _23672_, _43100_);
  and _44536_ (_00957_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _43100_);
  not _44537_ (_23702_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _44538_ (_23713_, _19977_, _23702_);
  and _44539_ (_23724_, _19655_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44540_ (_23735_, _23724_, _23713_);
  nor _44541_ (_23746_, _23735_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44542_ (_23757_, _19807_, _23702_);
  and _44543_ (_23767_, _20151_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _44544_ (_23778_, _23767_, _23757_);
  and _44545_ (_23789_, _23778_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44546_ (_23800_, _23789_, _23746_);
  nor _44547_ (_23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44548_ (_23822_, _23811_, _20325_);
  nor _44549_ (_23833_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor _44550_ (_23844_, _23833_, _23822_);
  not _44551_ (_23854_, _23844_);
  and _44552_ (_23865_, _18990_, _23702_);
  and _44553_ (_23876_, _18671_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44554_ (_23897_, _23876_, _23865_);
  nor _44555_ (_23898_, _23897_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44556_ (_23909_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44557_ (_23920_, _18836_, _23702_);
  and _44558_ (_23930_, _19166_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44559_ (_23941_, _23930_, _23920_);
  nor _44560_ (_23952_, _23941_, _23909_);
  nor _44561_ (_23963_, _23952_, _23898_);
  nor _44562_ (_23974_, _23963_, _23854_);
  and _44563_ (_23985_, _23963_, _23854_);
  nor _44564_ (_23996_, _23985_, _23974_);
  and _44565_ (_24007_, _23811_, _19481_);
  nor _44566_ (_24017_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor _44567_ (_24028_, _24017_, _24007_);
  not _44568_ (_24039_, _24028_);
  nor _44569_ (_24050_, _19977_, _23702_);
  nor _44570_ (_24061_, _24050_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44571_ (_24082_, _19655_, _23702_);
  and _44572_ (_24083_, _19807_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44573_ (_24094_, _24083_, _24082_);
  nor _44574_ (_24104_, _24094_, _23909_);
  nor _44575_ (_24115_, _24104_, _24061_);
  nor _44576_ (_24126_, _24115_, _24039_);
  and _44577_ (_24137_, _24115_, _24039_);
  nor _44578_ (_24148_, _24137_, _24126_);
  not _44579_ (_24159_, _24148_);
  nor _44580_ (_24170_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and _44581_ (_24181_, _23811_, _20521_);
  nor _44582_ (_24191_, _24181_, _24170_);
  not _44583_ (_24202_, _24191_);
  nor _44584_ (_24213_, _18990_, _23702_);
  nor _44585_ (_24224_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44586_ (_24235_, _18671_, _23702_);
  and _44587_ (_24246_, _18836_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44588_ (_24257_, _24246_, _24235_);
  nor _44589_ (_24267_, _24257_, _23909_);
  nor _44590_ (_24278_, _24267_, _24224_);
  nor _44591_ (_24289_, _24278_, _24202_);
  and _44592_ (_24300_, _24278_, _24202_);
  and _44593_ (_24311_, _23735_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44594_ (_24322_, _24311_);
  nor _44595_ (_24333_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and _44596_ (_24344_, _23811_, _20695_);
  nor _44597_ (_24354_, _24344_, _24333_);
  and _44598_ (_24365_, _24354_, _24322_);
  and _44599_ (_24377_, _23897_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44600_ (_24388_, _24377_);
  and _44601_ (_24399_, _23811_, _21054_);
  nor _44602_ (_24410_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor _44603_ (_24421_, _24410_, _24399_);
  and _44604_ (_24431_, _24421_, _24388_);
  nor _44605_ (_24442_, _24421_, _24388_);
  nor _44606_ (_24453_, _24442_, _24431_);
  not _44607_ (_24464_, _24453_);
  and _44608_ (_24475_, _24050_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44609_ (_24486_, _24475_);
  and _44610_ (_24497_, _23811_, _21555_);
  nor _44611_ (_24508_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor _44612_ (_24518_, _24508_, _24497_);
  and _44613_ (_24529_, _24518_, _24486_);
  and _44614_ (_24540_, _24213_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44615_ (_24551_, _24540_);
  and _44616_ (_24562_, _23811_, _21381_);
  nor _44617_ (_24573_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  nor _44618_ (_24584_, _24573_, _24562_);
  nor _44619_ (_24595_, _24584_, _24551_);
  not _44620_ (_24615_, _24595_);
  nor _44621_ (_24616_, _24518_, _24486_);
  nor _44622_ (_24627_, _24616_, _24529_);
  and _44623_ (_24638_, _24627_, _24615_);
  nor _44624_ (_24649_, _24638_, _24529_);
  nor _44625_ (_24660_, _24649_, _24464_);
  nor _44626_ (_24671_, _24660_, _24431_);
  nor _44627_ (_24681_, _24354_, _24322_);
  nor _44628_ (_24692_, _24681_, _24365_);
  not _44629_ (_24703_, _24692_);
  nor _44630_ (_24714_, _24703_, _24671_);
  nor _44631_ (_24725_, _24714_, _24365_);
  nor _44632_ (_24736_, _24725_, _24300_);
  nor _44633_ (_24747_, _24736_, _24289_);
  nor _44634_ (_24758_, _24747_, _24159_);
  nor _44635_ (_24768_, _24758_, _24126_);
  not _44636_ (_24779_, _24768_);
  and _44637_ (_24790_, _24779_, _23996_);
  or _44638_ (_24801_, _24790_, _23974_);
  and _44639_ (_24812_, _20151_, _19166_);
  or _44640_ (_24823_, _24812_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _44641_ (_24834_, _23941_);
  and _44642_ (_24845_, _23778_, _24834_);
  nor _44643_ (_24856_, _24257_, _24094_);
  and _44644_ (_24867_, _24856_, _24845_);
  or _44645_ (_24878_, _24867_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44646_ (_24889_, _24878_, _24823_);
  and _44647_ (_24900_, _24889_, _24801_);
  and _44648_ (_24911_, _24900_, _23800_);
  nor _44649_ (_24922_, _24779_, _23996_);
  or _44650_ (_24933_, _24922_, _24790_);
  and _44651_ (_24944_, _24933_, _24911_);
  nor _44652_ (_24955_, _24911_, _23844_);
  nor _44653_ (_24966_, _24955_, _24944_);
  not _44654_ (_24977_, _24966_);
  and _44655_ (_24988_, _24966_, _23800_);
  not _44656_ (_24999_, _23963_);
  nor _44657_ (_25010_, _24911_, _24039_);
  and _44658_ (_25021_, _24747_, _24159_);
  nor _44659_ (_25031_, _25021_, _24758_);
  and _44660_ (_25042_, _25031_, _24911_);
  or _44661_ (_25053_, _25042_, _25010_);
  and _44662_ (_25064_, _25053_, _24999_);
  nor _44663_ (_25075_, _25053_, _24999_);
  nor _44664_ (_25086_, _25075_, _25064_);
  not _44665_ (_25097_, _25086_);
  not _44666_ (_25108_, _24115_);
  nor _44667_ (_25119_, _24911_, _24202_);
  nor _44668_ (_25130_, _24300_, _24289_);
  nor _44669_ (_25141_, _25130_, _24725_);
  and _44670_ (_25162_, _25130_, _24725_);
  or _44671_ (_25163_, _25162_, _25141_);
  and _44672_ (_25174_, _25163_, _24911_);
  or _44673_ (_25185_, _25174_, _25119_);
  and _44674_ (_25196_, _25185_, _25108_);
  nor _44675_ (_25207_, _25185_, _25108_);
  not _44676_ (_25218_, _24278_);
  and _44677_ (_25229_, _24703_, _24671_);
  or _44678_ (_25240_, _25229_, _24714_);
  and _44679_ (_25251_, _25240_, _24911_);
  nor _44680_ (_25262_, _24911_, _24354_);
  nor _44681_ (_25273_, _25262_, _25251_);
  and _44682_ (_25284_, _25273_, _25218_);
  and _44683_ (_25295_, _24649_, _24464_);
  nor _44684_ (_25306_, _25295_, _24660_);
  not _44685_ (_25317_, _25306_);
  and _44686_ (_25328_, _25317_, _24911_);
  nor _44687_ (_25339_, _24911_, _24421_);
  nor _44688_ (_25350_, _25339_, _25328_);
  and _44689_ (_25361_, _25350_, _24322_);
  nor _44690_ (_25372_, _25350_, _24322_);
  nor _44691_ (_25383_, _25372_, _25361_);
  not _44692_ (_25394_, _25383_);
  nor _44693_ (_25404_, _24627_, _24615_);
  nor _44694_ (_25425_, _25404_, _24638_);
  not _44695_ (_25426_, _25425_);
  and _44696_ (_25437_, _25426_, _24911_);
  nor _44697_ (_25448_, _24911_, _24518_);
  nor _44698_ (_25459_, _25448_, _25437_);
  and _44699_ (_25470_, _25459_, _24388_);
  and _44700_ (_25481_, _24911_, _24540_);
  nor _44701_ (_25492_, _25481_, _24584_);
  and _44702_ (_25503_, _25481_, _24584_);
  nor _44703_ (_25514_, _25503_, _25492_);
  and _44704_ (_25525_, _25514_, _24486_);
  nor _44705_ (_25536_, _25514_, _24486_);
  nor _44706_ (_25547_, _25536_, _25525_);
  and _44707_ (_25558_, _23811_, _21925_);
  nor _44708_ (_25569_, _23811_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _44709_ (_25580_, _25569_, _25558_);
  nor _44710_ (_25591_, _25580_, _24551_);
  not _44711_ (_25602_, _25591_);
  and _44712_ (_25613_, _25602_, _25547_);
  nor _44713_ (_25624_, _25613_, _25525_);
  nor _44714_ (_25635_, _25459_, _24388_);
  nor _44715_ (_25646_, _25635_, _25470_);
  not _44716_ (_25657_, _25646_);
  nor _44717_ (_25668_, _25657_, _25624_);
  nor _44718_ (_25679_, _25668_, _25470_);
  nor _44719_ (_25690_, _25679_, _25394_);
  nor _44720_ (_25701_, _25690_, _25361_);
  nor _44721_ (_25712_, _25273_, _25218_);
  nor _44722_ (_25733_, _25712_, _25284_);
  not _44723_ (_25734_, _25733_);
  nor _44724_ (_25745_, _25734_, _25701_);
  nor _44725_ (_25755_, _25745_, _25284_);
  nor _44726_ (_25766_, _25755_, _25207_);
  nor _44727_ (_25777_, _25766_, _25196_);
  nor _44728_ (_25788_, _25777_, _25097_);
  or _44729_ (_25799_, _25788_, _25064_);
  or _44730_ (_25810_, _25799_, _24988_);
  and _44731_ (_25821_, _25810_, _24889_);
  nor _44732_ (_25832_, _25821_, _24977_);
  and _44733_ (_25843_, _24988_, _24889_);
  and _44734_ (_25854_, _25843_, _25799_);
  or _44735_ (_25865_, _25854_, _25832_);
  and _44736_ (_00976_, _25865_, _43100_);
  or _44737_ (_25886_, _24966_, _23800_);
  and _44738_ (_25897_, _25886_, _25821_);
  and _44739_ (_02839_, _25897_, _43100_);
  and _44740_ (_02851_, _24911_, _43100_);
  and _44741_ (_02873_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _43100_);
  and _44742_ (_02897_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _43100_);
  and _44743_ (_02919_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _43100_);
  or _44744_ (_25958_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44745_ (_25969_, _23639_, rst);
  and _44746_ (_02931_, _25969_, _25958_);
  and _44747_ (_25990_, _25897_, _24540_);
  or _44748_ (_26001_, _25990_, _25580_);
  nand _44749_ (_26012_, _25990_, _25580_);
  and _44750_ (_26023_, _26012_, _26001_);
  and _44751_ (_02944_, _26023_, _43100_);
  nor _44752_ (_26054_, _25602_, _25547_);
  or _44753_ (_26055_, _26054_, _25613_);
  nand _44754_ (_26066_, _26055_, _25897_);
  or _44755_ (_26077_, _25897_, _25514_);
  and _44756_ (_26088_, _26077_, _26066_);
  and _44757_ (_02957_, _26088_, _43100_);
  and _44758_ (_26108_, _25657_, _25624_);
  or _44759_ (_26119_, _26108_, _25668_);
  nand _44760_ (_26130_, _26119_, _25897_);
  or _44761_ (_26141_, _25897_, _25459_);
  and _44762_ (_26152_, _26141_, _26130_);
  and _44763_ (_02969_, _26152_, _43100_);
  and _44764_ (_26173_, _25679_, _25394_);
  or _44765_ (_26184_, _26173_, _25690_);
  nand _44766_ (_26195_, _26184_, _25897_);
  or _44767_ (_26206_, _25897_, _25350_);
  and _44768_ (_26217_, _26206_, _26195_);
  and _44769_ (_02980_, _26217_, _43100_);
  and _44770_ (_26238_, _25734_, _25701_);
  or _44771_ (_26249_, _26238_, _25745_);
  nand _44772_ (_26260_, _26249_, _25897_);
  or _44773_ (_26271_, _25897_, _25273_);
  and _44774_ (_26282_, _26271_, _26260_);
  and _44775_ (_02994_, _26282_, _43100_);
  or _44776_ (_26303_, _25207_, _25196_);
  and _44777_ (_26314_, _26303_, _25755_);
  nor _44778_ (_26325_, _26303_, _25755_);
  or _44779_ (_26336_, _26325_, _26314_);
  nand _44780_ (_26347_, _26336_, _25897_);
  or _44781_ (_26358_, _25897_, _25185_);
  and _44782_ (_26369_, _26358_, _26347_);
  and _44783_ (_03006_, _26369_, _43100_);
  and _44784_ (_26390_, _25777_, _25097_);
  or _44785_ (_26401_, _26390_, _25788_);
  nand _44786_ (_26412_, _26401_, _25897_);
  or _44787_ (_26423_, _25897_, _25053_);
  and _44788_ (_26433_, _26423_, _26412_);
  and _44789_ (_03020_, _26433_, _43100_);
  not _44790_ (_26454_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44791_ (_26465_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18201_);
  and _44792_ (_26476_, _26465_, _26454_);
  and _44793_ (_26487_, _26476_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _44794_ (_26498_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44795_ (_26509_, _26498_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44796_ (_26530_, _26498_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44797_ (_26531_, _26530_, _26509_);
  and _44798_ (_26542_, _26531_, _26487_);
  not _44799_ (_26553_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _44800_ (_26564_, _26476_, _26553_);
  and _44801_ (_26575_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _44802_ (_26586_, _26575_, _26542_);
  not _44803_ (_26597_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _44804_ (_26608_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18201_);
  and _44805_ (_26619_, _26608_, _26597_);
  and _44806_ (_26630_, _26619_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44807_ (_26641_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _44808_ (_26652_, _26619_, _26454_);
  and _44809_ (_26663_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or _44810_ (_26674_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44811_ (_26685_, _26674_, _18201_);
  nor _44812_ (_26696_, _26685_, _26608_);
  and _44813_ (_26707_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _44814_ (_26718_, _26707_, _26663_);
  nor _44815_ (_26729_, _26718_, _26641_);
  and _44816_ (_26740_, _26729_, _26586_);
  and _44817_ (_26761_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor _44818_ (_26762_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _44819_ (_26773_, _26762_, _26498_);
  and _44820_ (_26784_, _26773_, _26487_);
  nor _44821_ (_26794_, _26784_, _26761_);
  and _44822_ (_26805_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and _44823_ (_26816_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and _44824_ (_26827_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or _44825_ (_26838_, _26827_, _26816_);
  nor _44826_ (_26849_, _26838_, _26805_);
  and _44827_ (_26860_, _26849_, _26794_);
  and _44828_ (_26871_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and _44829_ (_26882_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _44830_ (_26893_, _26882_, _26871_);
  and _44831_ (_26904_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not _44832_ (_26915_, _26904_);
  not _44833_ (_26926_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44834_ (_26937_, _26487_, _26926_);
  and _44835_ (_26948_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _44836_ (_26959_, _26948_, _26937_);
  and _44837_ (_26970_, _26959_, _26915_);
  and _44838_ (_26981_, _26970_, _26893_);
  and _44839_ (_26992_, _26981_, _26860_);
  and _44840_ (_27003_, _26992_, _26740_);
  and _44841_ (_27014_, _26509_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _44842_ (_27025_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _44843_ (_27036_, _27025_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _44844_ (_27047_, _27036_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _44845_ (_27058_, _27047_);
  not _44846_ (_27069_, _26487_);
  nor _44847_ (_27080_, _27036_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _44848_ (_27091_, _27080_, _27069_);
  and _44849_ (_27102_, _27091_, _27058_);
  not _44850_ (_27113_, _27102_);
  and _44851_ (_27124_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44852_ (_27134_, _27124_, _26465_);
  and _44853_ (_27145_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _44854_ (_27156_, _27145_, _27134_);
  and _44855_ (_27167_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _44856_ (_27178_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _44857_ (_27189_, _27178_, _27167_);
  and _44858_ (_27200_, _27189_, _27156_);
  and _44859_ (_27211_, _27200_, _27113_);
  nor _44860_ (_27222_, _27025_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _44861_ (_27233_, _27222_);
  nor _44862_ (_27244_, _27036_, _27069_);
  and _44863_ (_27255_, _27244_, _27233_);
  not _44864_ (_27266_, _27255_);
  and _44865_ (_27277_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _44866_ (_27288_, _27277_, _27134_);
  and _44867_ (_27299_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _44868_ (_27310_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _44869_ (_27321_, _27310_, _27299_);
  and _44870_ (_27342_, _27321_, _27288_);
  and _44871_ (_27343_, _27342_, _27266_);
  nor _44872_ (_27354_, _27343_, _27211_);
  not _44873_ (_27365_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _44874_ (_27376_, _27047_, _27365_);
  and _44875_ (_27387_, _27047_, _27365_);
  nor _44876_ (_27398_, _27387_, _27376_);
  nor _44877_ (_27409_, _27398_, _27069_);
  not _44878_ (_27420_, _27409_);
  and _44879_ (_27431_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor _44880_ (_27442_, _27431_, _27134_);
  and _44881_ (_27453_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _44882_ (_27464_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor _44883_ (_27475_, _27464_, _27453_);
  and _44884_ (_27485_, _27475_, _27442_);
  and _44885_ (_27496_, _27485_, _27420_);
  not _44886_ (_27507_, _27496_);
  and _44887_ (_27518_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _44888_ (_27529_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _44889_ (_27540_, _27529_, _27518_);
  not _44890_ (_27551_, _27014_);
  nor _44891_ (_27562_, _26509_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _44892_ (_27573_, _27562_, _27069_);
  and _44893_ (_27584_, _27573_, _27551_);
  and _44894_ (_27595_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _44895_ (_27606_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _44896_ (_27617_, _27606_, _27595_);
  not _44897_ (_27628_, _27617_);
  nor _44898_ (_27639_, _27628_, _27584_);
  and _44899_ (_27650_, _27639_, _27540_);
  not _44900_ (_27661_, _27650_);
  and _44901_ (_27672_, _26564_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _44902_ (_27683_, _27672_, _27134_);
  and _44903_ (_27694_, _26630_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not _44904_ (_27705_, _27694_);
  and _44905_ (_27716_, _27705_, _27683_);
  nor _44906_ (_27727_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _44907_ (_27738_, _27727_);
  nor _44908_ (_27749_, _27025_, _27069_);
  and _44909_ (_27760_, _27749_, _27738_);
  and _44910_ (_27771_, _26652_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and _44911_ (_27782_, _26696_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor _44912_ (_27793_, _27782_, _27771_);
  not _44913_ (_27804_, _27793_);
  nor _44914_ (_27814_, _27804_, _27760_);
  and _44915_ (_27825_, _27814_, _27716_);
  nor _44916_ (_27836_, _27825_, _27661_);
  and _44917_ (_27847_, _27836_, _27507_);
  and _44918_ (_27858_, _27847_, _27354_);
  nand _44919_ (_27869_, _27858_, _27003_);
  and _44920_ (_27880_, _25865_, _23628_);
  not _44921_ (_27891_, _27880_);
  and _44922_ (_27902_, _23035_, _18267_);
  not _44923_ (_27913_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _44924_ (_27924_, _18212_, _27913_);
  and _44925_ (_27935_, _27924_, _18256_);
  not _44926_ (_27946_, _27935_);
  nor _44927_ (_27957_, _20325_, _20151_);
  and _44928_ (_27978_, _20325_, _20151_);
  nor _44929_ (_27979_, _27978_, _27957_);
  not _44930_ (_27990_, _19166_);
  nor _44931_ (_28001_, _19481_, _27990_);
  nor _44932_ (_28012_, _19481_, _19166_);
  and _44933_ (_28023_, _19481_, _19166_);
  nor _44934_ (_28034_, _28023_, _28012_);
  not _44935_ (_28045_, _19807_);
  nor _44936_ (_28056_, _20521_, _28045_);
  nor _44937_ (_28067_, _20521_, _19807_);
  and _44938_ (_28078_, _20521_, _19807_);
  nor _44939_ (_28089_, _28078_, _28067_);
  not _44940_ (_28100_, _18836_);
  and _44941_ (_28111_, _20695_, _28100_);
  nor _44942_ (_28122_, _28111_, _28089_);
  nor _44943_ (_28132_, _28122_, _28056_);
  nor _44944_ (_28143_, _28132_, _28034_);
  nor _44945_ (_28154_, _28143_, _28001_);
  and _44946_ (_28165_, _28132_, _28034_);
  nor _44947_ (_28176_, _28165_, _28143_);
  not _44948_ (_28187_, _28176_);
  and _44949_ (_28198_, _28111_, _28089_);
  nor _44950_ (_28209_, _28198_, _28122_);
  not _44951_ (_28220_, _28209_);
  nor _44952_ (_28231_, _20695_, _18836_);
  and _44953_ (_28242_, _20695_, _18836_);
  nor _44954_ (_28253_, _28242_, _28231_);
  not _44955_ (_28264_, _28253_);
  and _44956_ (_28285_, _21054_, _19655_);
  nor _44957_ (_28286_, _21054_, _19655_);
  nor _44958_ (_28297_, _28286_, _28285_);
  nor _44959_ (_28308_, _21555_, _18671_);
  and _44960_ (_28319_, _21555_, _18671_);
  nor _44961_ (_28330_, _28319_, _28308_);
  nor _44962_ (_28341_, _21381_, _19977_);
  and _44963_ (_28352_, _21381_, _19977_);
  nor _44964_ (_28363_, _28352_, _28341_);
  not _44965_ (_28374_, _18990_);
  and _44966_ (_28385_, _21925_, _28374_);
  nor _44967_ (_28396_, _28385_, _28363_);
  not _44968_ (_28407_, _19977_);
  nor _44969_ (_28418_, _21381_, _28407_);
  nor _44970_ (_28429_, _28418_, _28396_);
  nor _44971_ (_28440_, _28429_, _28330_);
  not _44972_ (_28450_, _18671_);
  nor _44973_ (_28461_, _21555_, _28450_);
  nor _44974_ (_28472_, _28461_, _28440_);
  nor _44975_ (_28483_, _28472_, _28297_);
  and _44976_ (_28494_, _28472_, _28297_);
  nor _44977_ (_28505_, _28494_, _28483_);
  not _44978_ (_28516_, _28505_);
  and _44979_ (_28527_, _28429_, _28330_);
  nor _44980_ (_28538_, _28527_, _28440_);
  not _44981_ (_28549_, _28538_);
  and _44982_ (_28560_, _28385_, _28363_);
  nor _44983_ (_28571_, _28560_, _28396_);
  not _44984_ (_28582_, _28571_);
  nor _44985_ (_28593_, _21925_, _18990_);
  and _44986_ (_28604_, _21925_, _18990_);
  nor _44987_ (_28615_, _28604_, _28593_);
  not _44988_ (_28636_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _44989_ (_28637_, _18475_, _28636_);
  not _44990_ (_28648_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _44991_ (_28659_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44992_ (_28670_, _28659_, _20043_);
  nor _44993_ (_28681_, _28670_, _28648_);
  nor _44994_ (_28692_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44995_ (_28703_, _28692_, _18716_);
  not _44996_ (_28714_, _28703_);
  not _44997_ (_28725_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44998_ (_28736_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _28725_);
  and _44999_ (_28746_, _28736_, _19699_);
  not _45000_ (_28757_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _45001_ (_28768_, _28757_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45002_ (_28779_, _28768_, _19056_);
  nor _45003_ (_28790_, _28779_, _28746_);
  and _45004_ (_28801_, _28790_, _28714_);
  and _45005_ (_28812_, _28801_, _28681_);
  and _45006_ (_28823_, _28659_, _19547_);
  nor _45007_ (_28834_, _28823_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _45008_ (_28845_, _28768_, _18518_);
  not _45009_ (_28856_, _28845_);
  and _45010_ (_28867_, _28736_, _19874_);
  and _45011_ (_28878_, _28692_, _18880_);
  nor _45012_ (_28889_, _28878_, _28867_);
  and _45013_ (_28900_, _28889_, _28856_);
  and _45014_ (_28911_, _28900_, _28834_);
  nor _45015_ (_28922_, _28911_, _28812_);
  nor _45016_ (_28933_, _28922_, _18475_);
  nor _45017_ (_28944_, _28933_, _28637_);
  and _45018_ (_28955_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _45019_ (_28966_, _28955_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _45020_ (_28977_, _28966_);
  and _45021_ (_28988_, _28977_, _28944_);
  and _45022_ (_29009_, _28977_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _45023_ (_29010_, _29009_, _28988_);
  nor _45024_ (_29021_, _29010_, _28615_);
  and _45025_ (_29032_, _29021_, _28582_);
  and _45026_ (_29043_, _29032_, _28549_);
  and _45027_ (_29054_, _29043_, _28516_);
  not _45028_ (_29064_, _19655_);
  or _45029_ (_29075_, _21054_, _29064_);
  and _45030_ (_29086_, _21054_, _29064_);
  or _45031_ (_29097_, _28472_, _29086_);
  and _45032_ (_29108_, _29097_, _29075_);
  or _45033_ (_29119_, _29108_, _29054_);
  and _45034_ (_29130_, _29119_, _28264_);
  and _45035_ (_29141_, _29130_, _28220_);
  and _45036_ (_29152_, _29141_, _28187_);
  nor _45037_ (_29163_, _29152_, _28154_);
  nor _45038_ (_29174_, _29163_, _27979_);
  and _45039_ (_29185_, _29163_, _27979_);
  nor _45040_ (_29196_, _29185_, _29174_);
  nor _45041_ (_29207_, _29196_, _27946_);
  not _45042_ (_29218_, _29207_);
  not _45043_ (_29229_, _27979_);
  not _45044_ (_29240_, _28034_);
  and _45045_ (_29251_, _28231_, _28089_);
  nor _45046_ (_29262_, _29251_, _28067_);
  nor _45047_ (_29273_, _29262_, _29240_);
  not _45048_ (_29284_, _28330_);
  and _45049_ (_29295_, _28593_, _28363_);
  nor _45050_ (_29306_, _29295_, _28341_);
  nor _45051_ (_29317_, _29306_, _29284_);
  nor _45052_ (_29328_, _29317_, _28308_);
  nor _45053_ (_29339_, _29328_, _28297_);
  and _45054_ (_29350_, _29328_, _28297_);
  nor _45055_ (_29361_, _29350_, _29339_);
  not _45056_ (_29371_, _28615_);
  nor _45057_ (_29382_, _29010_, _29371_);
  and _45058_ (_29393_, _29382_, _28363_);
  and _45059_ (_29404_, _29306_, _29284_);
  nor _45060_ (_29415_, _29404_, _29317_);
  and _45061_ (_29426_, _29415_, _29393_);
  not _45062_ (_29437_, _29426_);
  nor _45063_ (_29448_, _29437_, _29361_);
  nor _45064_ (_29459_, _29328_, _28285_);
  or _45065_ (_29470_, _29459_, _28286_);
  or _45066_ (_29481_, _29470_, _29448_);
  and _45067_ (_29492_, _29481_, _28253_);
  and _45068_ (_29503_, _29492_, _28089_);
  and _45069_ (_29514_, _29262_, _29240_);
  nor _45070_ (_29535_, _29514_, _29273_);
  and _45071_ (_29536_, _29535_, _29503_);
  or _45072_ (_29547_, _29536_, _29273_);
  nor _45073_ (_29558_, _29547_, _28012_);
  and _45074_ (_29569_, _29558_, _29229_);
  nor _45075_ (_29580_, _29558_, _29229_);
  not _45076_ (_29591_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _45077_ (_29602_, _23585_, _29591_);
  and _45078_ (_29613_, _29602_, _18256_);
  not _45079_ (_29624_, _29613_);
  or _45080_ (_29635_, _29624_, _29580_);
  nor _45081_ (_29646_, _29635_, _29569_);
  and _45082_ (_29657_, _18245_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _45083_ (_29668_, _29657_, _27924_);
  nor _45084_ (_29678_, _21925_, _21381_);
  and _45085_ (_29689_, _29678_, _21566_);
  and _45086_ (_29700_, _29689_, _21065_);
  and _45087_ (_29711_, _29700_, _20706_);
  and _45088_ (_29722_, _29711_, _20532_);
  and _45089_ (_29733_, _29722_, _19492_);
  and _45090_ (_29744_, _29733_, _29010_);
  not _45091_ (_29755_, _29010_);
  and _45092_ (_29766_, _19481_, _20521_);
  and _45093_ (_29777_, _21555_, _21381_);
  and _45094_ (_29788_, _29777_, _21925_);
  and _45095_ (_29808_, _29788_, _21054_);
  and _45096_ (_29809_, _29808_, _20695_);
  and _45097_ (_29820_, _29809_, _29766_);
  and _45098_ (_29831_, _29820_, _29755_);
  nor _45099_ (_29842_, _29831_, _29744_);
  and _45100_ (_29853_, _29842_, _20325_);
  nor _45101_ (_29864_, _29842_, _20325_);
  nor _45102_ (_29875_, _29864_, _29853_);
  and _45103_ (_29886_, _29875_, _29668_);
  not _45104_ (_29897_, _20151_);
  nor _45105_ (_29908_, _29010_, _29897_);
  not _45106_ (_29919_, _29908_);
  and _45107_ (_29930_, _29010_, _20325_);
  and _45108_ (_29941_, _29657_, _18223_);
  not _45109_ (_29951_, _29941_);
  nor _45110_ (_29962_, _29951_, _29930_);
  and _45111_ (_29973_, _29962_, _29919_);
  nor _45112_ (_29984_, _29973_, _29886_);
  and _45113_ (_29995_, _29602_, _23617_);
  nor _45114_ (_30006_, _29777_, _21054_);
  and _45115_ (_30017_, _30006_, _29995_);
  and _45116_ (_30028_, _30017_, _20706_);
  nor _45117_ (_30039_, _30028_, _20532_);
  and _45118_ (_30050_, _30039_, _19481_);
  nor _45119_ (_30061_, _29766_, _20325_);
  nor _45120_ (_30072_, _30061_, _30017_);
  and _45121_ (_30083_, _30072_, _29010_);
  nor _45122_ (_30093_, _30083_, _30050_);
  nor _45123_ (_30104_, _30093_, _20336_);
  and _45124_ (_30115_, _30093_, _20336_);
  nor _45125_ (_30126_, _30115_, _30104_);
  and _45126_ (_30137_, _30126_, _29995_);
  and _45127_ (_30148_, _29657_, _29602_);
  not _45128_ (_30159_, _30148_);
  nor _45129_ (_30170_, _30159_, _29010_);
  not _45130_ (_30181_, _30170_);
  not _45131_ (_30192_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _45132_ (_30203_, _18245_, _30192_);
  and _45133_ (_30214_, _30203_, _29602_);
  not _45134_ (_30225_, _30214_);
  nor _45135_ (_30235_, _30225_, _27978_);
  and _45136_ (_30246_, _30203_, _23596_);
  and _45137_ (_30257_, _30246_, _27979_);
  nor _45138_ (_30268_, _30257_, _30235_);
  and _45139_ (_30279_, _23617_, _18223_);
  and _45140_ (_30290_, _30279_, _27957_);
  and _45141_ (_30301_, _27924_, _23617_);
  and _45142_ (_30312_, _30301_, _20325_);
  nor _45143_ (_30323_, _30312_, _30290_);
  and _45144_ (_30334_, _30203_, _18212_);
  not _45145_ (_30345_, _30334_);
  nor _45146_ (_30356_, _30345_, _19481_);
  not _45147_ (_30367_, _30356_);
  and _45148_ (_30377_, _23596_, _18256_);
  not _45149_ (_30388_, _30377_);
  nor _45150_ (_30399_, _30388_, _20325_);
  and _45151_ (_30410_, _29657_, _23596_);
  and _45152_ (_30431_, _30410_, _21935_);
  nor _45153_ (_30432_, _30431_, _30399_);
  and _45154_ (_30443_, _30432_, _30367_);
  and _45155_ (_30454_, _30443_, _30323_);
  and _45156_ (_30465_, _30454_, _30268_);
  and _45157_ (_30476_, _30465_, _30181_);
  not _45158_ (_30487_, _30476_);
  nor _45159_ (_30498_, _30487_, _30137_);
  and _45160_ (_30509_, _30498_, _29984_);
  not _45161_ (_30519_, _30509_);
  nor _45162_ (_30530_, _30519_, _29646_);
  and _45163_ (_30541_, _30530_, _29218_);
  not _45164_ (_30552_, _30541_);
  nor _45165_ (_30563_, _30552_, _27902_);
  and _45166_ (_30574_, _30563_, _27891_);
  not _45167_ (_30585_, _30574_);
  or _45168_ (_30596_, _30585_, _27869_);
  not _45169_ (_30607_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _45170_ (_30618_, \oc8051_top_1.oc8051_decoder1.wr , _18201_);
  not _45171_ (_30629_, _30618_);
  nor _45172_ (_30640_, _30629_, _26476_);
  and _45173_ (_30651_, _30640_, _30607_);
  not _45174_ (_30661_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _45175_ (_30672_, _27869_, _30661_);
  and _45176_ (_30683_, _30672_, _30651_);
  and _45177_ (_30694_, _30683_, _30596_);
  nor _45178_ (_30705_, _30640_, _30661_);
  nor _45179_ (_30716_, _29580_, _27957_);
  nor _45180_ (_30727_, _30716_, _29624_);
  not _45181_ (_30738_, _30727_);
  and _45182_ (_30749_, _20325_, _29897_);
  nor _45183_ (_30759_, _30749_, _29174_);
  nor _45184_ (_30770_, _30759_, _27946_);
  and _45185_ (_30781_, _29010_, _19481_);
  and _45186_ (_30792_, _30781_, _30039_);
  nor _45187_ (_30803_, _30792_, _29930_);
  not _45188_ (_30814_, _29995_);
  nor _45189_ (_30825_, _29010_, _20325_);
  not _45190_ (_30836_, _30825_);
  nor _45191_ (_30847_, _30836_, _30050_);
  nor _45192_ (_30858_, _30847_, _30814_);
  and _45193_ (_30869_, _30858_, _30803_);
  not _45194_ (_30879_, _30869_);
  nor _45195_ (_30890_, _29009_, _28944_);
  not _45196_ (_30901_, _30246_);
  nor _45197_ (_30912_, _30901_, _28988_);
  nor _45198_ (_30923_, _30912_, _30214_);
  nor _45199_ (_30934_, _30923_, _30890_);
  not _45200_ (_30945_, _30934_);
  nor _45201_ (_30956_, _30388_, _29010_);
  not _45202_ (_30967_, _30956_);
  and _45203_ (_30978_, _28966_, _28944_);
  and _45204_ (_30988_, _30203_, _27924_);
  and _45205_ (_30999_, _30279_, _28944_);
  nor _45206_ (_31010_, _30999_, _30988_);
  nor _45207_ (_31021_, _31010_, _30978_);
  not _45208_ (_31032_, _31021_);
  not _45209_ (_31043_, _29009_);
  and _45210_ (_31054_, _30301_, _31043_);
  and _45211_ (_31065_, _30410_, _29009_);
  nor _45212_ (_31076_, _31065_, _31054_);
  nor _45213_ (_31087_, _31076_, _28988_);
  not _45214_ (_31097_, _31087_);
  nor _45215_ (_31108_, _30159_, _21925_);
  and _45216_ (_31119_, _30203_, _18223_);
  not _45217_ (_31141_, _31119_);
  nor _45218_ (_31142_, _31141_, _20325_);
  nor _45219_ (_31164_, _31142_, _31108_);
  not _45220_ (_31165_, _31164_);
  nor _45221_ (_31187_, _31165_, _30017_);
  and _45222_ (_31188_, _31187_, _31097_);
  and _45223_ (_31210_, _31188_, _31032_);
  and _45224_ (_31211_, _31210_, _30967_);
  and _45225_ (_31221_, _31211_, _30945_);
  and _45226_ (_31232_, _31221_, _30879_);
  not _45227_ (_31243_, _31232_);
  nor _45228_ (_31264_, _31243_, _30770_);
  and _45229_ (_31265_, _31264_, _30738_);
  not _45230_ (_31286_, _26740_);
  nor _45231_ (_31287_, _26981_, _26860_);
  and _45232_ (_31308_, _31287_, _31286_);
  and _45233_ (_31309_, _31308_, _27858_);
  nand _45234_ (_31329_, _31309_, _31265_);
  or _45235_ (_31330_, _31309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _45236_ (_31351_, _30640_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _45237_ (_31352_, _31351_, _31330_);
  and _45238_ (_31373_, _31352_, _31329_);
  or _45239_ (_31374_, _31373_, _30705_);
  or _45240_ (_31395_, _31374_, _30694_);
  and _45241_ (_06664_, _31395_, _43100_);
  and _45242_ (_31416_, _26023_, _23628_);
  not _45243_ (_31417_, _31416_);
  and _45244_ (_31437_, _23352_, _18267_);
  and _45245_ (_31438_, _29010_, _29371_);
  nor _45246_ (_31459_, _31438_, _29382_);
  not _45247_ (_31460_, _31459_);
  nor _45248_ (_31481_, _29613_, _27935_);
  nor _45249_ (_31482_, _31481_, _31460_);
  nor _45250_ (_31503_, _31141_, _29010_);
  not _45251_ (_31504_, _31503_);
  nor _45252_ (_31525_, _30901_, _28593_);
  nor _45253_ (_31526_, _31525_, _30214_);
  or _45254_ (_31546_, _31526_, _28604_);
  and _45255_ (_31547_, _29657_, _29591_);
  not _45256_ (_31568_, _31547_);
  nor _45257_ (_31569_, _31568_, _21381_);
  and _45258_ (_31590_, _30988_, _20336_);
  nor _45259_ (_31591_, _31590_, _31569_);
  and _45260_ (_31612_, _30279_, _28593_);
  and _45261_ (_31613_, _30301_, _21925_);
  nor _45262_ (_31634_, _31613_, _31612_);
  nor _45263_ (_31635_, _29951_, _18990_);
  and _45264_ (_31655_, _29668_, _21925_);
  nor _45265_ (_31656_, _31655_, _31635_);
  nor _45266_ (_31677_, _30377_, _29995_);
  nor _45267_ (_31678_, _31677_, _21925_);
  not _45268_ (_31699_, _31678_);
  and _45269_ (_31700_, _31699_, _31656_);
  and _45270_ (_31721_, _31700_, _31634_);
  and _45271_ (_31722_, _31721_, _31591_);
  and _45272_ (_31743_, _31722_, _31546_);
  and _45273_ (_31744_, _31743_, _31504_);
  not _45274_ (_31764_, _31744_);
  nor _45275_ (_31765_, _31764_, _31482_);
  not _45276_ (_31786_, _31765_);
  nor _45277_ (_31787_, _31786_, _31437_);
  and _45278_ (_31808_, _31787_, _31417_);
  not _45279_ (_31809_, _31808_);
  or _45280_ (_31830_, _31809_, _27869_);
  not _45281_ (_31831_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _45282_ (_31852_, _27869_, _31831_);
  and _45283_ (_31853_, _31852_, _30651_);
  and _45284_ (_31864_, _31853_, _31830_);
  nor _45285_ (_31874_, _30640_, _31831_);
  not _45286_ (_31885_, _31265_);
  or _45287_ (_31896_, _31885_, _27869_);
  and _45288_ (_31907_, _31852_, _31351_);
  and _45289_ (_31918_, _31907_, _31896_);
  or _45290_ (_31929_, _31918_, _31874_);
  or _45291_ (_31940_, _31929_, _31864_);
  and _45292_ (_08905_, _31940_, _43100_);
  and _45293_ (_31961_, _23384_, _18267_);
  not _45294_ (_31972_, _31961_);
  and _45295_ (_31982_, _26088_, _23628_);
  nor _45296_ (_31993_, _28593_, _28363_);
  or _45297_ (_32004_, _31993_, _29295_);
  and _45298_ (_32015_, _32004_, _29382_);
  nor _45299_ (_32026_, _32004_, _29382_);
  or _45300_ (_32037_, _32026_, _32015_);
  and _45301_ (_32048_, _32037_, _29613_);
  nor _45302_ (_32059_, _29021_, _28582_);
  nor _45303_ (_32070_, _32059_, _29032_);
  nor _45304_ (_32081_, _32070_, _27946_);
  not _45305_ (_32091_, _32081_);
  nor _45306_ (_32102_, _30006_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _45307_ (_32113_, _32102_, _21392_);
  nor _45308_ (_32124_, _32102_, _21392_);
  nor _45309_ (_32135_, _32124_, _32113_);
  nor _45310_ (_32146_, _32135_, _30814_);
  not _45311_ (_32157_, _32146_);
  and _45312_ (_32168_, _30246_, _28363_);
  nor _45313_ (_32179_, _30225_, _28352_);
  not _45314_ (_32190_, _32179_);
  and _45315_ (_32200_, _30279_, _28341_);
  and _45316_ (_32211_, _30301_, _21381_);
  nor _45317_ (_32222_, _32211_, _32200_);
  nand _45318_ (_32233_, _32222_, _32190_);
  nor _45319_ (_32244_, _32233_, _32168_);
  nor _45320_ (_32255_, _30345_, _21925_);
  not _45321_ (_32266_, _32255_);
  nor _45322_ (_32277_, _30388_, _21381_);
  nor _45323_ (_32288_, _31568_, _21555_);
  nor _45324_ (_32299_, _32288_, _32277_);
  and _45325_ (_32309_, _32299_, _32266_);
  and _45326_ (_32320_, _32309_, _32244_);
  and _45327_ (_32331_, _32320_, _32157_);
  and _45328_ (_32342_, _32331_, _32091_);
  nor _45329_ (_32353_, _29951_, _19977_);
  and _45330_ (_32364_, _21925_, _21381_);
  nor _45331_ (_32375_, _32364_, _29678_);
  not _45332_ (_32386_, _32375_);
  nor _45333_ (_32397_, _32386_, _29010_);
  and _45334_ (_32408_, _32386_, _29010_);
  nor _45335_ (_32418_, _32408_, _32397_);
  and _45336_ (_32429_, _32418_, _29668_);
  nor _45337_ (_32440_, _32429_, _32353_);
  nand _45338_ (_32451_, _32440_, _32342_);
  nor _45339_ (_32462_, _32451_, _32048_);
  not _45340_ (_32473_, _32462_);
  nor _45341_ (_32484_, _32473_, _31982_);
  and _45342_ (_32495_, _32484_, _31972_);
  not _45343_ (_32506_, _32495_);
  or _45344_ (_32517_, _32506_, _27869_);
  not _45345_ (_32527_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _45346_ (_32538_, _27869_, _32527_);
  and _45347_ (_32549_, _32538_, _30651_);
  and _45348_ (_32560_, _32549_, _32517_);
  nor _45349_ (_32571_, _30640_, _32527_);
  not _45350_ (_32582_, _26981_);
  and _45351_ (_32593_, _32582_, _26860_);
  and _45352_ (_32604_, _32593_, _26740_);
  and _45353_ (_32615_, _32604_, _27858_);
  nand _45354_ (_32626_, _32615_, _31265_);
  or _45355_ (_32636_, _32615_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _45356_ (_32647_, _32636_, _31351_);
  and _45357_ (_32658_, _32647_, _32626_);
  or _45358_ (_32669_, _32658_, _32571_);
  or _45359_ (_32680_, _32669_, _32560_);
  and _45360_ (_08916_, _32680_, _43100_);
  and _45361_ (_32701_, _26152_, _23628_);
  not _45362_ (_32712_, _32701_);
  and _45363_ (_32723_, _23415_, _18267_);
  nor _45364_ (_32734_, _29951_, _18671_);
  nor _45365_ (_32744_, _32364_, _29010_);
  nor _45366_ (_32755_, _29678_, _29755_);
  nor _45367_ (_32766_, _32755_, _32744_);
  and _45368_ (_32777_, _32766_, _21566_);
  not _45369_ (_32788_, _32777_);
  not _45370_ (_32799_, _29668_);
  nor _45371_ (_32810_, _32766_, _21566_);
  nor _45372_ (_32821_, _32810_, _32799_);
  and _45373_ (_32832_, _32821_, _32788_);
  nor _45374_ (_32843_, _32832_, _32734_);
  nor _45375_ (_32854_, _29032_, _28549_);
  nor _45376_ (_32864_, _32854_, _29043_);
  nor _45377_ (_32875_, _32864_, _27946_);
  and _45378_ (_32886_, _30246_, _28330_);
  nor _45379_ (_32897_, _30225_, _28319_);
  not _45380_ (_32908_, _32897_);
  and _45381_ (_32919_, _30279_, _28308_);
  and _45382_ (_32930_, _30301_, _21555_);
  nor _45383_ (_32941_, _32930_, _32919_);
  nand _45384_ (_32952_, _32941_, _32908_);
  nor _45385_ (_32963_, _32952_, _32886_);
  nor _45386_ (_32973_, _30345_, _21381_);
  not _45387_ (_32984_, _32973_);
  nor _45388_ (_32995_, _30388_, _21555_);
  nor _45389_ (_33006_, _31568_, _21054_);
  nor _45390_ (_33017_, _33006_, _32995_);
  and _45391_ (_33028_, _33017_, _32984_);
  and _45392_ (_33039_, _33028_, _32963_);
  not _45393_ (_33050_, _33039_);
  nor _45394_ (_33061_, _33050_, _32875_);
  nor _45395_ (_33071_, _29415_, _29393_);
  nor _45396_ (_33082_, _33071_, _29624_);
  and _45397_ (_33093_, _33082_, _29437_);
  and _45398_ (_33104_, _29777_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45399_ (_33115_, _32124_, _21555_);
  nor _45400_ (_33126_, _33115_, _33104_);
  nor _45401_ (_33137_, _33126_, _30814_);
  nor _45402_ (_33148_, _33137_, _33093_);
  and _45403_ (_33159_, _33148_, _33061_);
  and _45404_ (_33170_, _33159_, _32843_);
  not _45405_ (_33180_, _33170_);
  nor _45406_ (_33191_, _33180_, _32723_);
  and _45407_ (_33202_, _33191_, _32712_);
  not _45408_ (_33213_, _33202_);
  or _45409_ (_33224_, _33213_, _27869_);
  not _45410_ (_33235_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _45411_ (_33246_, _27869_, _33235_);
  and _45412_ (_33257_, _33246_, _30651_);
  and _45413_ (_33268_, _33257_, _33224_);
  nor _45414_ (_33279_, _30640_, _33235_);
  nand _45415_ (_33289_, _27858_, _26740_);
  or _45416_ (_33300_, _31287_, _33289_);
  and _45417_ (_33311_, _33300_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _45418_ (_33322_, _26860_);
  and _45419_ (_33333_, _26740_, _26981_);
  and _45420_ (_33344_, _33333_, _33322_);
  not _45421_ (_33355_, _33344_);
  nor _45422_ (_33366_, _33355_, _31265_);
  and _45423_ (_33377_, _26740_, _26860_);
  and _45424_ (_33388_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _45425_ (_33399_, _33388_, _33366_);
  and _45426_ (_33409_, _33399_, _27858_);
  or _45427_ (_33420_, _33409_, _33311_);
  and _45428_ (_33431_, _33420_, _31351_);
  or _45429_ (_33442_, _33431_, _33279_);
  or _45430_ (_33453_, _33442_, _33268_);
  and _45431_ (_08927_, _33453_, _43100_);
  and _45432_ (_33474_, _26217_, _23628_);
  not _45433_ (_33485_, _33474_);
  not _45434_ (_33496_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45435_ (_33507_, _29777_, _33496_);
  nor _45436_ (_33517_, _33507_, _21065_);
  nor _45437_ (_33528_, _30388_, _21054_);
  nor _45438_ (_33539_, _30006_, _30814_);
  nor _45439_ (_33550_, _33539_, _33528_);
  nor _45440_ (_33561_, _33550_, _33517_);
  not _45441_ (_33572_, _33561_);
  nor _45442_ (_33583_, _30225_, _28285_);
  and _45443_ (_33594_, _30246_, _28297_);
  nor _45444_ (_33605_, _33594_, _33583_);
  and _45445_ (_33616_, _30279_, _28286_);
  and _45446_ (_33626_, _30301_, _21054_);
  nor _45447_ (_33637_, _33626_, _33616_);
  nor _45448_ (_33648_, _31568_, _20695_);
  nor _45449_ (_33659_, _30345_, _21555_);
  nor _45450_ (_33670_, _33659_, _33648_);
  and _45451_ (_33681_, _33670_, _33637_);
  and _45452_ (_33692_, _33681_, _33605_);
  and _45453_ (_33703_, _33692_, _33572_);
  nor _45454_ (_33714_, _29043_, _28516_);
  nor _45455_ (_33725_, _33714_, _29054_);
  nor _45456_ (_33735_, _33725_, _27946_);
  and _45457_ (_33746_, _29437_, _29361_);
  or _45458_ (_33757_, _33746_, _29624_);
  nor _45459_ (_33768_, _33757_, _29448_);
  nor _45460_ (_33779_, _33768_, _33735_);
  and _45461_ (_33790_, _33779_, _33703_);
  and _45462_ (_33801_, _23468_, _18267_);
  not _45463_ (_33812_, _33801_);
  nor _45464_ (_33823_, _29951_, _19655_);
  and _45465_ (_33833_, _29689_, _29010_);
  and _45466_ (_33844_, _29788_, _29755_);
  nor _45467_ (_33855_, _33844_, _33833_);
  nor _45468_ (_33866_, _33855_, _21054_);
  not _45469_ (_33877_, _33866_);
  and _45470_ (_33888_, _33855_, _21054_);
  nor _45471_ (_33899_, _33888_, _32799_);
  and _45472_ (_33910_, _33899_, _33877_);
  nor _45473_ (_33921_, _33910_, _33823_);
  and _45474_ (_33932_, _33921_, _33812_);
  and _45475_ (_33943_, _33932_, _33790_);
  and _45476_ (_33953_, _33943_, _33485_);
  not _45477_ (_33964_, _33953_);
  or _45478_ (_33975_, _33964_, _27869_);
  not _45479_ (_33986_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _45480_ (_33997_, _27869_, _33986_);
  and _45481_ (_34008_, _33997_, _30651_);
  and _45482_ (_34019_, _34008_, _33975_);
  nor _45483_ (_34030_, _30640_, _33986_);
  and _45484_ (_34041_, _33289_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _45485_ (_34052_, _31287_, _26740_);
  and _45486_ (_34062_, _34052_, _31885_);
  nor _45487_ (_34073_, _33377_, _33333_);
  nor _45488_ (_34084_, _34073_, _33986_);
  or _45489_ (_34095_, _34084_, _34062_);
  and _45490_ (_34106_, _34095_, _27858_);
  or _45491_ (_34117_, _34106_, _34041_);
  and _45492_ (_34128_, _34117_, _31351_);
  or _45493_ (_34139_, _34128_, _34030_);
  or _45494_ (_34150_, _34139_, _34019_);
  and _45495_ (_08938_, _34150_, _43100_);
  and _45496_ (_34170_, _23490_, _18267_);
  not _45497_ (_34181_, _34170_);
  and _45498_ (_34192_, _26282_, _23628_);
  nor _45499_ (_34203_, _29010_, _18836_);
  and _45500_ (_34214_, _29010_, _20706_);
  nor _45501_ (_34225_, _34214_, _34203_);
  nor _45502_ (_34236_, _34225_, _29951_);
  and _45503_ (_34247_, _29700_, _29010_);
  and _45504_ (_34258_, _29808_, _29755_);
  nor _45505_ (_34269_, _34258_, _34247_);
  and _45506_ (_34281_, _34269_, _20695_);
  nor _45507_ (_34300_, _34269_, _20695_);
  nor _45508_ (_34311_, _34300_, _34281_);
  and _45509_ (_34322_, _34311_, _29668_);
  nor _45510_ (_34333_, _34322_, _34236_);
  and _45511_ (_34344_, _30279_, _28231_);
  and _45512_ (_34355_, _30301_, _20695_);
  nor _45513_ (_34366_, _34355_, _34344_);
  nor _45514_ (_34377_, _31568_, _20521_);
  not _45515_ (_34388_, _34377_);
  and _45516_ (_34398_, _34388_, _34366_);
  nor _45517_ (_34409_, _30017_, _20706_);
  not _45518_ (_34420_, _34409_);
  nor _45519_ (_34431_, _30028_, _30814_);
  and _45520_ (_34442_, _34431_, _34420_);
  nor _45521_ (_34453_, _30225_, _28242_);
  and _45522_ (_34464_, _30246_, _28253_);
  nor _45523_ (_34475_, _34464_, _34453_);
  nor _45524_ (_34486_, _30345_, _21054_);
  nor _45525_ (_34497_, _30388_, _20695_);
  nor _45526_ (_34507_, _34497_, _34486_);
  nand _45527_ (_34518_, _34507_, _34475_);
  nor _45528_ (_34529_, _34518_, _34442_);
  and _45529_ (_34540_, _34529_, _34398_);
  nor _45530_ (_34551_, _29119_, _28253_);
  and _45531_ (_34562_, _29119_, _28253_);
  nor _45532_ (_34573_, _34562_, _34551_);
  and _45533_ (_34584_, _34573_, _27935_);
  nor _45534_ (_34595_, _29481_, _28253_);
  not _45535_ (_34606_, _34595_);
  nor _45536_ (_34616_, _29624_, _29492_);
  and _45537_ (_34627_, _34616_, _34606_);
  nor _45538_ (_34638_, _34627_, _34584_);
  and _45539_ (_34649_, _34638_, _34540_);
  and _45540_ (_34660_, _34649_, _34333_);
  not _45541_ (_34671_, _34660_);
  nor _45542_ (_34682_, _34671_, _34192_);
  and _45543_ (_34693_, _34682_, _34181_);
  not _45544_ (_34704_, _34693_);
  or _45545_ (_34715_, _34704_, _27869_);
  not _45546_ (_34725_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _45547_ (_34736_, _27869_, _34725_);
  and _45548_ (_34747_, _34736_, _30651_);
  and _45549_ (_34758_, _34747_, _34715_);
  nor _45550_ (_34769_, _30640_, _34725_);
  not _45551_ (_34780_, _27858_);
  and _45552_ (_34791_, _26992_, _31286_);
  nor _45553_ (_34802_, _26992_, _31286_);
  nor _45554_ (_34813_, _34802_, _34791_);
  or _45555_ (_34824_, _34813_, _34780_);
  and _45556_ (_34834_, _34824_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _45557_ (_34845_, _34791_, _31885_);
  and _45558_ (_34856_, _34802_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _45559_ (_34867_, _34856_, _34845_);
  and _45560_ (_34878_, _34867_, _27858_);
  or _45561_ (_34889_, _34878_, _34834_);
  and _45562_ (_34900_, _34889_, _31351_);
  or _45563_ (_34911_, _34900_, _34769_);
  or _45564_ (_34922_, _34911_, _34758_);
  and _45565_ (_08949_, _34922_, _43100_);
  and _45566_ (_34942_, _26369_, _23628_);
  not _45567_ (_34953_, _34942_);
  and _45568_ (_34964_, _23532_, _18267_);
  nor _45569_ (_34975_, _28231_, _28089_);
  nor _45570_ (_34986_, _34975_, _29251_);
  nor _45571_ (_34997_, _34986_, _29492_);
  nor _45572_ (_35008_, _34997_, _29503_);
  and _45573_ (_35019_, _35008_, _29613_);
  not _45574_ (_35030_, _35019_);
  nor _45575_ (_35041_, _29130_, _28220_);
  nor _45576_ (_35051_, _35041_, _29141_);
  nor _45577_ (_35062_, _35051_, _27946_);
  nor _45578_ (_35073_, _29010_, _19807_);
  and _45579_ (_35084_, _29010_, _20532_);
  nor _45580_ (_35095_, _35084_, _35073_);
  nor _45581_ (_35106_, _35095_, _29951_);
  and _45582_ (_35117_, _29711_, _29010_);
  and _45583_ (_35128_, _29809_, _29755_);
  nor _45584_ (_35139_, _35128_, _35117_);
  nor _45585_ (_35150_, _35139_, _20521_);
  and _45586_ (_35160_, _35139_, _20521_);
  or _45587_ (_35171_, _35160_, _32799_);
  nor _45588_ (_35182_, _35171_, _35150_);
  nor _45589_ (_35193_, _35182_, _35106_);
  not _45590_ (_35204_, _30083_);
  and _45591_ (_35215_, _35204_, _30039_);
  nor _45592_ (_35226_, _30083_, _30028_);
  nor _45593_ (_35237_, _35226_, _20521_);
  nor _45594_ (_35248_, _35237_, _35215_);
  nor _45595_ (_35259_, _35248_, _30814_);
  and _45596_ (_35269_, _30246_, _28089_);
  nor _45597_ (_35280_, _30225_, _28078_);
  not _45598_ (_35291_, _35280_);
  and _45599_ (_35302_, _30279_, _28067_);
  and _45600_ (_35313_, _30301_, _20521_);
  nor _45601_ (_35324_, _35313_, _35302_);
  nand _45602_ (_35335_, _35324_, _35291_);
  nor _45603_ (_35346_, _35335_, _35269_);
  nor _45604_ (_35356_, _30388_, _20521_);
  not _45605_ (_35367_, _35356_);
  nor _45606_ (_35378_, _31568_, _19481_);
  nor _45607_ (_35389_, _30345_, _20695_);
  nor _45608_ (_35400_, _35389_, _35378_);
  and _45609_ (_35411_, _35400_, _35367_);
  and _45610_ (_35422_, _35411_, _35346_);
  not _45611_ (_35433_, _35422_);
  nor _45612_ (_35444_, _35433_, _35259_);
  and _45613_ (_35455_, _35444_, _35193_);
  not _45614_ (_35465_, _35455_);
  nor _45615_ (_35476_, _35465_, _35062_);
  and _45616_ (_35487_, _35476_, _35030_);
  not _45617_ (_35498_, _35487_);
  nor _45618_ (_35509_, _35498_, _34964_);
  and _45619_ (_35520_, _35509_, _34953_);
  not _45620_ (_35531_, _35520_);
  or _45621_ (_35542_, _35531_, _27869_);
  not _45622_ (_35553_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _45623_ (_35564_, _27869_, _35553_);
  and _45624_ (_35575_, _35564_, _30651_);
  and _45625_ (_35585_, _35575_, _35542_);
  nor _45626_ (_35596_, _30640_, _35553_);
  and _45627_ (_35607_, _32593_, _31286_);
  and _45628_ (_35618_, _35607_, _27858_);
  nand _45629_ (_35629_, _35618_, _31265_);
  or _45630_ (_35640_, _35618_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _45631_ (_35651_, _35640_, _31351_);
  and _45632_ (_35662_, _35651_, _35629_);
  or _45633_ (_35673_, _35662_, _35596_);
  or _45634_ (_35684_, _35673_, _35585_);
  and _45635_ (_08960_, _35684_, _43100_);
  and _45636_ (_35704_, _26433_, _23628_);
  not _45637_ (_35715_, _35704_);
  and _45638_ (_35726_, _23564_, _18267_);
  nor _45639_ (_35737_, _29141_, _28187_);
  nor _45640_ (_35748_, _35737_, _29152_);
  nor _45641_ (_35759_, _35748_, _27946_);
  not _45642_ (_35770_, _35759_);
  nor _45643_ (_35781_, _29535_, _29503_);
  not _45644_ (_35792_, _35781_);
  nor _45645_ (_35803_, _29624_, _29536_);
  and _45646_ (_35814_, _35803_, _35792_);
  nor _45647_ (_35825_, _29010_, _27990_);
  or _45648_ (_35835_, _35825_, _29951_);
  nor _45649_ (_35846_, _35835_, _30781_);
  or _45650_ (_35857_, _29010_, _20521_);
  or _45651_ (_35868_, _35128_, _29722_);
  and _45652_ (_35879_, _35868_, _35857_);
  nor _45653_ (_35890_, _35879_, _19492_);
  and _45654_ (_35901_, _35879_, _19492_);
  or _45655_ (_35912_, _35901_, _32799_);
  nor _45656_ (_35923_, _35912_, _35890_);
  nor _45657_ (_35934_, _35923_, _35846_);
  nor _45658_ (_35945_, _35215_, _19481_);
  and _45659_ (_35955_, _35215_, _19481_);
  nor _45660_ (_35966_, _35955_, _35945_);
  nor _45661_ (_35977_, _35966_, _30814_);
  and _45662_ (_35988_, _30246_, _28034_);
  nor _45663_ (_35999_, _30225_, _28023_);
  not _45664_ (_36010_, _35999_);
  and _45665_ (_36021_, _30279_, _28012_);
  and _45666_ (_36032_, _30301_, _19481_);
  nor _45667_ (_36043_, _36032_, _36021_);
  nand _45668_ (_36054_, _36043_, _36010_);
  nor _45669_ (_36065_, _36054_, _35988_);
  nor _45670_ (_36076_, _31568_, _20325_);
  not _45671_ (_36086_, _36076_);
  nor _45672_ (_36097_, _30388_, _19481_);
  nor _45673_ (_36108_, _30345_, _20521_);
  nor _45674_ (_36119_, _36108_, _36097_);
  and _45675_ (_36130_, _36119_, _36086_);
  and _45676_ (_36141_, _36130_, _36065_);
  not _45677_ (_36152_, _36141_);
  nor _45678_ (_36162_, _36152_, _35977_);
  and _45679_ (_36173_, _36162_, _35934_);
  not _45680_ (_36184_, _36173_);
  nor _45681_ (_36195_, _36184_, _35814_);
  and _45682_ (_36206_, _36195_, _35770_);
  not _45683_ (_36217_, _36206_);
  nor _45684_ (_36228_, _36217_, _35726_);
  and _45685_ (_36239_, _36228_, _35715_);
  not _45686_ (_36249_, _36239_);
  or _45687_ (_36260_, _36249_, _27869_);
  not _45688_ (_36271_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _45689_ (_36282_, _27869_, _36271_);
  and _45690_ (_36293_, _36282_, _30651_);
  and _45691_ (_36304_, _36293_, _36260_);
  nor _45692_ (_36315_, _30640_, _36271_);
  nor _45693_ (_36326_, _26740_, _26860_);
  and _45694_ (_36336_, _36326_, _26981_);
  and _45695_ (_36347_, _36336_, _27858_);
  nand _45696_ (_36358_, _36347_, _31265_);
  or _45697_ (_36369_, _36347_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _45698_ (_36380_, _36369_, _31351_);
  and _45699_ (_36391_, _36380_, _36358_);
  or _45700_ (_36402_, _36391_, _36315_);
  or _45701_ (_36413_, _36402_, _36304_);
  and _45702_ (_08971_, _36413_, _43100_);
  and _45703_ (_36433_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45704_ (_36444_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or _45705_ (_36455_, _36444_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _45706_ (_36466_, _36455_);
  not _45707_ (_36477_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _45708_ (_36488_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _45709_ (_36498_, _36488_, _36477_);
  and _45710_ (_36509_, _36444_, _18201_);
  and _45711_ (_36520_, _36509_, _36498_);
  not _45712_ (_36531_, _36520_);
  not _45713_ (_36542_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _45714_ (_36553_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _45715_ (_36564_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45716_ (_36575_, _36564_, _36553_);
  and _45717_ (_36585_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _45718_ (_36596_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45719_ (_36607_, _36596_, _36553_);
  and _45720_ (_36618_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not _45721_ (_36629_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45722_ (_36640_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _36629_);
  and _45723_ (_36651_, _36640_, _36553_);
  and _45724_ (_36662_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _45725_ (_36672_, _36662_, _36618_);
  or _45726_ (_36683_, _36672_, _36585_);
  and _45727_ (_36694_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _45728_ (_36705_, _36596_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _45729_ (_36716_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _45730_ (_36727_, _36716_, _36694_);
  nor _45731_ (_36738_, _36596_, _36553_);
  and _45732_ (_36749_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not _45733_ (_36760_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _45734_ (_36770_, _36760_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45735_ (_36781_, _36770_, _36553_);
  and _45736_ (_36792_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _45737_ (_36803_, _36792_, _36749_);
  or _45738_ (_36814_, _36803_, _36727_);
  nor _45739_ (_36825_, _36814_, _36683_);
  and _45740_ (_36836_, _36825_, _36542_);
  nor _45741_ (_36847_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _36542_);
  or _45742_ (_36858_, _36847_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45743_ (_36869_, _36858_, _36836_);
  and _45744_ (_36880_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _45745_ (_36890_, _36880_, _36869_);
  nor _45746_ (_36901_, _36890_, _36531_);
  not _45747_ (_36912_, _36901_);
  not _45748_ (_36923_, _36498_);
  nor _45749_ (_36934_, _36509_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _45750_ (_36945_, _36934_, _36923_);
  and _45751_ (_36956_, _36945_, _36912_);
  not _45752_ (_36967_, _36956_);
  and _45753_ (_36978_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45754_ (_36989_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45755_ (_37000_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and _45756_ (_37011_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _45757_ (_37022_, _37011_, _37000_);
  and _45758_ (_37033_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _45759_ (_37044_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _45760_ (_37055_, _37044_, _37033_);
  and _45761_ (_37066_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and _45762_ (_37077_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _45763_ (_37088_, _37077_, _37066_);
  and _45764_ (_37099_, _37088_, _37055_);
  and _45765_ (_37110_, _37099_, _37022_);
  nor _45766_ (_37121_, _37110_, _36694_);
  and _45767_ (_37132_, _37121_, _36542_);
  nor _45768_ (_37142_, _37132_, _36989_);
  nor _45769_ (_37153_, _37142_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45770_ (_37164_, _37153_, _36978_);
  and _45771_ (_37175_, _37164_, _36520_);
  not _45772_ (_37186_, _37175_);
  nor _45773_ (_37197_, _36509_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _45774_ (_37208_, _37197_, _36923_);
  and _45775_ (_37219_, _37208_, _37186_);
  and _45776_ (_37230_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not _45777_ (_37241_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45778_ (_37251_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  or _45779_ (_37262_, _36694_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45780_ (_37273_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _45781_ (_37284_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _45782_ (_37295_, _37284_, _37273_);
  and _45783_ (_37306_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and _45784_ (_37317_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _45785_ (_37328_, _37317_, _37306_);
  and _45786_ (_37339_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and _45787_ (_37350_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _45788_ (_37361_, _37350_, _37339_);
  and _45789_ (_37371_, _37361_, _37328_);
  and _45790_ (_37382_, _37371_, _37295_);
  nor _45791_ (_37393_, _37382_, _37262_);
  or _45792_ (_37404_, _37393_, _37251_);
  and _45793_ (_37415_, _37404_, _37241_);
  nor _45794_ (_37426_, _37415_, _37230_);
  nor _45795_ (_37437_, _37426_, _36531_);
  and _45796_ (_37448_, _36531_, \oc8051_top_1.oc8051_decoder1.op [7]);
  or _45797_ (_37459_, _37448_, _37437_);
  and _45798_ (_37470_, _37459_, _36498_);
  and _45799_ (_37480_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45800_ (_37491_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45801_ (_37502_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _45802_ (_37513_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _45803_ (_37524_, _37513_, _37502_);
  and _45804_ (_37535_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _45805_ (_37546_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _45806_ (_37557_, _37546_, _37535_);
  and _45807_ (_37568_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and _45808_ (_37579_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _45809_ (_37590_, _37579_, _37568_);
  and _45810_ (_37601_, _37590_, _37557_);
  and _45811_ (_37612_, _37601_, _37524_);
  nor _45812_ (_37623_, _37612_, _37262_);
  or _45813_ (_37634_, _37623_, _37491_);
  and _45814_ (_37645_, _37634_, _37241_);
  nor _45815_ (_37654_, _37645_, _37480_);
  and _45816_ (_37665_, _37654_, _36520_);
  not _45817_ (_37676_, _37665_);
  nor _45818_ (_37687_, _36509_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _45819_ (_37698_, _37687_, _36923_);
  and _45820_ (_37709_, _37698_, _37676_);
  not _45821_ (_37720_, _37709_);
  and _45822_ (_37731_, _37720_, _37470_);
  and _45823_ (_37742_, _37731_, _37219_);
  and _45824_ (_37753_, _37742_, _36967_);
  and _45825_ (_37764_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45826_ (_37775_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45827_ (_37786_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _45828_ (_37797_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _45829_ (_37808_, _37797_, _37786_);
  and _45830_ (_37819_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _45831_ (_37830_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _45832_ (_37841_, _37830_, _37819_);
  and _45833_ (_37852_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _45834_ (_37863_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _45835_ (_37874_, _37863_, _37852_);
  and _45836_ (_37885_, _37874_, _37841_);
  and _45837_ (_37896_, _37885_, _37808_);
  nor _45838_ (_37907_, _37896_, _36694_);
  and _45839_ (_37918_, _37907_, _36542_);
  nor _45840_ (_37929_, _37918_, _37775_);
  nor _45841_ (_37940_, _37929_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45842_ (_37951_, _37940_, _37764_);
  and _45843_ (_37962_, _37951_, _36520_);
  not _45844_ (_37973_, _37962_);
  nor _45845_ (_37984_, _36509_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _45846_ (_37995_, _37984_, _36923_);
  and _45847_ (_38006_, _37995_, _37973_);
  not _45848_ (_38017_, _36694_);
  and _45849_ (_38028_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _45850_ (_38039_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _45851_ (_38050_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _45852_ (_38061_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _45853_ (_38072_, _38061_, _38050_);
  and _45854_ (_38083_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and _45855_ (_38094_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _45856_ (_38105_, _38094_, _38083_);
  nand _45857_ (_38116_, _38105_, _38072_);
  or _45858_ (_38127_, _38116_, _38039_);
  nor _45859_ (_38138_, _38127_, _38028_);
  and _45860_ (_38149_, _38138_, _38017_);
  and _45861_ (_38160_, _38149_, _36542_);
  nor _45862_ (_38171_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _36542_);
  nor _45863_ (_38182_, _38171_, _38160_);
  nor _45864_ (_38193_, _38182_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45865_ (_38204_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _37241_);
  nor _45866_ (_38215_, _38204_, _38193_);
  nor _45867_ (_38226_, _38215_, _36531_);
  not _45868_ (_38237_, _38226_);
  nor _45869_ (_38248_, _36509_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _45870_ (_38259_, _38248_, _36923_);
  and _45871_ (_38270_, _38259_, _38237_);
  and _45872_ (_38281_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45873_ (_38292_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45874_ (_38302_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _45875_ (_38313_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _45876_ (_38324_, _38313_, _38302_);
  and _45877_ (_38335_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _45878_ (_38345_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _45879_ (_38356_, _38345_, _38335_);
  and _45880_ (_38367_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _45881_ (_38378_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _45882_ (_38389_, _38378_, _38367_);
  and _45883_ (_38400_, _38389_, _38356_);
  and _45884_ (_38406_, _38400_, _38324_);
  nor _45885_ (_38407_, _38406_, _37262_);
  nor _45886_ (_38408_, _38407_, _38292_);
  nor _45887_ (_38409_, _38408_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45888_ (_38410_, _38409_, _38281_);
  nor _45889_ (_38411_, _38410_, _36531_);
  and _45890_ (_38412_, _36531_, \oc8051_top_1.oc8051_decoder1.op [2]);
  or _45891_ (_38413_, _38412_, _38411_);
  and _45892_ (_38414_, _38413_, _36498_);
  and _45893_ (_38415_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45894_ (_38416_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45895_ (_38417_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and _45896_ (_38418_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _45897_ (_38419_, _38418_, _38417_);
  and _45898_ (_38420_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _45899_ (_38421_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _45900_ (_38422_, _38421_, _38420_);
  and _45901_ (_38423_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _45902_ (_38424_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _45903_ (_38425_, _38424_, _38423_);
  and _45904_ (_38426_, _38425_, _38422_);
  and _45905_ (_38427_, _38426_, _38419_);
  nor _45906_ (_38428_, _38427_, _36694_);
  and _45907_ (_38429_, _38428_, _36542_);
  or _45908_ (_38430_, _38429_, _38416_);
  and _45909_ (_38431_, _38430_, _37241_);
  nor _45910_ (_38432_, _38431_, _38415_);
  and _45911_ (_38433_, _38432_, _36520_);
  not _45912_ (_38434_, _38433_);
  nor _45913_ (_38435_, _36509_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _45914_ (_38436_, _38435_, _36923_);
  and _45915_ (_38437_, _38436_, _38434_);
  nor _45916_ (_38438_, _38437_, _38414_);
  and _45917_ (_38439_, _38438_, _38270_);
  and _45918_ (_38440_, _38439_, _38006_);
  and _45919_ (_38441_, _38440_, _37753_);
  not _45920_ (_38442_, _38441_);
  nor _45921_ (_38443_, _37720_, _37470_);
  and _45922_ (_38444_, _38443_, _37219_);
  and _45923_ (_38445_, _38444_, _36956_);
  and _45924_ (_38446_, _38440_, _38445_);
  nor _45925_ (_38447_, _37219_, _37709_);
  and _45926_ (_38448_, _38447_, _37470_);
  and _45927_ (_38449_, _38448_, _36956_);
  and _45928_ (_38450_, _38440_, _38449_);
  nor _45929_ (_38451_, _38450_, _38446_);
  and _45930_ (_38452_, _38451_, _38442_);
  and _45931_ (_38453_, _38448_, _36967_);
  not _45932_ (_38454_, _38437_);
  and _45933_ (_38455_, _38454_, _38414_);
  nor _45934_ (_38456_, _38006_, _38270_);
  and _45935_ (_38457_, _38456_, _38455_);
  and _45936_ (_38458_, _38457_, _38453_);
  and _45937_ (_38459_, _38457_, _37753_);
  nor _45938_ (_38460_, _38459_, _38458_);
  and _45939_ (_38461_, _38460_, _38452_);
  nor _45940_ (_38462_, _38461_, _36466_);
  not _45941_ (_38463_, _38462_);
  not _45942_ (_38464_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _45943_ (_38465_, _18201_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _45944_ (_38466_, _38465_, _38464_);
  and _45945_ (_38467_, _38456_, _38438_);
  and _45946_ (_38468_, _38467_, _38443_);
  and _45947_ (_38469_, _38468_, _38466_);
  and _45948_ (_38470_, _38459_, _18201_);
  and _45949_ (_38471_, _38458_, _18201_);
  nor _45950_ (_38472_, _38471_, _38470_);
  nor _45951_ (_38473_, _38472_, _36444_);
  nor _45952_ (_38474_, _38473_, _38469_);
  and _45953_ (_38475_, _38474_, _38463_);
  nor _45954_ (_38476_, _38475_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45955_ (_38477_, _38476_, _36433_);
  and _45956_ (_38478_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _45957_ (_38479_, _38006_);
  nor _45958_ (_38480_, _38479_, _38270_);
  and _45959_ (_38481_, _38480_, _38455_);
  and _45960_ (_38482_, _37709_, _37470_);
  and _45961_ (_38483_, _38482_, _37219_);
  and _45962_ (_38484_, _38483_, _36967_);
  and _45963_ (_38485_, _38484_, _38481_);
  not _45964_ (_38486_, _38485_);
  and _45965_ (_38487_, _38270_, _38455_);
  and _45966_ (_38488_, _38487_, _36967_);
  and _45967_ (_38489_, _38488_, _37742_);
  not _45968_ (_38490_, _38481_);
  and _45969_ (_38491_, _37742_, _36956_);
  nor _45970_ (_38492_, _38491_, _38449_);
  nor _45971_ (_38493_, _38492_, _38490_);
  nor _45972_ (_38494_, _38493_, _38489_);
  and _45973_ (_38495_, _38494_, _38486_);
  nor _45974_ (_38496_, _37709_, _37470_);
  and _45975_ (_38497_, _38496_, _37219_);
  not _45976_ (_38498_, _37219_);
  and _45977_ (_38499_, _38443_, _38498_);
  and _45978_ (_38500_, _38499_, _36956_);
  nor _45979_ (_38501_, _38500_, _38497_);
  nor _45980_ (_38502_, _38501_, _38490_);
  not _45981_ (_38503_, _38502_);
  and _45982_ (_38504_, _38439_, _38479_);
  and _45983_ (_38505_, _38504_, _38497_);
  not _45984_ (_38506_, _38505_);
  and _45985_ (_38507_, _38496_, _38498_);
  and _45986_ (_38508_, _38507_, _36967_);
  and _45987_ (_38509_, _38508_, _38481_);
  and _45988_ (_38510_, _37753_, _38437_);
  nor _45989_ (_38511_, _38510_, _38509_);
  and _45990_ (_38512_, _38511_, _38506_);
  and _45991_ (_38513_, _38512_, _38503_);
  and _45992_ (_38514_, _38444_, _36967_);
  and _45993_ (_38515_, _38514_, _38481_);
  and _45994_ (_38516_, _38482_, _38498_);
  and _45995_ (_38517_, _38516_, _36967_);
  and _45996_ (_38518_, _38517_, _38481_);
  nor _45997_ (_38519_, _38518_, _38515_);
  and _45998_ (_38520_, _38516_, _36956_);
  and _45999_ (_38521_, _38520_, _38504_);
  and _46000_ (_38522_, _37753_, _38504_);
  nor _46001_ (_38523_, _38522_, _38521_);
  and _46002_ (_38524_, _38523_, _38519_);
  and _46003_ (_38525_, _38524_, _38513_);
  and _46004_ (_38526_, _38525_, _38495_);
  and _46005_ (_38527_, _38499_, _36967_);
  and _46006_ (_38528_, _38527_, _38439_);
  not _46007_ (_38529_, _38528_);
  and _46008_ (_38530_, _38507_, _36956_);
  and _46009_ (_38531_, _38530_, _38481_);
  and _46010_ (_38532_, _38467_, _38491_);
  nor _46011_ (_38533_, _38532_, _38531_);
  and _46012_ (_38534_, _38533_, _38529_);
  and _46013_ (_38535_, _38445_, _38504_);
  and _46014_ (_38536_, _38520_, _38481_);
  nor _46015_ (_38537_, _38536_, _38535_);
  and _46016_ (_38538_, _38537_, _38534_);
  and _46017_ (_38539_, _38467_, _37753_);
  and _46018_ (_38540_, _38527_, _38481_);
  nor _46019_ (_38541_, _38540_, _38539_);
  and _46020_ (_38542_, _38504_, _38491_);
  and _46021_ (_38543_, _38517_, _38504_);
  nor _46022_ (_38544_, _38543_, _38542_);
  and _46023_ (_38545_, _38544_, _38541_);
  and _46024_ (_38546_, _38545_, _38538_);
  and _46025_ (_38547_, _38453_, _38504_);
  and _46026_ (_38548_, _38439_, _38500_);
  nor _46027_ (_38549_, _38548_, _38547_);
  and _46028_ (_38550_, _38504_, _38449_);
  and _46029_ (_38551_, _38453_, _38481_);
  nor _46030_ (_38552_, _38551_, _38550_);
  and _46031_ (_38553_, _38552_, _38549_);
  and _46032_ (_38554_, _38497_, _36956_);
  and _46033_ (_38555_, _38554_, _38467_);
  not _46034_ (_38556_, _38555_);
  and _46035_ (_38557_, _38497_, _36967_);
  and _46036_ (_38558_, _38557_, _38467_);
  and _46037_ (_38559_, _38467_, _38530_);
  nor _46038_ (_38560_, _38559_, _38558_);
  and _46039_ (_38561_, _38560_, _38556_);
  and _46040_ (_38562_, _38467_, _38516_);
  and _46041_ (_38563_, _38514_, _38439_);
  nor _46042_ (_38564_, _38563_, _38562_);
  and _46043_ (_38565_, _38564_, _38561_);
  and _46044_ (_38566_, _38565_, _38553_);
  and _46045_ (_38567_, _38566_, _38546_);
  and _46046_ (_38568_, _38567_, _38526_);
  nor _46047_ (_38569_, _38568_, _36466_);
  and _46048_ (_38570_, \oc8051_top_1.oc8051_decoder1.state [0], _18201_);
  and _46049_ (_38571_, _38570_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _46050_ (_38572_, _38571_, _38505_);
  nor _46051_ (_38573_, _38572_, _38469_);
  not _46052_ (_38574_, _38573_);
  nor _46053_ (_38575_, _38574_, _38569_);
  nor _46054_ (_38576_, _38575_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46055_ (_38577_, _38576_, _38478_);
  and _46056_ (_38578_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _46057_ (_38579_, _38270_, _38414_);
  nor _46058_ (_38580_, _36967_, _38437_);
  and _46059_ (_38581_, _38580_, _38579_);
  and _46060_ (_38582_, _38581_, _38499_);
  and _46061_ (_38583_, _38497_, _38487_);
  or _46062_ (_38584_, _38583_, _38582_);
  not _46063_ (_38585_, _38584_);
  and _46064_ (_38586_, _38453_, _38487_);
  nor _46065_ (_38587_, _38586_, _38505_);
  and _46066_ (_38588_, _38581_, _37742_);
  and _46067_ (_38589_, _38507_, _38487_);
  nor _46068_ (_38590_, _38589_, _38588_);
  not _46069_ (_38591_, _38590_);
  or _46070_ (_38592_, _38499_, _38483_);
  and _46071_ (_38593_, _38592_, _38488_);
  nor _46072_ (_38594_, _38593_, _38591_);
  and _46073_ (_38595_, _38594_, _38587_);
  and _46074_ (_38596_, _38595_, _38585_);
  and _46075_ (_38597_, _38562_, _36956_);
  not _46076_ (_38598_, _38597_);
  and _46077_ (_38599_, _38516_, _38487_);
  and _46078_ (_38600_, _38581_, _38448_);
  nor _46079_ (_38601_, _38600_, _38599_);
  not _46080_ (_38602_, _38601_);
  and _46081_ (_38603_, _38514_, _38487_);
  nor _46082_ (_38604_, _38603_, _38602_);
  and _46083_ (_38605_, _38604_, _38598_);
  and _46084_ (_38606_, _38605_, _38452_);
  and _46085_ (_38607_, _38606_, _38596_);
  nor _46086_ (_38608_, _38607_, _36466_);
  and _46087_ (_38609_, _38466_, _38444_);
  and _46088_ (_38610_, _38609_, _38467_);
  or _46089_ (_38611_, _38610_, _38572_);
  nor _46090_ (_38612_, _38611_, _38608_);
  nor _46091_ (_38613_, _38612_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46092_ (_38614_, _38613_, _38578_);
  nor _46093_ (_38615_, _38614_, _38577_);
  and _46094_ (_38616_, _38615_, _38477_);
  and _46095_ (_09521_, _38616_, _43100_);
  and _46096_ (_38617_, _30651_, _27650_);
  and _46097_ (_38618_, _27825_, _27343_);
  and _46098_ (_38619_, _27211_, _27507_);
  and _46099_ (_38620_, _38619_, _38618_);
  and _46100_ (_38621_, _38620_, _32593_);
  and _46101_ (_38622_, _38621_, _26740_);
  and _46102_ (_38623_, _38622_, _38617_);
  not _46103_ (_38624_, _38623_);
  and _46104_ (_38625_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _46105_ (_38626_, _23628_, _18267_);
  and _46106_ (_38627_, _29602_, _23606_);
  nor _46107_ (_38628_, _30377_, _38627_);
  and _46108_ (_38629_, _38628_, _30345_);
  and _46109_ (_38630_, _38629_, _38626_);
  and _46110_ (_38631_, _38630_, _31568_);
  nor _46111_ (_38632_, _38631_, _19481_);
  not _46112_ (_38633_, _38632_);
  and _46113_ (_38634_, _38633_, _36065_);
  and _46114_ (_38635_, _38634_, _35934_);
  nor _46115_ (_38636_, _38635_, _38624_);
  nor _46116_ (_38637_, _38636_, _38625_);
  and _46117_ (_38638_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _46118_ (_38639_, _38631_, _20521_);
  not _46119_ (_38640_, _38639_);
  and _46120_ (_38641_, _38640_, _35346_);
  and _46121_ (_38642_, _38641_, _35193_);
  nor _46122_ (_38643_, _38642_, _38624_);
  nor _46123_ (_38644_, _38643_, _38638_);
  and _46124_ (_38645_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _46125_ (_38646_, _38631_, _20695_);
  not _46126_ (_38647_, _38646_);
  and _46127_ (_38648_, _38647_, _34366_);
  and _46128_ (_38649_, _38648_, _34475_);
  and _46129_ (_38650_, _38649_, _34333_);
  nor _46130_ (_38651_, _38650_, _38624_);
  nor _46131_ (_38652_, _38651_, _38645_);
  and _46132_ (_38653_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _46133_ (_38654_, _38631_, _21054_);
  not _46134_ (_38655_, _38654_);
  and _46135_ (_38656_, _38655_, _33637_);
  and _46136_ (_38657_, _38656_, _33605_);
  and _46137_ (_38658_, _38657_, _33921_);
  nor _46138_ (_38659_, _38658_, _38624_);
  nor _46139_ (_38660_, _38659_, _38653_);
  and _46140_ (_38661_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _46141_ (_38662_, _38631_, _21555_);
  not _46142_ (_38663_, _38662_);
  and _46143_ (_38664_, _38663_, _32963_);
  and _46144_ (_38665_, _38664_, _32843_);
  nor _46145_ (_38666_, _38665_, _38624_);
  nor _46146_ (_38667_, _38666_, _38661_);
  and _46147_ (_38668_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _46148_ (_38669_, _38631_, _21381_);
  not _46149_ (_38670_, _38669_);
  and _46150_ (_38671_, _38670_, _32244_);
  and _46151_ (_38672_, _38671_, _32440_);
  nor _46152_ (_38673_, _38672_, _38624_);
  nor _46153_ (_38674_, _38673_, _38668_);
  and _46154_ (_38675_, _38617_, _26740_);
  and _46155_ (_38676_, _38675_, _38621_);
  nor _46156_ (_38677_, _38676_, _26926_);
  nor _46157_ (_38678_, _38631_, _21925_);
  not _46158_ (_38679_, _38678_);
  and _46159_ (_38680_, _38679_, _31656_);
  and _46160_ (_38681_, _38680_, _31634_);
  and _46161_ (_38682_, _38681_, _31546_);
  not _46162_ (_38683_, _38682_);
  and _46163_ (_38684_, _38683_, _38623_);
  nor _46164_ (_38685_, _38684_, _38677_);
  and _46165_ (_38686_, _38685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _46166_ (_38687_, _38686_, _38674_);
  and _46167_ (_38688_, _38687_, _38667_);
  and _46168_ (_38689_, _38688_, _38660_);
  and _46169_ (_38690_, _38689_, _38652_);
  and _46170_ (_38691_, _38690_, _38644_);
  and _46171_ (_38692_, _38691_, _38637_);
  nor _46172_ (_38693_, _38676_, _27365_);
  nand _46173_ (_38694_, _38693_, _38692_);
  or _46174_ (_38695_, _38693_, _38692_);
  and _46175_ (_38696_, _38695_, _27069_);
  and _46176_ (_38697_, _38696_, _38694_);
  or _46177_ (_38698_, _38676_, _27409_);
  or _46178_ (_38699_, _38698_, _38697_);
  nor _46179_ (_38700_, _38631_, _20325_);
  not _46180_ (_38701_, _38700_);
  and _46181_ (_38702_, _38701_, _30323_);
  and _46182_ (_38703_, _38702_, _30268_);
  and _46183_ (_38704_, _38703_, _29984_);
  nand _46184_ (_38705_, _38704_, _38676_);
  and _46185_ (_38706_, _38705_, _38699_);
  and _46186_ (_09542_, _38706_, _43100_);
  not _46187_ (_38707_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _46188_ (_38708_, _38685_, _38707_);
  nor _46189_ (_38709_, _38685_, _38707_);
  nor _46190_ (_38710_, _38709_, _38708_);
  and _46191_ (_38711_, _38710_, _27069_);
  nor _46192_ (_38712_, _38711_, _26937_);
  nor _46193_ (_38713_, _38712_, _38623_);
  nor _46194_ (_38714_, _38713_, _38684_);
  nand _46195_ (_10698_, _38714_, _43100_);
  nor _46196_ (_38715_, _38686_, _38674_);
  nor _46197_ (_38716_, _38715_, _38687_);
  nor _46198_ (_38717_, _38716_, _26487_);
  nor _46199_ (_38718_, _38717_, _26784_);
  nor _46200_ (_38719_, _38718_, _38623_);
  nor _46201_ (_38720_, _38719_, _38673_);
  nand _46202_ (_10709_, _38720_, _43100_);
  nor _46203_ (_38721_, _38687_, _38667_);
  nor _46204_ (_38722_, _38721_, _38688_);
  nor _46205_ (_38723_, _38722_, _26487_);
  nor _46206_ (_38724_, _38723_, _26542_);
  nor _46207_ (_38725_, _38724_, _38623_);
  nor _46208_ (_38726_, _38725_, _38666_);
  nand _46209_ (_10720_, _38726_, _43100_);
  nor _46210_ (_38727_, _38688_, _38660_);
  nor _46211_ (_38728_, _38727_, _38689_);
  nor _46212_ (_38729_, _38728_, _26487_);
  nor _46213_ (_38730_, _38729_, _27584_);
  nor _46214_ (_38731_, _38730_, _38623_);
  nor _46215_ (_38732_, _38731_, _38659_);
  nor _46216_ (_10731_, _38732_, rst);
  nor _46217_ (_38733_, _38689_, _38652_);
  nor _46218_ (_38734_, _38733_, _38690_);
  nor _46219_ (_38735_, _38734_, _26487_);
  nor _46220_ (_38736_, _38735_, _27760_);
  nor _46221_ (_38737_, _38736_, _38623_);
  nor _46222_ (_38738_, _38737_, _38651_);
  nor _46223_ (_10742_, _38738_, rst);
  nor _46224_ (_38739_, _38690_, _38644_);
  nor _46225_ (_38740_, _38739_, _38691_);
  nor _46226_ (_38741_, _38740_, _26487_);
  nor _46227_ (_38742_, _38741_, _27255_);
  nor _46228_ (_38743_, _38742_, _38623_);
  nor _46229_ (_38744_, _38743_, _38643_);
  nor _46230_ (_10753_, _38744_, rst);
  nor _46231_ (_38745_, _38691_, _38637_);
  nor _46232_ (_38746_, _38745_, _38692_);
  nor _46233_ (_38747_, _38746_, _26487_);
  nor _46234_ (_38748_, _38747_, _27102_);
  nor _46235_ (_38749_, _38748_, _38623_);
  nor _46236_ (_38750_, _38749_, _38636_);
  nor _46237_ (_10764_, _38750_, rst);
  and _46238_ (_38751_, _38620_, _34052_);
  nand _46239_ (_38752_, _38751_, _38617_);
  nor _46240_ (_38753_, _38752_, _30574_);
  and _46241_ (_38754_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18201_);
  and _46242_ (_38755_, _38754_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46243_ (_38756_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _46244_ (_38757_, _38756_, _38755_);
  or _46245_ (_38758_, _38757_, _38753_);
  nor _46246_ (_38759_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _46247_ (_38760_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _46248_ (_38761_, _38760_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46249_ (_38762_, _38761_, _38759_);
  nor _46250_ (_38763_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _46251_ (_38764_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _46252_ (_38765_, _38764_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46253_ (_38766_, _38765_, _38763_);
  nor _46254_ (_38767_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _46255_ (_38768_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _46256_ (_38769_, _38768_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46257_ (_38770_, _38769_, _38767_);
  nor _46258_ (_38771_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not _46259_ (_38772_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _46260_ (_38773_, _38772_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46261_ (_38774_, _38773_, _38771_);
  nor _46262_ (_38775_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _46263_ (_38776_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _46264_ (_38777_, _38776_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46265_ (_38778_, _38777_, _38775_);
  not _46266_ (_38779_, _38778_);
  nor _46267_ (_38780_, _38779_, _30716_);
  nor _46268_ (_38781_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not _46269_ (_38782_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _46270_ (_38783_, _38782_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46271_ (_38784_, _38783_, _38781_);
  and _46272_ (_38785_, _38784_, _38780_);
  nor _46273_ (_38786_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not _46274_ (_38787_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _46275_ (_38788_, _38787_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46276_ (_38789_, _38788_, _38786_);
  and _46277_ (_38790_, _38789_, _38785_);
  and _46278_ (_38791_, _38790_, _38774_);
  nor _46279_ (_38792_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not _46280_ (_38793_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _46281_ (_38794_, _38793_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46282_ (_38795_, _38794_, _38792_);
  and _46283_ (_38796_, _38795_, _38791_);
  and _46284_ (_38797_, _38796_, _38770_);
  and _46285_ (_38798_, _38797_, _38766_);
  or _46286_ (_38799_, _38798_, _38762_);
  nand _46287_ (_38800_, _38798_, _38762_);
  and _46288_ (_38801_, _38800_, _38799_);
  and _46289_ (_38802_, _38801_, _29613_);
  not _46290_ (_38803_, _38802_);
  and _46291_ (_38804_, _23320_, _18267_);
  and _46292_ (_38805_, _29733_, _20336_);
  and _46293_ (_38806_, _38805_, _28374_);
  and _46294_ (_38807_, _38806_, _28407_);
  and _46295_ (_38808_, _38807_, _28450_);
  and _46296_ (_38809_, _38808_, _29064_);
  nor _46297_ (_38810_, _38809_, _29755_);
  and _46298_ (_38811_, _29010_, _18836_);
  nor _46299_ (_38812_, _38811_, _38810_);
  and _46300_ (_38813_, _29820_, _20325_);
  and _46301_ (_38814_, _19655_, _18671_);
  and _46302_ (_38815_, _19977_, _18990_);
  and _46303_ (_38816_, _38815_, _38814_);
  and _46304_ (_38817_, _38816_, _38813_);
  and _46305_ (_38818_, _19807_, _18836_);
  and _46306_ (_38819_, _38818_, _38817_);
  nor _46307_ (_38820_, _38819_, _29010_);
  and _46308_ (_38821_, _29010_, _19807_);
  nor _46309_ (_38822_, _38821_, _38820_);
  and _46310_ (_38823_, _38822_, _38812_);
  nor _46311_ (_38824_, _29010_, _19166_);
  and _46312_ (_38825_, _29010_, _19166_);
  nor _46313_ (_38826_, _38825_, _38824_);
  and _46314_ (_38827_, _38826_, _38823_);
  and _46315_ (_38828_, _38827_, _29897_);
  nor _46316_ (_38829_, _38827_, _29897_);
  nor _46317_ (_38830_, _38829_, _38828_);
  and _46318_ (_38831_, _38830_, _29668_);
  and _46319_ (_38832_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and _46320_ (_38833_, _29010_, _29897_);
  nor _46321_ (_38834_, _38833_, _30825_);
  nor _46322_ (_38835_, _38834_, _29951_);
  nor _46323_ (_38836_, _31141_, _21054_);
  nor _46324_ (_38837_, _30388_, _20151_);
  or _46325_ (_38838_, _38837_, _38836_);
  or _46326_ (_38839_, _38838_, _38835_);
  nor _46327_ (_38840_, _38839_, _38832_);
  not _46328_ (_38841_, _38840_);
  nor _46329_ (_38842_, _38841_, _38831_);
  not _46330_ (_38843_, _38842_);
  nor _46331_ (_38844_, _38843_, _38804_);
  and _46332_ (_38845_, _38844_, _38803_);
  nand _46333_ (_38846_, _38845_, _38755_);
  and _46334_ (_38847_, _38846_, _43100_);
  and _46335_ (_12715_, _38847_, _38758_);
  and _46336_ (_38848_, _38620_, _33344_);
  and _46337_ (_38849_, _38848_, _38617_);
  nor _46338_ (_38850_, _38849_, _38755_);
  not _46339_ (_38851_, _38850_);
  nand _46340_ (_38852_, _38851_, _30574_);
  or _46341_ (_38853_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _46342_ (_38854_, _38853_, _43100_);
  and _46343_ (_12736_, _38854_, _38852_);
  nor _46344_ (_38855_, _38752_, _31808_);
  and _46345_ (_38856_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _46346_ (_38857_, _38856_, _38755_);
  or _46347_ (_38858_, _38857_, _38855_);
  and _46348_ (_38859_, _25897_, _23628_);
  not _46349_ (_38860_, _38859_);
  and _46350_ (_38861_, _38779_, _30716_);
  nor _46351_ (_38862_, _38861_, _38780_);
  and _46352_ (_38863_, _38862_, _29613_);
  nor _46353_ (_38864_, _30825_, _29930_);
  not _46354_ (_38865_, _38864_);
  nor _46355_ (_38866_, _38865_, _29842_);
  nor _46356_ (_38867_, _38866_, _28374_);
  and _46357_ (_38868_, _38866_, _28374_);
  or _46358_ (_38869_, _38868_, _32799_);
  nor _46359_ (_38870_, _38869_, _38867_);
  nor _46360_ (_38871_, _30388_, _18990_);
  and _46361_ (_38872_, _23098_, _18267_);
  nor _46362_ (_38873_, _31141_, _20695_);
  nor _46363_ (_38874_, _29951_, _21925_);
  or _46364_ (_38875_, _38874_, _38873_);
  or _46365_ (_38876_, _38875_, _38872_);
  nor _46366_ (_38877_, _38876_, _38871_);
  not _46367_ (_38878_, _38877_);
  nor _46368_ (_38879_, _38878_, _38870_);
  not _46369_ (_38880_, _38879_);
  nor _46370_ (_38881_, _38880_, _38863_);
  and _46371_ (_38882_, _38881_, _38860_);
  nand _46372_ (_38883_, _38882_, _38755_);
  and _46373_ (_38884_, _38883_, _43100_);
  and _46374_ (_13649_, _38884_, _38858_);
  nor _46375_ (_38885_, _38752_, _32495_);
  and _46376_ (_38886_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _46377_ (_38887_, _38886_, _38755_);
  or _46378_ (_38888_, _38887_, _38885_);
  nor _46379_ (_38889_, _38784_, _38780_);
  not _46380_ (_38890_, _38889_);
  nor _46381_ (_38891_, _38785_, _29624_);
  and _46382_ (_38892_, _38891_, _38890_);
  not _46383_ (_38893_, _38892_);
  and _46384_ (_38894_, _24911_, _23628_);
  nor _46385_ (_38895_, _20325_, _18990_);
  and _46386_ (_38896_, _38895_, _29733_);
  and _46387_ (_38897_, _38896_, _29010_);
  and _46388_ (_38898_, _38813_, _18990_);
  and _46389_ (_38899_, _38898_, _29755_);
  nor _46390_ (_38900_, _38899_, _38897_);
  nor _46391_ (_38901_, _38900_, _28407_);
  and _46392_ (_38902_, _38900_, _28407_);
  nor _46393_ (_38903_, _38902_, _38901_);
  nor _46394_ (_38904_, _38903_, _32799_);
  nor _46395_ (_38905_, _30388_, _19977_);
  and _46396_ (_38906_, _23130_, _18267_);
  nor _46397_ (_38907_, _31141_, _20521_);
  nor _46398_ (_38908_, _29951_, _21381_);
  or _46399_ (_38909_, _38908_, _38907_);
  or _46400_ (_38910_, _38909_, _38906_);
  nor _46401_ (_38911_, _38910_, _38905_);
  not _46402_ (_38912_, _38911_);
  nor _46403_ (_38913_, _38912_, _38904_);
  not _46404_ (_38914_, _38913_);
  nor _46405_ (_38915_, _38914_, _38894_);
  and _46406_ (_38916_, _38915_, _38893_);
  nand _46407_ (_38917_, _38916_, _38755_);
  and _46408_ (_38918_, _38917_, _43100_);
  and _46409_ (_13660_, _38918_, _38888_);
  nor _46410_ (_38919_, _38752_, _33202_);
  and _46411_ (_38920_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _46412_ (_38921_, _38920_, _38755_);
  or _46413_ (_38922_, _38921_, _38919_);
  nor _46414_ (_38923_, _38789_, _38785_);
  nor _46415_ (_38924_, _38923_, _38790_);
  and _46416_ (_38925_, _38924_, _29613_);
  not _46417_ (_38926_, _38925_);
  and _46418_ (_38927_, _38898_, _19977_);
  and _46419_ (_38928_, _38927_, _29755_);
  and _46420_ (_38929_, _38896_, _28407_);
  and _46421_ (_38930_, _38929_, _29010_);
  nor _46422_ (_38931_, _38930_, _38928_);
  and _46423_ (_38932_, _38931_, _18671_);
  nor _46424_ (_38933_, _38931_, _18671_);
  nor _46425_ (_38934_, _38933_, _38932_);
  and _46426_ (_38935_, _38934_, _29668_);
  not _46427_ (_38936_, _38935_);
  nor _46428_ (_38937_, _29951_, _21555_);
  and _46429_ (_38938_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _46430_ (_38939_, _38938_, _38937_);
  and _46431_ (_38940_, _23162_, _18267_);
  nor _46432_ (_38941_, _31141_, _19481_);
  nor _46433_ (_38942_, _30388_, _18671_);
  or _46434_ (_38943_, _38942_, _38941_);
  nor _46435_ (_38944_, _38943_, _38940_);
  and _46436_ (_38945_, _38944_, _38939_);
  and _46437_ (_38946_, _38945_, _38936_);
  and _46438_ (_38947_, _38946_, _38926_);
  nand _46439_ (_38948_, _38947_, _38755_);
  and _46440_ (_38949_, _38948_, _43100_);
  and _46441_ (_13671_, _38949_, _38922_);
  nor _46442_ (_38950_, _38752_, _33953_);
  and _46443_ (_38951_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _46444_ (_38952_, _38951_, _38755_);
  or _46445_ (_38953_, _38952_, _38950_);
  nor _46446_ (_38954_, _38790_, _38774_);
  nor _46447_ (_38955_, _38954_, _38791_);
  and _46448_ (_38956_, _38955_, _29613_);
  not _46449_ (_38957_, _38956_);
  nor _46450_ (_38958_, _38808_, _29064_);
  not _46451_ (_38959_, _38958_);
  and _46452_ (_38960_, _38959_, _38810_);
  and _46453_ (_38961_, _38927_, _18671_);
  nor _46454_ (_38962_, _38961_, _19655_);
  nor _46455_ (_38963_, _38962_, _38817_);
  nor _46456_ (_38964_, _38963_, _29010_);
  nor _46457_ (_38965_, _38964_, _38960_);
  nor _46458_ (_38966_, _38965_, _32799_);
  nor _46459_ (_38967_, _30388_, _19655_);
  or _46460_ (_38968_, _38967_, _31142_);
  nor _46461_ (_38969_, _38968_, _38966_);
  and _46462_ (_38970_, _23193_, _18267_);
  nor _46463_ (_38971_, _29951_, _21054_);
  and _46464_ (_38972_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _46465_ (_38973_, _38972_, _38971_);
  nor _46466_ (_38974_, _38973_, _38970_);
  and _46467_ (_38975_, _38974_, _38969_);
  and _46468_ (_38976_, _38975_, _38957_);
  nand _46469_ (_38977_, _38976_, _38755_);
  and _46470_ (_38978_, _38977_, _43100_);
  and _46471_ (_13682_, _38978_, _38953_);
  nor _46472_ (_38979_, _38752_, _34693_);
  and _46473_ (_38980_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _46474_ (_38981_, _38980_, _38755_);
  or _46475_ (_38982_, _38981_, _38979_);
  nor _46476_ (_38983_, _38795_, _38791_);
  nor _46477_ (_38984_, _38983_, _38796_);
  and _46478_ (_38985_, _38984_, _29613_);
  not _46479_ (_38986_, _38985_);
  and _46480_ (_38987_, _23225_, _18267_);
  nor _46481_ (_38988_, _38817_, _29010_);
  nor _46482_ (_38989_, _38988_, _38810_);
  nor _46483_ (_38990_, _38989_, _28100_);
  and _46484_ (_38991_, _38989_, _28100_);
  nor _46485_ (_38992_, _38991_, _38990_);
  and _46486_ (_38993_, _38992_, _29668_);
  and _46487_ (_38994_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _46488_ (_38995_, _29010_, _20706_);
  or _46489_ (_38996_, _38995_, _29951_);
  nor _46490_ (_38997_, _38996_, _38811_);
  nor _46491_ (_38998_, _31141_, _21925_);
  nor _46492_ (_38999_, _30388_, _18836_);
  or _46493_ (_39000_, _38999_, _38998_);
  or _46494_ (_39001_, _39000_, _38997_);
  nor _46495_ (_39002_, _39001_, _38994_);
  not _46496_ (_39003_, _39002_);
  nor _46497_ (_39004_, _39003_, _38993_);
  not _46498_ (_39005_, _39004_);
  nor _46499_ (_39006_, _39005_, _38987_);
  and _46500_ (_39007_, _39006_, _38986_);
  nand _46501_ (_39008_, _39007_, _38755_);
  and _46502_ (_39009_, _39008_, _43100_);
  and _46503_ (_13693_, _39009_, _38982_);
  nor _46504_ (_39010_, _38752_, _35520_);
  and _46505_ (_39011_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _46506_ (_39012_, _39011_, _38755_);
  or _46507_ (_39013_, _39012_, _39010_);
  nor _46508_ (_39014_, _38796_, _38770_);
  not _46509_ (_39015_, _39014_);
  nor _46510_ (_39016_, _38797_, _29624_);
  and _46511_ (_39017_, _39016_, _39015_);
  not _46512_ (_39018_, _39017_);
  and _46513_ (_39019_, _23257_, _18267_);
  and _46514_ (_39020_, _38817_, _18836_);
  nor _46515_ (_39021_, _39020_, _29010_);
  not _46516_ (_39022_, _39021_);
  and _46517_ (_39023_, _39022_, _38812_);
  and _46518_ (_39024_, _39023_, _19807_);
  nor _46519_ (_39025_, _39023_, _19807_);
  nor _46520_ (_39026_, _39025_, _39024_);
  nor _46521_ (_39027_, _39026_, _32799_);
  and _46522_ (_39028_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _46523_ (_39029_, _29010_, _20532_);
  or _46524_ (_39030_, _39029_, _29951_);
  nor _46525_ (_39031_, _39030_, _38821_);
  nor _46526_ (_39032_, _31141_, _21381_);
  nor _46527_ (_39033_, _30388_, _19807_);
  or _46528_ (_39034_, _39033_, _39032_);
  or _46529_ (_39035_, _39034_, _39031_);
  nor _46530_ (_39036_, _39035_, _39028_);
  not _46531_ (_39037_, _39036_);
  nor _46532_ (_39038_, _39037_, _39027_);
  not _46533_ (_39039_, _39038_);
  nor _46534_ (_39040_, _39039_, _39019_);
  and _46535_ (_39041_, _39040_, _39018_);
  nand _46536_ (_39042_, _39041_, _38755_);
  and _46537_ (_39043_, _39042_, _43100_);
  and _46538_ (_13704_, _39043_, _39013_);
  nor _46539_ (_39044_, _38752_, _36239_);
  and _46540_ (_39045_, _38752_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _46541_ (_39046_, _39045_, _38755_);
  or _46542_ (_39047_, _39046_, _39044_);
  nor _46543_ (_39048_, _38797_, _38766_);
  not _46544_ (_39049_, _39048_);
  nor _46545_ (_39050_, _38798_, _29624_);
  and _46546_ (_39051_, _39050_, _39049_);
  not _46547_ (_39052_, _39051_);
  and _46548_ (_39053_, _23288_, _18267_);
  and _46549_ (_39054_, _38823_, _19166_);
  nor _46550_ (_39055_, _38823_, _19166_);
  nor _46551_ (_39056_, _39055_, _39054_);
  nor _46552_ (_39057_, _39056_, _32799_);
  and _46553_ (_39058_, _23628_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _46554_ (_39059_, _29010_, _19492_);
  or _46555_ (_39060_, _39059_, _29951_);
  nor _46556_ (_39061_, _39060_, _38825_);
  nor _46557_ (_39062_, _31141_, _21555_);
  nor _46558_ (_39063_, _30388_, _19166_);
  or _46559_ (_39064_, _39063_, _39062_);
  or _46560_ (_39065_, _39064_, _39061_);
  nor _46561_ (_39066_, _39065_, _39058_);
  not _46562_ (_39067_, _39066_);
  nor _46563_ (_39068_, _39067_, _39057_);
  not _46564_ (_39069_, _39068_);
  nor _46565_ (_39070_, _39069_, _39053_);
  and _46566_ (_39071_, _39070_, _39052_);
  nand _46567_ (_39072_, _39071_, _38755_);
  and _46568_ (_39073_, _39072_, _43100_);
  and _46569_ (_13715_, _39073_, _39047_);
  nand _46570_ (_39074_, _38851_, _31808_);
  or _46571_ (_39075_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _46572_ (_39076_, _39075_, _43100_);
  and _46573_ (_13726_, _39076_, _39074_);
  nand _46574_ (_39077_, _38851_, _32495_);
  or _46575_ (_39078_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _46576_ (_39079_, _39078_, _43100_);
  and _46577_ (_13737_, _39079_, _39077_);
  nand _46578_ (_39080_, _38851_, _33202_);
  or _46579_ (_39081_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _46580_ (_39082_, _39081_, _43100_);
  and _46581_ (_13748_, _39082_, _39080_);
  nand _46582_ (_39083_, _38851_, _33953_);
  or _46583_ (_39084_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _46584_ (_39085_, _39084_, _43100_);
  and _46585_ (_13758_, _39085_, _39083_);
  nand _46586_ (_39086_, _38851_, _34693_);
  or _46587_ (_39087_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _46588_ (_39088_, _39087_, _43100_);
  and _46589_ (_13769_, _39088_, _39086_);
  nand _46590_ (_39089_, _38851_, _35520_);
  or _46591_ (_39090_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _46592_ (_39091_, _39090_, _43100_);
  and _46593_ (_13780_, _39091_, _39089_);
  nand _46594_ (_39092_, _38851_, _36239_);
  or _46595_ (_39093_, _38851_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _46596_ (_39094_, _39093_, _43100_);
  and _46597_ (_13791_, _39094_, _39092_);
  not _46598_ (_39095_, _27343_);
  nor _46599_ (_39096_, _39095_, _27211_);
  and _46600_ (_39097_, _39096_, _31351_);
  and _46601_ (_39098_, _39097_, _27847_);
  not _46602_ (_39099_, _31308_);
  nor _46603_ (_39100_, _39099_, _31265_);
  not _46604_ (_39101_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _46605_ (_39102_, _31308_, _39101_);
  or _46606_ (_39103_, _39102_, _39100_);
  and _46607_ (_39104_, _39103_, _39098_);
  nor _46608_ (_39105_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _46609_ (_39106_, _39105_);
  nand _46610_ (_39107_, _39106_, _31265_);
  and _46611_ (_39108_, _39105_, _39101_);
  nor _46612_ (_39109_, _39108_, _39098_);
  and _46613_ (_39110_, _39109_, _39107_);
  nor _46614_ (_39111_, _27825_, _39095_);
  nor _46615_ (_39112_, _27211_, _27496_);
  and _46616_ (_39113_, _38617_, _27003_);
  and _46617_ (_39114_, _39113_, _39112_);
  and _46618_ (_39115_, _39114_, _39111_);
  or _46619_ (_39116_, _39115_, _39110_);
  or _46620_ (_39117_, _39116_, _39104_);
  nand _46621_ (_39118_, _39115_, _38704_);
  and _46622_ (_39119_, _39118_, _43100_);
  and _46623_ (_15195_, _39119_, _39117_);
  and _46624_ (_39120_, _39098_, _32604_);
  nand _46625_ (_39121_, _39120_, _31265_);
  not _46626_ (_39122_, _39115_);
  or _46627_ (_39123_, _39120_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _46628_ (_39124_, _39123_, _39122_);
  and _46629_ (_39125_, _39124_, _39121_);
  nor _46630_ (_39126_, _39122_, _38672_);
  or _46631_ (_39127_, _39126_, _39125_);
  and _46632_ (_17376_, _39127_, _43100_);
  or _46633_ (_39128_, _23384_, _23352_);
  or _46634_ (_39129_, _39128_, _23415_);
  or _46635_ (_39130_, _39129_, _23468_);
  or _46636_ (_39131_, _39130_, _23490_);
  or _46637_ (_39132_, _39131_, _23532_);
  and _46638_ (_39133_, _39132_, _18267_);
  or _46639_ (_39134_, _30759_, _29163_);
  not _46640_ (_39135_, _30749_);
  nand _46641_ (_39136_, _39135_, _29163_);
  and _46642_ (_39137_, _39136_, _27935_);
  and _46643_ (_39138_, _39137_, _39134_);
  not _46644_ (_39139_, _27957_);
  nand _46645_ (_39140_, _29558_, _39139_);
  or _46646_ (_39141_, _29558_, _27978_);
  and _46647_ (_39142_, _29613_, _39141_);
  and _46648_ (_39143_, _39142_, _39140_);
  and _46649_ (_39144_, _38818_, _24812_);
  and _46650_ (_39145_, _38816_, _23628_);
  nand _46651_ (_39146_, _39145_, _39144_);
  nand _46652_ (_39147_, _39146_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _46653_ (_39148_, _39147_, _39143_);
  or _46654_ (_39149_, _39148_, _39138_);
  or _46655_ (_39150_, _39149_, _35726_);
  or _46656_ (_39151_, _39150_, _39133_);
  or _46657_ (_39152_, _39151_, _27902_);
  nor _46658_ (_39153_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _46659_ (_39154_, _39153_, _39098_);
  and _46660_ (_39155_, _39154_, _39152_);
  and _46661_ (_39156_, _33355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _46662_ (_39157_, _39156_, _33366_);
  and _46663_ (_39158_, _39157_, _39098_);
  or _46664_ (_39159_, _39158_, _39115_);
  or _46665_ (_39160_, _39159_, _39155_);
  nand _46666_ (_39161_, _39115_, _38665_);
  and _46667_ (_39162_, _39161_, _43100_);
  and _46668_ (_17387_, _39162_, _39160_);
  and _46669_ (_39163_, _39098_, _34052_);
  nand _46670_ (_39164_, _39163_, _31265_);
  or _46671_ (_39165_, _39163_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _46672_ (_39166_, _39165_, _39122_);
  and _46673_ (_39167_, _39166_, _39164_);
  nor _46674_ (_39168_, _39122_, _38658_);
  or _46675_ (_39169_, _39168_, _39167_);
  and _46676_ (_17398_, _39169_, _43100_);
  not _46677_ (_39170_, _39098_);
  or _46678_ (_39171_, _39170_, _34813_);
  and _46679_ (_39172_, _39171_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _46680_ (_39175_, _34802_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _46681_ (_39177_, _39175_, _34845_);
  and _46682_ (_39178_, _39177_, _39098_);
  or _46683_ (_39179_, _39178_, _39172_);
  and _46684_ (_39180_, _39179_, _39122_);
  nor _46685_ (_39181_, _39122_, _38650_);
  or _46686_ (_39182_, _39181_, _39180_);
  and _46687_ (_17409_, _39182_, _43100_);
  and _46688_ (_39183_, _39098_, _35607_);
  nand _46689_ (_39184_, _39183_, _31265_);
  or _46690_ (_39185_, _39183_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _46691_ (_39187_, _39185_, _39122_);
  and _46692_ (_39196_, _39187_, _39184_);
  nor _46693_ (_39202_, _39122_, _38642_);
  or _46694_ (_39208_, _39202_, _39196_);
  and _46695_ (_17420_, _39208_, _43100_);
  and _46696_ (_39211_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _46697_ (_39212_, _39211_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _46698_ (_39213_, _29119_, _27935_);
  and _46699_ (_39214_, _29613_, _29481_);
  nand _46700_ (_39215_, _30377_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _46701_ (_39216_, _39215_, _39211_);
  or _46702_ (_39217_, _39216_, _39214_);
  or _46703_ (_39218_, _39217_, _39213_);
  and _46704_ (_39219_, _39218_, _39212_);
  or _46705_ (_39220_, _39219_, _39098_);
  not _46706_ (_39221_, _36336_);
  nor _46707_ (_39222_, _39221_, _31265_);
  or _46708_ (_39223_, _36336_, _33496_);
  nand _46709_ (_39224_, _39223_, _39098_);
  or _46710_ (_39225_, _39224_, _39222_);
  and _46711_ (_39226_, _39225_, _39220_);
  or _46712_ (_39227_, _39226_, _39115_);
  nand _46713_ (_39228_, _39115_, _38635_);
  and _46714_ (_39229_, _39228_, _43100_);
  and _46715_ (_17431_, _39229_, _39227_);
  not _46716_ (_39230_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46717_ (_39231_, _38754_, _39230_);
  not _46718_ (_39232_, _39231_);
  nor _46719_ (_39233_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _46720_ (_39236_, _39233_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46721_ (_39237_, _27003_, _27650_);
  and _46722_ (_39238_, _27825_, _39095_);
  and _46723_ (_39239_, _39238_, _39112_);
  and _46724_ (_39240_, _39239_, _39237_);
  and _46725_ (_39241_, _39240_, _30651_);
  nor _46726_ (_39242_, _39241_, _39236_);
  nor _46727_ (_39243_, _39242_, _30574_);
  and _46728_ (_39244_, _27825_, _27650_);
  and _46729_ (_39245_, _39244_, _27354_);
  not _46730_ (_39246_, _31351_);
  nor _46731_ (_39247_, _39246_, _27496_);
  and _46732_ (_39248_, _39247_, _39245_);
  and _46733_ (_39249_, _39248_, _31308_);
  and _46734_ (_39250_, _39249_, _31265_);
  nor _46735_ (_39251_, _39249_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _46736_ (_39252_, _39251_);
  and _46737_ (_39253_, _39242_, _39232_);
  and _46738_ (_39254_, _39253_, _39252_);
  not _46739_ (_39255_, _39254_);
  nor _46740_ (_39256_, _39255_, _39250_);
  or _46741_ (_39257_, _39256_, _39243_);
  and _46742_ (_39258_, _39257_, _39232_);
  nor _46743_ (_39259_, _39232_, _38845_);
  or _46744_ (_39260_, _39259_, _39258_);
  and _46745_ (_18000_, _39260_, _43100_);
  nor _46746_ (_39261_, _39232_, _38882_);
  not _46747_ (_39262_, _39242_);
  and _46748_ (_39263_, _39262_, _31808_);
  not _46749_ (_39264_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _46750_ (_39265_, _39248_, _39264_);
  nor _46751_ (_39266_, _39265_, _39262_);
  not _46752_ (_39267_, _39266_);
  and _46753_ (_39268_, _31885_, _27003_);
  nor _46754_ (_39269_, _27003_, _39264_);
  nor _46755_ (_39270_, _39269_, _39268_);
  and _46756_ (_39271_, _39244_, _27507_);
  and _46757_ (_39272_, _31351_, _27354_);
  and _46758_ (_39274_, _39272_, _39271_);
  and _46759_ (_39278_, _39253_, _39274_);
  not _46760_ (_39284_, _39278_);
  nor _46761_ (_39289_, _39284_, _39270_);
  nor _46762_ (_39296_, _39289_, _39267_);
  nor _46763_ (_39304_, _39296_, _39231_);
  not _46764_ (_39312_, _39304_);
  nor _46765_ (_39313_, _39312_, _39263_);
  nor _46766_ (_39314_, _39313_, _39261_);
  nor _46767_ (_19851_, _39314_, rst);
  nor _46768_ (_39315_, _39242_, _32495_);
  and _46769_ (_39316_, _39248_, _32604_);
  and _46770_ (_39317_, _39316_, _31265_);
  nor _46771_ (_39318_, _39316_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not _46772_ (_39319_, _39318_);
  and _46773_ (_39320_, _39319_, _39253_);
  not _46774_ (_39321_, _39320_);
  nor _46775_ (_39322_, _39321_, _39317_);
  or _46776_ (_39323_, _39322_, _39315_);
  and _46777_ (_39324_, _39323_, _39232_);
  nor _46778_ (_39325_, _39232_, _38916_);
  or _46779_ (_39326_, _39325_, _39324_);
  and _46780_ (_19863_, _39326_, _43100_);
  nor _46781_ (_39327_, _39242_, _33202_);
  and _46782_ (_39328_, _39248_, _33344_);
  and _46783_ (_39329_, _39328_, _31265_);
  nor _46784_ (_39330_, _39328_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not _46785_ (_39331_, _39330_);
  and _46786_ (_39332_, _39331_, _39253_);
  not _46787_ (_39333_, _39332_);
  nor _46788_ (_39334_, _39333_, _39329_);
  or _46789_ (_39335_, _39334_, _39327_);
  and _46790_ (_39336_, _39335_, _39232_);
  nor _46791_ (_39337_, _39232_, _38947_);
  or _46792_ (_39338_, _39337_, _39336_);
  and _46793_ (_19875_, _39338_, _43100_);
  nor _46794_ (_39339_, _39232_, _38976_);
  and _46795_ (_39340_, _39262_, _33953_);
  not _46796_ (_39341_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _46797_ (_39342_, _39248_, _39341_);
  not _46798_ (_39343_, _39342_);
  not _46799_ (_39344_, _39248_);
  nor _46800_ (_39345_, _34052_, _39341_);
  nor _46801_ (_39346_, _39345_, _34062_);
  or _46802_ (_39352_, _39346_, _39344_);
  and _46803_ (_39363_, _39352_, _39242_);
  and _46804_ (_39364_, _39363_, _39343_);
  nor _46805_ (_39365_, _39364_, _39231_);
  not _46806_ (_39366_, _39365_);
  nor _46807_ (_39377_, _39366_, _39340_);
  nor _46808_ (_39383_, _39377_, _39339_);
  nor _46809_ (_19886_, _39383_, rst);
  nor _46810_ (_39384_, _39242_, _34693_);
  and _46811_ (_39385_, _39248_, _34791_);
  and _46812_ (_39386_, _39385_, _31265_);
  nor _46813_ (_39387_, _39385_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not _46814_ (_39388_, _39387_);
  and _46815_ (_39389_, _39388_, _39253_);
  not _46816_ (_39390_, _39389_);
  nor _46817_ (_39391_, _39390_, _39386_);
  or _46818_ (_39392_, _39391_, _39384_);
  and _46819_ (_39393_, _39392_, _39232_);
  nor _46820_ (_39394_, _39232_, _39007_);
  or _46821_ (_39395_, _39394_, _39393_);
  and _46822_ (_19898_, _39395_, _43100_);
  nor _46823_ (_39396_, _39242_, _35520_);
  and _46824_ (_39397_, _39248_, _35607_);
  and _46825_ (_39398_, _39397_, _31265_);
  nor _46826_ (_39399_, _39397_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not _46827_ (_39400_, _39399_);
  and _46828_ (_39401_, _39400_, _39253_);
  not _46829_ (_39402_, _39401_);
  nor _46830_ (_39403_, _39402_, _39398_);
  or _46831_ (_39404_, _39403_, _39396_);
  and _46832_ (_39405_, _39404_, _39232_);
  nor _46833_ (_39406_, _39232_, _39041_);
  or _46834_ (_39407_, _39406_, _39405_);
  and _46835_ (_19910_, _39407_, _43100_);
  nor _46836_ (_39408_, _39242_, _36239_);
  and _46837_ (_39409_, _39253_, _39344_);
  and _46838_ (_39410_, _39409_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _46839_ (_39411_, _39221_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _46840_ (_39412_, _39411_, _39222_);
  nor _46841_ (_39413_, _39412_, _39284_);
  nor _46842_ (_39414_, _39413_, _39410_);
  and _46843_ (_39415_, _39414_, _39232_);
  not _46844_ (_39416_, _39415_);
  nor _46845_ (_39417_, _39416_, _39408_);
  and _46846_ (_39418_, _39231_, _39071_);
  or _46847_ (_39419_, _39418_, _39417_);
  nor _46848_ (_19922_, _39419_, rst);
  and _46849_ (_39420_, _27343_, _27211_);
  and _46850_ (_39421_, _39271_, _39420_);
  and _46851_ (_39422_, _39421_, _31308_);
  nand _46852_ (_39423_, _39422_, _31265_);
  or _46853_ (_39424_, _39422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46854_ (_39425_, _39424_, _31351_);
  and _46855_ (_39426_, _39425_, _39423_);
  and _46856_ (_39427_, _38620_, _39237_);
  nand _46857_ (_39428_, _39427_, _38704_);
  or _46858_ (_39429_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46859_ (_39430_, _39429_, _30651_);
  and _46860_ (_39431_, _39430_, _39428_);
  not _46861_ (_39432_, _30640_);
  and _46862_ (_39433_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _46863_ (_39434_, _39433_, rst);
  or _46864_ (_39435_, _39434_, _39431_);
  or _46865_ (_31130_, _39435_, _39426_);
  and _46866_ (_39436_, _39420_, _27847_);
  and _46867_ (_39437_, _39436_, _31308_);
  nand _46868_ (_39438_, _39437_, _31265_);
  or _46869_ (_39439_, _39437_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _46870_ (_39440_, _39439_, _31351_);
  and _46871_ (_39441_, _39440_, _39438_);
  and _46872_ (_39442_, _39111_, _38619_);
  and _46873_ (_39443_, _39442_, _39237_);
  nand _46874_ (_39444_, _39443_, _38704_);
  or _46875_ (_39445_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _46876_ (_39446_, _39445_, _30651_);
  and _46877_ (_39447_, _39446_, _39444_);
  and _46878_ (_39448_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _46879_ (_39449_, _39448_, rst);
  or _46880_ (_39450_, _39449_, _39447_);
  or _46881_ (_31153_, _39450_, _39441_);
  and _46882_ (_39451_, _39095_, _27211_);
  and _46883_ (_39452_, _39451_, _39271_);
  and _46884_ (_39453_, _39452_, _31308_);
  nand _46885_ (_39454_, _39453_, _31265_);
  or _46886_ (_39455_, _39453_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _46887_ (_39456_, _39455_, _31351_);
  and _46888_ (_39457_, _39456_, _39454_);
  and _46889_ (_39458_, _39238_, _38619_);
  and _46890_ (_39459_, _39458_, _39237_);
  not _46891_ (_39460_, _39459_);
  nor _46892_ (_39461_, _39460_, _38704_);
  and _46893_ (_39462_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _46894_ (_39463_, _39462_, _39461_);
  and _46895_ (_39464_, _39463_, _30651_);
  and _46896_ (_39465_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _46897_ (_39466_, _39465_, rst);
  or _46898_ (_39467_, _39466_, _39464_);
  or _46899_ (_31176_, _39467_, _39457_);
  and _46900_ (_39468_, _39451_, _27847_);
  and _46901_ (_39469_, _39468_, _31308_);
  nand _46902_ (_39470_, _39469_, _31265_);
  or _46903_ (_39471_, _39469_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _46904_ (_39472_, _39471_, _31351_);
  and _46905_ (_39473_, _39472_, _39470_);
  nor _46906_ (_39474_, _27825_, _27343_);
  and _46907_ (_39475_, _38619_, _39474_);
  and _46908_ (_39476_, _39475_, _39237_);
  not _46909_ (_39477_, _39476_);
  nor _46910_ (_39478_, _39477_, _38704_);
  and _46911_ (_39479_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _46912_ (_39480_, _39479_, _39478_);
  and _46913_ (_39481_, _39480_, _30651_);
  and _46914_ (_39482_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _46915_ (_39483_, _39482_, rst);
  or _46916_ (_39484_, _39483_, _39481_);
  or _46917_ (_31199_, _39484_, _39473_);
  or _46918_ (_39485_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _46919_ (_39486_, _39485_, _31351_);
  and _46920_ (_39487_, _39421_, _27003_);
  nand _46921_ (_39488_, _39487_, _31265_);
  and _46922_ (_39489_, _39488_, _39486_);
  nand _46923_ (_39490_, _39427_, _38682_);
  and _46924_ (_39491_, _39490_, _30651_);
  and _46925_ (_39492_, _39491_, _39485_);
  not _46926_ (_39493_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _46927_ (_39494_, _30640_, _39493_);
  or _46928_ (_39495_, _39494_, rst);
  or _46929_ (_39496_, _39495_, _39492_);
  or _46930_ (_40808_, _39496_, _39489_);
  and _46931_ (_39497_, _32604_, _27650_);
  and _46932_ (_39498_, _39497_, _38620_);
  nand _46933_ (_39499_, _39498_, _31265_);
  or _46934_ (_39500_, _39498_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46935_ (_39501_, _39500_, _31351_);
  and _46936_ (_39502_, _39501_, _39499_);
  nand _46937_ (_39503_, _39427_, _38672_);
  or _46938_ (_39504_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46939_ (_39505_, _39504_, _30651_);
  and _46940_ (_39506_, _39505_, _39503_);
  and _46941_ (_39507_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _46942_ (_39508_, _39507_, rst);
  or _46943_ (_39509_, _39508_, _39506_);
  or _46944_ (_40810_, _39509_, _39502_);
  not _46945_ (_39510_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  not _46946_ (_39511_, _34073_);
  and _46947_ (_39512_, _39421_, _39511_);
  nor _46948_ (_39513_, _39512_, _39510_);
  and _46949_ (_39514_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _46950_ (_39515_, _39514_, _33366_);
  and _46951_ (_39516_, _39515_, _39421_);
  or _46952_ (_39517_, _39516_, _39513_);
  and _46953_ (_39518_, _39517_, _31351_);
  nand _46954_ (_39519_, _39427_, _38665_);
  or _46955_ (_39520_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _46956_ (_39521_, _39520_, _30651_);
  and _46957_ (_39522_, _39521_, _39519_);
  nor _46958_ (_39523_, _30640_, _39510_);
  or _46959_ (_39524_, _39523_, rst);
  or _46960_ (_39525_, _39524_, _39522_);
  or _46961_ (_40812_, _39525_, _39518_);
  and _46962_ (_39526_, _39421_, _34052_);
  nand _46963_ (_39527_, _39526_, _31265_);
  or _46964_ (_39528_, _39526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _46965_ (_39529_, _39528_, _31351_);
  and _46966_ (_39530_, _39529_, _39527_);
  nand _46967_ (_39531_, _39427_, _38658_);
  or _46968_ (_39532_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _46969_ (_39533_, _39532_, _30651_);
  and _46970_ (_39534_, _39533_, _39531_);
  and _46971_ (_39535_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _46972_ (_39536_, _39535_, rst);
  or _46973_ (_39537_, _39536_, _39534_);
  or _46974_ (_40814_, _39537_, _39530_);
  not _46975_ (_39538_, _39421_);
  or _46976_ (_39539_, _39538_, _34813_);
  and _46977_ (_39540_, _39539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46978_ (_39541_, _34802_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _46979_ (_39542_, _39541_, _34845_);
  and _46980_ (_39543_, _39542_, _39421_);
  or _46981_ (_39544_, _39543_, _39540_);
  and _46982_ (_39545_, _39544_, _31351_);
  nand _46983_ (_39546_, _39427_, _38650_);
  or _46984_ (_39547_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46985_ (_39548_, _39547_, _30651_);
  and _46986_ (_39549_, _39548_, _39546_);
  and _46987_ (_39550_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _46988_ (_39551_, _39550_, rst);
  or _46989_ (_39552_, _39551_, _39549_);
  or _46990_ (_40816_, _39552_, _39545_);
  and _46991_ (_39553_, _39421_, _35607_);
  nand _46992_ (_39554_, _39553_, _31265_);
  or _46993_ (_39555_, _39553_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _46994_ (_39556_, _39555_, _31351_);
  and _46995_ (_39557_, _39556_, _39554_);
  nand _46996_ (_39566_, _39427_, _38642_);
  or _46997_ (_39577_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _46998_ (_39588_, _39577_, _30651_);
  and _46999_ (_39597_, _39588_, _39566_);
  and _47000_ (_39603_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _47001_ (_39614_, _39603_, rst);
  or _47002_ (_39625_, _39614_, _39597_);
  or _47003_ (_40818_, _39625_, _39557_);
  and _47004_ (_39646_, _39421_, _36336_);
  nand _47005_ (_39657_, _39646_, _31265_);
  or _47006_ (_39668_, _39646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _47007_ (_39679_, _39668_, _31351_);
  and _47008_ (_39690_, _39679_, _39657_);
  nand _47009_ (_39701_, _39427_, _38635_);
  or _47010_ (_39712_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _47011_ (_39723_, _39712_, _30651_);
  and _47012_ (_39734_, _39723_, _39701_);
  and _47013_ (_39745_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _47014_ (_39756_, _39745_, rst);
  or _47015_ (_39767_, _39756_, _39734_);
  or _47016_ (_40820_, _39767_, _39690_);
  and _47017_ (_39771_, _39436_, _27003_);
  nand _47018_ (_39772_, _39771_, _31265_);
  or _47019_ (_39773_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _47020_ (_39774_, _39773_, _31351_);
  and _47021_ (_39775_, _39774_, _39772_);
  nand _47022_ (_39776_, _39443_, _38682_);
  and _47023_ (_39777_, _39776_, _30651_);
  and _47024_ (_39778_, _39777_, _39773_);
  not _47025_ (_39779_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _47026_ (_39780_, _30640_, _39779_);
  or _47027_ (_39781_, _39780_, rst);
  or _47028_ (_39782_, _39781_, _39778_);
  or _47029_ (_40821_, _39782_, _39775_);
  and _47030_ (_39783_, _39436_, _32604_);
  nand _47031_ (_39784_, _39783_, _31265_);
  or _47032_ (_39785_, _39783_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _47033_ (_39786_, _39785_, _31351_);
  and _47034_ (_39787_, _39786_, _39784_);
  nand _47035_ (_39788_, _39443_, _38672_);
  or _47036_ (_39789_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _47037_ (_39790_, _39789_, _30651_);
  and _47038_ (_39791_, _39790_, _39788_);
  and _47039_ (_39792_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _47040_ (_39793_, _39792_, rst);
  or _47041_ (_39794_, _39793_, _39791_);
  or _47042_ (_40823_, _39794_, _39787_);
  and _47043_ (_39795_, _39436_, _33344_);
  nand _47044_ (_39796_, _39795_, _31265_);
  or _47045_ (_39797_, _39795_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _47046_ (_39798_, _39797_, _31351_);
  and _47047_ (_39799_, _39798_, _39796_);
  nand _47048_ (_39800_, _39443_, _38665_);
  or _47049_ (_39801_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _47050_ (_39802_, _39801_, _30651_);
  and _47051_ (_39803_, _39802_, _39800_);
  and _47052_ (_39804_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _47053_ (_39805_, _39804_, rst);
  or _47054_ (_39806_, _39805_, _39803_);
  or _47055_ (_40825_, _39806_, _39799_);
  and _47056_ (_39807_, _39436_, _34052_);
  nand _47057_ (_39808_, _39807_, _31265_);
  or _47058_ (_39809_, _39807_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _47059_ (_39810_, _39809_, _31351_);
  and _47060_ (_39811_, _39810_, _39808_);
  nand _47061_ (_39812_, _39443_, _38658_);
  or _47062_ (_39813_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _47063_ (_39814_, _39813_, _30651_);
  and _47064_ (_39815_, _39814_, _39812_);
  and _47065_ (_39816_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _47066_ (_39817_, _39816_, rst);
  or _47067_ (_39818_, _39817_, _39815_);
  or _47068_ (_40827_, _39818_, _39811_);
  and _47069_ (_39819_, _39436_, _34791_);
  nand _47070_ (_39820_, _39819_, _31265_);
  or _47071_ (_39821_, _39819_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47072_ (_39822_, _39821_, _31351_);
  and _47073_ (_39823_, _39822_, _39820_);
  nand _47074_ (_39824_, _39443_, _38650_);
  or _47075_ (_39825_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47076_ (_39826_, _39825_, _30651_);
  and _47077_ (_39827_, _39826_, _39824_);
  and _47078_ (_39828_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _47079_ (_39829_, _39828_, rst);
  or _47080_ (_39830_, _39829_, _39827_);
  or _47081_ (_40829_, _39830_, _39823_);
  and _47082_ (_39831_, _39436_, _35607_);
  nand _47083_ (_39832_, _39831_, _31265_);
  or _47084_ (_39833_, _39831_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _47085_ (_39834_, _39833_, _31351_);
  and _47086_ (_39835_, _39834_, _39832_);
  nand _47087_ (_39836_, _39443_, _38642_);
  or _47088_ (_39837_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _47089_ (_39838_, _39837_, _30651_);
  and _47090_ (_39839_, _39838_, _39836_);
  and _47091_ (_39840_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _47092_ (_39841_, _39840_, rst);
  or _47093_ (_39842_, _39841_, _39839_);
  or _47094_ (_40831_, _39842_, _39835_);
  and _47095_ (_39843_, _39436_, _36336_);
  nand _47096_ (_39844_, _39843_, _31265_);
  or _47097_ (_39845_, _39843_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _47098_ (_39846_, _39845_, _31351_);
  and _47099_ (_39847_, _39846_, _39844_);
  nand _47100_ (_39848_, _39443_, _38635_);
  or _47101_ (_39849_, _39443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _47102_ (_39850_, _39849_, _30651_);
  and _47103_ (_39851_, _39850_, _39848_);
  and _47104_ (_39852_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _47105_ (_39853_, _39852_, rst);
  or _47106_ (_39854_, _39853_, _39851_);
  or _47107_ (_40833_, _39854_, _39847_);
  nand _47108_ (_39855_, _39459_, _31265_);
  or _47109_ (_39856_, _39459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _47110_ (_39857_, _39856_, _31351_);
  and _47111_ (_39858_, _39857_, _39855_);
  and _47112_ (_39859_, _39459_, _38683_);
  not _47113_ (_39860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _47114_ (_39861_, _39459_, _39860_);
  or _47115_ (_39862_, _39861_, _39859_);
  and _47116_ (_39863_, _39862_, _30651_);
  nor _47117_ (_39864_, _30640_, _39860_);
  or _47118_ (_39865_, _39864_, rst);
  or _47119_ (_39866_, _39865_, _39863_);
  or _47120_ (_40835_, _39866_, _39858_);
  and _47121_ (_39867_, _39452_, _32604_);
  nand _47122_ (_39868_, _39867_, _31265_);
  or _47123_ (_39869_, _39867_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _47124_ (_39870_, _39869_, _31351_);
  and _47125_ (_39871_, _39870_, _39868_);
  nor _47126_ (_39872_, _39460_, _38672_);
  and _47127_ (_39873_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _47128_ (_39874_, _39873_, _39872_);
  and _47129_ (_39875_, _39874_, _30651_);
  and _47130_ (_39876_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _47131_ (_39877_, _39876_, rst);
  or _47132_ (_39878_, _39877_, _39875_);
  or _47133_ (_40837_, _39878_, _39871_);
  and _47134_ (_39879_, _39452_, _33344_);
  nand _47135_ (_39880_, _39879_, _31265_);
  or _47136_ (_39881_, _39879_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _47137_ (_39882_, _39881_, _31351_);
  and _47138_ (_39883_, _39882_, _39880_);
  nor _47139_ (_39884_, _39460_, _38665_);
  and _47140_ (_39885_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _47141_ (_39886_, _39885_, _39884_);
  and _47142_ (_39887_, _39886_, _30651_);
  and _47143_ (_39888_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _47144_ (_39889_, _39888_, rst);
  or _47145_ (_39890_, _39889_, _39887_);
  or _47146_ (_40839_, _39890_, _39883_);
  and _47147_ (_39891_, _39452_, _34052_);
  nand _47148_ (_39892_, _39891_, _31265_);
  or _47149_ (_39893_, _39891_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _47150_ (_39894_, _39893_, _31351_);
  and _47151_ (_39895_, _39894_, _39892_);
  nor _47152_ (_39896_, _39460_, _38658_);
  and _47153_ (_39897_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _47154_ (_39898_, _39897_, _39896_);
  and _47155_ (_39899_, _39898_, _30651_);
  and _47156_ (_39900_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _47157_ (_39901_, _39900_, rst);
  or _47158_ (_39902_, _39901_, _39899_);
  or _47159_ (_40841_, _39902_, _39895_);
  and _47160_ (_39903_, _39452_, _34791_);
  nand _47161_ (_39904_, _39903_, _31265_);
  or _47162_ (_39905_, _39903_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _47163_ (_39906_, _39905_, _31351_);
  and _47164_ (_39907_, _39906_, _39904_);
  nor _47165_ (_39908_, _39460_, _38650_);
  and _47166_ (_39909_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _47167_ (_39910_, _39909_, _39908_);
  and _47168_ (_39911_, _39910_, _30651_);
  and _47169_ (_39912_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _47170_ (_39913_, _39912_, rst);
  or _47171_ (_39914_, _39913_, _39911_);
  or _47172_ (_40843_, _39914_, _39907_);
  and _47173_ (_39915_, _39452_, _35607_);
  nand _47174_ (_39916_, _39915_, _31265_);
  or _47175_ (_39917_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _47176_ (_39918_, _39917_, _31351_);
  and _47177_ (_39919_, _39918_, _39916_);
  nor _47178_ (_39920_, _39460_, _38642_);
  and _47179_ (_39921_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _47180_ (_39922_, _39921_, _39920_);
  and _47181_ (_39923_, _39922_, _30651_);
  and _47182_ (_39924_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _47183_ (_39925_, _39924_, rst);
  or _47184_ (_39926_, _39925_, _39923_);
  or _47185_ (_40845_, _39926_, _39919_);
  and _47186_ (_39927_, _39452_, _36336_);
  nand _47187_ (_39928_, _39927_, _31265_);
  or _47188_ (_39929_, _39927_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _47189_ (_39930_, _39929_, _31351_);
  and _47190_ (_39931_, _39930_, _39928_);
  nor _47191_ (_39932_, _39460_, _38635_);
  and _47192_ (_39933_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _47193_ (_39934_, _39933_, _39932_);
  and _47194_ (_39935_, _39934_, _30651_);
  and _47195_ (_39936_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _47196_ (_39937_, _39936_, rst);
  or _47197_ (_39938_, _39937_, _39935_);
  or _47198_ (_40847_, _39938_, _39931_);
  and _47199_ (_39939_, _39468_, _27003_);
  nand _47200_ (_39940_, _39939_, _31265_);
  or _47201_ (_39941_, _39476_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _47202_ (_39942_, _39941_, _31351_);
  and _47203_ (_39943_, _39942_, _39940_);
  nand _47204_ (_39944_, _39476_, _38682_);
  and _47205_ (_39945_, _39941_, _30651_);
  and _47206_ (_39946_, _39945_, _39944_);
  not _47207_ (_39947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _47208_ (_39948_, _30640_, _39947_);
  or _47209_ (_39949_, _39948_, rst);
  or _47210_ (_39950_, _39949_, _39946_);
  or _47211_ (_40849_, _39950_, _39943_);
  and _47212_ (_39951_, _39468_, _32604_);
  nand _47213_ (_39952_, _39951_, _31265_);
  or _47214_ (_39953_, _39951_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _47215_ (_39954_, _39953_, _31351_);
  and _47216_ (_39955_, _39954_, _39952_);
  nor _47217_ (_39956_, _39477_, _38672_);
  and _47218_ (_39957_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _47219_ (_39958_, _39957_, _39956_);
  and _47220_ (_39959_, _39958_, _30651_);
  and _47221_ (_39960_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _47222_ (_39961_, _39960_, rst);
  or _47223_ (_39962_, _39961_, _39959_);
  or _47224_ (_40851_, _39962_, _39955_);
  and _47225_ (_39963_, _39468_, _33344_);
  nand _47226_ (_39964_, _39963_, _31265_);
  or _47227_ (_39965_, _39963_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _47228_ (_39966_, _39965_, _31351_);
  and _47229_ (_39967_, _39966_, _39964_);
  nor _47230_ (_39968_, _39477_, _38665_);
  and _47231_ (_39969_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _47232_ (_39970_, _39969_, _39968_);
  and _47233_ (_39971_, _39970_, _30651_);
  and _47234_ (_39972_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _47235_ (_39973_, _39972_, rst);
  or _47236_ (_39974_, _39973_, _39971_);
  or _47237_ (_40852_, _39974_, _39967_);
  and _47238_ (_39975_, _39468_, _34052_);
  nand _47239_ (_39976_, _39975_, _31265_);
  or _47240_ (_39977_, _39975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _47241_ (_39978_, _39977_, _31351_);
  and _47242_ (_39979_, _39978_, _39976_);
  nor _47243_ (_39984_, _39477_, _38658_);
  and _47244_ (_39986_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _47245_ (_39987_, _39986_, _39984_);
  and _47246_ (_39988_, _39987_, _30651_);
  and _47247_ (_39989_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _47248_ (_39990_, _39989_, rst);
  or _47249_ (_39991_, _39990_, _39988_);
  or _47250_ (_40854_, _39991_, _39979_);
  and _47251_ (_39992_, _39468_, _34791_);
  nand _47252_ (_39993_, _39992_, _31265_);
  or _47253_ (_39994_, _39992_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47254_ (_39995_, _39994_, _31351_);
  and _47255_ (_39996_, _39995_, _39993_);
  nor _47256_ (_39997_, _39477_, _38650_);
  and _47257_ (_39998_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _47258_ (_39999_, _39998_, _39997_);
  and _47259_ (_40000_, _39999_, _30651_);
  and _47260_ (_40001_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _47261_ (_40002_, _40001_, rst);
  or _47262_ (_40003_, _40002_, _40000_);
  or _47263_ (_40856_, _40003_, _39996_);
  and _47264_ (_40004_, _39468_, _35607_);
  nand _47265_ (_40005_, _40004_, _31265_);
  or _47266_ (_40006_, _40004_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _47267_ (_40007_, _40006_, _31351_);
  and _47268_ (_40008_, _40007_, _40005_);
  nor _47269_ (_40009_, _39477_, _38642_);
  and _47270_ (_40010_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _47271_ (_40011_, _40010_, _40009_);
  and _47272_ (_40012_, _40011_, _30651_);
  and _47273_ (_40020_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _47274_ (_40031_, _40020_, rst);
  or _47275_ (_40042_, _40031_, _40012_);
  or _47276_ (_40858_, _40042_, _40008_);
  and _47277_ (_40044_, _39468_, _36336_);
  nand _47278_ (_40045_, _40044_, _31265_);
  or _47279_ (_40046_, _40044_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _47280_ (_40047_, _40046_, _31351_);
  and _47281_ (_40048_, _40047_, _40045_);
  nor _47282_ (_40049_, _39477_, _38635_);
  and _47283_ (_40050_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _47284_ (_40051_, _40050_, _40049_);
  and _47285_ (_40052_, _40051_, _30651_);
  and _47286_ (_40053_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _47287_ (_40054_, _40053_, rst);
  or _47288_ (_40055_, _40054_, _40052_);
  or _47289_ (_40860_, _40055_, _40048_);
  and _47290_ (_41311_, t0_i, _43100_);
  and _47291_ (_41314_, t1_i, _43100_);
  nor _47292_ (_40056_, _26740_, _27650_);
  and _47293_ (_40057_, _40056_, _38621_);
  and _47294_ (_40058_, _40057_, _30651_);
  not _47295_ (_40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _47296_ (_40060_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _47297_ (_40061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _47298_ (_40062_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _40061_);
  nor _47299_ (_40063_, _40062_, _40060_);
  or _47300_ (_40064_, _40063_, _40058_);
  and _47301_ (_40065_, _40064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _47302_ (_40066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _47303_ (_40067_, t1_i);
  and _47304_ (_40068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _40067_);
  nor _47305_ (_40069_, _40068_, _40066_);
  not _47306_ (_40071_, _40069_);
  not _47307_ (_40077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _47308_ (_40078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _40077_);
  nor _47309_ (_40079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _47310_ (_40080_, _40079_);
  and _47311_ (_40081_, _40080_, _40078_);
  and _47312_ (_40082_, _40081_, _40071_);
  not _47313_ (_40083_, _40082_);
  nand _47314_ (_40084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _47315_ (_40085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or _47316_ (_40086_, _40085_, _40084_);
  nor _47317_ (_40087_, _40086_, _40083_);
  and _47318_ (_40088_, _40087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _47319_ (_40089_, _40088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _47320_ (_40090_, _40089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _47321_ (_40091_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _47322_ (_40092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _47323_ (_40093_, _40086_, _40092_);
  and _47324_ (_40094_, _40093_, _40082_);
  and _47325_ (_40095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _47326_ (_40096_, _40095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _47327_ (_40097_, _40096_, _40094_);
  nor _47328_ (_40098_, _40097_, _40063_);
  and _47329_ (_40099_, _40098_, _40091_);
  and _47330_ (_40100_, _40097_, _40060_);
  and _47331_ (_40101_, _40100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47332_ (_40102_, _40101_, _40099_);
  nor _47333_ (_40103_, _40102_, _40058_);
  or _47334_ (_40104_, _40103_, _40065_);
  and _47335_ (_40105_, _34052_, _27661_);
  and _47336_ (_40106_, _40105_, _38620_);
  and _47337_ (_40107_, _40106_, _30651_);
  not _47338_ (_40108_, _40107_);
  and _47339_ (_40109_, _40108_, _40104_);
  nor _47340_ (_40110_, _40108_, _38704_);
  or _47341_ (_40111_, _40110_, _40109_);
  and _47342_ (_41317_, _40111_, _43100_);
  not _47343_ (_40112_, _30651_);
  nor _47344_ (_40113_, _40112_, _27650_);
  and _47345_ (_40114_, _40113_, _38751_);
  and _47346_ (_40115_, _40114_, _43100_);
  and _47347_ (_40116_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _47348_ (_40117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47349_ (_40118_, _40117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47350_ (_40119_, _40096_, _40093_);
  and _47351_ (_40120_, _40119_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47352_ (_40121_, _40120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _47353_ (_40122_, _40121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47354_ (_40123_, _40122_, _40082_);
  and _47355_ (_40124_, _40123_, _40118_);
  and _47356_ (_40125_, _40124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47357_ (_40126_, _40125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47358_ (_40127_, _40125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47359_ (_40128_, _40127_, _40126_);
  and _47360_ (_40129_, _40128_, _40062_);
  and _47361_ (_40130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _47362_ (_40131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47363_ (_40132_, _40131_, _40093_);
  and _47364_ (_40133_, _40132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47365_ (_40134_, _40133_, _40082_);
  and _47366_ (_40135_, _40134_, _40118_);
  and _47367_ (_40136_, _40135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47368_ (_40137_, _40136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47369_ (_40138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _47370_ (_40139_, _40136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _47371_ (_40140_, _40139_, _40138_);
  nor _47372_ (_40141_, _40140_, _40137_);
  or _47373_ (_40142_, _40141_, _40130_);
  nor _47374_ (_40143_, _40142_, _40129_);
  nor _47375_ (_40144_, _40143_, _40058_);
  not _47376_ (_40145_, _38704_);
  and _47377_ (_40146_, _40058_, _40145_);
  or _47378_ (_40147_, _40146_, _40144_);
  nor _47379_ (_40148_, _40114_, rst);
  and _47380_ (_40149_, _40148_, _40147_);
  or _47381_ (_41320_, _40149_, _40116_);
  and _47382_ (_40150_, _40083_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or _47383_ (_40151_, _40150_, _40126_);
  and _47384_ (_40152_, _40151_, _40062_);
  or _47385_ (_40153_, _40150_, _40137_);
  and _47386_ (_40154_, _40153_, _40138_);
  nand _47387_ (_40155_, _40082_, _40059_);
  and _47388_ (_40160_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _47389_ (_40167_, _40160_, _40155_);
  or _47390_ (_40168_, _40167_, _40100_);
  or _47391_ (_40169_, _40168_, _40154_);
  nor _47392_ (_40170_, _40169_, _40152_);
  nor _47393_ (_40171_, _40170_, _40058_);
  and _47394_ (_41323_, _40171_, _40148_);
  and _47395_ (_40172_, _40113_, _34791_);
  and _47396_ (_40173_, _40172_, _38620_);
  nor _47397_ (_40174_, _40173_, rst);
  and _47398_ (_40175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47399_ (_40176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _47400_ (_40177_, _40176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47401_ (_40178_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47402_ (_40179_, _40178_, _40175_);
  and _47403_ (_40180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _47404_ (_40181_, _40180_, _40179_);
  or _47405_ (_40182_, _40181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _47406_ (_40183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _47407_ (_40184_, _40183_);
  and _47408_ (_40185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _47409_ (_40186_, _40185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _47410_ (_40187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _47411_ (_40188_, t0_i);
  and _47412_ (_40189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _40188_);
  nor _47413_ (_40190_, _40189_, _40187_);
  not _47414_ (_40191_, _40190_);
  not _47415_ (_40192_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _47416_ (_40193_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _47417_ (_40194_, _40193_, _40192_);
  and _47418_ (_40195_, _40194_, _40191_);
  and _47419_ (_40196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _47420_ (_40197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47421_ (_40198_, _40197_, _40196_);
  and _47422_ (_40199_, _40198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _47423_ (_40200_, _40199_, _40195_);
  and _47424_ (_40201_, _40200_, _40186_);
  and _47425_ (_40202_, _40201_, _40184_);
  and _47426_ (_40203_, _40202_, _40182_);
  not _47427_ (_40204_, _40195_);
  and _47428_ (_40205_, _40204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and _47429_ (_40206_, _40200_, _40179_);
  and _47430_ (_40207_, _40206_, _40180_);
  and _47431_ (_40208_, _40207_, _40183_);
  or _47432_ (_40209_, _40208_, _40205_);
  nor _47433_ (_40210_, _40209_, _40203_);
  and _47434_ (_40211_, _40113_, _33344_);
  and _47435_ (_40212_, _40211_, _38620_);
  nor _47436_ (_40213_, _40212_, _40210_);
  and _47437_ (_41326_, _40213_, _40174_);
  and _47438_ (_40214_, _40113_, _38848_);
  nand _47439_ (_40215_, _40214_, _38704_);
  and _47440_ (_40216_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _47441_ (_40217_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47442_ (_40218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40217_);
  not _47443_ (_40219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47444_ (_40220_, _40219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _47445_ (_40221_, _40220_, _40218_);
  not _47446_ (_40222_, _40201_);
  and _47447_ (_40223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47448_ (_40224_, _40223_, _40222_);
  or _47449_ (_40225_, _40224_, _40221_);
  nand _47450_ (_40226_, _40220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _47451_ (_40227_, _40226_, _40201_);
  and _47452_ (_40228_, _40227_, _40225_);
  or _47453_ (_40229_, _40228_, _40216_);
  or _47454_ (_40230_, _40229_, _40173_);
  and _47455_ (_40231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _47456_ (_40232_, _40231_, _40200_);
  nor _47457_ (_40233_, _40232_, _40173_);
  or _47458_ (_40234_, _40233_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _47459_ (_40235_, _40234_, _40230_);
  or _47460_ (_40236_, _40235_, _40214_);
  and _47461_ (_40238_, _40236_, _43100_);
  and _47462_ (_41329_, _40238_, _40215_);
  nand _47463_ (_40242_, _40173_, _38704_);
  not _47464_ (_40243_, _40212_);
  not _47465_ (_40244_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _47466_ (_40245_, _40199_, _40186_);
  and _47467_ (_40246_, _40195_, _40217_);
  and _47468_ (_40247_, _40246_, _40245_);
  and _47469_ (_40248_, _40247_, _40179_);
  and _47470_ (_40249_, _40248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _47471_ (_40250_, _40249_, _40244_);
  and _47472_ (_40251_, _40249_, _40244_);
  or _47473_ (_40252_, _40251_, _40250_);
  and _47474_ (_40253_, _40252_, _40221_);
  and _47475_ (_40254_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _47476_ (_40255_, _40254_, _40178_);
  and _47477_ (_40256_, _40255_, _40175_);
  and _47478_ (_40257_, _40256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _47479_ (_40267_, _40257_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _47480_ (_40268_, _40254_, _40181_);
  and _47481_ (_40269_, _40268_, _40267_);
  and _47482_ (_40270_, _40269_, _40223_);
  and _47483_ (_40271_, _40206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _47484_ (_40272_, _40271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _47485_ (_40273_, _40207_, _40184_);
  and _47486_ (_40274_, _40273_, _40272_);
  or _47487_ (_40275_, _40274_, _40270_);
  or _47488_ (_40276_, _40275_, _40253_);
  or _47489_ (_40277_, _40276_, _40173_);
  and _47490_ (_40278_, _40277_, _40243_);
  and _47491_ (_40279_, _40278_, _40242_);
  and _47492_ (_40280_, _40212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _47493_ (_40281_, _40280_, _40279_);
  and _47494_ (_41332_, _40281_, _43100_);
  or _47495_ (_40282_, _40254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _47496_ (_40283_, _40223_, _43100_);
  nand _47497_ (_40284_, _40283_, _40282_);
  nor _47498_ (_40285_, _40284_, _40173_);
  not _47499_ (_40286_, _40254_);
  nor _47500_ (_40287_, _40286_, _40181_);
  nor _47501_ (_40288_, _40287_, _40212_);
  and _47502_ (_41335_, _40288_, _40285_);
  and _47503_ (_40289_, _40113_, _38622_);
  or _47504_ (_40290_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _47505_ (_40291_, _40290_, _43100_);
  nand _47506_ (_40292_, _40289_, _38704_);
  and _47507_ (_41338_, _40292_, _40291_);
  and _47508_ (_40293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _47509_ (_40294_, _40293_, _40058_);
  and _47510_ (_40295_, _40294_, _40082_);
  or _47511_ (_40296_, _40295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  not _47512_ (_40297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _47513_ (_40298_, _40060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _47514_ (_40299_, _40298_, _40119_);
  nor _47515_ (_40300_, _40299_, _40058_);
  nor _47516_ (_40301_, _40300_, _40297_);
  nand _47517_ (_40302_, _40301_, _40295_);
  and _47518_ (_40303_, _40302_, _40148_);
  and _47519_ (_40304_, _40303_, _40296_);
  and _47520_ (_40305_, _40115_, _38683_);
  or _47521_ (_41820_, _40305_, _40304_);
  not _47522_ (_40306_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _47523_ (_40307_, _40294_, _40306_);
  not _47524_ (_40308_, _40293_);
  and _47525_ (_40309_, _40082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _47526_ (_40310_, _40309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _47527_ (_40311_, _40309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _47528_ (_40312_, _40311_, _40310_);
  and _47529_ (_40313_, _40312_, _40308_);
  and _47530_ (_40314_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _47531_ (_40315_, _40314_, _40060_);
  and _47532_ (_40316_, _40315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _47533_ (_40317_, _40316_, _40313_);
  nor _47534_ (_40318_, _40317_, _40058_);
  or _47535_ (_40319_, _40318_, _40307_);
  and _47536_ (_40320_, _40319_, _40108_);
  nor _47537_ (_40321_, _40108_, _38672_);
  or _47538_ (_40322_, _40321_, _40320_);
  and _47539_ (_41822_, _40322_, _43100_);
  not _47540_ (_40323_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _47541_ (_40324_, _40294_, _40323_);
  nor _47542_ (_40325_, _40310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _47543_ (_40326_, _40310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _47544_ (_40327_, _40326_, _40325_);
  and _47545_ (_40328_, _40327_, _40308_);
  and _47546_ (_40329_, _40100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _47547_ (_40330_, _40329_, _40328_);
  nor _47548_ (_40331_, _40330_, _40058_);
  or _47549_ (_40332_, _40331_, _40324_);
  and _47550_ (_40333_, _40332_, _40148_);
  not _47551_ (_40334_, _38665_);
  and _47552_ (_40335_, _40115_, _40334_);
  or _47553_ (_41823_, _40335_, _40333_);
  not _47554_ (_40336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _47555_ (_40337_, _40294_, _40336_);
  or _47556_ (_40338_, _40326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _47557_ (_40339_, _40293_, _40087_);
  and _47558_ (_40340_, _40339_, _40338_);
  and _47559_ (_40341_, _40100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _47560_ (_40342_, _40341_, _40340_);
  nor _47561_ (_40343_, _40342_, _40058_);
  or _47562_ (_40344_, _40343_, _40337_);
  and _47563_ (_40345_, _40344_, _40148_);
  not _47564_ (_40346_, _38658_);
  and _47565_ (_40347_, _40115_, _40346_);
  or _47566_ (_41825_, _40347_, _40345_);
  nor _47567_ (_40348_, _40294_, _40092_);
  or _47568_ (_40349_, _40087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _47569_ (_40350_, _40293_, _40094_);
  and _47570_ (_40351_, _40350_, _40349_);
  and _47571_ (_40352_, _40100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _47572_ (_40353_, _40352_, _40351_);
  nor _47573_ (_40354_, _40353_, _40058_);
  or _47574_ (_40355_, _40354_, _40348_);
  and _47575_ (_40356_, _40355_, _40148_);
  not _47576_ (_40357_, _38650_);
  and _47577_ (_40358_, _40115_, _40357_);
  or _47578_ (_41827_, _40358_, _40356_);
  and _47579_ (_40359_, _40064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _47580_ (_40360_, _40315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _47581_ (_40361_, _40063_);
  and _47582_ (_40362_, _40094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _47583_ (_40363_, _40094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _47584_ (_40364_, _40363_, _40362_);
  and _47585_ (_40365_, _40364_, _40361_);
  nor _47586_ (_40366_, _40365_, _40360_);
  nor _47587_ (_40367_, _40366_, _40058_);
  or _47588_ (_40368_, _40367_, _40359_);
  and _47589_ (_40369_, _40368_, _40148_);
  not _47590_ (_40370_, _38642_);
  and _47591_ (_40371_, _40115_, _40370_);
  or _47592_ (_41829_, _40371_, _40369_);
  and _47593_ (_40372_, _40064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _47594_ (_40373_, _40060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47595_ (_40374_, _40373_, _40082_);
  and _47596_ (_40375_, _40374_, _40119_);
  or _47597_ (_40376_, _40362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _47598_ (_40377_, _40376_, _40361_);
  nor _47599_ (_40378_, _40377_, _40090_);
  nor _47600_ (_40379_, _40378_, _40375_);
  nor _47601_ (_40380_, _40379_, _40058_);
  or _47602_ (_40381_, _40380_, _40372_);
  and _47603_ (_40382_, _40381_, _40148_);
  not _47604_ (_40383_, _38635_);
  and _47605_ (_40384_, _40115_, _40383_);
  or _47606_ (_41831_, _40384_, _40382_);
  not _47607_ (_40385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47608_ (_40386_, _40094_, _40061_);
  nor _47609_ (_40387_, _40096_, _40059_);
  not _47610_ (_40388_, _40387_);
  and _47611_ (_40389_, _40388_, _40386_);
  nor _47612_ (_40390_, _40389_, _40385_);
  and _47613_ (_40391_, _40389_, _40385_);
  or _47614_ (_40392_, _40391_, _40390_);
  or _47615_ (_40393_, _40392_, _40058_);
  nand _47616_ (_40394_, _40058_, _38682_);
  and _47617_ (_40395_, _40394_, _40148_);
  and _47618_ (_40396_, _40395_, _40393_);
  and _47619_ (_40397_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or _47620_ (_41833_, _40397_, _40396_);
  nand _47621_ (_40398_, _40058_, _38672_);
  not _47622_ (_40399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not _47623_ (_40400_, _40062_);
  nor _47624_ (_40401_, _40097_, _40400_);
  not _47625_ (_40402_, _40401_);
  nor _47626_ (_40403_, _40386_, _40062_);
  nor _47627_ (_40404_, _40403_, _40385_);
  and _47628_ (_40405_, _40404_, _40402_);
  nor _47629_ (_40406_, _40405_, _40399_);
  and _47630_ (_40407_, _40405_, _40399_);
  or _47631_ (_40408_, _40407_, _40406_);
  or _47632_ (_40409_, _40408_, _40058_);
  and _47633_ (_40410_, _40409_, _40148_);
  and _47634_ (_40411_, _40410_, _40398_);
  and _47635_ (_40412_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _47636_ (_41835_, _40412_, _40411_);
  and _47637_ (_40413_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _47638_ (_40414_, _40058_, _38665_);
  and _47639_ (_40415_, _40131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47640_ (_40416_, _40415_, _40094_);
  nand _47641_ (_40417_, _40416_, _40061_);
  or _47642_ (_40418_, _40417_, _40387_);
  and _47643_ (_40419_, _40418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _47644_ (_40420_, _40387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _47645_ (_40421_, _40420_);
  not _47646_ (_40422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47647_ (_40423_, _40131_, _40422_);
  and _47648_ (_40424_, _40423_, _40094_);
  and _47649_ (_40425_, _40424_, _40421_);
  or _47650_ (_40426_, _40425_, _40419_);
  or _47651_ (_40427_, _40426_, _40058_);
  and _47652_ (_40428_, _40427_, _40148_);
  and _47653_ (_40429_, _40428_, _40414_);
  or _47654_ (_41837_, _40429_, _40413_);
  and _47655_ (_40430_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _47656_ (_40431_, _40058_, _38658_);
  and _47657_ (_40432_, _40416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _47658_ (_40433_, _40432_, _40096_);
  or _47659_ (_40434_, _40123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _47660_ (_40435_, _40434_, _40062_);
  nor _47661_ (_40436_, _40435_, _40433_);
  and _47662_ (_40437_, _40417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _47663_ (_40438_, _40417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _47664_ (_40439_, _40438_, _40437_);
  and _47665_ (_40440_, _40439_, _40400_);
  or _47666_ (_40441_, _40440_, _40436_);
  or _47667_ (_40442_, _40441_, _40058_);
  and _47668_ (_40443_, _40442_, _40148_);
  and _47669_ (_40444_, _40443_, _40431_);
  or _47670_ (_41839_, _40444_, _40430_);
  nand _47671_ (_40445_, _40058_, _38650_);
  or _47672_ (_40446_, _40433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _47673_ (_40447_, _40446_, _40062_);
  and _47674_ (_40448_, _40433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _47675_ (_40449_, _40448_, _40447_);
  and _47676_ (_40450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47677_ (_40451_, _40134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _47678_ (_40452_, _40451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _47679_ (_40453_, _40451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47680_ (_40454_, _40453_, _40452_);
  and _47681_ (_40455_, _40454_, _40138_);
  or _47682_ (_40456_, _40455_, _40450_);
  or _47683_ (_40457_, _40456_, _40449_);
  or _47684_ (_40458_, _40457_, _40058_);
  and _47685_ (_40459_, _40458_, _40148_);
  and _47686_ (_40460_, _40459_, _40445_);
  and _47687_ (_40461_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _47688_ (_41840_, _40461_, _40460_);
  nand _47689_ (_40462_, _40058_, _38642_);
  and _47690_ (_40463_, _40432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47691_ (_40464_, _40463_, _40138_);
  and _47692_ (_40465_, _40448_, _40062_);
  nor _47693_ (_40466_, _40465_, _40464_);
  and _47694_ (_40467_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _47695_ (_40468_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _47696_ (_40469_, _40468_, _40467_);
  or _47697_ (_40470_, _40469_, _40058_);
  and _47698_ (_40471_, _40470_, _40148_);
  and _47699_ (_40472_, _40471_, _40462_);
  and _47700_ (_40473_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _47701_ (_41842_, _40473_, _40472_);
  nand _47702_ (_40474_, _40058_, _38635_);
  and _47703_ (_40475_, _40463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47704_ (_40476_, _40421_, _40475_);
  or _47705_ (_40477_, _40476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _47706_ (_40478_, _40476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47707_ (_40479_, _40478_, _40477_);
  or _47708_ (_40480_, _40479_, _40058_);
  and _47709_ (_40481_, _40480_, _40148_);
  and _47710_ (_40482_, _40481_, _40474_);
  and _47711_ (_40483_, _40115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _47712_ (_41844_, _40483_, _40482_);
  nor _47713_ (_40484_, _40204_, _40173_);
  or _47714_ (_40485_, _40484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47715_ (_40486_, _40195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47716_ (_40487_, _40220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47717_ (_40488_, _40487_, _40245_);
  nand _47718_ (_40489_, _40488_, _40486_);
  or _47719_ (_40490_, _40489_, _40173_);
  and _47720_ (_40491_, _40490_, _40485_);
  or _47721_ (_40492_, _40491_, _40212_);
  nand _47722_ (_40493_, _40212_, _38682_);
  and _47723_ (_40494_, _40493_, _43100_);
  and _47724_ (_41846_, _40494_, _40492_);
  not _47725_ (_40495_, _40214_);
  nor _47726_ (_40496_, _40486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _47727_ (_40497_, _40486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _47728_ (_40498_, _40497_, _40496_);
  and _47729_ (_40499_, _40220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _47730_ (_40500_, _40499_, _40201_);
  nor _47731_ (_40501_, _40500_, _40498_);
  nor _47732_ (_40502_, _40501_, _40173_);
  and _47733_ (_40503_, _40173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _47734_ (_40504_, _40503_, _40502_);
  and _47735_ (_40505_, _40504_, _40495_);
  nor _47736_ (_40506_, _40243_, _38672_);
  or _47737_ (_40507_, _40506_, _40505_);
  and _47738_ (_41848_, _40507_, _43100_);
  nor _47739_ (_40508_, _40497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _47740_ (_40509_, _40486_, _40196_);
  nor _47741_ (_40510_, _40509_, _40508_);
  and _47742_ (_40511_, _40220_, _40201_);
  and _47743_ (_40512_, _40511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _47744_ (_40513_, _40512_, _40510_);
  nor _47745_ (_40514_, _40513_, _40173_);
  and _47746_ (_40515_, _40173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _47747_ (_40516_, _40515_, _40514_);
  and _47748_ (_40517_, _40516_, _40495_);
  nor _47749_ (_40518_, _40243_, _38665_);
  or _47750_ (_40519_, _40518_, _40517_);
  and _47751_ (_41850_, _40519_, _43100_);
  and _47752_ (_40520_, _40198_, _40195_);
  nor _47753_ (_40521_, _40509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _47754_ (_40522_, _40521_, _40520_);
  and _47755_ (_40523_, _40511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _47756_ (_40524_, _40523_, _40522_);
  nor _47757_ (_40525_, _40524_, _40173_);
  and _47758_ (_40526_, _40173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _47759_ (_40527_, _40526_, _40525_);
  and _47760_ (_40528_, _40527_, _40495_);
  nor _47761_ (_40529_, _40243_, _38658_);
  or _47762_ (_40530_, _40529_, _40528_);
  and _47763_ (_41852_, _40530_, _43100_);
  nor _47764_ (_40531_, _40520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _47765_ (_40532_, _40531_, _40200_);
  and _47766_ (_40533_, _40511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _47767_ (_40534_, _40533_, _40532_);
  or _47768_ (_40535_, _40534_, _40173_);
  not _47769_ (_40536_, _40173_);
  or _47770_ (_40537_, _40536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _47771_ (_40538_, _40537_, _40243_);
  and _47772_ (_40539_, _40538_, _40535_);
  nor _47773_ (_40540_, _40243_, _38650_);
  or _47774_ (_40541_, _40540_, _40539_);
  and _47775_ (_41854_, _40541_, _43100_);
  nand _47776_ (_40542_, _40214_, _38642_);
  or _47777_ (_40543_, _40536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _47778_ (_40544_, _40511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47779_ (_40545_, _40200_, _40184_);
  or _47780_ (_40546_, _40545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _47781_ (_40547_, _40545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _47782_ (_40548_, _40547_);
  or _47783_ (_40549_, _40548_, _40173_);
  and _47784_ (_40550_, _40549_, _40546_);
  or _47785_ (_40551_, _40550_, _40544_);
  and _47786_ (_40552_, _40551_, _40543_);
  or _47787_ (_40553_, _40552_, _40214_);
  and _47788_ (_40554_, _40553_, _43100_);
  and _47789_ (_41855_, _40554_, _40542_);
  and _47790_ (_40555_, _40220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _47791_ (_40556_, _40555_, _40195_);
  and _47792_ (_40557_, _40556_, _40245_);
  nor _47793_ (_40558_, _40548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _47794_ (_40559_, _40558_, _40557_);
  nor _47795_ (_40560_, _40559_, _40173_);
  and _47796_ (_40561_, _40549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _47797_ (_40562_, _40561_, _40560_);
  and _47798_ (_40563_, _40562_, _40495_);
  nor _47799_ (_40564_, _40243_, _38635_);
  or _47800_ (_40565_, _40564_, _40563_);
  and _47801_ (_41857_, _40565_, _43100_);
  or _47802_ (_40566_, _40247_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47803_ (_40567_, _40566_, _40221_);
  and _47804_ (_40568_, _40247_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _47805_ (_40569_, _40568_, _40567_);
  and _47806_ (_40570_, _40254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _47807_ (_40571_, _40254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47808_ (_40572_, _40571_, _40223_);
  nor _47809_ (_40573_, _40572_, _40570_);
  and _47810_ (_40574_, _40200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _47811_ (_40575_, _40200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47812_ (_40576_, _40575_, _40183_);
  nor _47813_ (_40577_, _40576_, _40574_);
  or _47814_ (_40578_, _40577_, _40573_);
  or _47815_ (_40579_, _40578_, _40569_);
  or _47816_ (_40580_, _40579_, _40173_);
  nand _47817_ (_40581_, _40173_, _38682_);
  and _47818_ (_40582_, _40581_, _40580_);
  or _47819_ (_40583_, _40582_, _40214_);
  or _47820_ (_40584_, _40495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _47821_ (_40585_, _40584_, _43100_);
  and _47822_ (_41859_, _40585_, _40583_);
  nand _47823_ (_40586_, _40173_, _38672_);
  or _47824_ (_40587_, _40568_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _47825_ (_40588_, _40245_, _40195_);
  and _47826_ (_40589_, _40588_, _40176_);
  not _47827_ (_40590_, _40589_);
  or _47828_ (_40591_, _40590_, _40220_);
  and _47829_ (_40592_, _40591_, _40221_);
  and _47830_ (_40593_, _40592_, _40587_);
  not _47831_ (_40594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _47832_ (_40595_, _40570_, _40594_);
  and _47833_ (_40596_, _40570_, _40594_);
  or _47834_ (_40597_, _40596_, _40595_);
  and _47835_ (_40598_, _40597_, _40223_);
  and _47836_ (_40599_, _40574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _47837_ (_40600_, _40574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _47838_ (_40601_, _40600_, _40183_);
  nor _47839_ (_40602_, _40601_, _40599_);
  or _47840_ (_40603_, _40602_, _40598_);
  or _47841_ (_40604_, _40603_, _40593_);
  or _47842_ (_40605_, _40604_, _40173_);
  and _47843_ (_40606_, _40605_, _40243_);
  and _47844_ (_40607_, _40606_, _40586_);
  and _47845_ (_40608_, _40212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _47846_ (_40609_, _40608_, _40607_);
  and _47847_ (_41861_, _40609_, _43100_);
  nor _47848_ (_40610_, _40536_, _38665_);
  or _47849_ (_40611_, _40589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47850_ (_40612_, _40588_, _40177_);
  not _47851_ (_40613_, _40612_);
  and _47852_ (_40614_, _40613_, _40218_);
  and _47853_ (_40615_, _40614_, _40611_);
  or _47854_ (_40616_, _40599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47855_ (_40617_, _40200_, _40177_);
  nor _47856_ (_40618_, _40617_, _40184_);
  and _47857_ (_40619_, _40618_, _40616_);
  and _47858_ (_40620_, _40176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47859_ (_40621_, _40620_, _40254_);
  or _47860_ (_40622_, _40621_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47861_ (_40623_, _40254_, _40177_);
  nand _47862_ (_40624_, _40623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47863_ (_40625_, _40624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47864_ (_40626_, _40625_, _40622_);
  or _47865_ (_40627_, _40626_, _40619_);
  nor _47866_ (_40628_, _40627_, _40615_);
  nor _47867_ (_40629_, _40628_, _40173_);
  or _47868_ (_40630_, _40629_, _40214_);
  or _47869_ (_40631_, _40630_, _40610_);
  or _47870_ (_40632_, _40495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47871_ (_40633_, _40632_, _43100_);
  and _47872_ (_41863_, _40633_, _40631_);
  nor _47873_ (_40634_, _40536_, _38658_);
  not _47874_ (_40635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47875_ (_40636_, _40612_, _40217_);
  nor _47876_ (_40637_, _40636_, _40635_);
  and _47877_ (_40638_, _40636_, _40635_);
  or _47878_ (_40639_, _40638_, _40637_);
  and _47879_ (_40640_, _40639_, _40221_);
  or _47880_ (_40641_, _40623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _47881_ (_40642_, _40255_);
  and _47882_ (_40643_, _40642_, _40223_);
  and _47883_ (_40644_, _40643_, _40641_);
  or _47884_ (_40645_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47885_ (_40646_, _40200_, _40178_);
  nor _47886_ (_40647_, _40646_, _40184_);
  and _47887_ (_40648_, _40647_, _40645_);
  or _47888_ (_40649_, _40648_, _40644_);
  nor _47889_ (_40650_, _40649_, _40640_);
  nor _47890_ (_40651_, _40650_, _40173_);
  or _47891_ (_40652_, _40651_, _40214_);
  or _47892_ (_40653_, _40652_, _40634_);
  nand _47893_ (_40654_, _40214_, _40635_);
  and _47894_ (_40655_, _40654_, _43100_);
  and _47895_ (_41865_, _40655_, _40653_);
  nand _47896_ (_40656_, _40173_, _38650_);
  or _47897_ (_40657_, _40646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47898_ (_40658_, _40599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47899_ (_40659_, _40658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47900_ (_40660_, _40659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _47901_ (_40661_, _40660_, _40184_);
  and _47902_ (_40662_, _40661_, _40657_);
  and _47903_ (_40663_, _40588_, _40178_);
  or _47904_ (_40664_, _40663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _47905_ (_40665_, _40663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47906_ (_40666_, _40665_, _40218_);
  and _47907_ (_40667_, _40666_, _40664_);
  and _47908_ (_40668_, _40255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _47909_ (_40669_, _40668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47910_ (_40670_, _40669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47911_ (_40671_, _40255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _47912_ (_40672_, _40671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47913_ (_40673_, _40672_, _40670_);
  or _47914_ (_40674_, _40673_, _40667_);
  or _47915_ (_40675_, _40674_, _40662_);
  or _47916_ (_40676_, _40675_, _40173_);
  and _47917_ (_40677_, _40676_, _40243_);
  and _47918_ (_40678_, _40677_, _40656_);
  and _47919_ (_40679_, _40212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _47920_ (_40680_, _40679_, _40678_);
  and _47921_ (_41867_, _40680_, _43100_);
  nor _47922_ (_40681_, _40536_, _38642_);
  not _47923_ (_40682_, _40660_);
  nor _47924_ (_40683_, _40682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47925_ (_40684_, _40682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _47926_ (_40685_, _40684_, _40683_);
  and _47927_ (_40686_, _40685_, _40183_);
  nor _47928_ (_40687_, _40665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _47929_ (_40688_, _40687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _47930_ (_40689_, _40687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47931_ (_40690_, _40689_, _40221_);
  and _47932_ (_40691_, _40690_, _40688_);
  not _47933_ (_40692_, _40256_);
  and _47934_ (_40693_, _40692_, _40223_);
  or _47935_ (_40694_, _40671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47936_ (_40695_, _40694_, _40693_);
  or _47937_ (_40696_, _40695_, _40691_);
  or _47938_ (_40697_, _40696_, _40686_);
  and _47939_ (_40698_, _40697_, _40536_);
  or _47940_ (_40699_, _40698_, _40214_);
  or _47941_ (_40700_, _40699_, _40681_);
  or _47942_ (_40701_, _40495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47943_ (_40702_, _40701_, _43100_);
  and _47944_ (_41869_, _40702_, _40700_);
  nand _47945_ (_40703_, _40173_, _38635_);
  or _47946_ (_40704_, _40248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _47947_ (_40705_, _40704_, _40221_);
  nor _47948_ (_40706_, _40705_, _40249_);
  or _47949_ (_40707_, _40256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _47950_ (_40708_, _40257_);
  and _47951_ (_40709_, _40708_, _40223_);
  and _47952_ (_40710_, _40709_, _40707_);
  or _47953_ (_40711_, _40206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _47954_ (_40712_, _40271_, _40184_);
  and _47955_ (_40713_, _40712_, _40711_);
  or _47956_ (_40714_, _40713_, _40710_);
  or _47957_ (_40715_, _40714_, _40706_);
  or _47958_ (_40716_, _40715_, _40173_);
  and _47959_ (_40717_, _40716_, _40243_);
  and _47960_ (_40718_, _40717_, _40703_);
  and _47961_ (_40719_, _40212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _47962_ (_40720_, _40719_, _40718_);
  and _47963_ (_41870_, _40720_, _43100_);
  nor _47964_ (_40721_, _40289_, _40219_);
  and _47965_ (_40722_, _40289_, _38683_);
  or _47966_ (_40723_, _40722_, _40721_);
  and _47967_ (_41872_, _40723_, _43100_);
  or _47968_ (_40724_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47969_ (_40725_, _40724_, _43100_);
  nand _47970_ (_40726_, _40289_, _38672_);
  and _47971_ (_41874_, _40726_, _40725_);
  or _47972_ (_40727_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _47973_ (_40728_, _40727_, _43100_);
  nand _47974_ (_40729_, _40289_, _38665_);
  and _47975_ (_41876_, _40729_, _40728_);
  or _47976_ (_40730_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _47977_ (_40731_, _40730_, _43100_);
  nand _47978_ (_40732_, _40289_, _38658_);
  and _47979_ (_41877_, _40732_, _40731_);
  or _47980_ (_40733_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _47981_ (_40734_, _40733_, _43100_);
  nand _47982_ (_40735_, _40289_, _38650_);
  and _47983_ (_41879_, _40735_, _40734_);
  or _47984_ (_40736_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _47985_ (_40737_, _40736_, _43100_);
  nand _47986_ (_40738_, _40289_, _38642_);
  and _47987_ (_41881_, _40738_, _40737_);
  or _47988_ (_40739_, _40289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _47989_ (_40740_, _40739_, _43100_);
  nand _47990_ (_40741_, _40289_, _38635_);
  and _47991_ (_41883_, _40741_, _40740_);
  not _47992_ (_40742_, _27825_);
  nor _47993_ (_40743_, _39246_, _27650_);
  nand _47994_ (_40744_, _40743_, _40742_);
  nor _47995_ (_40745_, _40744_, _27496_);
  and _47996_ (_40746_, _40745_, _39451_);
  and _47997_ (_40747_, _40746_, _31308_);
  nand _47998_ (_40748_, _40747_, _31265_);
  and _47999_ (_40749_, _38617_, _31308_);
  and _48000_ (_40750_, _40749_, _39475_);
  nor _48001_ (_40751_, _40747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nor _48002_ (_40752_, _40751_, _40750_);
  and _48003_ (_40753_, _40752_, _40748_);
  and _48004_ (_40754_, _39469_, _30651_);
  and _48005_ (_40755_, _40754_, _40145_);
  or _48006_ (_40756_, _40755_, _40753_);
  and _48007_ (_43045_, _40756_, _43100_);
  and _48008_ (_40757_, _40113_, _27003_);
  and _48009_ (_40758_, _40757_, _39458_);
  not _48010_ (_40759_, _40758_);
  and _48011_ (_40760_, _27825_, _27661_);
  and _48012_ (_40761_, _40760_, _39247_);
  and _48013_ (_40762_, _40761_, _39451_);
  and _48014_ (_40763_, _40762_, _31308_);
  or _48015_ (_40764_, _40763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _48016_ (_40765_, _40764_, _40759_);
  nand _48017_ (_40766_, _40763_, _31265_);
  and _48018_ (_40767_, _40766_, _40765_);
  nor _48019_ (_40768_, _40759_, _38704_);
  or _48020_ (_40769_, _40768_, _40767_);
  and _48021_ (_43048_, _40769_, _43100_);
  and _48022_ (_40770_, _40757_, _38620_);
  and _48023_ (_40771_, _40743_, _27825_);
  and _48024_ (_40772_, _40771_, _27507_);
  and _48025_ (_40773_, _40772_, _39420_);
  nand _48026_ (_40774_, _40773_, _26981_);
  and _48027_ (_40775_, _40774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _48028_ (_40776_, _40775_, _40770_);
  or _48029_ (_40777_, _26992_, _33333_);
  and _48030_ (_40778_, _40777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _48031_ (_40779_, _40778_, _39222_);
  and _48032_ (_40780_, _40779_, _40773_);
  or _48033_ (_40781_, _40780_, _40776_);
  nand _48034_ (_40782_, _40770_, _38635_);
  and _48035_ (_40783_, _40782_, _43100_);
  and _48036_ (_43050_, _40783_, _40781_);
  not _48037_ (_40784_, _40770_);
  nor _48038_ (_40785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _48039_ (_40786_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _48040_ (_40787_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _48041_ (_40788_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _48042_ (_40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _48043_ (_40790_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40789_);
  and _48044_ (_40791_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48045_ (_40792_, _40791_, _40790_);
  nor _48046_ (_40793_, _40792_, _40788_);
  or _48047_ (_40794_, _40793_, _40787_);
  and _48048_ (_40795_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _48049_ (_40796_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _48050_ (_40797_, _40796_, _40795_);
  nor _48051_ (_40798_, _40797_, _40788_);
  and _48052_ (_40799_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40789_);
  and _48053_ (_40800_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48054_ (_40801_, _40800_, _40799_);
  nand _48055_ (_40802_, _40801_, _40798_);
  or _48056_ (_40803_, _40802_, _40794_);
  and _48057_ (_40804_, _40803_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _48058_ (_40805_, _40804_, _40786_);
  and _48059_ (_40806_, _38620_, _31308_);
  and _48060_ (_40807_, _40806_, _40743_);
  or _48061_ (_40809_, _40807_, _40805_);
  and _48062_ (_40811_, _40809_, _40784_);
  nand _48063_ (_40813_, _40807_, _31265_);
  and _48064_ (_40815_, _40813_, _40811_);
  nor _48065_ (_40817_, _40784_, _38704_);
  or _48066_ (_40819_, _40817_, _40815_);
  and _48067_ (_43052_, _40819_, _43100_);
  and _48068_ (_40822_, _40057_, _31351_);
  nand _48069_ (_40824_, _40822_, _31265_);
  not _48070_ (_40826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _48071_ (_40828_, _40826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _48072_ (_40830_, _40801_, _40788_);
  not _48073_ (_40832_, _40830_);
  or _48074_ (_40834_, _40832_, _40798_);
  or _48075_ (_40836_, _40834_, _40794_);
  and _48076_ (_40838_, _40836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _48077_ (_40840_, _40838_, _40828_);
  or _48078_ (_40842_, _40840_, _40822_);
  and _48079_ (_40844_, _40842_, _40784_);
  and _48080_ (_40846_, _40844_, _40824_);
  nor _48081_ (_40848_, _40784_, _38642_);
  or _48082_ (_40850_, _40848_, _40846_);
  and _48083_ (_43054_, _40850_, _43100_);
  not _48084_ (_40853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _48085_ (_40855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40853_);
  nand _48086_ (_40857_, _40793_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _48087_ (_40859_, _40830_, _40798_);
  or _48088_ (_40861_, _40859_, _40857_);
  and _48089_ (_40862_, _40861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _48090_ (_40863_, _40862_, _40855_);
  and _48091_ (_40864_, _40743_, _38622_);
  or _48092_ (_40865_, _40864_, _40863_);
  and _48093_ (_40866_, _40865_, _40784_);
  nand _48094_ (_40867_, _40864_, _31265_);
  and _48095_ (_40868_, _40867_, _40866_);
  nor _48096_ (_40869_, _40784_, _38672_);
  or _48097_ (_40870_, _40869_, _40868_);
  and _48098_ (_43056_, _40870_, _43100_);
  and _48099_ (_40871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _48100_ (_40872_, _40857_, _40834_);
  and _48101_ (_40873_, _40872_, _40871_);
  and _48102_ (_40874_, _40743_, _38751_);
  or _48103_ (_40875_, _40874_, _40873_);
  and _48104_ (_40876_, _40875_, _40784_);
  nand _48105_ (_40877_, _40874_, _31265_);
  and _48106_ (_40878_, _40877_, _40876_);
  nor _48107_ (_40879_, _40784_, _38658_);
  or _48108_ (_40880_, _40879_, _40878_);
  and _48109_ (_43058_, _40880_, _43100_);
  and _48110_ (_40881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _48111_ (_40882_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40789_);
  nor _48112_ (_40883_, _40882_, _40881_);
  and _48113_ (_40884_, _40883_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _48114_ (_40885_, _40884_, _40788_);
  and _48115_ (_40886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _48116_ (_40887_, _40886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _48117_ (_40888_, _40887_);
  and _48118_ (_40889_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _48119_ (_40890_, _40889_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _48120_ (_40891_, _40890_);
  and _48121_ (_40892_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _48122_ (_40893_, _40892_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _48123_ (_40894_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _48124_ (_40895_, _40894_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _48125_ (_40896_, _40895_, _40893_);
  and _48126_ (_40897_, _40896_, _40891_);
  and _48127_ (_40898_, _40897_, _40888_);
  not _48128_ (_40899_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _48129_ (_40900_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _48130_ (_40901_, _40900_, _40899_);
  nand _48131_ (_40902_, _40901_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _48132_ (_40903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _48133_ (_40904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _48134_ (_40905_, _40904_, _40903_);
  and _48135_ (_40906_, _40905_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _48136_ (_40907_, _40906_);
  and _48137_ (_40908_, _40907_, _40902_);
  and _48138_ (_40909_, _40908_, _40898_);
  nor _48139_ (_40910_, _40909_, _40885_);
  and _48140_ (_40911_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _48141_ (_40912_, _40911_, _40789_);
  and _48142_ (_40913_, _40912_, _40910_);
  not _48143_ (_40914_, _40913_);
  not _48144_ (_40915_, _40912_);
  and _48145_ (_40916_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40788_);
  not _48146_ (_40917_, _40916_);
  not _48147_ (_40918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _48148_ (_40919_, _40889_, _40918_);
  not _48149_ (_40920_, _40919_);
  not _48150_ (_40921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _48151_ (_40922_, _40892_, _40921_);
  not _48152_ (_40923_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _48153_ (_40924_, _40894_, _40923_);
  nor _48154_ (_40925_, _40924_, _40922_);
  and _48155_ (_40926_, _40925_, _40920_);
  nor _48156_ (_40927_, _40926_, _40917_);
  not _48157_ (_40928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _48158_ (_40929_, _40901_, _40928_);
  not _48159_ (_40930_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _48160_ (_40931_, _40905_, _40930_);
  nor _48161_ (_40932_, _40931_, _40929_);
  not _48162_ (_40933_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _48163_ (_40934_, _40886_, _40933_);
  not _48164_ (_40935_, _40934_);
  and _48165_ (_40936_, _40935_, _40932_);
  nor _48166_ (_40937_, _40936_, _40917_);
  nor _48167_ (_40938_, _40937_, _40927_);
  or _48168_ (_40939_, _40938_, _40915_);
  and _48169_ (_40940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _43100_);
  and _48170_ (_40941_, _40940_, _40939_);
  and _48171_ (_43087_, _40941_, _40914_);
  nor _48172_ (_40942_, _40911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _48173_ (_40943_, _40942_);
  not _48174_ (_40944_, _40910_);
  and _48175_ (_40945_, _40938_, _40944_);
  nor _48176_ (_40946_, _40945_, _40943_);
  nand _48177_ (_40947_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _43100_);
  nor _48178_ (_43089_, _40947_, _40946_);
  and _48179_ (_40948_, _40908_, _40888_);
  nand _48180_ (_40949_, _40948_, _40910_);
  or _48181_ (_40950_, _40937_, _40910_);
  and _48182_ (_40951_, _40950_, _40912_);
  and _48183_ (_40952_, _40951_, _40949_);
  or _48184_ (_40953_, _40952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _48185_ (_40954_, _40914_, _40897_);
  nor _48186_ (_40955_, _40915_, _40910_);
  nand _48187_ (_40956_, _40955_, _40927_);
  and _48188_ (_40957_, _40956_, _43100_);
  and _48189_ (_40958_, _40957_, _40954_);
  and _48190_ (_43091_, _40958_, _40953_);
  and _48191_ (_40959_, _40949_, _40942_);
  or _48192_ (_40960_, _40959_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _48193_ (_40961_, _40942_, _40910_);
  not _48194_ (_40962_, _40961_);
  or _48195_ (_40963_, _40962_, _40897_);
  or _48196_ (_40964_, _40937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand _48197_ (_40965_, _40942_, _40927_);
  and _48198_ (_40966_, _40965_, _40964_);
  or _48199_ (_40967_, _40966_, _40910_);
  and _48200_ (_40968_, _40967_, _43100_);
  and _48201_ (_40969_, _40968_, _40963_);
  and _48202_ (_43093_, _40969_, _40960_);
  nand _48203_ (_40970_, _40945_, _40788_);
  nor _48204_ (_40971_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _48205_ (_40972_, _40971_, _40911_);
  and _48206_ (_40973_, _40972_, _43100_);
  and _48207_ (_43094_, _40973_, _40970_);
  and _48208_ (_40974_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _48209_ (_40975_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _48210_ (_40976_, _40975_, _40971_);
  nor _48211_ (_40977_, _40976_, _40944_);
  or _48212_ (_40978_, _40977_, _40911_);
  or _48213_ (_40984_, _40978_, _40974_);
  not _48214_ (_40990_, _40911_);
  or _48215_ (_40996_, _40976_, _40990_);
  and _48216_ (_41002_, _40996_, _43100_);
  and _48217_ (_43096_, _41002_, _40984_);
  and _48218_ (_41006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _43100_);
  and _48219_ (_43098_, _41006_, _40911_);
  nor _48220_ (_43102_, _40785_, rst);
  and _48221_ (_43104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _43100_);
  nor _48222_ (_41007_, _40945_, _40911_);
  and _48223_ (_41008_, _40911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _48224_ (_41009_, _41008_, _41007_);
  and _48225_ (_00131_, _41009_, _43100_);
  and _48226_ (_41010_, _40911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _48227_ (_41011_, _41010_, _41007_);
  and _48228_ (_00133_, _41011_, _43100_);
  and _48229_ (_41012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _43100_);
  and _48230_ (_00135_, _41012_, _40911_);
  not _48231_ (_41015_, _40924_);
  nor _48232_ (_41019_, _40931_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _48233_ (_41023_, _41019_, _40929_);
  or _48234_ (_41024_, _41023_, _40934_);
  and _48235_ (_41025_, _41024_, _41015_);
  or _48236_ (_41026_, _41025_, _40922_);
  nor _48237_ (_41032_, _40938_, _40910_);
  and _48238_ (_41036_, _41032_, _40920_);
  and _48239_ (_41037_, _41036_, _41026_);
  not _48240_ (_41039_, _40895_);
  or _48241_ (_41040_, _40906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _48242_ (_41046_, _41040_, _40902_);
  or _48243_ (_41049_, _41046_, _40887_);
  and _48244_ (_41050_, _41049_, _41039_);
  or _48245_ (_41051_, _41050_, _40893_);
  and _48246_ (_41057_, _40910_, _40891_);
  and _48247_ (_41061_, _41057_, _41051_);
  or _48248_ (_41062_, _41061_, _40911_);
  or _48249_ (_41064_, _41062_, _41037_);
  or _48250_ (_41065_, _40990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _48251_ (_41073_, _41065_, _43100_);
  and _48252_ (_00137_, _41073_, _41064_);
  not _48253_ (_41074_, _40893_);
  or _48254_ (_41076_, _40895_, _40887_);
  and _48255_ (_41082_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _48256_ (_41085_, _41082_, _41076_);
  and _48257_ (_41086_, _41085_, _41074_);
  and _48258_ (_41087_, _41086_, _41057_);
  nor _48259_ (_41093_, _40922_, _40919_);
  or _48260_ (_41097_, _40934_, _40924_);
  and _48261_ (_41098_, _40932_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _48262_ (_41099_, _41098_, _41097_);
  and _48263_ (_41105_, _41099_, _41093_);
  and _48264_ (_41109_, _41105_, _41032_);
  or _48265_ (_41110_, _41109_, _40911_);
  or _48266_ (_41111_, _41110_, _41087_);
  or _48267_ (_41113_, _40990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _48268_ (_41119_, _41113_, _43100_);
  and _48269_ (_00139_, _41119_, _41111_);
  and _48270_ (_41122_, _40935_, _40916_);
  nand _48271_ (_41129_, _41122_, _40926_);
  nor _48272_ (_41130_, _41129_, _40932_);
  nor _48273_ (_41133_, _40908_, _40885_);
  or _48274_ (_41134_, _41133_, _41130_);
  or _48275_ (_41135_, _40898_, _40885_);
  and _48276_ (_41141_, _41135_, _41134_);
  or _48277_ (_41145_, _41141_, _40911_);
  or _48278_ (_41146_, _40990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _48279_ (_41147_, _41146_, _43100_);
  and _48280_ (_00140_, _41147_, _41145_);
  and _48281_ (_41156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _43100_);
  and _48282_ (_00142_, _41156_, _40911_);
  and _48283_ (_41157_, _40911_, _40789_);
  or _48284_ (_41161_, _41157_, _40946_);
  or _48285_ (_41167_, _41161_, _40955_);
  and _48286_ (_00144_, _41167_, _43100_);
  not _48287_ (_41168_, _41007_);
  and _48288_ (_41172_, _41168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _48289_ (_41178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _48290_ (_41179_, _40906_, _40789_);
  or _48291_ (_41180_, _41179_, _41178_);
  nor _48292_ (_41183_, _40902_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48293_ (_41189_, _41183_, _40887_);
  nand _48294_ (_41191_, _41189_, _41180_);
  or _48295_ (_41192_, _40888_, _40791_);
  and _48296_ (_41195_, _41192_, _41191_);
  or _48297_ (_41201_, _41195_, _40895_);
  or _48298_ (_41202_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40789_);
  or _48299_ (_41203_, _41202_, _41039_);
  and _48300_ (_41204_, _41203_, _41074_);
  and _48301_ (_41205_, _41204_, _41201_);
  and _48302_ (_41206_, _40893_, _40791_);
  or _48303_ (_41207_, _41206_, _40890_);
  or _48304_ (_41208_, _41207_, _41205_);
  or _48305_ (_41209_, _41202_, _40891_);
  and _48306_ (_41210_, _41209_, _40910_);
  and _48307_ (_41211_, _41210_, _41208_);
  and _48308_ (_41212_, _40931_, _40789_);
  or _48309_ (_41213_, _41212_, _41178_);
  and _48310_ (_41214_, _40929_, _40789_);
  nor _48311_ (_41215_, _41214_, _40934_);
  nand _48312_ (_41216_, _41215_, _41213_);
  or _48313_ (_41217_, _40935_, _40791_);
  and _48314_ (_41218_, _41217_, _41216_);
  or _48315_ (_41219_, _41218_, _40924_);
  not _48316_ (_41220_, _40922_);
  or _48317_ (_41221_, _41202_, _41015_);
  and _48318_ (_41222_, _41221_, _41220_);
  and _48319_ (_41223_, _41222_, _41219_);
  and _48320_ (_41224_, _40922_, _40791_);
  or _48321_ (_41225_, _41224_, _40919_);
  or _48322_ (_41226_, _41225_, _41223_);
  and _48323_ (_41227_, _41202_, _41032_);
  or _48324_ (_41228_, _41227_, _41036_);
  and _48325_ (_41229_, _41228_, _41226_);
  or _48326_ (_41230_, _41229_, _41211_);
  and _48327_ (_41231_, _41230_, _40990_);
  or _48328_ (_41232_, _41231_, _41172_);
  and _48329_ (_00146_, _41232_, _43100_);
  and _48330_ (_41233_, _41168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _48331_ (_41234_, _41179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _48332_ (_41235_, _41234_, _41189_);
  and _48333_ (_41236_, _40887_, _40800_);
  or _48334_ (_41237_, _41236_, _41235_);
  and _48335_ (_41238_, _41237_, _40896_);
  not _48336_ (_41239_, _40896_);
  or _48337_ (_41240_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40789_);
  and _48338_ (_41241_, _41240_, _41239_);
  or _48339_ (_41242_, _41241_, _40890_);
  or _48340_ (_41243_, _41242_, _41238_);
  or _48341_ (_41244_, _40891_, _40800_);
  and _48342_ (_41245_, _41244_, _40910_);
  and _48343_ (_41246_, _41245_, _41243_);
  and _48344_ (_41247_, _40919_, _40800_);
  and _48345_ (_41248_, _41240_, _40920_);
  or _48346_ (_41249_, _41248_, _40926_);
  and _48347_ (_41250_, _40934_, _40800_);
  not _48348_ (_41251_, _40925_);
  or _48349_ (_41252_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _48350_ (_41253_, _41252_, _41215_);
  or _48351_ (_41254_, _41253_, _41251_);
  or _48352_ (_41255_, _41254_, _41250_);
  and _48353_ (_41256_, _41255_, _41249_);
  or _48354_ (_41257_, _41256_, _41247_);
  and _48355_ (_41258_, _41257_, _41032_);
  or _48356_ (_41259_, _41258_, _41246_);
  and _48357_ (_41260_, _41259_, _40990_);
  or _48358_ (_41261_, _41260_, _41233_);
  and _48359_ (_00148_, _41261_, _43100_);
  and _48360_ (_41262_, _41168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _48361_ (_41263_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48362_ (_41264_, _41263_, _40891_);
  and _48363_ (_41265_, _41264_, _40910_);
  not _48364_ (_41266_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _48365_ (_41267_, _40906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48366_ (_41268_, _41267_, _41266_);
  nor _48367_ (_41269_, _40902_, _40789_);
  nor _48368_ (_41270_, _41269_, _40887_);
  nand _48369_ (_41271_, _41270_, _41268_);
  or _48370_ (_41272_, _40888_, _40790_);
  and _48371_ (_41273_, _41272_, _41271_);
  or _48372_ (_41274_, _41273_, _40895_);
  or _48373_ (_41275_, _41263_, _41039_);
  and _48374_ (_41276_, _41275_, _41074_);
  and _48375_ (_41277_, _41276_, _41274_);
  and _48376_ (_41278_, _40893_, _40790_);
  or _48377_ (_41279_, _41278_, _40890_);
  or _48378_ (_41280_, _41279_, _41277_);
  and _48379_ (_41281_, _41280_, _41265_);
  or _48380_ (_41282_, _41263_, _40920_);
  and _48381_ (_41283_, _40931_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48382_ (_41284_, _41283_, _41266_);
  and _48383_ (_41285_, _40929_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48384_ (_41286_, _41285_, _40934_);
  nand _48385_ (_41287_, _41286_, _41284_);
  or _48386_ (_41288_, _40935_, _40790_);
  and _48387_ (_41289_, _41288_, _41287_);
  or _48388_ (_41290_, _41289_, _40924_);
  or _48389_ (_41291_, _41263_, _41015_);
  and _48390_ (_41292_, _41291_, _41220_);
  and _48391_ (_41293_, _41292_, _41290_);
  and _48392_ (_41294_, _40922_, _40790_);
  or _48393_ (_41295_, _41294_, _40919_);
  or _48394_ (_41296_, _41295_, _41293_);
  and _48395_ (_41297_, _41296_, _41032_);
  and _48396_ (_41298_, _41297_, _41282_);
  or _48397_ (_41299_, _41298_, _41281_);
  and _48398_ (_41300_, _41299_, _40990_);
  or _48399_ (_41301_, _41300_, _41262_);
  and _48400_ (_00150_, _41301_, _43100_);
  and _48401_ (_41302_, _41168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _48402_ (_41303_, _41267_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _48403_ (_41304_, _41303_, _41270_);
  and _48404_ (_41305_, _40887_, _40799_);
  or _48405_ (_41306_, _41305_, _41304_);
  and _48406_ (_41307_, _41306_, _40896_);
  or _48407_ (_41308_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _48408_ (_41309_, _41308_, _41239_);
  or _48409_ (_41310_, _41309_, _40890_);
  or _48410_ (_41312_, _41310_, _41307_);
  or _48411_ (_41313_, _40891_, _40799_);
  and _48412_ (_41315_, _41313_, _40910_);
  and _48413_ (_41316_, _41315_, _41312_);
  and _48414_ (_41318_, _40919_, _40799_);
  and _48415_ (_41319_, _41308_, _40920_);
  or _48416_ (_41321_, _41319_, _40926_);
  and _48417_ (_41322_, _40934_, _40799_);
  or _48418_ (_41324_, _41283_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _48419_ (_41325_, _41324_, _41286_);
  or _48420_ (_41327_, _41325_, _41251_);
  or _48421_ (_41328_, _41327_, _41322_);
  and _48422_ (_41330_, _41328_, _41321_);
  or _48423_ (_41331_, _41330_, _41318_);
  and _48424_ (_41333_, _41331_, _41032_);
  or _48425_ (_41334_, _41333_, _41316_);
  and _48426_ (_41336_, _41334_, _40990_);
  or _48427_ (_41337_, _41336_, _41302_);
  and _48428_ (_00151_, _41337_, _43100_);
  or _48429_ (_41339_, _40943_, _40938_);
  and _48430_ (_41340_, _41339_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _48431_ (_41341_, _41340_, _40961_);
  and _48432_ (_00153_, _41341_, _43100_);
  and _48433_ (_41342_, _40939_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _48434_ (_41343_, _41342_, _40913_);
  and _48435_ (_00155_, _41343_, _43100_);
  and _48436_ (_41344_, _40773_, _27003_);
  or _48437_ (_41345_, _41344_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _48438_ (_41346_, _41345_, _40784_);
  nand _48439_ (_41347_, _41344_, _31265_);
  and _48440_ (_41348_, _41347_, _41346_);
  and _48441_ (_41349_, _40770_, _38683_);
  or _48442_ (_41350_, _41349_, _41348_);
  and _48443_ (_00157_, _41350_, _43100_);
  and _48444_ (_41351_, _40773_, _33344_);
  or _48445_ (_41352_, _41351_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _48446_ (_41353_, _41352_, _40784_);
  nand _48447_ (_41354_, _41351_, _31265_);
  and _48448_ (_41355_, _41354_, _41353_);
  nor _48449_ (_41356_, _40784_, _38665_);
  or _48450_ (_41357_, _41356_, _41355_);
  and _48451_ (_00159_, _41357_, _43100_);
  and _48452_ (_41358_, _40773_, _34791_);
  or _48453_ (_41359_, _41358_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _48454_ (_41360_, _41359_, _40784_);
  nand _48455_ (_41361_, _41358_, _31265_);
  and _48456_ (_41362_, _41361_, _41360_);
  nor _48457_ (_41363_, _40784_, _38650_);
  or _48458_ (_41364_, _41363_, _41362_);
  and _48459_ (_00161_, _41364_, _43100_);
  and _48460_ (_41365_, _40762_, _27003_);
  or _48461_ (_41366_, _41365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _48462_ (_41367_, _41366_, _40759_);
  nand _48463_ (_41368_, _41365_, _31265_);
  and _48464_ (_41369_, _41368_, _41367_);
  and _48465_ (_41370_, _40758_, _38683_);
  or _48466_ (_41371_, _41370_, _41369_);
  and _48467_ (_00162_, _41371_, _43100_);
  and _48468_ (_41372_, _40762_, _32604_);
  or _48469_ (_41373_, _41372_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _48470_ (_41374_, _41373_, _40759_);
  nand _48471_ (_41375_, _41372_, _31265_);
  and _48472_ (_41376_, _41375_, _41374_);
  nor _48473_ (_41377_, _40759_, _38672_);
  or _48474_ (_41378_, _41377_, _41376_);
  and _48475_ (_00164_, _41378_, _43100_);
  nand _48476_ (_41379_, _40762_, _39511_);
  and _48477_ (_41380_, _41379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _48478_ (_41381_, _41380_, _40758_);
  and _48479_ (_41382_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _48480_ (_41383_, _41382_, _33366_);
  and _48481_ (_41384_, _41383_, _40762_);
  or _48482_ (_41385_, _41384_, _41381_);
  nand _48483_ (_41386_, _40758_, _38665_);
  and _48484_ (_41387_, _41386_, _43100_);
  and _48485_ (_00166_, _41387_, _41385_);
  and _48486_ (_41388_, _40762_, _34052_);
  or _48487_ (_41389_, _41388_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _48488_ (_41390_, _41389_, _40759_);
  nand _48489_ (_41391_, _41388_, _31265_);
  and _48490_ (_41392_, _41391_, _41390_);
  nor _48491_ (_41393_, _40759_, _38658_);
  or _48492_ (_41394_, _41393_, _41392_);
  and _48493_ (_00168_, _41394_, _43100_);
  and _48494_ (_41395_, _40762_, _34791_);
  or _48495_ (_41396_, _41395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _48496_ (_41397_, _41396_, _40759_);
  nand _48497_ (_41398_, _41395_, _31265_);
  and _48498_ (_41399_, _41398_, _41397_);
  nor _48499_ (_41400_, _40759_, _38650_);
  or _48500_ (_41401_, _41400_, _41399_);
  and _48501_ (_00170_, _41401_, _43100_);
  and _48502_ (_41402_, _40762_, _35607_);
  or _48503_ (_41403_, _41402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _48504_ (_41404_, _41403_, _40759_);
  nand _48505_ (_41405_, _41402_, _31265_);
  and _48506_ (_41406_, _41405_, _41404_);
  nor _48507_ (_41407_, _40759_, _38642_);
  or _48508_ (_41408_, _41407_, _41406_);
  and _48509_ (_00172_, _41408_, _43100_);
  and _48510_ (_41409_, _40762_, _36336_);
  or _48511_ (_41410_, _41409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _48512_ (_41411_, _41410_, _40759_);
  nand _48513_ (_41412_, _41409_, _31265_);
  and _48514_ (_41413_, _41412_, _41411_);
  nor _48515_ (_41414_, _40759_, _38635_);
  or _48516_ (_41415_, _41414_, _41413_);
  and _48517_ (_00173_, _41415_, _43100_);
  and _48518_ (_41416_, _40746_, _27003_);
  nand _48519_ (_41417_, _41416_, _31265_);
  nor _48520_ (_41418_, _41416_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor _48521_ (_41419_, _41418_, _40750_);
  and _48522_ (_41420_, _41419_, _41417_);
  and _48523_ (_41421_, _40754_, _38683_);
  or _48524_ (_41422_, _41421_, _41420_);
  and _48525_ (_00175_, _41422_, _43100_);
  and _48526_ (_41423_, _40746_, _32604_);
  nand _48527_ (_41424_, _41423_, _31265_);
  nor _48528_ (_41425_, _41423_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _48529_ (_41426_, _41425_, _40750_);
  and _48530_ (_41427_, _41426_, _41424_);
  not _48531_ (_41428_, _38672_);
  and _48532_ (_41429_, _40754_, _41428_);
  or _48533_ (_41430_, _41429_, _41427_);
  and _48534_ (_00177_, _41430_, _43100_);
  and _48535_ (_41431_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _48536_ (_41432_, _41431_, _33366_);
  and _48537_ (_41433_, _41432_, _40746_);
  nand _48538_ (_41434_, _40746_, _39511_);
  and _48539_ (_41435_, _41434_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _48540_ (_41436_, _41435_, _40750_);
  or _48541_ (_41437_, _41436_, _41433_);
  nand _48542_ (_41438_, _40750_, _38665_);
  and _48543_ (_41439_, _41438_, _43100_);
  and _48544_ (_00179_, _41439_, _41437_);
  and _48545_ (_41440_, _40746_, _34052_);
  nand _48546_ (_41441_, _41440_, _31265_);
  nor _48547_ (_41442_, _41440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor _48548_ (_41443_, _41442_, _40750_);
  and _48549_ (_41444_, _41443_, _41441_);
  and _48550_ (_41445_, _40754_, _40346_);
  or _48551_ (_41446_, _41445_, _41444_);
  and _48552_ (_00181_, _41446_, _43100_);
  and _48553_ (_41447_, _40746_, _34791_);
  nand _48554_ (_41448_, _41447_, _31265_);
  nor _48555_ (_41449_, _41447_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor _48556_ (_41450_, _41449_, _40750_);
  and _48557_ (_41451_, _41450_, _41448_);
  and _48558_ (_41452_, _40754_, _40357_);
  or _48559_ (_41453_, _41452_, _41451_);
  and _48560_ (_00183_, _41453_, _43100_);
  not _48561_ (_41454_, _40750_);
  and _48562_ (_41455_, _40746_, _35607_);
  and _48563_ (_41456_, _41455_, _31265_);
  nor _48564_ (_41457_, _41455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _48565_ (_41458_, _41457_, _41456_);
  nand _48566_ (_41459_, _41458_, _41454_);
  nand _48567_ (_41460_, _40750_, _38642_);
  and _48568_ (_41461_, _41460_, _43100_);
  and _48569_ (_00184_, _41461_, _41459_);
  and _48570_ (_41462_, _40746_, _36336_);
  nand _48571_ (_41463_, _41462_, _31265_);
  nor _48572_ (_41464_, _41462_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor _48573_ (_41465_, _41464_, _40750_);
  and _48574_ (_41466_, _41465_, _41463_);
  and _48575_ (_41467_, _40754_, _40383_);
  or _48576_ (_41468_, _41467_, _41466_);
  and _48577_ (_00186_, _41468_, _43100_);
  and _48578_ (_41469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _48579_ (_41470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _48580_ (_41471_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _48581_ (_41472_, _41471_, _41470_);
  not _48582_ (_41473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _48583_ (_41474_, _41473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _48584_ (_41475_, _41474_, _41472_);
  nor _48585_ (_41476_, _41475_, _41469_);
  or _48586_ (_41477_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _48587_ (_41478_, _41477_, _43100_);
  nor _48588_ (_00546_, _41478_, _41476_);
  nor _48589_ (_41479_, _41476_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _48590_ (_41480_, _41479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _48591_ (_41481_, _41479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _48592_ (_41482_, _41481_, _43100_);
  and _48593_ (_00549_, _41482_, _41480_);
  not _48594_ (_41483_, rxd_i);
  and _48595_ (_41484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _41483_);
  nor _48596_ (_41485_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _48597_ (_41486_, _41485_);
  and _48598_ (_41487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _48599_ (_41488_, _41487_, _41486_);
  and _48600_ (_41489_, _41488_, _41484_);
  not _48601_ (_41490_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _48602_ (_41491_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _41490_);
  and _48603_ (_41492_, _41491_, _41485_);
  or _48604_ (_41493_, _41492_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or _48605_ (_41494_, _41493_, _41489_);
  and _48606_ (_41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _43100_);
  and _48607_ (_00552_, _41495_, _41494_);
  and _48608_ (_41496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _48609_ (_41497_, _41496_, _41486_);
  not _48610_ (_41498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _48611_ (_41499_, _41485_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48612_ (_41500_, _41499_, _41498_);
  nor _48613_ (_41501_, _41500_, _41497_);
  not _48614_ (_41502_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _48615_ (_41503_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _41502_);
  not _48616_ (_41504_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _48617_ (_41505_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _41504_);
  and _48618_ (_41506_, _41505_, _41503_);
  not _48619_ (_41507_, _41506_);
  or _48620_ (_41508_, _41507_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and _48621_ (_41509_, _41506_, _41497_);
  and _48622_ (_41510_, _41497_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48623_ (_41511_, _41510_, _41509_);
  and _48624_ (_41512_, _41511_, _41508_);
  or _48625_ (_41513_, _41512_, _41501_);
  not _48626_ (_41514_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand _48627_ (_41515_, _41485_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor _48628_ (_41516_, _41515_, _41514_);
  not _48629_ (_41517_, _41516_);
  or _48630_ (_41518_, _41517_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _48631_ (_41519_, _41518_, _41513_);
  nand _48632_ (_00554_, _41519_, _41495_);
  not _48633_ (_41520_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _48634_ (_41521_, _41497_);
  nor _48635_ (_41522_, _41498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _48636_ (_41523_, _41522_);
  not _48637_ (_41524_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48638_ (_41525_, _41485_, _41524_);
  and _48639_ (_41526_, _41525_, _41523_);
  and _48640_ (_41527_, _41526_, _41521_);
  nor _48641_ (_41528_, _41527_, _41520_);
  and _48642_ (_41529_, _41527_, rxd_i);
  or _48643_ (_41530_, _41529_, rst);
  or _48644_ (_00557_, _41530_, _41528_);
  nor _48645_ (_41531_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48646_ (_41532_, _41531_, _41503_);
  and _48647_ (_41533_, _41532_, _41510_);
  nand _48648_ (_41534_, _41533_, _41483_);
  or _48649_ (_41535_, _41533_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _48650_ (_41536_, _41535_, _43100_);
  and _48651_ (_00560_, _41536_, _41534_);
  and _48652_ (_41537_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48653_ (_41538_, _41537_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _48654_ (_41539_, _41538_, _41502_);
  and _48655_ (_41540_, _41539_, _41510_);
  and _48656_ (_41541_, _41488_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48657_ (_41542_, _41541_, _41510_);
  nor _48658_ (_41543_, _41538_, _41521_);
  or _48659_ (_41544_, _41543_, _41542_);
  and _48660_ (_41545_, _41544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _48661_ (_41546_, _41545_, _41540_);
  and _48662_ (_00562_, _41546_, _43100_);
  and _48663_ (_41547_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _43100_);
  nand _48664_ (_41548_, _41547_, _41524_);
  nand _48665_ (_41549_, _41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _48666_ (_00565_, _41549_, _41548_);
  and _48667_ (_41550_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41524_);
  not _48668_ (_41551_, _41488_);
  nand _48669_ (_41552_, _41492_, _41514_);
  and _48670_ (_41553_, _41552_, _41551_);
  nand _48671_ (_41554_, _41553_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _48672_ (_41555_, _41554_, _41521_);
  or _48673_ (_41556_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor _48674_ (_41557_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _48675_ (_41558_, _41557_, _41509_);
  and _48676_ (_41559_, _41558_, _41556_);
  and _48677_ (_41560_, _41559_, _41555_);
  or _48678_ (_41561_, _41560_, _41516_);
  nand _48679_ (_41562_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _48680_ (_41563_, _41562_, _41497_);
  or _48681_ (_41564_, _41563_, _41507_);
  and _48682_ (_41565_, _41564_, _41517_);
  or _48683_ (_41566_, _41565_, rxd_i);
  and _48684_ (_41567_, _41566_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48685_ (_41568_, _41567_, _41561_);
  or _48686_ (_41569_, _41568_, _41550_);
  and _48687_ (_00568_, _41569_, _43100_);
  and _48688_ (_41570_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _48689_ (_41571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _48690_ (_41572_, _41471_, _41571_);
  or _48691_ (_41573_, _41572_, _41474_);
  nor _48692_ (_41574_, _41573_, _41570_);
  or _48693_ (_41575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _48694_ (_41576_, _41575_, _43100_);
  nor _48695_ (_00571_, _41576_, _41574_);
  nor _48696_ (_41577_, _41574_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _48697_ (_41578_, _41577_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _48698_ (_41579_, _41577_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _48699_ (_41580_, _41579_, _43100_);
  and _48700_ (_00573_, _41580_, _41578_);
  not _48701_ (_41581_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _48702_ (_41582_, _32604_, _27661_);
  and _48703_ (_41583_, _41582_, _30651_);
  and _48704_ (_41584_, _41583_, _39442_);
  and _48705_ (_41585_, _41584_, _43100_);
  nand _48706_ (_41586_, _41585_, _41581_);
  not _48707_ (_41587_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _48708_ (_41588_, _41515_, _41587_);
  nor _48709_ (_41589_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not _48710_ (_41590_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _48711_ (_41591_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _48712_ (_41592_, _41591_, _41590_);
  and _48713_ (_41593_, _41592_, _41589_);
  not _48714_ (_41594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _48715_ (_41595_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _48716_ (_41596_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _48717_ (_41597_, _41596_, _41595_);
  and _48718_ (_41598_, _41597_, _41594_);
  and _48719_ (_41599_, _41598_, _41593_);
  or _48720_ (_41600_, _41599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _48721_ (_41601_, _41599_, _41581_);
  nand _48722_ (_41602_, _41601_, _41600_);
  nand _48723_ (_41603_, _41602_, _41588_);
  nor _48724_ (_41604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _48725_ (_41605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _48726_ (_41606_, _41605_, _41604_);
  and _48727_ (_41607_, _41486_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _48728_ (_41608_, _41607_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _48729_ (_41609_, _41608_, _41606_);
  not _48730_ (_41610_, _41609_);
  or _48731_ (_41611_, _41610_, _41600_);
  and _48732_ (_41612_, _41606_, _41607_);
  or _48733_ (_41613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _41587_);
  or _48734_ (_41614_, _41613_, _41612_);
  or _48735_ (_41615_, _41614_, _41588_);
  and _48736_ (_41616_, _41615_, _41611_);
  nand _48737_ (_41617_, _41616_, _41603_);
  nor _48738_ (_41618_, _41584_, rst);
  nand _48739_ (_41619_, _41618_, _41617_);
  and _48740_ (_00576_, _41619_, _41586_);
  not _48741_ (_41620_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and _48742_ (_41621_, _41599_, _41620_);
  nand _48743_ (_41622_, _41612_, _41621_);
  and _48744_ (_41623_, _41599_, _41588_);
  or _48745_ (_41624_, _41587_, rst);
  nor _48746_ (_41625_, _41624_, _41623_);
  and _48747_ (_41626_, _41625_, _41622_);
  or _48748_ (_00579_, _41626_, _41585_);
  or _48749_ (_41627_, _41610_, _41621_);
  or _48750_ (_41628_, _41612_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _48751_ (_41629_, _41515_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _48752_ (_41630_, _41629_, _41628_);
  and _48753_ (_41631_, _41630_, _41627_);
  or _48754_ (_41632_, _41631_, _41623_);
  and _48755_ (_00581_, _41632_, _41618_);
  and _48756_ (_41633_, _41608_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _48757_ (_41634_, _41633_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _48758_ (_41635_, _41634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or _48759_ (_41636_, _41635_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _48760_ (_41637_, _41635_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _48761_ (_41638_, _41637_, _41636_);
  and _48762_ (_00584_, _41638_, _41618_);
  nor _48763_ (_41639_, _41609_, _41588_);
  and _48764_ (_41640_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _48765_ (_41641_, _41640_, _41618_);
  and _48766_ (_41642_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _48767_ (_00587_, _41642_, _41641_);
  and _48768_ (_41643_, _40749_, _38620_);
  or _48769_ (_41644_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _48770_ (_41645_, _41644_, _43100_);
  nand _48771_ (_41646_, _41643_, _38704_);
  and _48772_ (_00589_, _41646_, _41645_);
  and _48773_ (_41647_, _40745_, _39420_);
  and _48774_ (_41648_, _41647_, _31308_);
  nand _48775_ (_41649_, _41648_, _31265_);
  and _48776_ (_41650_, _40757_, _39442_);
  nor _48777_ (_41651_, _41648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _48778_ (_41652_, _41651_, _41650_);
  and _48779_ (_41653_, _41652_, _41649_);
  not _48780_ (_41654_, _41650_);
  nor _48781_ (_41655_, _41654_, _38704_);
  or _48782_ (_41656_, _41655_, _41653_);
  and _48783_ (_00592_, _41656_, _43100_);
  nor _48784_ (_41657_, _41516_, _41509_);
  not _48785_ (_41658_, _41657_);
  nor _48786_ (_41659_, _41553_, _41497_);
  nor _48787_ (_41660_, _41659_, _41658_);
  nor _48788_ (_41661_, _41660_, _41524_);
  or _48789_ (_41662_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _48790_ (_41663_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _41524_);
  or _48791_ (_41664_, _41663_, _41657_);
  and _48792_ (_41665_, _41664_, _43100_);
  and _48793_ (_01211_, _41665_, _41662_);
  or _48794_ (_41666_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _48795_ (_41667_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _41524_);
  or _48796_ (_41668_, _41667_, _41657_);
  and _48797_ (_41669_, _41668_, _43100_);
  and _48798_ (_01213_, _41669_, _41666_);
  or _48799_ (_41670_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _48800_ (_41671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41524_);
  or _48801_ (_41672_, _41671_, _41657_);
  and _48802_ (_41673_, _41672_, _43100_);
  and _48803_ (_01215_, _41673_, _41670_);
  or _48804_ (_41674_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _48805_ (_41675_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41524_);
  or _48806_ (_41676_, _41675_, _41657_);
  and _48807_ (_41677_, _41676_, _43100_);
  and _48808_ (_01217_, _41677_, _41674_);
  or _48809_ (_41678_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _48810_ (_41679_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41524_);
  or _48811_ (_41680_, _41679_, _41657_);
  and _48812_ (_41681_, _41680_, _43100_);
  and _48813_ (_01219_, _41681_, _41678_);
  or _48814_ (_41682_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _48815_ (_41683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41524_);
  or _48816_ (_41684_, _41683_, _41657_);
  and _48817_ (_41685_, _41684_, _43100_);
  and _48818_ (_01221_, _41685_, _41682_);
  or _48819_ (_41686_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _48820_ (_41687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41524_);
  or _48821_ (_41688_, _41687_, _41657_);
  and _48822_ (_41689_, _41688_, _43100_);
  and _48823_ (_01223_, _41689_, _41686_);
  or _48824_ (_41690_, _41661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _48825_ (_41691_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _41524_);
  or _48826_ (_41692_, _41691_, _41657_);
  and _48827_ (_41693_, _41692_, _43100_);
  and _48828_ (_01224_, _41693_, _41690_);
  nor _48829_ (_41694_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _48830_ (_41695_, _41694_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _48831_ (_41696_, _41507_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or _48832_ (_41697_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _48833_ (_41698_, _41697_, _41497_);
  and _48834_ (_41699_, _41698_, _41696_);
  or _48835_ (_41700_, _41488_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _48836_ (_41701_, _41700_, _41552_);
  and _48837_ (_41702_, _41701_, _41521_);
  or _48838_ (_41703_, _41702_, _41699_);
  or _48839_ (_41704_, _41703_, _41516_);
  or _48840_ (_41705_, _41517_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _48841_ (_41706_, _41705_, _41495_);
  and _48842_ (_41707_, _41706_, _41704_);
  or _48843_ (_01226_, _41707_, _41695_);
  and _48844_ (_41708_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _48845_ (_41709_, _41708_, _41553_);
  or _48846_ (_41710_, _41709_, _41660_);
  and _48847_ (_41711_, _41710_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _48848_ (_41712_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _41524_);
  nand _48849_ (_41713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48850_ (_41714_, _41713_, _41657_);
  or _48851_ (_41715_, _41714_, _41712_);
  or _48852_ (_41716_, _41715_, _41711_);
  and _48853_ (_01228_, _41716_, _43100_);
  not _48854_ (_41717_, _41661_);
  and _48855_ (_41718_, _41717_, _41547_);
  or _48856_ (_41719_, _41709_, _41658_);
  and _48857_ (_41720_, _41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _48858_ (_41721_, _41720_, _41719_);
  or _48859_ (_01230_, _41721_, _41718_);
  or _48860_ (_41722_, _41540_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _48861_ (_41723_, _41540_, _41483_);
  and _48862_ (_41724_, _41723_, _43100_);
  and _48863_ (_01232_, _41724_, _41722_);
  or _48864_ (_41725_, _41542_, _41504_);
  or _48865_ (_41726_, _41510_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48866_ (_41727_, _41726_, _43100_);
  and _48867_ (_01234_, _41727_, _41725_);
  and _48868_ (_41728_, _41542_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _48869_ (_41729_, _41531_, _41537_);
  and _48870_ (_41730_, _41729_, _41510_);
  or _48871_ (_41731_, _41730_, _41728_);
  and _48872_ (_01236_, _41731_, _43100_);
  and _48873_ (_41732_, _41544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _48874_ (_41733_, _41537_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48875_ (_41734_, _41733_, _41543_);
  or _48876_ (_41735_, _41734_, _41732_);
  and _48877_ (_01238_, _41735_, _43100_);
  and _48878_ (_41736_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41524_);
  and _48879_ (_41737_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48880_ (_41738_, _41737_, _41736_);
  and _48881_ (_01240_, _41738_, _43100_);
  and _48882_ (_41739_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41524_);
  and _48883_ (_41740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48884_ (_41741_, _41740_, _41739_);
  and _48885_ (_01242_, _41741_, _43100_);
  and _48886_ (_41742_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41524_);
  and _48887_ (_41743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48888_ (_41744_, _41743_, _41742_);
  and _48889_ (_01244_, _41744_, _43100_);
  and _48890_ (_41745_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41524_);
  and _48891_ (_41746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48892_ (_41747_, _41746_, _41745_);
  and _48893_ (_01246_, _41747_, _43100_);
  and _48894_ (_41748_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41524_);
  and _48895_ (_41749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48896_ (_41750_, _41749_, _41748_);
  and _48897_ (_01248_, _41750_, _43100_);
  and _48898_ (_41751_, _41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _48899_ (_01250_, _41751_, _41695_);
  and _48900_ (_41752_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48901_ (_41753_, _41752_, _41712_);
  and _48902_ (_01252_, _41753_, _43100_);
  nor _48903_ (_41754_, _41608_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _48904_ (_41755_, _41754_, _41633_);
  and _48905_ (_01254_, _41755_, _41618_);
  nor _48906_ (_41756_, _41633_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _48907_ (_41757_, _41756_, _41634_);
  and _48908_ (_01256_, _41757_, _41618_);
  nor _48909_ (_41758_, _41634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _48910_ (_41759_, _41758_, _41635_);
  and _48911_ (_01258_, _41759_, _41618_);
  and _48912_ (_41760_, _41609_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _48913_ (_41761_, _41588_, _41620_);
  nor _48914_ (_41762_, _41761_, _41609_);
  or _48915_ (_41763_, _41762_, _41760_);
  and _48916_ (_41764_, _41599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _48917_ (_41765_, _41764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _48918_ (_41766_, _41765_, _41588_);
  nor _48919_ (_41767_, _41766_, _41763_);
  nor _48920_ (_41768_, _41767_, _41584_);
  nor _48921_ (_41769_, _41486_, _38682_);
  and _48922_ (_41770_, _41769_, _41584_);
  or _48923_ (_41771_, _41770_, _41768_);
  and _48924_ (_01259_, _41771_, _43100_);
  not _48925_ (_41772_, _41639_);
  and _48926_ (_41773_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _48927_ (_41774_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _48928_ (_41775_, _41774_, _41773_);
  and _48929_ (_41776_, _41775_, _41618_);
  nand _48930_ (_41777_, _41485_, _38672_);
  nand _48931_ (_41778_, _41486_, _38682_);
  and _48932_ (_41779_, _41778_, _41585_);
  and _48933_ (_41780_, _41779_, _41777_);
  or _48934_ (_01261_, _41780_, _41776_);
  nor _48935_ (_41781_, _41639_, _41594_);
  and _48936_ (_41782_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or _48937_ (_41783_, _41782_, _41781_);
  and _48938_ (_41784_, _41783_, _41618_);
  nand _48939_ (_41785_, _41485_, _38665_);
  nand _48940_ (_41786_, _41486_, _38672_);
  and _48941_ (_41787_, _41786_, _41585_);
  and _48942_ (_41788_, _41787_, _41785_);
  or _48943_ (_01263_, _41788_, _41784_);
  nor _48944_ (_41789_, _41639_, _41590_);
  and _48945_ (_41790_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _48946_ (_41791_, _41790_, _41789_);
  and _48947_ (_41792_, _41791_, _41618_);
  nand _48948_ (_41793_, _41486_, _38665_);
  nand _48949_ (_41794_, _41485_, _38658_);
  and _48950_ (_41795_, _41794_, _41585_);
  and _48951_ (_41796_, _41795_, _41793_);
  or _48952_ (_01265_, _41796_, _41792_);
  and _48953_ (_41797_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _48954_ (_41798_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or _48955_ (_41799_, _41798_, _41797_);
  and _48956_ (_41800_, _41799_, _41618_);
  nand _48957_ (_41801_, _41485_, _38650_);
  nand _48958_ (_41802_, _41486_, _38658_);
  and _48959_ (_41803_, _41802_, _41585_);
  and _48960_ (_41804_, _41803_, _41801_);
  or _48961_ (_01267_, _41804_, _41800_);
  and _48962_ (_41805_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _48963_ (_41806_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _48964_ (_41807_, _41806_, _41805_);
  and _48965_ (_41808_, _41807_, _41618_);
  nand _48966_ (_41809_, _41486_, _38650_);
  nand _48967_ (_41810_, _41485_, _38642_);
  and _48968_ (_41811_, _41810_, _41585_);
  and _48969_ (_41812_, _41811_, _41809_);
  or _48970_ (_01269_, _41812_, _41808_);
  and _48971_ (_41813_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _48972_ (_41814_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or _48973_ (_41815_, _41814_, _41813_);
  and _48974_ (_41816_, _41815_, _41618_);
  nand _48975_ (_41817_, _41485_, _38635_);
  nand _48976_ (_41818_, _41486_, _38642_);
  and _48977_ (_41819_, _41818_, _41585_);
  and _48978_ (_41821_, _41819_, _41817_);
  or _48979_ (_01271_, _41821_, _41816_);
  and _48980_ (_41824_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _48981_ (_41826_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _48982_ (_41828_, _41826_, _41824_);
  and _48983_ (_41830_, _41828_, _41618_);
  nand _48984_ (_41832_, _41485_, _38704_);
  nand _48985_ (_41834_, _41486_, _38635_);
  and _48986_ (_41836_, _41834_, _41585_);
  and _48987_ (_41838_, _41836_, _41832_);
  or _48988_ (_01273_, _41838_, _41830_);
  and _48989_ (_41841_, _41584_, _41486_);
  nand _48990_ (_41843_, _41841_, _38704_);
  or _48991_ (_41845_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _48992_ (_41847_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _48993_ (_41849_, _41847_, _41845_);
  or _48994_ (_41851_, _41849_, _41584_);
  and _48995_ (_41853_, _41851_, _43100_);
  and _48996_ (_01275_, _41853_, _41843_);
  and _48997_ (_41856_, _41772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _48998_ (_41858_, _41639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _48999_ (_41860_, _41858_, _41856_);
  and _49000_ (_41862_, _41860_, _41618_);
  or _49001_ (_41864_, _41473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _49002_ (_41866_, _41864_, _41486_);
  and _49003_ (_41868_, _41866_, _41585_);
  or _49004_ (_01277_, _41868_, _41862_);
  nand _49005_ (_41871_, _41643_, _38682_);
  or _49006_ (_41873_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _49007_ (_41875_, _41873_, _43100_);
  and _49008_ (_01279_, _41875_, _41871_);
  or _49009_ (_41878_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _49010_ (_41880_, _41878_, _43100_);
  nand _49011_ (_41882_, _41643_, _38672_);
  and _49012_ (_01281_, _41882_, _41880_);
  or _49013_ (_41884_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _49014_ (_41885_, _41884_, _43100_);
  nand _49015_ (_41886_, _41643_, _38665_);
  and _49016_ (_01283_, _41886_, _41885_);
  or _49017_ (_41887_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _49018_ (_41888_, _41887_, _43100_);
  nand _49019_ (_41889_, _41643_, _38658_);
  and _49020_ (_01285_, _41889_, _41888_);
  or _49021_ (_41890_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _49022_ (_41891_, _41890_, _43100_);
  nand _49023_ (_41892_, _41643_, _38650_);
  and _49024_ (_01287_, _41892_, _41891_);
  or _49025_ (_41893_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _49026_ (_41894_, _41893_, _43100_);
  nand _49027_ (_41895_, _41643_, _38642_);
  and _49028_ (_01289_, _41895_, _41894_);
  or _49029_ (_41896_, _41643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _49030_ (_41897_, _41896_, _43100_);
  nand _49031_ (_41898_, _41643_, _38635_);
  and _49032_ (_01291_, _41898_, _41897_);
  not _49033_ (_41899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _49034_ (_41900_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41899_);
  or _49035_ (_41901_, _41900_, _41485_);
  nor _49036_ (_41902_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _49037_ (_41903_, _41902_, _41901_);
  or _49038_ (_41904_, _41903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _49039_ (_41905_, _41904_, _41647_);
  or _49040_ (_41906_, _27003_, _41490_);
  nand _49041_ (_41907_, _41906_, _41647_);
  or _49042_ (_41908_, _41907_, _39268_);
  and _49043_ (_41909_, _41908_, _41905_);
  or _49044_ (_41910_, _41909_, _41650_);
  nand _49045_ (_41911_, _41650_, _38682_);
  and _49046_ (_41912_, _41911_, _43100_);
  and _49047_ (_01293_, _41912_, _41910_);
  or _49048_ (_41913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _49049_ (_41914_, _41913_, _41647_);
  not _49050_ (_41915_, _32604_);
  nor _49051_ (_41916_, _41915_, _31265_);
  nand _49052_ (_41917_, _41915_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _49053_ (_41918_, _41917_, _41647_);
  or _49054_ (_41919_, _41918_, _41916_);
  and _49055_ (_41920_, _41919_, _41914_);
  or _49056_ (_41921_, _41920_, _41650_);
  nand _49057_ (_41922_, _41650_, _38672_);
  and _49058_ (_41923_, _41922_, _43100_);
  and _49059_ (_01294_, _41923_, _41921_);
  not _49060_ (_41924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not _49061_ (_41925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _49062_ (_41926_, _41499_, _41925_);
  nor _49063_ (_41927_, _41926_, _41924_);
  and _49064_ (_41928_, _41926_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _49065_ (_41929_, _41928_, _41927_);
  or _49066_ (_41930_, _41929_, _41647_);
  or _49067_ (_41931_, _33344_, _41924_);
  nand _49068_ (_41932_, _41931_, _41647_);
  or _49069_ (_41933_, _41932_, _33366_);
  and _49070_ (_41934_, _41933_, _41930_);
  or _49071_ (_41935_, _41934_, _41650_);
  nand _49072_ (_41936_, _41650_, _38665_);
  and _49073_ (_41937_, _41936_, _43100_);
  and _49074_ (_01296_, _41937_, _41935_);
  and _49075_ (_41938_, _41647_, _34052_);
  nand _49076_ (_41939_, _41938_, _31265_);
  nor _49077_ (_41940_, _41938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor _49078_ (_41941_, _41940_, _41650_);
  and _49079_ (_41942_, _41941_, _41939_);
  nor _49080_ (_41943_, _41654_, _38658_);
  or _49081_ (_41944_, _41943_, _41942_);
  and _49082_ (_01298_, _41944_, _43100_);
  and _49083_ (_41945_, _41647_, _34791_);
  nand _49084_ (_41946_, _41945_, _31265_);
  nor _49085_ (_41947_, _41945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _49086_ (_41948_, _41947_, _41650_);
  and _49087_ (_41949_, _41948_, _41946_);
  nor _49088_ (_41950_, _41654_, _38650_);
  or _49089_ (_41951_, _41950_, _41949_);
  and _49090_ (_01300_, _41951_, _43100_);
  and _49091_ (_41952_, _41647_, _35607_);
  nand _49092_ (_41953_, _41952_, _31265_);
  nor _49093_ (_41954_, _41952_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nor _49094_ (_41955_, _41954_, _41650_);
  and _49095_ (_41956_, _41955_, _41953_);
  nor _49096_ (_41957_, _41654_, _38642_);
  or _49097_ (_41958_, _41957_, _41956_);
  and _49098_ (_01302_, _41958_, _43100_);
  and _49099_ (_41959_, _41647_, _36336_);
  nand _49100_ (_41960_, _41959_, _31265_);
  nor _49101_ (_41961_, _41959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nor _49102_ (_41962_, _41961_, _41650_);
  and _49103_ (_41963_, _41962_, _41960_);
  nor _49104_ (_41964_, _41654_, _38635_);
  or _49105_ (_41965_, _41964_, _41963_);
  and _49106_ (_01304_, _41965_, _43100_);
  and _49107_ (_01630_, t2_i, _43100_);
  nor _49108_ (_41966_, t2_i, rst);
  and _49109_ (_01633_, _41966_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand _49110_ (_41967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _43100_);
  nor _49111_ (_01636_, _41967_, t2ex_i);
  and _49112_ (_01639_, t2ex_i, _43100_);
  and _49113_ (_41968_, _38618_, _39112_);
  and _49114_ (_41969_, _41968_, _40211_);
  nand _49115_ (_41970_, _41969_, _38704_);
  and _49116_ (_41971_, _40113_, _34052_);
  and _49117_ (_41972_, _41968_, _41971_);
  not _49118_ (_41973_, _41972_);
  and _49119_ (_41974_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _49120_ (_41975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _49121_ (_41976_, _41975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _49122_ (_41977_, _41976_, _41974_);
  not _49123_ (_41978_, _41977_);
  and _49124_ (_41979_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _49125_ (_41980_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _49126_ (_41981_, _41980_, _41979_);
  or _49127_ (_41982_, _41969_, _41981_);
  and _49128_ (_41983_, _41982_, _41973_);
  and _49129_ (_41984_, _41983_, _41970_);
  and _49130_ (_41985_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _49131_ (_41986_, _41985_, _41984_);
  and _49132_ (_01642_, _41986_, _43100_);
  nand _49133_ (_41987_, _41972_, _38704_);
  nor _49134_ (_41988_, _41969_, _41978_);
  or _49135_ (_41989_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not _49136_ (_41990_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _49137_ (_41991_, _41988_, _41990_);
  and _49138_ (_41992_, _41991_, _41989_);
  or _49139_ (_41993_, _41992_, _41972_);
  and _49140_ (_41994_, _41993_, _43100_);
  and _49141_ (_01645_, _41994_, _41987_);
  and _49142_ (_41995_, _41968_, _35607_);
  and _49143_ (_41996_, _41995_, _40113_);
  and _49144_ (_41997_, _41968_, _40172_);
  nor _49145_ (_41998_, _41997_, _41996_);
  not _49146_ (_41999_, _41975_);
  or _49147_ (_42000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _49148_ (_42001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _49149_ (_42002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _42001_);
  and _49150_ (_42003_, _42002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _49151_ (_42004_, _42003_, _42000_);
  and _49152_ (_42005_, _42004_, _41999_);
  and _49153_ (_42006_, _42005_, _41998_);
  and _49154_ (_42007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49155_ (_42008_, _42007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _49156_ (_42009_, _42008_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _49157_ (_42010_, _42009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _49158_ (_42011_, _42010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _49159_ (_42012_, _42011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _49160_ (_42013_, _42012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _49161_ (_42014_, _42013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _49162_ (_42015_, _42014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _49163_ (_42016_, _42015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _49164_ (_42017_, _42016_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _49165_ (_42018_, _42017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _49166_ (_42019_, _42018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _49167_ (_42020_, _42019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _49168_ (_42021_, _42020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not _49169_ (_42022_, _42021_);
  nand _49170_ (_42023_, _42022_, _42006_);
  or _49171_ (_42024_, _42006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _49172_ (_42025_, _42024_, _43100_);
  and _49173_ (_01648_, _42025_, _42023_);
  nand _49174_ (_42026_, _41997_, _38704_);
  not _49175_ (_42027_, _41996_);
  not _49176_ (_42028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _49177_ (_42029_, _41974_, _42028_);
  and _49178_ (_42030_, _42029_, _41975_);
  and _49179_ (_42031_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not _49180_ (_42032_, _42030_);
  not _49181_ (_42033_, _41976_);
  and _49182_ (_42034_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _49183_ (_42035_, _42021_, _42004_);
  and _49184_ (_42036_, _42035_, _42034_);
  and _49185_ (_42037_, _42012_, _42004_);
  or _49186_ (_42038_, _42037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _49187_ (_42039_, _42037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _49188_ (_42040_, _42039_, _42038_);
  or _49189_ (_42041_, _42040_, _42036_);
  and _49190_ (_42042_, _42041_, _42032_);
  or _49191_ (_42043_, _42042_, _42031_);
  or _49192_ (_42044_, _42043_, _41997_);
  and _49193_ (_42045_, _42044_, _42027_);
  and _49194_ (_42046_, _42045_, _42026_);
  and _49195_ (_42047_, _41996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _49196_ (_42048_, _42047_, _42046_);
  and _49197_ (_01651_, _42048_, _43100_);
  nand _49198_ (_42049_, _41996_, _38704_);
  nor _49199_ (_42050_, _42030_, _41990_);
  and _49200_ (_42051_, _42032_, _42004_);
  and _49201_ (_42052_, _42051_, _42020_);
  or _49202_ (_42053_, _42052_, _42050_);
  nand _49203_ (_42054_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _49204_ (_42055_, _42054_, _42035_);
  and _49205_ (_42056_, _42055_, _42053_);
  nand _49206_ (_42057_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _49207_ (_42058_, _42057_, _41998_);
  or _49208_ (_42059_, _42058_, _42056_);
  nand _49209_ (_42060_, _41997_, _41990_);
  and _49210_ (_42061_, _42060_, _43100_);
  and _49211_ (_42062_, _42061_, _42059_);
  and _49212_ (_01654_, _42062_, _42049_);
  and _49213_ (_42063_, _41975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _49214_ (_42064_, _42063_, _42052_);
  nand _49215_ (_42065_, _42064_, _41998_);
  or _49216_ (_42066_, _41998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49217_ (_42067_, _42066_, _43100_);
  and _49218_ (_01657_, _42067_, _42065_);
  or _49219_ (_42068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49220_ (_42069_, _40761_, _39096_);
  or _49221_ (_42070_, _42069_, _42068_);
  nand _49222_ (_42071_, _39099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _49223_ (_42072_, _42071_, _42069_);
  or _49224_ (_42073_, _42072_, _39100_);
  and _49225_ (_42074_, _42073_, _42070_);
  and _49226_ (_42075_, _41968_, _40757_);
  or _49227_ (_42076_, _42075_, _42074_);
  nand _49228_ (_42077_, _42075_, _38704_);
  and _49229_ (_42078_, _42077_, _43100_);
  and _49230_ (_01660_, _42078_, _42076_);
  not _49231_ (_42079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor _49232_ (_42080_, _41977_, _42079_);
  and _49233_ (_42081_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _49234_ (_42082_, _42081_, _42080_);
  or _49235_ (_42083_, _42082_, _41969_);
  nand _49236_ (_42084_, _41969_, _38682_);
  and _49237_ (_42085_, _42084_, _42083_);
  or _49238_ (_42086_, _42085_, _41972_);
  nand _49239_ (_42087_, _41972_, _42079_);
  and _49240_ (_42088_, _42087_, _43100_);
  and _49241_ (_02112_, _42088_, _42086_);
  nand _49242_ (_42089_, _41969_, _38672_);
  and _49243_ (_42090_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _49244_ (_42091_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _49245_ (_42092_, _42091_, _42090_);
  or _49246_ (_42093_, _42092_, _41969_);
  and _49247_ (_42094_, _42093_, _41973_);
  and _49248_ (_42095_, _42094_, _42089_);
  and _49249_ (_42096_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _49250_ (_42097_, _42096_, _42095_);
  and _49251_ (_02114_, _42097_, _43100_);
  nand _49252_ (_42098_, _41969_, _38665_);
  and _49253_ (_42099_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _49254_ (_42100_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _49255_ (_42101_, _42100_, _42099_);
  or _49256_ (_42102_, _42101_, _41969_);
  and _49257_ (_42103_, _42102_, _41973_);
  and _49258_ (_42104_, _42103_, _42098_);
  and _49259_ (_42105_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _49260_ (_42106_, _42105_, _42104_);
  and _49261_ (_02116_, _42106_, _43100_);
  not _49262_ (_42107_, _41969_);
  nor _49263_ (_42108_, _42107_, _38658_);
  and _49264_ (_42109_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49265_ (_42110_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _49266_ (_42111_, _42110_, _42109_);
  nor _49267_ (_42112_, _42111_, _41969_);
  or _49268_ (_42113_, _42112_, _41972_);
  or _49269_ (_42114_, _42113_, _42108_);
  or _49270_ (_42115_, _41973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49271_ (_42116_, _42115_, _43100_);
  and _49272_ (_02117_, _42116_, _42114_);
  nand _49273_ (_42117_, _41969_, _38650_);
  and _49274_ (_42118_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49275_ (_42119_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _49276_ (_42120_, _42119_, _42118_);
  or _49277_ (_42121_, _42120_, _41969_);
  and _49278_ (_42122_, _42121_, _41973_);
  and _49279_ (_42123_, _42122_, _42117_);
  and _49280_ (_42124_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _49281_ (_42125_, _42124_, _42123_);
  and _49282_ (_02119_, _42125_, _43100_);
  nand _49283_ (_42126_, _41969_, _38642_);
  and _49284_ (_42127_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _49285_ (_42128_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _49286_ (_42129_, _42128_, _42127_);
  or _49287_ (_42130_, _42129_, _41969_);
  and _49288_ (_42131_, _42130_, _41973_);
  and _49289_ (_42132_, _42131_, _42126_);
  and _49290_ (_42133_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _49291_ (_42134_, _42133_, _42132_);
  and _49292_ (_02121_, _42134_, _43100_);
  nand _49293_ (_42135_, _41969_, _38635_);
  and _49294_ (_42136_, _41978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _49295_ (_42137_, _41977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _49296_ (_42138_, _42137_, _42136_);
  or _49297_ (_42139_, _42138_, _41969_);
  and _49298_ (_42140_, _42139_, _41973_);
  and _49299_ (_42141_, _42140_, _42135_);
  and _49300_ (_42142_, _41972_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _49301_ (_42143_, _42142_, _42141_);
  and _49302_ (_02123_, _42143_, _43100_);
  or _49303_ (_42144_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not _49304_ (_42145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _49305_ (_42146_, _41988_, _42145_);
  and _49306_ (_42147_, _42146_, _42144_);
  or _49307_ (_42148_, _42147_, _41972_);
  nand _49308_ (_42149_, _41972_, _38682_);
  and _49309_ (_42150_, _42149_, _43100_);
  and _49310_ (_02124_, _42150_, _42148_);
  not _49311_ (_42151_, _41988_);
  and _49312_ (_42152_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _49313_ (_42153_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _49314_ (_42154_, _42153_, _42152_);
  or _49315_ (_42155_, _42154_, _41972_);
  nand _49316_ (_42156_, _41972_, _38672_);
  and _49317_ (_42157_, _42156_, _43100_);
  and _49318_ (_02126_, _42157_, _42155_);
  nand _49319_ (_42158_, _41972_, _38665_);
  and _49320_ (_42159_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _49321_ (_42160_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _49322_ (_42161_, _42160_, _42159_);
  or _49323_ (_42162_, _42161_, _41972_);
  and _49324_ (_42163_, _42162_, _43100_);
  and _49325_ (_02128_, _42163_, _42158_);
  nand _49326_ (_42164_, _41972_, _38658_);
  and _49327_ (_42165_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _49328_ (_42166_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49329_ (_42167_, _42166_, _42165_);
  or _49330_ (_42168_, _42167_, _41972_);
  and _49331_ (_42169_, _42168_, _43100_);
  and _49332_ (_02130_, _42169_, _42164_);
  nand _49333_ (_42170_, _41972_, _38650_);
  and _49334_ (_42171_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _49335_ (_42172_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _49336_ (_42173_, _42172_, _42171_);
  or _49337_ (_42174_, _42173_, _41972_);
  and _49338_ (_42175_, _42174_, _43100_);
  and _49339_ (_02131_, _42175_, _42170_);
  nand _49340_ (_42176_, _41972_, _38642_);
  and _49341_ (_42177_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _49342_ (_42178_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _49343_ (_42179_, _42178_, _42177_);
  or _49344_ (_42180_, _42179_, _41972_);
  and _49345_ (_42181_, _42180_, _43100_);
  and _49346_ (_02133_, _42181_, _42176_);
  nand _49347_ (_42182_, _41972_, _38635_);
  and _49348_ (_42183_, _42151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _49349_ (_42184_, _41988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _49350_ (_42185_, _42184_, _42183_);
  or _49351_ (_42186_, _42185_, _41972_);
  and _49352_ (_42187_, _42186_, _43100_);
  and _49353_ (_02135_, _42187_, _42182_);
  and _49354_ (_42188_, _42004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _49355_ (_42189_, _41976_, _42079_);
  nand _49356_ (_42190_, _42189_, _42021_);
  nand _49357_ (_42191_, _42190_, _42188_);
  or _49358_ (_42192_, _42004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49359_ (_42193_, _42192_, _42032_);
  and _49360_ (_42194_, _42193_, _42191_);
  and _49361_ (_42195_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _49362_ (_42196_, _42195_, _41997_);
  or _49363_ (_42197_, _42196_, _42194_);
  and _49364_ (_42198_, _41997_, _38682_);
  nor _49365_ (_42199_, _42198_, _41996_);
  and _49366_ (_42200_, _42199_, _42197_);
  and _49367_ (_42201_, _41996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _49368_ (_42202_, _42201_, _42200_);
  and _49369_ (_02137_, _42202_, _43100_);
  and _49370_ (_42203_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _49371_ (_42204_, _42203_, _42051_);
  and _49372_ (_42205_, _42204_, _42021_);
  and _49373_ (_42206_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _49374_ (_42207_, _42188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _49375_ (_42208_, _42007_, _42004_);
  nor _49376_ (_42209_, _42208_, _42030_);
  and _49377_ (_42210_, _42209_, _42207_);
  nor _49378_ (_42211_, _42210_, _42206_);
  nand _49379_ (_42212_, _42211_, _41998_);
  or _49380_ (_42213_, _42212_, _42205_);
  nand _49381_ (_42214_, _41997_, _38672_);
  or _49382_ (_42215_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _49383_ (_42216_, _42215_, _43100_);
  and _49384_ (_42217_, _42216_, _42214_);
  and _49385_ (_02138_, _42217_, _42213_);
  and _49386_ (_42218_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _49387_ (_42219_, _42218_, _42035_);
  not _49388_ (_42220_, _42208_);
  nor _49389_ (_42221_, _42220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _49390_ (_42222_, _42220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _49391_ (_42223_, _42222_, _42221_);
  or _49392_ (_42224_, _42223_, _42219_);
  and _49393_ (_42225_, _42224_, _42032_);
  nand _49394_ (_42226_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand _49395_ (_42227_, _42226_, _41998_);
  or _49396_ (_42228_, _42227_, _42225_);
  nand _49397_ (_42229_, _41997_, _38665_);
  or _49398_ (_42230_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _49399_ (_42231_, _42230_, _43100_);
  and _49400_ (_42232_, _42231_, _42229_);
  and _49401_ (_02140_, _42232_, _42228_);
  not _49402_ (_42233_, _41997_);
  and _49403_ (_42234_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49404_ (_42235_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49405_ (_42236_, _42235_, _42035_);
  nand _49406_ (_42237_, _42008_, _42004_);
  nor _49407_ (_42238_, _42237_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _49408_ (_42239_, _42237_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _49409_ (_42240_, _42239_, _42238_);
  or _49410_ (_42241_, _42240_, _42236_);
  and _49411_ (_42242_, _42241_, _42032_);
  or _49412_ (_42243_, _42242_, _42234_);
  and _49413_ (_42244_, _42243_, _42233_);
  nor _49414_ (_42245_, _42233_, _38658_);
  or _49415_ (_42246_, _42245_, _42244_);
  and _49416_ (_42247_, _42246_, _42027_);
  and _49417_ (_42248_, _41996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _49418_ (_42249_, _42248_, _42247_);
  and _49419_ (_02142_, _42249_, _43100_);
  and _49420_ (_42250_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49421_ (_42251_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49422_ (_42252_, _42251_, _42035_);
  nand _49423_ (_42253_, _42009_, _42004_);
  nor _49424_ (_42254_, _42253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _49425_ (_42255_, _42253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _49426_ (_42256_, _42255_, _42254_);
  or _49427_ (_42257_, _42256_, _42252_);
  and _49428_ (_42258_, _42257_, _42032_);
  or _49429_ (_42259_, _42258_, _42250_);
  and _49430_ (_42260_, _42259_, _42233_);
  nor _49431_ (_42261_, _42233_, _38650_);
  or _49432_ (_42262_, _42261_, _41996_);
  or _49433_ (_42263_, _42262_, _42260_);
  or _49434_ (_42264_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _49435_ (_42265_, _42264_, _43100_);
  and _49436_ (_02144_, _42265_, _42263_);
  and _49437_ (_42266_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _49438_ (_42267_, _42266_, _42035_);
  nand _49439_ (_42268_, _42010_, _42004_);
  nor _49440_ (_42269_, _42268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _49441_ (_42270_, _42268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _49442_ (_42271_, _42270_, _42269_);
  or _49443_ (_42272_, _42271_, _42267_);
  and _49444_ (_42273_, _42272_, _42032_);
  nand _49445_ (_42274_, _42030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand _49446_ (_42275_, _42274_, _41998_);
  or _49447_ (_42276_, _42275_, _42273_);
  nand _49448_ (_42277_, _41997_, _38642_);
  or _49449_ (_42278_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _49450_ (_42279_, _42278_, _43100_);
  and _49451_ (_42280_, _42279_, _42277_);
  and _49452_ (_02145_, _42280_, _42276_);
  nor _49453_ (_42281_, _42233_, _38635_);
  and _49454_ (_42282_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _49455_ (_42283_, _42282_, _42035_);
  and _49456_ (_42284_, _42011_, _42004_);
  nor _49457_ (_42285_, _42284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _49458_ (_42286_, _42285_, _42037_);
  or _49459_ (_42287_, _42286_, _42030_);
  or _49460_ (_42288_, _42287_, _42283_);
  or _49461_ (_42289_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _49462_ (_42290_, _42289_, _41998_);
  and _49463_ (_42291_, _42290_, _42288_);
  and _49464_ (_42292_, _41996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _49465_ (_42293_, _42292_, _42291_);
  or _49466_ (_42294_, _42293_, _42281_);
  and _49467_ (_02147_, _42294_, _43100_);
  not _49468_ (_42295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _49469_ (_42296_, _41976_, _42295_);
  and _49470_ (_42297_, _42296_, _42035_);
  and _49471_ (_42298_, _42013_, _42004_);
  or _49472_ (_42299_, _42298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _49473_ (_42300_, _42298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _49474_ (_42301_, _42300_, _42299_);
  or _49475_ (_42302_, _42301_, _42030_);
  or _49476_ (_42303_, _42302_, _42297_);
  nand _49477_ (_42304_, _42030_, _42295_);
  and _49478_ (_42305_, _42304_, _41998_);
  and _49479_ (_42306_, _42305_, _42303_);
  and _49480_ (_42307_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _49481_ (_42308_, _41996_, _38683_);
  or _49482_ (_42309_, _42308_, _42307_);
  or _49483_ (_42310_, _42309_, _42306_);
  and _49484_ (_02149_, _42310_, _43100_);
  and _49485_ (_42311_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _49486_ (_42312_, _42311_, _42035_);
  and _49487_ (_42313_, _42014_, _42004_);
  or _49488_ (_42314_, _42313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _49489_ (_42315_, _42313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _49490_ (_42316_, _42315_, _42314_);
  or _49491_ (_42317_, _42316_, _42030_);
  or _49492_ (_42318_, _42317_, _42312_);
  not _49493_ (_42319_, _41998_);
  nor _49494_ (_42320_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _49495_ (_42321_, _42320_, _42319_);
  and _49496_ (_42322_, _42321_, _42318_);
  and _49497_ (_42323_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _49498_ (_42324_, _42027_, _38672_);
  or _49499_ (_42325_, _42324_, _42323_);
  or _49500_ (_42326_, _42325_, _42322_);
  and _49501_ (_02151_, _42326_, _43100_);
  and _49502_ (_42327_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _49503_ (_42328_, _42327_, _42035_);
  and _49504_ (_42329_, _42015_, _42004_);
  or _49505_ (_42330_, _42329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand _49506_ (_42331_, _42329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _49507_ (_42332_, _42331_, _42330_);
  or _49508_ (_42333_, _42332_, _42030_);
  or _49509_ (_42334_, _42333_, _42328_);
  nor _49510_ (_42335_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _49511_ (_42336_, _42335_, _42319_);
  and _49512_ (_42337_, _42336_, _42334_);
  nor _49513_ (_42338_, _42027_, _38665_);
  and _49514_ (_42339_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _49515_ (_42340_, _42339_, _42338_);
  or _49516_ (_42341_, _42340_, _42337_);
  and _49517_ (_02152_, _42341_, _43100_);
  and _49518_ (_42342_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _49519_ (_42343_, _42342_, _42035_);
  nand _49520_ (_42344_, _42016_, _42004_);
  nor _49521_ (_42345_, _42344_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _49522_ (_42346_, _42344_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49523_ (_42347_, _42346_, _42030_);
  or _49524_ (_42348_, _42347_, _42345_);
  or _49525_ (_42349_, _42348_, _42343_);
  or _49526_ (_42350_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _49527_ (_42351_, _42350_, _41998_);
  and _49528_ (_42352_, _42351_, _42349_);
  and _49529_ (_42353_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49530_ (_42354_, _42353_, _42352_);
  nor _49531_ (_42355_, _42027_, _38658_);
  or _49532_ (_42356_, _42355_, _42354_);
  and _49533_ (_02154_, _42356_, _43100_);
  and _49534_ (_42357_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _49535_ (_42358_, _42357_, _42035_);
  nand _49536_ (_42359_, _42017_, _42004_);
  nor _49537_ (_42360_, _42359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _49538_ (_42361_, _42359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _49539_ (_42362_, _42361_, _42030_);
  or _49540_ (_42363_, _42362_, _42360_);
  or _49541_ (_42364_, _42363_, _42358_);
  or _49542_ (_42365_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _49543_ (_42366_, _42365_, _41998_);
  and _49544_ (_42367_, _42366_, _42364_);
  and _49545_ (_42368_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _49546_ (_42369_, _42368_, _42367_);
  nor _49547_ (_42370_, _42027_, _38650_);
  or _49548_ (_42371_, _42370_, _42369_);
  and _49549_ (_02156_, _42371_, _43100_);
  and _49550_ (_42372_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _49551_ (_42373_, _42372_, _42035_);
  nand _49552_ (_42374_, _42018_, _42004_);
  and _49553_ (_42375_, _42374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _49554_ (_42376_, _42374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _49555_ (_42377_, _42376_, _42030_);
  or _49556_ (_42378_, _42377_, _42375_);
  or _49557_ (_42379_, _42378_, _42373_);
  or _49558_ (_42380_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _49559_ (_42381_, _42380_, _41998_);
  and _49560_ (_42382_, _42381_, _42379_);
  and _49561_ (_42383_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _49562_ (_42384_, _42027_, _38642_);
  or _49563_ (_42385_, _42384_, _42383_);
  or _49564_ (_42386_, _42385_, _42382_);
  and _49565_ (_02158_, _42386_, _43100_);
  and _49566_ (_42387_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _49567_ (_42388_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _49568_ (_42389_, _42388_, _42035_);
  nand _49569_ (_42390_, _42019_, _42004_);
  and _49570_ (_42391_, _42390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _49571_ (_42392_, _42390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _49572_ (_42393_, _42392_, _42030_);
  or _49573_ (_42394_, _42393_, _42391_);
  or _49574_ (_42395_, _42394_, _42389_);
  or _49575_ (_42396_, _42032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _49576_ (_42397_, _42396_, _41998_);
  and _49577_ (_42398_, _42397_, _42395_);
  or _49578_ (_42399_, _42398_, _42387_);
  nor _49579_ (_42400_, _42027_, _38635_);
  or _49580_ (_42401_, _42400_, _42399_);
  and _49581_ (_02159_, _42401_, _43100_);
  not _49582_ (_42402_, _42075_);
  and _49583_ (_42403_, _42069_, _27003_);
  or _49584_ (_42404_, _42403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _49585_ (_42405_, _42404_, _42402_);
  nand _49586_ (_42406_, _42403_, _31265_);
  and _49587_ (_42407_, _42406_, _42405_);
  and _49588_ (_42408_, _42075_, _38683_);
  or _49589_ (_42409_, _42408_, _42407_);
  and _49590_ (_02161_, _42409_, _43100_);
  and _49591_ (_42410_, _42069_, _32604_);
  or _49592_ (_42411_, _42410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _49593_ (_42412_, _42411_, _42402_);
  nand _49594_ (_42413_, _42410_, _31265_);
  and _49595_ (_42414_, _42413_, _42412_);
  nor _49596_ (_42415_, _42402_, _38672_);
  or _49597_ (_42416_, _42415_, _42414_);
  and _49598_ (_02163_, _42416_, _43100_);
  nand _49599_ (_42417_, _42069_, _39511_);
  and _49600_ (_42418_, _42417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _49601_ (_42419_, _42418_, _42075_);
  and _49602_ (_42420_, _33377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _49603_ (_42421_, _42420_, _33366_);
  and _49604_ (_42422_, _42421_, _42069_);
  or _49605_ (_42423_, _42422_, _42419_);
  nand _49606_ (_42424_, _42075_, _38665_);
  and _49607_ (_42425_, _42424_, _43100_);
  and _49608_ (_02165_, _42425_, _42423_);
  and _49609_ (_42426_, _42069_, _34052_);
  or _49610_ (_42427_, _42426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _49611_ (_42428_, _42427_, _42402_);
  nand _49612_ (_42429_, _42426_, _31265_);
  and _49613_ (_42430_, _42429_, _42428_);
  nor _49614_ (_42431_, _42402_, _38658_);
  or _49615_ (_42432_, _42431_, _42430_);
  and _49616_ (_02166_, _42432_, _43100_);
  and _49617_ (_42433_, _42069_, _34791_);
  or _49618_ (_42434_, _42433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _49619_ (_42435_, _42434_, _42402_);
  nand _49620_ (_42436_, _42433_, _31265_);
  and _49621_ (_42437_, _42436_, _42435_);
  nor _49622_ (_42438_, _42402_, _38650_);
  or _49623_ (_42439_, _42438_, _42437_);
  and _49624_ (_02167_, _42439_, _43100_);
  and _49625_ (_42440_, _42069_, _35607_);
  or _49626_ (_42441_, _42440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _49627_ (_42442_, _42441_, _42402_);
  nand _49628_ (_42443_, _42440_, _31265_);
  and _49629_ (_42444_, _42443_, _42442_);
  nor _49630_ (_42445_, _42402_, _38642_);
  or _49631_ (_42446_, _42445_, _42444_);
  and _49632_ (_02168_, _42446_, _43100_);
  not _49633_ (_42447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49634_ (_42448_, _41974_, _42447_);
  or _49635_ (_42449_, _42448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _49636_ (_42450_, _42449_, _42069_);
  nand _49637_ (_42451_, _39221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _49638_ (_42452_, _42451_, _42069_);
  or _49639_ (_42453_, _42452_, _39222_);
  and _49640_ (_42454_, _42453_, _42450_);
  or _49641_ (_42455_, _42454_, _42075_);
  nand _49642_ (_42456_, _42075_, _38635_);
  and _49643_ (_42457_, _42456_, _43100_);
  and _49644_ (_02169_, _42457_, _42455_);
  nor _49645_ (_42458_, _27496_, _26476_);
  nor _49646_ (_42459_, _42458_, _30629_);
  and _49647_ (_42460_, _38706_, _38615_);
  not _49648_ (_42461_, _42460_);
  not _49649_ (_42462_, _38614_);
  and _49650_ (_42463_, _42462_, _38577_);
  nand _49651_ (_42464_, _38006_, _26981_);
  or _49652_ (_42465_, _38006_, _26981_);
  not _49653_ (_42466_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _49654_ (_42467_, _30618_, _42466_);
  and _49655_ (_42468_, _42467_, _33377_);
  and _49656_ (_42469_, _42468_, _27496_);
  and _49657_ (_42470_, _42469_, _42465_);
  and _49658_ (_42471_, _42470_, _42464_);
  and _49659_ (_42472_, _39111_, _39112_);
  and _49660_ (_42473_, _42472_, _39113_);
  not _49661_ (_42474_, _42473_);
  and _49662_ (_42475_, _42474_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _49663_ (_42476_, _42475_, _39168_);
  and _49664_ (_42477_, _42476_, _27661_);
  nor _49665_ (_42478_, _42476_, _27661_);
  nor _49666_ (_42479_, _42478_, _42477_);
  and _49667_ (_42480_, _42479_, _42471_);
  not _49668_ (_42481_, _42480_);
  and _49669_ (_42482_, _42476_, _38479_);
  and _49670_ (_42483_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor _49671_ (_42484_, _42476_, _38006_);
  and _49672_ (_42485_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _49673_ (_42486_, _42485_, _42483_);
  nor _49674_ (_42487_, _42476_, _38479_);
  and _49675_ (_42488_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _49676_ (_42489_, _42476_, _38006_);
  and _49677_ (_42490_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor _49678_ (_42491_, _42490_, _42488_);
  and _49679_ (_42492_, _42491_, _42486_);
  and _49680_ (_42493_, _42492_, _42481_);
  and _49681_ (_42494_, _42480_, _38704_);
  nor _49682_ (_42495_, _42494_, _42493_);
  and _49683_ (_42496_, _42495_, _42463_);
  not _49684_ (_42497_, _42496_);
  not _49685_ (_42498_, _38477_);
  nor _49686_ (_42499_, _42462_, _38577_);
  not _49687_ (_42500_, _36509_);
  and _49688_ (_42501_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and _49689_ (_42502_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _49690_ (_42503_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _49691_ (_42504_, _42503_, _42502_);
  and _49692_ (_42505_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _49693_ (_42506_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _49694_ (_42507_, _42506_, _42505_);
  and _49695_ (_42508_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _49696_ (_42509_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _49697_ (_42510_, _42509_, _42508_);
  and _49698_ (_42511_, _42510_, _42507_);
  and _49699_ (_42512_, _42511_, _42504_);
  and _49700_ (_42513_, _38017_, _36509_);
  not _49701_ (_42514_, _42513_);
  nor _49702_ (_42515_, _42514_, _42512_);
  nor _49703_ (_42516_, _42515_, _42501_);
  not _49704_ (_42517_, _42516_);
  and _49705_ (_42518_, _42517_, _42499_);
  nor _49706_ (_42519_, _42518_, _42498_);
  and _49707_ (_42520_, _42519_, _42497_);
  and _49708_ (_42521_, _42520_, _42461_);
  not _49709_ (_42522_, _38550_);
  and _49710_ (_42523_, _42522_, _38544_);
  nor _49711_ (_42524_, _38539_, _38535_);
  nor _49712_ (_42525_, _38547_, _38532_);
  and _49713_ (_42526_, _42525_, _42524_);
  and _49714_ (_42527_, _38561_, _38523_);
  and _49715_ (_42528_, _42527_, _42526_);
  and _49716_ (_42529_, _42528_, _42523_);
  nor _49717_ (_42530_, _42529_, _36466_);
  nor _49718_ (_42531_, _38559_, _38555_);
  not _49719_ (_42532_, _38466_);
  nor _49720_ (_42533_, _42532_, _42531_);
  nor _49721_ (_42534_, _42533_, _42530_);
  not _49722_ (_42535_, _42534_);
  and _49723_ (_42536_, _42535_, _42521_);
  and _49724_ (_42537_, _42499_, _38477_);
  and _49725_ (_42538_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and _49726_ (_42539_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _49727_ (_42540_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _49728_ (_42541_, _42540_, _42539_);
  and _49729_ (_42542_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _49730_ (_42543_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _49731_ (_42544_, _42543_, _42542_);
  and _49732_ (_42545_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _49733_ (_42546_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _49734_ (_42547_, _42546_, _42545_);
  and _49735_ (_42548_, _42547_, _42544_);
  and _49736_ (_42549_, _42548_, _42541_);
  nor _49737_ (_42550_, _42549_, _42514_);
  nor _49738_ (_42551_, _42550_, _42538_);
  not _49739_ (_42552_, _42551_);
  and _49740_ (_42553_, _42552_, _42537_);
  not _49741_ (_42554_, _42553_);
  and _49742_ (_42555_, _42498_, _38614_);
  and _49743_ (_42556_, _38614_, _38577_);
  and _49744_ (_42557_, _42556_, _38477_);
  and _49745_ (_42558_, _42474_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _49746_ (_42559_, _42558_, _39181_);
  and _49747_ (_42560_, _42559_, _42557_);
  nor _49748_ (_42561_, _42560_, _42555_);
  and _49749_ (_42562_, _42561_, _42554_);
  not _49750_ (_42563_, _38738_);
  and _49751_ (_42564_, _42563_, _38616_);
  and _49752_ (_42565_, _42463_, _38477_);
  and _49753_ (_42566_, _42480_, _40357_);
  and _49754_ (_42567_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _49755_ (_42568_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _49756_ (_42569_, _42568_, _42567_);
  and _49757_ (_42570_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _49758_ (_42571_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _49759_ (_42572_, _42571_, _42570_);
  and _49760_ (_42573_, _42572_, _42569_);
  nor _49761_ (_42574_, _42573_, _42480_);
  nor _49762_ (_42575_, _42574_, _42566_);
  not _49763_ (_42576_, _42575_);
  and _49764_ (_42577_, _42576_, _42565_);
  nor _49765_ (_42578_, _42577_, _42564_);
  and _49766_ (_42579_, _42578_, _42562_);
  not _49767_ (_42580_, _42579_);
  and _49768_ (_42581_, _42580_, _42536_);
  and _49769_ (_42582_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _49770_ (_42583_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _49771_ (_42584_, _42583_, _42582_);
  and _49772_ (_42585_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _49773_ (_42586_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _49774_ (_42587_, _42586_, _42585_);
  and _49775_ (_42588_, _42587_, _42584_);
  nor _49776_ (_42589_, _42588_, _42480_);
  and _49777_ (_42590_, _42480_, _41428_);
  nor _49778_ (_42591_, _42590_, _42589_);
  not _49779_ (_42592_, _42591_);
  and _49780_ (_42593_, _42592_, _42565_);
  and _49781_ (_42594_, _42463_, _42498_);
  not _49782_ (_42595_, _38720_);
  and _49783_ (_42596_, _42595_, _38616_);
  or _49784_ (_42597_, _42596_, _42594_);
  and _49785_ (_42598_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _49786_ (_42599_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _49787_ (_42600_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _49788_ (_42601_, _42600_, _42599_);
  and _49789_ (_42602_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _49790_ (_42603_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _49791_ (_42604_, _42603_, _42602_);
  and _49792_ (_42605_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _49793_ (_42606_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _49794_ (_42607_, _42606_, _42605_);
  and _49795_ (_42608_, _42607_, _42604_);
  and _49796_ (_42609_, _42608_, _42601_);
  nor _49797_ (_42610_, _42609_, _42514_);
  nor _49798_ (_42611_, _42610_, _42598_);
  not _49799_ (_42612_, _42611_);
  and _49800_ (_42613_, _42612_, _42537_);
  and _49801_ (_42614_, _42557_, _38270_);
  or _49802_ (_42615_, _42614_, _42613_);
  or _49803_ (_42616_, _42615_, _42597_);
  nor _49804_ (_42617_, _42616_, _42593_);
  nor _49805_ (_42618_, _42617_, _42535_);
  nor _49806_ (_42619_, _42618_, _42581_);
  and _49807_ (_42620_, _27496_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49808_ (_42621_, _42620_, _40742_);
  nor _49809_ (_42622_, _26860_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _49810_ (_42623_, _42622_, _42621_);
  nand _49811_ (_42624_, _42623_, _42619_);
  or _49812_ (_42625_, _42623_, _42619_);
  and _49813_ (_42626_, _42625_, _42624_);
  and _49814_ (_42627_, _42620_, _27661_);
  nor _49815_ (_42628_, _26981_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _49816_ (_42629_, _42628_, _42627_);
  not _49817_ (_42630_, _42629_);
  not _49818_ (_42631_, _42476_);
  and _49819_ (_42632_, _42557_, _42631_);
  and _49820_ (_42633_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _49821_ (_42634_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _49822_ (_42635_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _49823_ (_42636_, _42635_, _42634_);
  and _49824_ (_42637_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _49825_ (_42638_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _49826_ (_42639_, _42638_, _42637_);
  and _49827_ (_42640_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _49828_ (_42641_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _49829_ (_42642_, _42641_, _42640_);
  and _49830_ (_42643_, _42642_, _42639_);
  and _49831_ (_42644_, _42643_, _42636_);
  nor _49832_ (_42645_, _42644_, _42514_);
  nor _49833_ (_42646_, _42645_, _42633_);
  not _49834_ (_42647_, _42646_);
  and _49835_ (_42648_, _42647_, _42537_);
  nor _49836_ (_42649_, _42648_, _42632_);
  not _49837_ (_42650_, _38732_);
  and _49838_ (_42651_, _42650_, _38616_);
  and _49839_ (_42652_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _49840_ (_42653_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _49841_ (_42654_, _42653_, _42652_);
  and _49842_ (_42655_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _49843_ (_42656_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _49844_ (_42657_, _42656_, _42655_);
  and _49845_ (_42658_, _42657_, _42654_);
  nor _49846_ (_42659_, _42658_, _42480_);
  and _49847_ (_42660_, _42480_, _40346_);
  nor _49848_ (_42661_, _42660_, _42659_);
  not _49849_ (_42662_, _42661_);
  and _49850_ (_42663_, _42662_, _42565_);
  nor _49851_ (_42664_, _42663_, _42651_);
  and _49852_ (_42665_, _42664_, _42649_);
  not _49853_ (_42666_, _42665_);
  and _49854_ (_42667_, _42666_, _42536_);
  and _49855_ (_42668_, _42557_, _38006_);
  and _49856_ (_42669_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _49857_ (_42670_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _49858_ (_42671_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _49859_ (_42672_, _42671_, _42670_);
  and _49860_ (_42673_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _49861_ (_42674_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _49862_ (_42675_, _42674_, _42673_);
  and _49863_ (_42676_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _49864_ (_42677_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _49865_ (_42678_, _42677_, _42676_);
  and _49866_ (_42679_, _42678_, _42675_);
  and _49867_ (_42680_, _42679_, _42672_);
  nor _49868_ (_42681_, _42680_, _42514_);
  nor _49869_ (_42682_, _42681_, _42669_);
  not _49870_ (_42683_, _42682_);
  and _49871_ (_42684_, _42683_, _42537_);
  nor _49872_ (_42685_, _42684_, _42668_);
  not _49873_ (_42686_, _38714_);
  and _49874_ (_42687_, _42686_, _38616_);
  and _49875_ (_42688_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _49876_ (_42689_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _49877_ (_42690_, _42689_, _42688_);
  and _49878_ (_42691_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _49879_ (_42692_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _49880_ (_42693_, _42692_, _42691_);
  and _49881_ (_42694_, _42693_, _42690_);
  nor _49882_ (_42695_, _42694_, _42480_);
  and _49883_ (_42696_, _42480_, _38683_);
  nor _49884_ (_42697_, _42696_, _42695_);
  not _49885_ (_42698_, _42697_);
  and _49886_ (_42699_, _42698_, _42565_);
  nor _49887_ (_42700_, _42699_, _42687_);
  and _49888_ (_42701_, _42700_, _42685_);
  nor _49889_ (_42702_, _42701_, _42535_);
  nor _49890_ (_42703_, _42702_, _42667_);
  and _49891_ (_42704_, _42703_, _42630_);
  nor _49892_ (_42705_, _42703_, _42630_);
  nor _49893_ (_42706_, _42705_, _42704_);
  not _49894_ (_42707_, _42706_);
  nor _49895_ (_42708_, _42707_, _42626_);
  nor _49896_ (_42709_, _42666_, _42536_);
  nor _49897_ (_42710_, _42463_, _38477_);
  and _49898_ (_42711_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _49899_ (_42712_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _49900_ (_42713_, _42712_, _42711_);
  and _49901_ (_42714_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _49902_ (_42715_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _49903_ (_42716_, _42715_, _42714_);
  and _49904_ (_42717_, _42716_, _42713_);
  nor _49905_ (_42718_, _42717_, _42480_);
  and _49906_ (_42719_, _42480_, _40383_);
  nor _49907_ (_42720_, _42719_, _42718_);
  not _49908_ (_42721_, _42720_);
  and _49909_ (_42722_, _42721_, _42565_);
  nor _49910_ (_42723_, _42722_, _42710_);
  not _49911_ (_42724_, _38750_);
  and _49912_ (_42725_, _42724_, _38616_);
  and _49913_ (_42726_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _49914_ (_42727_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _49915_ (_42728_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _49916_ (_42729_, _42728_, _42727_);
  and _49917_ (_42730_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _49918_ (_42731_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _49919_ (_42732_, _42731_, _42730_);
  and _49920_ (_42733_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _49921_ (_42734_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _49922_ (_42735_, _42734_, _42733_);
  and _49923_ (_42736_, _42735_, _42732_);
  and _49924_ (_42737_, _42736_, _42729_);
  nor _49925_ (_42738_, _42737_, _42514_);
  nor _49926_ (_42739_, _42738_, _42726_);
  not _49927_ (_42740_, _42739_);
  and _49928_ (_42741_, _42740_, _42537_);
  nor _49929_ (_42742_, _42741_, _42725_);
  and _49930_ (_42743_, _42742_, _42723_);
  and _49931_ (_42744_, _42743_, _42536_);
  nor _49932_ (_42745_, _42744_, _42709_);
  nor _49933_ (_42746_, _42620_, _27661_);
  and _49934_ (_42747_, _42620_, _27211_);
  nor _49935_ (_42748_, _42747_, _42746_);
  not _49936_ (_42749_, _42748_);
  and _49937_ (_42750_, _42749_, _42745_);
  nor _49938_ (_42751_, _42749_, _42745_);
  nor _49939_ (_42752_, _42751_, _42750_);
  and _49940_ (_42753_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _49941_ (_42754_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _49942_ (_42755_, _42754_, _42753_);
  and _49943_ (_42756_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _49944_ (_42757_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _49945_ (_42758_, _42757_, _42756_);
  and _49946_ (_42759_, _42758_, _42755_);
  and _49947_ (_42760_, _42759_, _42481_);
  and _49948_ (_42761_, _42480_, _38642_);
  nor _49949_ (_42762_, _42761_, _42760_);
  and _49950_ (_42763_, _42762_, _42565_);
  and _49951_ (_42764_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and _49952_ (_42765_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _49953_ (_42766_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _49954_ (_42767_, _42766_, _42765_);
  and _49955_ (_42768_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _49956_ (_42769_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _49957_ (_42770_, _42769_, _42768_);
  and _49958_ (_42771_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _49959_ (_42772_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _49960_ (_42773_, _42772_, _42771_);
  and _49961_ (_42774_, _42773_, _42770_);
  and _49962_ (_42775_, _42774_, _42767_);
  nor _49963_ (_42776_, _42775_, _42514_);
  nor _49964_ (_42777_, _42776_, _42764_);
  not _49965_ (_42778_, _42777_);
  and _49966_ (_42779_, _42778_, _42537_);
  nor _49967_ (_42780_, _42779_, _42763_);
  nor _49968_ (_42781_, _38744_, _38614_);
  nor _49969_ (_42782_, _42781_, _42498_);
  or _49970_ (_42783_, _42556_, _38615_);
  not _49971_ (_42784_, _42783_);
  nor _49972_ (_42785_, _42784_, _42782_);
  not _49973_ (_42786_, _42785_);
  and _49974_ (_42787_, _42786_, _42780_);
  not _49975_ (_42788_, _42787_);
  and _49976_ (_42789_, _42788_, _42536_);
  and _49977_ (_42790_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _49978_ (_42791_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _49979_ (_42792_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _49980_ (_42793_, _42792_, _42791_);
  and _49981_ (_42794_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _49982_ (_42795_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _49983_ (_42796_, _42795_, _42794_);
  and _49984_ (_42797_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _49985_ (_42798_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _49986_ (_42799_, _42798_, _42797_);
  and _49987_ (_42800_, _42799_, _42796_);
  and _49988_ (_42801_, _42800_, _42793_);
  nor _49989_ (_42802_, _42801_, _42514_);
  nor _49990_ (_42803_, _42802_, _42790_);
  not _49991_ (_42804_, _42803_);
  and _49992_ (_42805_, _42804_, _42537_);
  and _49993_ (_42806_, _42489_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _49994_ (_42807_, _42484_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _49995_ (_42808_, _42807_, _42806_);
  and _49996_ (_42809_, _42487_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _49997_ (_42810_, _42482_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _49998_ (_42811_, _42810_, _42809_);
  and _49999_ (_42812_, _42811_, _42808_);
  nor _50000_ (_42813_, _42812_, _42480_);
  and _50001_ (_42814_, _42480_, _40334_);
  nor _50002_ (_42815_, _42814_, _42813_);
  not _50003_ (_42816_, _42815_);
  and _50004_ (_42817_, _42816_, _42565_);
  nor _50005_ (_42818_, _42817_, _42805_);
  not _50006_ (_42819_, _38726_);
  and _50007_ (_42820_, _42819_, _38616_);
  and _50008_ (_42821_, _42557_, _38414_);
  nor _50009_ (_42822_, _42821_, _42820_);
  and _50010_ (_42823_, _42822_, _42818_);
  nor _50011_ (_42824_, _42823_, _42535_);
  nor _50012_ (_42825_, _42824_, _42789_);
  and _50013_ (_42826_, _42620_, _39095_);
  nor _50014_ (_42827_, _26740_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _50015_ (_42828_, _42827_, _42826_);
  not _50016_ (_42829_, _42828_);
  nor _50017_ (_42830_, _42829_, _42825_);
  and _50018_ (_42831_, _42829_, _42825_);
  nor _50019_ (_42832_, _42831_, _42830_);
  and _50020_ (_42833_, _42832_, _42752_);
  and _50021_ (_42834_, _42833_, _42708_);
  and _50022_ (_42835_, _42834_, _42459_);
  nor _50023_ (_42836_, _42788_, _42536_);
  nor _50024_ (_42837_, _42620_, _39095_);
  not _50025_ (_42838_, _42837_);
  nor _50026_ (_42839_, _42838_, _42836_);
  and _50027_ (_42840_, _42838_, _42836_);
  nor _50028_ (_42841_, _42840_, _42839_);
  nor _50029_ (_42842_, _42579_, _42536_);
  nor _50030_ (_42843_, _42620_, _27825_);
  not _50031_ (_42844_, _42843_);
  nor _50032_ (_42845_, _42844_, _42842_);
  and _50033_ (_42846_, _42844_, _42842_);
  nor _50034_ (_42847_, _42846_, _42845_);
  and _50035_ (_42848_, _42847_, _42841_);
  nor _50036_ (_42849_, _42743_, _42536_);
  nor _50037_ (_42850_, _42620_, _27211_);
  not _50038_ (_42851_, _42850_);
  nor _50039_ (_42852_, _42851_, _42849_);
  and _50040_ (_42853_, _42851_, _42849_);
  nor _50041_ (_42854_, _42853_, _42852_);
  nor _50042_ (_42855_, _42521_, _27496_);
  and _50043_ (_42856_, _42521_, _27496_);
  nor _50044_ (_42857_, _42856_, _42855_);
  not _50045_ (_42858_, _42857_);
  and _50046_ (_42859_, _42858_, _42854_);
  and _50047_ (_42860_, _42859_, _42848_);
  and _50048_ (_42861_, _42860_, _42835_);
  not _50049_ (_42862_, _42825_);
  not _50050_ (_42863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _50051_ (_42864_, _42703_, _42863_);
  and _50052_ (_42865_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _50053_ (_42866_, _42865_, _42619_);
  or _50054_ (_42867_, _42866_, _42864_);
  and _50055_ (_42868_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not _50056_ (_42869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _50057_ (_42870_, _42703_, _42869_);
  nand _50058_ (_42871_, _42870_, _42619_);
  or _50059_ (_42872_, _42871_, _42868_);
  and _50060_ (_42873_, _42872_, _42867_);
  or _50061_ (_42874_, _42873_, _42862_);
  not _50062_ (_42875_, _42745_);
  not _50063_ (_42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _50064_ (_42877_, _42703_, _42876_);
  and _50065_ (_42878_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _50066_ (_42879_, _42878_, _42619_);
  or _50067_ (_42880_, _42879_, _42877_);
  and _50068_ (_42881_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not _50069_ (_42882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _50070_ (_42883_, _42703_, _42882_);
  nand _50071_ (_42884_, _42883_, _42619_);
  or _50072_ (_42885_, _42884_, _42881_);
  and _50073_ (_42886_, _42885_, _42880_);
  or _50074_ (_42887_, _42886_, _42825_);
  and _50075_ (_42888_, _42887_, _42875_);
  and _50076_ (_42889_, _42888_, _42874_);
  not _50077_ (_42890_, _42619_);
  not _50078_ (_42891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand _50079_ (_42892_, _42703_, _42891_);
  or _50080_ (_42893_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _50081_ (_42894_, _42893_, _42892_);
  or _50082_ (_42895_, _42894_, _42890_);
  or _50083_ (_42896_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not _50084_ (_42897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand _50085_ (_42898_, _42703_, _42897_);
  and _50086_ (_42899_, _42898_, _42896_);
  or _50087_ (_42900_, _42899_, _42619_);
  and _50088_ (_42901_, _42900_, _42895_);
  or _50089_ (_42902_, _42901_, _42862_);
  not _50090_ (_42903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand _50091_ (_42904_, _42703_, _42903_);
  or _50092_ (_42905_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _50093_ (_42906_, _42905_, _42904_);
  or _50094_ (_42907_, _42906_, _42890_);
  or _50095_ (_42908_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not _50096_ (_42909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand _50097_ (_42910_, _42703_, _42909_);
  and _50098_ (_42911_, _42910_, _42908_);
  or _50099_ (_42912_, _42911_, _42619_);
  and _50100_ (_42913_, _42912_, _42907_);
  or _50101_ (_42914_, _42913_, _42825_);
  and _50102_ (_42915_, _42914_, _42745_);
  and _50103_ (_42916_, _42915_, _42902_);
  or _50104_ (_42917_, _42916_, _42889_);
  or _50105_ (_42918_, _42917_, _42861_);
  not _50106_ (_42919_, _42861_);
  or _50107_ (_42920_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not _50108_ (_42921_, _42835_);
  nor _50109_ (_42922_, _42861_, _42921_);
  nor _50110_ (_42923_, _42922_, rst);
  and _50111_ (_42924_, _42923_, _42920_);
  and _50112_ (_42925_, _42924_, _42918_);
  and _50113_ (_42926_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _50114_ (_42927_, _42926_, _28659_);
  nor _50115_ (_42928_, _42927_, _31265_);
  nand _50116_ (_42929_, _28659_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50117_ (_42930_, _20043_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50118_ (_42931_, _42930_, _42929_);
  nor _50119_ (_42932_, _38704_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _50120_ (_42933_, _42932_, _42931_);
  or _50121_ (_42934_, _42933_, _42928_);
  and _50122_ (_40239_, _42934_, _43100_);
  and _50123_ (_42935_, _40239_, _42922_);
  or _50124_ (_02567_, _42935_, _42925_);
  not _50125_ (_42936_, _42459_);
  nor _50126_ (_42937_, _42629_, _42936_);
  nor _50127_ (_42938_, _42936_, _42623_);
  and _50128_ (_42939_, _42938_, _42937_);
  and _50129_ (_42940_, _42748_, _42459_);
  nor _50130_ (_42941_, _42936_, _42828_);
  and _50131_ (_42942_, _42941_, _42940_);
  and _50132_ (_42943_, _42942_, _42939_);
  and _50133_ (_42944_, _42934_, _42459_);
  and _50134_ (_42945_, _42944_, _42943_);
  not _50135_ (_42946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor _50136_ (_42947_, _42943_, _42946_);
  or _50137_ (_02578_, _42947_, _42945_);
  nor _50138_ (_42948_, _42941_, _42940_);
  nor _50139_ (_42949_, _42938_, _42937_);
  and _50140_ (_42950_, _42949_, _42459_);
  and _50141_ (_42951_, _42950_, _42948_);
  and _50142_ (_42952_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _28648_);
  and _50143_ (_42953_, _42952_, _28692_);
  nand _50144_ (_42954_, _42953_, _31265_);
  not _50145_ (_42955_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50146_ (_42956_, _38682_, _42955_);
  or _50147_ (_42957_, _18880_, _42955_);
  and _50148_ (_42958_, _42957_, _42956_);
  or _50149_ (_42959_, _42958_, _42953_);
  and _50150_ (_42960_, _42959_, _42954_);
  and _50151_ (_42961_, _42960_, _42951_);
  not _50152_ (_42962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _50153_ (_42963_, _42951_, _42962_);
  or _50154_ (_02802_, _42963_, _42961_);
  not _50155_ (_42964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _50156_ (_42965_, _42951_, _42964_);
  nand _50157_ (_42966_, _42952_, _28736_);
  nor _50158_ (_42967_, _42966_, _31265_);
  nor _50159_ (_42968_, _38672_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50160_ (_42969_, _42952_, _28757_);
  and _50161_ (_42970_, _42952_, _28659_);
  or _50162_ (_42971_, _42970_, _42926_);
  or _50163_ (_42972_, _42971_, _42969_);
  and _50164_ (_42973_, _42972_, _19874_);
  or _50165_ (_42974_, _42973_, _42968_);
  or _50166_ (_42975_, _42974_, _42967_);
  and _50167_ (_42976_, _42975_, _42951_);
  or _50168_ (_02807_, _42976_, _42965_);
  not _50169_ (_42977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _50170_ (_42978_, _42951_, _42977_);
  nand _50171_ (_42979_, _42952_, _28768_);
  nor _50172_ (_42980_, _42979_, _31265_);
  nor _50173_ (_42981_, _38665_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50174_ (_42982_, _42952_, _28725_);
  or _50175_ (_42983_, _42982_, _42971_);
  and _50176_ (_42984_, _42983_, _18518_);
  or _50177_ (_42985_, _42984_, _42981_);
  or _50178_ (_42986_, _42985_, _42980_);
  and _50179_ (_42987_, _42986_, _42951_);
  or _50180_ (_02812_, _42987_, _42978_);
  and _50181_ (_42988_, _42970_, _31885_);
  nor _50182_ (_42989_, _38658_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _50183_ (_42990_, _42969_, _42926_);
  or _50184_ (_42991_, _42990_, _42982_);
  and _50185_ (_42992_, _42991_, _19547_);
  or _50186_ (_42993_, _42992_, _42989_);
  or _50187_ (_42994_, _42993_, _42988_);
  and _50188_ (_42995_, _42994_, _42951_);
  not _50189_ (_42996_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _50190_ (_42997_, _42951_, _42996_);
  or _50191_ (_02817_, _42997_, _42995_);
  nand _50192_ (_42998_, _42926_, _28692_);
  nor _50193_ (_42999_, _42998_, _31265_);
  nor _50194_ (_43000_, _38650_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50195_ (_43001_, _28692_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50196_ (_43002_, _18716_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50197_ (_43003_, _43002_, _43001_);
  or _50198_ (_43004_, _43003_, _43000_);
  or _50199_ (_43005_, _43004_, _42999_);
  and _50200_ (_43006_, _43005_, _42951_);
  not _50201_ (_43007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _50202_ (_43008_, _42951_, _43007_);
  or _50203_ (_02822_, _43008_, _43006_);
  nand _50204_ (_43009_, _42926_, _28736_);
  nor _50205_ (_43010_, _43009_, _31265_);
  nor _50206_ (_43011_, _38642_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50207_ (_43012_, _28736_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50208_ (_43013_, _19699_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50209_ (_43014_, _43013_, _43012_);
  or _50210_ (_43015_, _43014_, _43011_);
  or _50211_ (_43016_, _43015_, _43010_);
  and _50212_ (_43017_, _43016_, _42951_);
  not _50213_ (_43018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _50214_ (_43019_, _42951_, _43018_);
  or _50215_ (_02827_, _43019_, _43017_);
  nand _50216_ (_43020_, _42926_, _28768_);
  nor _50217_ (_43021_, _43020_, _31265_);
  nor _50218_ (_43022_, _38635_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50219_ (_43023_, _28768_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50220_ (_43024_, _19056_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50221_ (_43025_, _43024_, _43023_);
  or _50222_ (_43026_, _43025_, _43022_);
  or _50223_ (_43027_, _43026_, _43021_);
  and _50224_ (_43028_, _43027_, _42951_);
  not _50225_ (_43029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _50226_ (_43030_, _42951_, _43029_);
  or _50227_ (_02832_, _43030_, _43028_);
  not _50228_ (_43031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _50229_ (_43032_, _42951_, _43031_);
  and _50230_ (_43033_, _42951_, _42934_);
  or _50231_ (_02834_, _43033_, _43032_);
  and _50232_ (_43034_, _42960_, _42459_);
  and _50233_ (_43035_, _42937_, _42623_);
  and _50234_ (_43036_, _43035_, _42948_);
  and _50235_ (_43037_, _43036_, _43034_);
  not _50236_ (_43038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _50237_ (_43039_, _43036_, _43038_);
  or _50238_ (_02842_, _43039_, _43037_);
  and _50239_ (_43040_, _42975_, _42459_);
  and _50240_ (_43041_, _43036_, _43040_);
  not _50241_ (_43042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _50242_ (_43043_, _43036_, _43042_);
  or _50243_ (_02845_, _43043_, _43041_);
  and _50244_ (_43044_, _42986_, _42459_);
  and _50245_ (_43046_, _43036_, _43044_);
  not _50246_ (_43047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _50247_ (_43049_, _43036_, _43047_);
  or _50248_ (_02848_, _43049_, _43046_);
  and _50249_ (_43051_, _42994_, _42459_);
  and _50250_ (_43053_, _43036_, _43051_);
  not _50251_ (_43055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _50252_ (_43057_, _43036_, _43055_);
  or _50253_ (_02853_, _43057_, _43053_);
  and _50254_ (_43059_, _43005_, _42459_);
  and _50255_ (_43060_, _43036_, _43059_);
  not _50256_ (_43061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _50257_ (_43062_, _43036_, _43061_);
  or _50258_ (_02856_, _43062_, _43060_);
  and _50259_ (_43063_, _43016_, _42459_);
  and _50260_ (_43064_, _43036_, _43063_);
  not _50261_ (_43065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _50262_ (_43066_, _43036_, _43065_);
  or _50263_ (_02859_, _43066_, _43064_);
  and _50264_ (_43067_, _43027_, _42459_);
  and _50265_ (_43068_, _43036_, _43067_);
  not _50266_ (_43069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _50267_ (_43070_, _43036_, _43069_);
  or _50268_ (_02862_, _43070_, _43068_);
  and _50269_ (_43071_, _43036_, _42944_);
  nor _50270_ (_43072_, _43036_, _42869_);
  or _50271_ (_02865_, _43072_, _43071_);
  and _50272_ (_43073_, _42938_, _42629_);
  and _50273_ (_43074_, _43073_, _42948_);
  and _50274_ (_43075_, _43074_, _43034_);
  not _50275_ (_43076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor _50276_ (_43077_, _43074_, _43076_);
  or _50277_ (_02871_, _43077_, _43075_);
  and _50278_ (_43078_, _43074_, _43040_);
  not _50279_ (_43079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor _50280_ (_43080_, _43074_, _43079_);
  or _50281_ (_02875_, _43080_, _43078_);
  and _50282_ (_43081_, _43074_, _43044_);
  not _50283_ (_43082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _50284_ (_43083_, _43074_, _43082_);
  or _50285_ (_02879_, _43083_, _43081_);
  and _50286_ (_43084_, _43074_, _43051_);
  not _50287_ (_43085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor _50288_ (_43086_, _43074_, _43085_);
  or _50289_ (_02882_, _43086_, _43084_);
  and _50290_ (_43088_, _43074_, _43059_);
  not _50291_ (_43090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _50292_ (_43092_, _43074_, _43090_);
  or _50293_ (_02886_, _43092_, _43088_);
  and _50294_ (_43095_, _43074_, _43063_);
  not _50295_ (_43097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _50296_ (_43099_, _43074_, _43097_);
  or _50297_ (_02889_, _43099_, _43095_);
  and _50298_ (_43101_, _43074_, _43067_);
  not _50299_ (_43103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _50300_ (_43105_, _43074_, _43103_);
  or _50301_ (_02893_, _43105_, _43101_);
  and _50302_ (_43106_, _43074_, _42944_);
  not _50303_ (_43107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _50304_ (_43108_, _43074_, _43107_);
  or _50305_ (_02895_, _43108_, _43106_);
  and _50306_ (_43109_, _42948_, _42939_);
  and _50307_ (_43110_, _43109_, _43034_);
  not _50308_ (_43111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _50309_ (_43112_, _43109_, _43111_);
  or _50310_ (_02901_, _43112_, _43110_);
  and _50311_ (_43113_, _43109_, _43040_);
  not _50312_ (_43114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _50313_ (_43115_, _43109_, _43114_);
  or _50314_ (_02904_, _43115_, _43113_);
  and _50315_ (_43116_, _43109_, _43044_);
  not _50316_ (_43117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _50317_ (_43118_, _43109_, _43117_);
  or _50318_ (_02907_, _43118_, _43116_);
  and _50319_ (_43119_, _43109_, _43051_);
  not _50320_ (_43120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _50321_ (_43121_, _43109_, _43120_);
  or _50322_ (_02910_, _43121_, _43119_);
  and _50323_ (_43122_, _43109_, _43059_);
  not _50324_ (_43123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor _50325_ (_43124_, _43109_, _43123_);
  or _50326_ (_02914_, _43124_, _43122_);
  and _50327_ (_43125_, _43109_, _43063_);
  not _50328_ (_43126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _50329_ (_43127_, _43109_, _43126_);
  or _50330_ (_02917_, _43127_, _43125_);
  and _50331_ (_43128_, _43109_, _43067_);
  not _50332_ (_43129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor _50333_ (_43130_, _43109_, _43129_);
  or _50334_ (_02922_, _43130_, _43128_);
  and _50335_ (_43131_, _43109_, _42944_);
  nor _50336_ (_43132_, _43109_, _42863_);
  or _50337_ (_02925_, _43132_, _43131_);
  and _50338_ (_43133_, _42941_, _42749_);
  and _50339_ (_43134_, _43133_, _42949_);
  and _50340_ (_43135_, _43134_, _43034_);
  not _50341_ (_43136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _50342_ (_43137_, _43134_, _43136_);
  or _50343_ (_02933_, _43137_, _43135_);
  and _50344_ (_43138_, _43134_, _43040_);
  not _50345_ (_43139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _50346_ (_43140_, _43134_, _43139_);
  or _50347_ (_02937_, _43140_, _43138_);
  and _50348_ (_43141_, _43134_, _43044_);
  not _50349_ (_43142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _50350_ (_43143_, _43134_, _43142_);
  or _50351_ (_02940_, _43143_, _43141_);
  and _50352_ (_43144_, _43134_, _43051_);
  not _50353_ (_43145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _50354_ (_43146_, _43134_, _43145_);
  or _50355_ (_02945_, _43146_, _43144_);
  and _50356_ (_43147_, _43134_, _43059_);
  not _50357_ (_43148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _50358_ (_43149_, _43134_, _43148_);
  or _50359_ (_02949_, _43149_, _43147_);
  and _50360_ (_43150_, _43134_, _43063_);
  not _50361_ (_43151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _50362_ (_43152_, _43134_, _43151_);
  or _50363_ (_02952_, _43152_, _43150_);
  and _50364_ (_43153_, _43134_, _43067_);
  not _50365_ (_43154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _50366_ (_43155_, _43134_, _43154_);
  or _50367_ (_02956_, _43155_, _43153_);
  and _50368_ (_43156_, _43134_, _42944_);
  not _50369_ (_43157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor _50370_ (_43158_, _43134_, _43157_);
  or _50371_ (_02959_, _43158_, _43156_);
  and _50372_ (_43159_, _43133_, _43035_);
  and _50373_ (_43160_, _43159_, _43034_);
  not _50374_ (_43161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _50375_ (_43162_, _43159_, _43161_);
  or _50376_ (_02963_, _43162_, _43160_);
  and _50377_ (_43163_, _43159_, _43040_);
  not _50378_ (_43164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor _50379_ (_43165_, _43159_, _43164_);
  or _50380_ (_02966_, _43165_, _43163_);
  and _50381_ (_43166_, _43159_, _43044_);
  not _50382_ (_43167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor _50383_ (_43168_, _43159_, _43167_);
  or _50384_ (_02971_, _43168_, _43166_);
  and _50385_ (_43169_, _43159_, _43051_);
  not _50386_ (_43170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _50387_ (_43171_, _43159_, _43170_);
  or _50388_ (_02974_, _43171_, _43169_);
  and _50389_ (_43172_, _43159_, _43059_);
  not _50390_ (_43173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _50391_ (_43174_, _43159_, _43173_);
  or _50392_ (_02977_, _43174_, _43172_);
  and _50393_ (_43175_, _43159_, _43063_);
  not _50394_ (_43176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor _50395_ (_43177_, _43159_, _43176_);
  or _50396_ (_02981_, _43177_, _43175_);
  and _50397_ (_43178_, _43159_, _43067_);
  not _50398_ (_43179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor _50399_ (_43180_, _43159_, _43179_);
  or _50400_ (_02985_, _43180_, _43178_);
  and _50401_ (_43181_, _43159_, _42944_);
  nor _50402_ (_43182_, _43159_, _42882_);
  or _50403_ (_02987_, _43182_, _43181_);
  and _50404_ (_43183_, _43133_, _43073_);
  and _50405_ (_43184_, _43183_, _43034_);
  not _50406_ (_43185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor _50407_ (_43186_, _43183_, _43185_);
  or _50408_ (_02992_, _43186_, _43184_);
  and _50409_ (_43187_, _43183_, _43040_);
  not _50410_ (_43188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor _50411_ (_43189_, _43183_, _43188_);
  or _50412_ (_02996_, _43189_, _43187_);
  and _50413_ (_43190_, _43183_, _43044_);
  not _50414_ (_43191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _50415_ (_43192_, _43183_, _43191_);
  or _50416_ (_03000_, _43192_, _43190_);
  and _50417_ (_43193_, _43183_, _43051_);
  not _50418_ (_43194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor _50419_ (_43195_, _43183_, _43194_);
  or _50420_ (_03003_, _43195_, _43193_);
  and _50421_ (_43196_, _43183_, _43059_);
  not _50422_ (_43197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor _50423_ (_43198_, _43183_, _43197_);
  or _50424_ (_03008_, _43198_, _43196_);
  and _50425_ (_43199_, _43183_, _43063_);
  not _50426_ (_43200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor _50427_ (_43201_, _43183_, _43200_);
  or _50428_ (_03012_, _43201_, _43199_);
  and _50429_ (_43202_, _43183_, _43067_);
  not _50430_ (_43203_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _50431_ (_43204_, _43183_, _43203_);
  or _50432_ (_03015_, _43204_, _43202_);
  and _50433_ (_43205_, _43183_, _42944_);
  not _50434_ (_43206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _50435_ (_43207_, _43183_, _43206_);
  or _50436_ (_03018_, _43207_, _43205_);
  and _50437_ (_43208_, _43133_, _42939_);
  and _50438_ (_43209_, _43208_, _43034_);
  not _50439_ (_43210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _50440_ (_43211_, _43208_, _43210_);
  or _50441_ (_03023_, _43211_, _43209_);
  and _50442_ (_43212_, _43208_, _43040_);
  not _50443_ (_43213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor _50444_ (_43214_, _43208_, _43213_);
  or _50445_ (_03027_, _43214_, _43212_);
  and _50446_ (_43215_, _43208_, _43044_);
  not _50447_ (_43216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor _50448_ (_43217_, _43208_, _43216_);
  or _50449_ (_03030_, _43217_, _43215_);
  and _50450_ (_43218_, _43208_, _43051_);
  not _50451_ (_43219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor _50452_ (_43220_, _43208_, _43219_);
  or _50453_ (_03034_, _43220_, _43218_);
  and _50454_ (_43221_, _43208_, _43059_);
  not _50455_ (_43222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor _50456_ (_43223_, _43208_, _43222_);
  or _50457_ (_03038_, _43223_, _43221_);
  and _50458_ (_43224_, _43208_, _43063_);
  not _50459_ (_43225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor _50460_ (_43226_, _43208_, _43225_);
  or _50461_ (_03041_, _43226_, _43224_);
  and _50462_ (_43227_, _43208_, _43067_);
  not _50463_ (_43228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor _50464_ (_43229_, _43208_, _43228_);
  or _50465_ (_03045_, _43229_, _43227_);
  and _50466_ (_43230_, _43208_, _42944_);
  nor _50467_ (_43231_, _43208_, _42876_);
  or _50468_ (_03047_, _43231_, _43230_);
  and _50469_ (_43232_, _42940_, _42828_);
  and _50470_ (_43233_, _43232_, _42949_);
  and _50471_ (_43234_, _43233_, _43034_);
  not _50472_ (_43235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _50473_ (_43236_, _43233_, _43235_);
  or _50474_ (_03054_, _43236_, _43234_);
  and _50475_ (_43237_, _43233_, _43040_);
  not _50476_ (_43238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _50477_ (_43239_, _43233_, _43238_);
  or _50478_ (_03058_, _43239_, _43237_);
  and _50479_ (_43240_, _43233_, _43044_);
  not _50480_ (_43241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _50481_ (_43242_, _43233_, _43241_);
  or _50482_ (_03062_, _43242_, _43240_);
  and _50483_ (_43243_, _43233_, _43051_);
  not _50484_ (_43244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _50485_ (_43245_, _43233_, _43244_);
  or _50486_ (_03065_, _43245_, _43243_);
  and _50487_ (_43246_, _43233_, _43059_);
  not _50488_ (_43247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _50489_ (_43248_, _43233_, _43247_);
  or _50490_ (_03069_, _43248_, _43246_);
  and _50491_ (_43249_, _43233_, _43063_);
  not _50492_ (_43250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _50493_ (_43251_, _43233_, _43250_);
  or _50494_ (_03072_, _43251_, _43249_);
  and _50495_ (_43252_, _43233_, _43067_);
  not _50496_ (_43253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _50497_ (_43254_, _43233_, _43253_);
  or _50498_ (_03076_, _43254_, _43252_);
  and _50499_ (_43255_, _43233_, _42944_);
  nor _50500_ (_43256_, _43233_, _42891_);
  or _50501_ (_03078_, _43256_, _43255_);
  and _50502_ (_43257_, _43232_, _43035_);
  and _50503_ (_43258_, _43257_, _43034_);
  not _50504_ (_43259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _50505_ (_43260_, _43257_, _43259_);
  or _50506_ (_03083_, _43260_, _43258_);
  and _50507_ (_43261_, _43257_, _43040_);
  not _50508_ (_43262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor _50509_ (_43263_, _43257_, _43262_);
  or _50510_ (_03086_, _43263_, _43261_);
  and _50511_ (_43264_, _43257_, _43044_);
  not _50512_ (_43265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor _50513_ (_43266_, _43257_, _43265_);
  or _50514_ (_03090_, _43266_, _43264_);
  and _50515_ (_43267_, _43257_, _43051_);
  not _50516_ (_43268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor _50517_ (_43269_, _43257_, _43268_);
  or _50518_ (_03094_, _43269_, _43267_);
  and _50519_ (_43270_, _43257_, _43059_);
  not _50520_ (_43271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _50521_ (_43272_, _43257_, _43271_);
  or _50522_ (_03097_, _43272_, _43270_);
  and _50523_ (_43273_, _43257_, _43063_);
  not _50524_ (_43274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor _50525_ (_43275_, _43257_, _43274_);
  or _50526_ (_03101_, _43275_, _43273_);
  and _50527_ (_43276_, _43257_, _43067_);
  not _50528_ (_43277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor _50529_ (_43278_, _43257_, _43277_);
  or _50530_ (_03104_, _43278_, _43276_);
  and _50531_ (_43279_, _43257_, _42944_);
  not _50532_ (_43280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor _50533_ (_43281_, _43257_, _43280_);
  or _50534_ (_03107_, _43281_, _43279_);
  and _50535_ (_43282_, _43232_, _43073_);
  and _50536_ (_43283_, _43282_, _43034_);
  not _50537_ (_43284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _50538_ (_43285_, _43282_, _43284_);
  or _50539_ (_03111_, _43285_, _43283_);
  and _50540_ (_43286_, _43282_, _43040_);
  not _50541_ (_43287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _50542_ (_43288_, _43282_, _43287_);
  or _50543_ (_03115_, _43288_, _43286_);
  and _50544_ (_43289_, _43282_, _43044_);
  not _50545_ (_43290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor _50546_ (_43291_, _43282_, _43290_);
  or _50547_ (_03119_, _43291_, _43289_);
  and _50548_ (_43292_, _43282_, _43051_);
  not _50549_ (_43293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor _50550_ (_43294_, _43282_, _43293_);
  or _50551_ (_03122_, _43294_, _43292_);
  and _50552_ (_43295_, _43282_, _43059_);
  not _50553_ (_43296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor _50554_ (_43297_, _43282_, _43296_);
  or _50555_ (_03127_, _43297_, _43295_);
  and _50556_ (_43298_, _43282_, _43063_);
  not _50557_ (_43299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor _50558_ (_43300_, _43282_, _43299_);
  or _50559_ (_03130_, _43300_, _43298_);
  and _50560_ (_43301_, _43282_, _43067_);
  not _50561_ (_43302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _50562_ (_43303_, _43282_, _43302_);
  or _50563_ (_03134_, _43303_, _43301_);
  and _50564_ (_43304_, _43282_, _42944_);
  nor _50565_ (_43305_, _43282_, _42897_);
  or _50566_ (_03137_, _43305_, _43304_);
  and _50567_ (_43306_, _43232_, _42939_);
  and _50568_ (_43307_, _43306_, _43034_);
  not _50569_ (_43308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _50570_ (_43309_, _43306_, _43308_);
  or _50571_ (_03141_, _43309_, _43307_);
  and _50572_ (_43310_, _43306_, _43040_);
  not _50573_ (_43311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _50574_ (_43312_, _43306_, _43311_);
  or _50575_ (_03145_, _43312_, _43310_);
  and _50576_ (_43313_, _43306_, _43044_);
  not _50577_ (_43314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _50578_ (_43315_, _43306_, _43314_);
  or _50579_ (_03148_, _43315_, _43313_);
  and _50580_ (_43316_, _43306_, _43051_);
  not _50581_ (_43317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor _50582_ (_43318_, _43306_, _43317_);
  or _50583_ (_03152_, _43318_, _43316_);
  and _50584_ (_43319_, _43306_, _43059_);
  not _50585_ (_43320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _50586_ (_43321_, _43306_, _43320_);
  or _50587_ (_03155_, _43321_, _43319_);
  and _50588_ (_43322_, _43306_, _43063_);
  not _50589_ (_43323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _50590_ (_43324_, _43306_, _43323_);
  or _50591_ (_03159_, _43324_, _43322_);
  and _50592_ (_43325_, _43306_, _43067_);
  not _50593_ (_43326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _50594_ (_43327_, _43306_, _43326_);
  or _50595_ (_03162_, _43327_, _43325_);
  and _50596_ (_43328_, _43306_, _42944_);
  not _50597_ (_43329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor _50598_ (_43330_, _43306_, _43329_);
  or _50599_ (_03165_, _43330_, _43328_);
  and _50600_ (_43331_, _42949_, _42942_);
  and _50601_ (_43332_, _43331_, _43034_);
  not _50602_ (_43333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _50603_ (_43334_, _43331_, _43333_);
  or _50604_ (_03170_, _43334_, _43332_);
  and _50605_ (_43335_, _43331_, _43040_);
  not _50606_ (_43336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _50607_ (_43337_, _43331_, _43336_);
  or _50608_ (_03173_, _43337_, _43335_);
  and _50609_ (_43338_, _43331_, _43044_);
  not _50610_ (_43339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor _50611_ (_43340_, _43331_, _43339_);
  or _50612_ (_03177_, _43340_, _43338_);
  and _50613_ (_43341_, _43331_, _43051_);
  not _50614_ (_43342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _50615_ (_43343_, _43331_, _43342_);
  or _50616_ (_03181_, _43343_, _43341_);
  and _50617_ (_43344_, _43331_, _43059_);
  not _50618_ (_43345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _50619_ (_43346_, _43331_, _43345_);
  or _50620_ (_03185_, _43346_, _43344_);
  and _50621_ (_43347_, _43331_, _43063_);
  not _50622_ (_43348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor _50623_ (_43349_, _43331_, _43348_);
  or _50624_ (_03189_, _43349_, _43347_);
  and _50625_ (_43350_, _43331_, _43067_);
  not _50626_ (_43351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _50627_ (_43352_, _43331_, _43351_);
  or _50628_ (_03193_, _43352_, _43350_);
  and _50629_ (_43353_, _43331_, _42944_);
  nor _50630_ (_43354_, _43331_, _42903_);
  or _50631_ (_03196_, _43354_, _43353_);
  and _50632_ (_43355_, _43035_, _42942_);
  and _50633_ (_43356_, _43355_, _43034_);
  not _50634_ (_43357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor _50635_ (_43358_, _43355_, _43357_);
  or _50636_ (_03201_, _43358_, _43356_);
  and _50637_ (_43359_, _43355_, _43040_);
  not _50638_ (_43360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor _50639_ (_43361_, _43355_, _43360_);
  or _50640_ (_03205_, _43361_, _43359_);
  and _50641_ (_43362_, _43355_, _43044_);
  not _50642_ (_43363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor _50643_ (_43364_, _43355_, _43363_);
  or _50644_ (_03209_, _43364_, _43362_);
  and _50645_ (_43365_, _43355_, _43051_);
  not _50646_ (_43366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor _50647_ (_43367_, _43355_, _43366_);
  or _50648_ (_03213_, _43367_, _43365_);
  and _50649_ (_43368_, _43355_, _43059_);
  not _50650_ (_43369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _50651_ (_43370_, _43355_, _43369_);
  or _50652_ (_03217_, _43370_, _43368_);
  and _50653_ (_43371_, _43355_, _43063_);
  not _50654_ (_43372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor _50655_ (_43373_, _43355_, _43372_);
  or _50656_ (_03221_, _43373_, _43371_);
  and _50657_ (_43374_, _43355_, _43067_);
  not _50658_ (_43375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor _50659_ (_43376_, _43355_, _43375_);
  or _50660_ (_03225_, _43376_, _43374_);
  and _50661_ (_43377_, _43355_, _42944_);
  not _50662_ (_43378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor _50663_ (_43379_, _43355_, _43378_);
  or _50664_ (_03228_, _43379_, _43377_);
  and _50665_ (_43380_, _43073_, _42942_);
  and _50666_ (_43381_, _43380_, _43034_);
  not _50667_ (_43382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor _50668_ (_43383_, _43380_, _43382_);
  or _50669_ (_03233_, _43383_, _43381_);
  and _50670_ (_43384_, _43380_, _43040_);
  not _50671_ (_43385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor _50672_ (_43386_, _43380_, _43385_);
  or _50673_ (_03237_, _43386_, _43384_);
  and _50674_ (_43387_, _43380_, _43044_);
  not _50675_ (_43388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor _50676_ (_43389_, _43380_, _43388_);
  or _50677_ (_03241_, _43389_, _43387_);
  and _50678_ (_43390_, _43380_, _43051_);
  not _50679_ (_43391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor _50680_ (_43392_, _43380_, _43391_);
  or _50681_ (_03245_, _43392_, _43390_);
  and _50682_ (_43393_, _43380_, _43059_);
  not _50683_ (_43394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _50684_ (_43395_, _43380_, _43394_);
  or _50685_ (_03249_, _43395_, _43393_);
  and _50686_ (_43396_, _43380_, _43063_);
  not _50687_ (_43397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _50688_ (_43398_, _43380_, _43397_);
  or _50689_ (_03253_, _43398_, _43396_);
  and _50690_ (_43399_, _43380_, _43067_);
  not _50691_ (_43400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor _50692_ (_43401_, _43380_, _43400_);
  or _50693_ (_03257_, _43401_, _43399_);
  and _50694_ (_43402_, _43380_, _42944_);
  nor _50695_ (_43403_, _43380_, _42909_);
  or _50696_ (_03260_, _43403_, _43402_);
  and _50697_ (_43404_, _43034_, _42943_);
  not _50698_ (_43405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor _50699_ (_43406_, _42943_, _43405_);
  or _50700_ (_03265_, _43406_, _43404_);
  and _50701_ (_43407_, _43040_, _42943_);
  not _50702_ (_43408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor _50703_ (_43409_, _42943_, _43408_);
  or _50704_ (_03269_, _43409_, _43407_);
  and _50705_ (_43410_, _43044_, _42943_);
  not _50706_ (_43411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor _50707_ (_43412_, _42943_, _43411_);
  or _50708_ (_03273_, _43412_, _43410_);
  and _50709_ (_43413_, _43051_, _42943_);
  not _50710_ (_43414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor _50711_ (_43415_, _42943_, _43414_);
  or _50712_ (_03277_, _43415_, _43413_);
  and _50713_ (_43416_, _43059_, _42943_);
  not _50714_ (_43417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor _50715_ (_43418_, _42943_, _43417_);
  or _50716_ (_03281_, _43418_, _43416_);
  and _50717_ (_43419_, _43063_, _42943_);
  not _50718_ (_43420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor _50719_ (_43421_, _42943_, _43420_);
  or _50720_ (_03285_, _43421_, _43419_);
  and _50721_ (_43422_, _43067_, _42943_);
  not _50722_ (_43423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor _50723_ (_43424_, _42943_, _43423_);
  or _50724_ (_03289_, _43424_, _43422_);
  nor _50725_ (_43425_, _42703_, _43111_);
  and _50726_ (_43426_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _50727_ (_43427_, _43426_, _42619_);
  or _50728_ (_43428_, _43427_, _43425_);
  and _50729_ (_43429_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _50730_ (_43430_, _42703_, _43038_);
  nand _50731_ (_43431_, _43430_, _42619_);
  or _50732_ (_43432_, _43431_, _43429_);
  and _50733_ (_43433_, _43432_, _43428_);
  or _50734_ (_43434_, _43433_, _42862_);
  nor _50735_ (_43435_, _42703_, _43210_);
  and _50736_ (_43436_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _50737_ (_43437_, _43436_, _42619_);
  or _50738_ (_43438_, _43437_, _43435_);
  and _50739_ (_43439_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _50740_ (_43440_, _42703_, _43161_);
  nand _50741_ (_43441_, _43440_, _42619_);
  or _50742_ (_43442_, _43441_, _43439_);
  and _50743_ (_43443_, _43442_, _43438_);
  or _50744_ (_43444_, _43443_, _42825_);
  and _50745_ (_43445_, _43444_, _42875_);
  and _50746_ (_43446_, _43445_, _43434_);
  nand _50747_ (_43447_, _42703_, _43235_);
  or _50748_ (_43448_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _50749_ (_43449_, _43448_, _43447_);
  or _50750_ (_43450_, _43449_, _42890_);
  or _50751_ (_43451_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand _50752_ (_43452_, _42703_, _43284_);
  and _50753_ (_43453_, _43452_, _43451_);
  or _50754_ (_43454_, _43453_, _42619_);
  and _50755_ (_43455_, _43454_, _43450_);
  or _50756_ (_43456_, _43455_, _42862_);
  nand _50757_ (_43457_, _42703_, _43333_);
  or _50758_ (_43458_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _50759_ (_43459_, _43458_, _43457_);
  or _50760_ (_43460_, _43459_, _42890_);
  or _50761_ (_43461_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand _50762_ (_43462_, _42703_, _43382_);
  and _50763_ (_43463_, _43462_, _43461_);
  or _50764_ (_43464_, _43463_, _42619_);
  and _50765_ (_43465_, _43464_, _43460_);
  or _50766_ (_43466_, _43465_, _42825_);
  and _50767_ (_43467_, _43466_, _42745_);
  and _50768_ (_43468_, _43467_, _43456_);
  or _50769_ (_43469_, _43468_, _43446_);
  or _50770_ (_43470_, _43469_, _42861_);
  or _50771_ (_43471_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _50772_ (_43472_, _43471_, _42923_);
  and _50773_ (_43473_, _43472_, _43470_);
  and _50774_ (_40258_, _42960_, _43100_);
  and _50775_ (_43474_, _40258_, _42922_);
  or _50776_ (_05085_, _43474_, _43473_);
  nor _50777_ (_43475_, _42703_, _43114_);
  and _50778_ (_43476_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _50779_ (_43477_, _43476_, _42619_);
  or _50780_ (_43478_, _43477_, _43475_);
  and _50781_ (_43479_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or _50782_ (_43480_, _42703_, _43042_);
  nand _50783_ (_43481_, _43480_, _42619_);
  or _50784_ (_43482_, _43481_, _43479_);
  and _50785_ (_43483_, _43482_, _43478_);
  or _50786_ (_43484_, _43483_, _42862_);
  nor _50787_ (_43485_, _42703_, _43213_);
  and _50788_ (_43486_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _50789_ (_43487_, _43486_, _42619_);
  or _50790_ (_43488_, _43487_, _43485_);
  and _50791_ (_43489_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _50792_ (_43490_, _42703_, _43164_);
  nand _50793_ (_43491_, _43490_, _42619_);
  or _50794_ (_43492_, _43491_, _43489_);
  and _50795_ (_43493_, _43492_, _43488_);
  or _50796_ (_43494_, _43493_, _42825_);
  and _50797_ (_43495_, _43494_, _42875_);
  and _50798_ (_43496_, _43495_, _43484_);
  nand _50799_ (_43497_, _42703_, _43238_);
  or _50800_ (_43498_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _50801_ (_43499_, _43498_, _43497_);
  or _50802_ (_43500_, _43499_, _42890_);
  or _50803_ (_43501_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand _50804_ (_43502_, _42703_, _43287_);
  and _50805_ (_43503_, _43502_, _43501_);
  or _50806_ (_43504_, _43503_, _42619_);
  and _50807_ (_43505_, _43504_, _43500_);
  or _50808_ (_43506_, _43505_, _42862_);
  nand _50809_ (_43507_, _42703_, _43336_);
  or _50810_ (_43508_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _50811_ (_43509_, _43508_, _43507_);
  or _50812_ (_43510_, _43509_, _42890_);
  or _50813_ (_43511_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand _50814_ (_43512_, _42703_, _43385_);
  and _50815_ (_43513_, _43512_, _43511_);
  or _50816_ (_43514_, _43513_, _42619_);
  and _50817_ (_43515_, _43514_, _43510_);
  or _50818_ (_43516_, _43515_, _42825_);
  and _50819_ (_43517_, _43516_, _42745_);
  and _50820_ (_43518_, _43517_, _43506_);
  or _50821_ (_43519_, _43518_, _43496_);
  or _50822_ (_43520_, _43519_, _42861_);
  or _50823_ (_43521_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _50824_ (_43522_, _43521_, _42923_);
  and _50825_ (_43523_, _43522_, _43520_);
  and _50826_ (_40259_, _42975_, _43100_);
  and _50827_ (_43524_, _40259_, _42922_);
  or _50828_ (_05087_, _43524_, _43523_);
  nor _50829_ (_43525_, _42703_, _43117_);
  and _50830_ (_43526_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _50831_ (_43527_, _43526_, _42619_);
  or _50832_ (_43528_, _43527_, _43525_);
  and _50833_ (_43529_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or _50834_ (_43530_, _42703_, _43047_);
  nand _50835_ (_43531_, _43530_, _42619_);
  or _50836_ (_43532_, _43531_, _43529_);
  and _50837_ (_43533_, _43532_, _43528_);
  or _50838_ (_43534_, _43533_, _42862_);
  nor _50839_ (_43535_, _42703_, _43216_);
  and _50840_ (_43536_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _50841_ (_43537_, _43536_, _42619_);
  or _50842_ (_43538_, _43537_, _43535_);
  and _50843_ (_43539_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _50844_ (_43540_, _42703_, _43167_);
  nand _50845_ (_43541_, _43540_, _42619_);
  or _50846_ (_43542_, _43541_, _43539_);
  and _50847_ (_43543_, _43542_, _43538_);
  or _50848_ (_43544_, _43543_, _42825_);
  and _50849_ (_43545_, _43544_, _42875_);
  and _50850_ (_43546_, _43545_, _43534_);
  nand _50851_ (_43547_, _42703_, _43241_);
  or _50852_ (_43548_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _50853_ (_43549_, _43548_, _43547_);
  or _50854_ (_43550_, _43549_, _42890_);
  or _50855_ (_43551_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand _50856_ (_43552_, _42703_, _43290_);
  and _50857_ (_43553_, _43552_, _43551_);
  or _50858_ (_43554_, _43553_, _42619_);
  and _50859_ (_43555_, _43554_, _43550_);
  or _50860_ (_43556_, _43555_, _42862_);
  nand _50861_ (_43557_, _42703_, _43339_);
  or _50862_ (_43558_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _50863_ (_43559_, _43558_, _43557_);
  or _50864_ (_43560_, _43559_, _42890_);
  or _50865_ (_43561_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand _50866_ (_43562_, _42703_, _43388_);
  and _50867_ (_43563_, _43562_, _43561_);
  or _50868_ (_43564_, _43563_, _42619_);
  and _50869_ (_43565_, _43564_, _43560_);
  or _50870_ (_43566_, _43565_, _42825_);
  and _50871_ (_43567_, _43566_, _42745_);
  and _50872_ (_43568_, _43567_, _43556_);
  or _50873_ (_43569_, _43568_, _43546_);
  or _50874_ (_43570_, _43569_, _42861_);
  or _50875_ (_43571_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _50876_ (_43572_, _43571_, _42923_);
  and _50877_ (_43573_, _43572_, _43570_);
  and _50878_ (_40260_, _42986_, _43100_);
  and _50879_ (_43574_, _40260_, _42922_);
  or _50880_ (_05089_, _43574_, _43573_);
  nor _50881_ (_43575_, _42703_, _43120_);
  and _50882_ (_43576_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _50883_ (_43577_, _43576_, _42619_);
  or _50884_ (_43578_, _43577_, _43575_);
  and _50885_ (_43579_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or _50886_ (_43580_, _42703_, _43055_);
  nand _50887_ (_43581_, _43580_, _42619_);
  or _50888_ (_43582_, _43581_, _43579_);
  and _50889_ (_43583_, _43582_, _43578_);
  or _50890_ (_43584_, _43583_, _42862_);
  nor _50891_ (_43585_, _42703_, _43219_);
  and _50892_ (_43586_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _50893_ (_43587_, _43586_, _42619_);
  or _50894_ (_43588_, _43587_, _43585_);
  and _50895_ (_43589_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _50896_ (_43590_, _42703_, _43170_);
  nand _50897_ (_43591_, _43590_, _42619_);
  or _50898_ (_43592_, _43591_, _43589_);
  and _50899_ (_43593_, _43592_, _43588_);
  or _50900_ (_43597_, _43593_, _42825_);
  and _50901_ (_43602_, _43597_, _42875_);
  and _50902_ (_43610_, _43602_, _43584_);
  nand _50903_ (_43616_, _42703_, _43244_);
  or _50904_ (_43620_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _50905_ (_43627_, _43620_, _43616_);
  or _50906_ (_43635_, _43627_, _42890_);
  or _50907_ (_43639_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand _50908_ (_43644_, _42703_, _43293_);
  and _50909_ (_43652_, _43644_, _43639_);
  or _50910_ (_43658_, _43652_, _42619_);
  and _50911_ (_43662_, _43658_, _43635_);
  or _50912_ (_43669_, _43662_, _42862_);
  nand _50913_ (_43677_, _42703_, _43342_);
  or _50914_ (_43681_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _50915_ (_43686_, _43681_, _43677_);
  or _50916_ (_43688_, _43686_, _42890_);
  or _50917_ (_43699_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand _50918_ (_43704_, _42703_, _43391_);
  and _50919_ (_43712_, _43704_, _43699_);
  or _50920_ (_43718_, _43712_, _42619_);
  and _50921_ (_43722_, _43718_, _43688_);
  or _50922_ (_43729_, _43722_, _42825_);
  and _50923_ (_43737_, _43729_, _42745_);
  and _50924_ (_43741_, _43737_, _43669_);
  or _50925_ (_43746_, _43741_, _43610_);
  or _50926_ (_43754_, _43746_, _42861_);
  or _50927_ (_43760_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and _50928_ (_43764_, _43760_, _42923_);
  and _50929_ (_43771_, _43764_, _43754_);
  and _50930_ (_40261_, _42994_, _43100_);
  and _50931_ (_43782_, _40261_, _42922_);
  or _50932_ (_05091_, _43782_, _43771_);
  and _50933_ (_43787_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _50934_ (_43788_, _42703_, _43061_);
  nand _50935_ (_43789_, _43788_, _42619_);
  or _50936_ (_43790_, _43789_, _43787_);
  nor _50937_ (_43791_, _42703_, _43123_);
  and _50938_ (_43792_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _50939_ (_43793_, _43792_, _42619_);
  or _50940_ (_43794_, _43793_, _43791_);
  and _50941_ (_43795_, _43794_, _43790_);
  or _50942_ (_43796_, _43795_, _42862_);
  nor _50943_ (_43797_, _42703_, _43222_);
  and _50944_ (_43798_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _50945_ (_43799_, _43798_, _42619_);
  or _50946_ (_43800_, _43799_, _43797_);
  and _50947_ (_43801_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _50948_ (_43802_, _42703_, _43173_);
  nand _50949_ (_43803_, _43802_, _42619_);
  or _50950_ (_43804_, _43803_, _43801_);
  and _50951_ (_43805_, _43804_, _43800_);
  or _50952_ (_43806_, _43805_, _42825_);
  and _50953_ (_43807_, _43806_, _42875_);
  and _50954_ (_43808_, _43807_, _43796_);
  nor _50955_ (_43809_, _42703_, _43320_);
  and _50956_ (_43810_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _50957_ (_43811_, _43810_, _42619_);
  or _50958_ (_43812_, _43811_, _43809_);
  and _50959_ (_43813_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _50960_ (_43814_, _42703_, _43271_);
  nand _50961_ (_43815_, _43814_, _42619_);
  or _50962_ (_43816_, _43815_, _43813_);
  and _50963_ (_43817_, _43816_, _43812_);
  or _50964_ (_43818_, _43817_, _42862_);
  nor _50965_ (_43819_, _42703_, _43417_);
  and _50966_ (_43820_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _50967_ (_43821_, _43820_, _42619_);
  or _50968_ (_43822_, _43821_, _43819_);
  and _50969_ (_43823_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or _50970_ (_43824_, _42703_, _43369_);
  nand _50971_ (_43825_, _43824_, _42619_);
  or _50972_ (_43826_, _43825_, _43823_);
  and _50973_ (_43827_, _43826_, _43822_);
  or _50974_ (_43828_, _43827_, _42825_);
  and _50975_ (_43829_, _43828_, _42745_);
  and _50976_ (_43830_, _43829_, _43818_);
  or _50977_ (_43831_, _43830_, _43808_);
  and _50978_ (_43832_, _43831_, _42921_);
  and _50979_ (_43833_, _43005_, _42922_);
  and _50980_ (_43834_, _42861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or _50981_ (_43835_, _43834_, _43833_);
  or _50982_ (_43836_, _43835_, _43832_);
  and _50983_ (_05093_, _43836_, _43100_);
  or _50984_ (_43837_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand _50985_ (_43838_, _42703_, _43397_);
  and _50986_ (_43839_, _43838_, _43837_);
  or _50987_ (_43840_, _43839_, _42619_);
  nand _50988_ (_43841_, _42703_, _43348_);
  or _50989_ (_43842_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _50990_ (_43843_, _43842_, _43841_);
  or _50991_ (_43844_, _43843_, _42890_);
  and _50992_ (_43845_, _43844_, _42745_);
  and _50993_ (_43846_, _43845_, _43840_);
  and _50994_ (_43847_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _50995_ (_43848_, _42703_, _43176_);
  nand _50996_ (_43849_, _43848_, _42619_);
  or _50997_ (_43850_, _43849_, _43847_);
  nor _50998_ (_43851_, _42703_, _43225_);
  and _50999_ (_43852_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _51000_ (_43853_, _43852_, _42619_);
  or _51001_ (_43854_, _43853_, _43851_);
  and _51002_ (_43855_, _43854_, _42875_);
  and _51003_ (_43856_, _43855_, _43850_);
  or _51004_ (_43857_, _43856_, _43846_);
  and _51005_ (_43858_, _43857_, _42862_);
  or _51006_ (_43859_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand _51007_ (_43860_, _42703_, _43299_);
  and _51008_ (_43861_, _43860_, _43859_);
  or _51009_ (_43862_, _43861_, _42619_);
  nand _51010_ (_43863_, _42703_, _43250_);
  or _51011_ (_43864_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _51012_ (_43865_, _43864_, _43863_);
  or _51013_ (_43866_, _43865_, _42890_);
  and _51014_ (_43867_, _43866_, _42745_);
  and _51015_ (_43868_, _43867_, _43862_);
  and _51016_ (_43869_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _51017_ (_43870_, _42703_, _43065_);
  nand _51018_ (_43871_, _43870_, _42619_);
  or _51019_ (_43872_, _43871_, _43869_);
  nor _51020_ (_43873_, _42703_, _43126_);
  and _51021_ (_43874_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _51022_ (_43875_, _43874_, _42619_);
  or _51023_ (_43876_, _43875_, _43873_);
  and _51024_ (_43877_, _43876_, _42875_);
  and _51025_ (_43878_, _43877_, _43872_);
  or _51026_ (_43879_, _43878_, _43868_);
  and _51027_ (_43880_, _43879_, _42825_);
  or _51028_ (_43881_, _43880_, _42835_);
  or _51029_ (_43882_, _43881_, _43858_);
  or _51030_ (_43883_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _51031_ (_40263_, _43016_, _43100_);
  or _51032_ (_43884_, _40263_, _42923_);
  and _51033_ (_43885_, _43884_, _43883_);
  and _51034_ (_05095_, _43885_, _43882_);
  nor _51035_ (_43886_, _42703_, _43129_);
  and _51036_ (_43887_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _51037_ (_43888_, _43887_, _42619_);
  or _51038_ (_43889_, _43888_, _43886_);
  and _51039_ (_43890_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _51040_ (_43891_, _42703_, _43069_);
  nand _51041_ (_43892_, _43891_, _42619_);
  or _51042_ (_43893_, _43892_, _43890_);
  and _51043_ (_43894_, _43893_, _43889_);
  or _51044_ (_43895_, _43894_, _42862_);
  nor _51045_ (_43896_, _42703_, _43228_);
  and _51046_ (_43897_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _51047_ (_43898_, _43897_, _42619_);
  or _51048_ (_43899_, _43898_, _43896_);
  and _51049_ (_43900_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _51050_ (_43901_, _42703_, _43179_);
  nand _51051_ (_43902_, _43901_, _42619_);
  or _51052_ (_43903_, _43902_, _43900_);
  and _51053_ (_43904_, _43903_, _43899_);
  or _51054_ (_43905_, _43904_, _42825_);
  and _51055_ (_43906_, _43905_, _42875_);
  and _51056_ (_43907_, _43906_, _43895_);
  nand _51057_ (_43908_, _42703_, _43253_);
  or _51058_ (_43909_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _51059_ (_43910_, _43909_, _43908_);
  or _51060_ (_43911_, _43910_, _42890_);
  or _51061_ (_43912_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand _51062_ (_43913_, _42703_, _43302_);
  and _51063_ (_43914_, _43913_, _43912_);
  or _51064_ (_43915_, _43914_, _42619_);
  and _51065_ (_43916_, _43915_, _43911_);
  or _51066_ (_43917_, _43916_, _42862_);
  nand _51067_ (_43918_, _42703_, _43351_);
  or _51068_ (_43919_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _51069_ (_43920_, _43919_, _43918_);
  or _51070_ (_43921_, _43920_, _42890_);
  or _51071_ (_43922_, _42703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand _51072_ (_43923_, _42703_, _43400_);
  and _51073_ (_43924_, _43923_, _43922_);
  or _51074_ (_43925_, _43924_, _42619_);
  and _51075_ (_43926_, _43925_, _43921_);
  or _51076_ (_43927_, _43926_, _42825_);
  and _51077_ (_43928_, _43927_, _42745_);
  and _51078_ (_43929_, _43928_, _43917_);
  or _51079_ (_43930_, _43929_, _43907_);
  or _51080_ (_43931_, _43930_, _42861_);
  or _51081_ (_43932_, _42919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _51082_ (_43933_, _43932_, _42923_);
  and _51083_ (_43934_, _43933_, _43931_);
  and _51084_ (_40264_, _43027_, _43100_);
  and _51085_ (_43935_, _40264_, _42922_);
  or _51086_ (_05097_, _43935_, _43934_);
  or _51087_ (_43936_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not _51088_ (_43937_, \oc8051_gm_cxrom_1.cell0.valid );
  or _51089_ (_43938_, _43937_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand _51090_ (_43939_, _43938_, _43936_);
  nand _51091_ (_43940_, _43939_, _43100_);
  or _51092_ (_43941_, \oc8051_gm_cxrom_1.cell0.data [7], _43100_);
  and _51093_ (_05105_, _43941_, _43940_);
  or _51094_ (_43942_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or _51095_ (_43943_, \oc8051_gm_cxrom_1.cell0.data [0], _43937_);
  nand _51096_ (_43944_, _43943_, _43942_);
  nand _51097_ (_43945_, _43944_, _43100_);
  or _51098_ (_43946_, \oc8051_gm_cxrom_1.cell0.data [0], _43100_);
  and _51099_ (_05111_, _43946_, _43945_);
  or _51100_ (_43947_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or _51101_ (_43948_, \oc8051_gm_cxrom_1.cell0.data [1], _43937_);
  nand _51102_ (_43949_, _43948_, _43947_);
  nand _51103_ (_43950_, _43949_, _43100_);
  or _51104_ (_43951_, \oc8051_gm_cxrom_1.cell0.data [1], _43100_);
  and _51105_ (_05115_, _43951_, _43950_);
  or _51106_ (_43952_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or _51107_ (_43953_, \oc8051_gm_cxrom_1.cell0.data [2], _43937_);
  nand _51108_ (_43954_, _43953_, _43952_);
  nand _51109_ (_43955_, _43954_, _43100_);
  or _51110_ (_43956_, \oc8051_gm_cxrom_1.cell0.data [2], _43100_);
  and _51111_ (_05119_, _43956_, _43955_);
  or _51112_ (_43957_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or _51113_ (_43958_, \oc8051_gm_cxrom_1.cell0.data [3], _43937_);
  nand _51114_ (_43959_, _43958_, _43957_);
  nand _51115_ (_43960_, _43959_, _43100_);
  or _51116_ (_43961_, \oc8051_gm_cxrom_1.cell0.data [3], _43100_);
  and _51117_ (_05123_, _43961_, _43960_);
  or _51118_ (_43962_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or _51119_ (_43963_, \oc8051_gm_cxrom_1.cell0.data [4], _43937_);
  nand _51120_ (_43964_, _43963_, _43962_);
  nand _51121_ (_43965_, _43964_, _43100_);
  or _51122_ (_43966_, \oc8051_gm_cxrom_1.cell0.data [4], _43100_);
  and _51123_ (_05127_, _43966_, _43965_);
  or _51124_ (_43967_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or _51125_ (_43968_, \oc8051_gm_cxrom_1.cell0.data [5], _43937_);
  nand _51126_ (_43969_, _43968_, _43967_);
  nand _51127_ (_43970_, _43969_, _43100_);
  or _51128_ (_43971_, \oc8051_gm_cxrom_1.cell0.data [5], _43100_);
  and _51129_ (_05131_, _43971_, _43970_);
  or _51130_ (_43972_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or _51131_ (_43973_, \oc8051_gm_cxrom_1.cell0.data [6], _43937_);
  nand _51132_ (_43974_, _43973_, _43972_);
  nand _51133_ (_43975_, _43974_, _43100_);
  or _51134_ (_43976_, \oc8051_gm_cxrom_1.cell0.data [6], _43100_);
  and _51135_ (_05135_, _43976_, _43975_);
  or _51136_ (_43977_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not _51137_ (_43978_, \oc8051_gm_cxrom_1.cell1.valid );
  or _51138_ (_43979_, _43978_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand _51139_ (_43980_, _43979_, _43977_);
  nand _51140_ (_43981_, _43980_, _43100_);
  or _51141_ (_43982_, \oc8051_gm_cxrom_1.cell1.data [7], _43100_);
  and _51142_ (_05156_, _43982_, _43981_);
  or _51143_ (_43983_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or _51144_ (_43984_, \oc8051_gm_cxrom_1.cell1.data [0], _43978_);
  nand _51145_ (_43985_, _43984_, _43983_);
  nand _51146_ (_43986_, _43985_, _43100_);
  or _51147_ (_43987_, \oc8051_gm_cxrom_1.cell1.data [0], _43100_);
  and _51148_ (_05163_, _43987_, _43986_);
  or _51149_ (_43988_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or _51150_ (_43989_, \oc8051_gm_cxrom_1.cell1.data [1], _43978_);
  nand _51151_ (_43990_, _43989_, _43988_);
  nand _51152_ (_43991_, _43990_, _43100_);
  or _51153_ (_43992_, \oc8051_gm_cxrom_1.cell1.data [1], _43100_);
  and _51154_ (_05167_, _43992_, _43991_);
  or _51155_ (_43993_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or _51156_ (_43994_, \oc8051_gm_cxrom_1.cell1.data [2], _43978_);
  nand _51157_ (_43995_, _43994_, _43993_);
  nand _51158_ (_43996_, _43995_, _43100_);
  or _51159_ (_43997_, \oc8051_gm_cxrom_1.cell1.data [2], _43100_);
  and _51160_ (_05171_, _43997_, _43996_);
  or _51161_ (_43998_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or _51162_ (_43999_, \oc8051_gm_cxrom_1.cell1.data [3], _43978_);
  nand _51163_ (_44000_, _43999_, _43998_);
  nand _51164_ (_44001_, _44000_, _43100_);
  or _51165_ (_44002_, \oc8051_gm_cxrom_1.cell1.data [3], _43100_);
  and _51166_ (_05175_, _44002_, _44001_);
  or _51167_ (_44003_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or _51168_ (_44004_, \oc8051_gm_cxrom_1.cell1.data [4], _43978_);
  nand _51169_ (_44005_, _44004_, _44003_);
  nand _51170_ (_44006_, _44005_, _43100_);
  or _51171_ (_44007_, \oc8051_gm_cxrom_1.cell1.data [4], _43100_);
  and _51172_ (_05179_, _44007_, _44006_);
  or _51173_ (_44008_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or _51174_ (_44009_, \oc8051_gm_cxrom_1.cell1.data [5], _43978_);
  nand _51175_ (_44010_, _44009_, _44008_);
  nand _51176_ (_44011_, _44010_, _43100_);
  or _51177_ (_44012_, \oc8051_gm_cxrom_1.cell1.data [5], _43100_);
  and _51178_ (_05183_, _44012_, _44011_);
  or _51179_ (_44013_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or _51180_ (_44014_, \oc8051_gm_cxrom_1.cell1.data [6], _43978_);
  nand _51181_ (_44015_, _44014_, _44013_);
  nand _51182_ (_44016_, _44015_, _43100_);
  or _51183_ (_44017_, \oc8051_gm_cxrom_1.cell1.data [6], _43100_);
  and _51184_ (_05186_, _44017_, _44016_);
  or _51185_ (_44018_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not _51186_ (_44019_, \oc8051_gm_cxrom_1.cell2.valid );
  or _51187_ (_44020_, _44019_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand _51188_ (_44021_, _44020_, _44018_);
  nand _51189_ (_44022_, _44021_, _43100_);
  or _51190_ (_44023_, \oc8051_gm_cxrom_1.cell2.data [7], _43100_);
  and _51191_ (_05208_, _44023_, _44022_);
  or _51192_ (_44024_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or _51193_ (_44025_, \oc8051_gm_cxrom_1.cell2.data [0], _44019_);
  nand _51194_ (_44026_, _44025_, _44024_);
  nand _51195_ (_44027_, _44026_, _43100_);
  or _51196_ (_44028_, \oc8051_gm_cxrom_1.cell2.data [0], _43100_);
  and _51197_ (_05215_, _44028_, _44027_);
  or _51198_ (_00002_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or _51199_ (_00003_, \oc8051_gm_cxrom_1.cell2.data [1], _44019_);
  nand _51200_ (_00004_, _00003_, _00002_);
  nand _51201_ (_00005_, _00004_, _43100_);
  or _51202_ (_00006_, \oc8051_gm_cxrom_1.cell2.data [1], _43100_);
  and _51203_ (_05219_, _00006_, _00005_);
  or _51204_ (_00007_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or _51205_ (_00008_, \oc8051_gm_cxrom_1.cell2.data [2], _44019_);
  nand _51206_ (_00009_, _00008_, _00007_);
  nand _51207_ (_00010_, _00009_, _43100_);
  or _51208_ (_00011_, \oc8051_gm_cxrom_1.cell2.data [2], _43100_);
  and _51209_ (_05222_, _00011_, _00010_);
  or _51210_ (_00012_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or _51211_ (_00013_, \oc8051_gm_cxrom_1.cell2.data [3], _44019_);
  nand _51212_ (_00014_, _00013_, _00012_);
  nand _51213_ (_00015_, _00014_, _43100_);
  or _51214_ (_00016_, \oc8051_gm_cxrom_1.cell2.data [3], _43100_);
  and _51215_ (_05226_, _00016_, _00015_);
  or _51216_ (_00017_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or _51217_ (_00018_, \oc8051_gm_cxrom_1.cell2.data [4], _44019_);
  nand _51218_ (_00019_, _00018_, _00017_);
  nand _51219_ (_00020_, _00019_, _43100_);
  or _51220_ (_00021_, \oc8051_gm_cxrom_1.cell2.data [4], _43100_);
  and _51221_ (_05230_, _00021_, _00020_);
  or _51222_ (_00022_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or _51223_ (_00023_, \oc8051_gm_cxrom_1.cell2.data [5], _44019_);
  nand _51224_ (_00024_, _00023_, _00022_);
  nand _51225_ (_00025_, _00024_, _43100_);
  or _51226_ (_00026_, \oc8051_gm_cxrom_1.cell2.data [5], _43100_);
  and _51227_ (_05234_, _00026_, _00025_);
  or _51228_ (_00027_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or _51229_ (_00028_, \oc8051_gm_cxrom_1.cell2.data [6], _44019_);
  nand _51230_ (_00029_, _00028_, _00027_);
  nand _51231_ (_00030_, _00029_, _43100_);
  or _51232_ (_00031_, \oc8051_gm_cxrom_1.cell2.data [6], _43100_);
  and _51233_ (_05238_, _00031_, _00030_);
  or _51234_ (_00032_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not _51235_ (_00033_, \oc8051_gm_cxrom_1.cell3.valid );
  or _51236_ (_00034_, _00033_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand _51237_ (_00035_, _00034_, _00032_);
  nand _51238_ (_00036_, _00035_, _43100_);
  or _51239_ (_00037_, \oc8051_gm_cxrom_1.cell3.data [7], _43100_);
  and _51240_ (_05259_, _00037_, _00036_);
  or _51241_ (_00038_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or _51242_ (_00039_, \oc8051_gm_cxrom_1.cell3.data [0], _00033_);
  nand _51243_ (_00040_, _00039_, _00038_);
  nand _51244_ (_00041_, _00040_, _43100_);
  or _51245_ (_00042_, \oc8051_gm_cxrom_1.cell3.data [0], _43100_);
  and _51246_ (_05266_, _00042_, _00041_);
  or _51247_ (_00043_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or _51248_ (_00044_, \oc8051_gm_cxrom_1.cell3.data [1], _00033_);
  nand _51249_ (_00045_, _00044_, _00043_);
  nand _51250_ (_00046_, _00045_, _43100_);
  or _51251_ (_00047_, \oc8051_gm_cxrom_1.cell3.data [1], _43100_);
  and _51252_ (_05270_, _00047_, _00046_);
  or _51253_ (_00048_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or _51254_ (_00049_, \oc8051_gm_cxrom_1.cell3.data [2], _00033_);
  nand _51255_ (_00050_, _00049_, _00048_);
  nand _51256_ (_00051_, _00050_, _43100_);
  or _51257_ (_00052_, \oc8051_gm_cxrom_1.cell3.data [2], _43100_);
  and _51258_ (_05274_, _00052_, _00051_);
  or _51259_ (_00053_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or _51260_ (_00054_, \oc8051_gm_cxrom_1.cell3.data [3], _00033_);
  nand _51261_ (_00055_, _00054_, _00053_);
  nand _51262_ (_00056_, _00055_, _43100_);
  or _51263_ (_00057_, \oc8051_gm_cxrom_1.cell3.data [3], _43100_);
  and _51264_ (_05278_, _00057_, _00056_);
  or _51265_ (_00058_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or _51266_ (_00059_, \oc8051_gm_cxrom_1.cell3.data [4], _00033_);
  nand _51267_ (_00060_, _00059_, _00058_);
  nand _51268_ (_00061_, _00060_, _43100_);
  or _51269_ (_00062_, \oc8051_gm_cxrom_1.cell3.data [4], _43100_);
  and _51270_ (_05282_, _00062_, _00061_);
  or _51271_ (_00063_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or _51272_ (_00064_, \oc8051_gm_cxrom_1.cell3.data [5], _00033_);
  nand _51273_ (_00065_, _00064_, _00063_);
  nand _51274_ (_00066_, _00065_, _43100_);
  or _51275_ (_00067_, \oc8051_gm_cxrom_1.cell3.data [5], _43100_);
  and _51276_ (_05286_, _00067_, _00066_);
  or _51277_ (_00068_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or _51278_ (_00069_, \oc8051_gm_cxrom_1.cell3.data [6], _00033_);
  nand _51279_ (_00070_, _00069_, _00068_);
  nand _51280_ (_00071_, _00070_, _43100_);
  or _51281_ (_00072_, \oc8051_gm_cxrom_1.cell3.data [6], _43100_);
  and _51282_ (_05290_, _00072_, _00071_);
  or _51283_ (_00073_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not _51284_ (_00074_, \oc8051_gm_cxrom_1.cell4.valid );
  or _51285_ (_00075_, _00074_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand _51286_ (_00076_, _00075_, _00073_);
  nand _51287_ (_00077_, _00076_, _43100_);
  or _51288_ (_00078_, \oc8051_gm_cxrom_1.cell4.data [7], _43100_);
  and _51289_ (_05311_, _00078_, _00077_);
  or _51290_ (_00079_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or _51291_ (_00080_, \oc8051_gm_cxrom_1.cell4.data [0], _00074_);
  nand _51292_ (_00081_, _00080_, _00079_);
  nand _51293_ (_00082_, _00081_, _43100_);
  or _51294_ (_00083_, \oc8051_gm_cxrom_1.cell4.data [0], _43100_);
  and _51295_ (_05318_, _00083_, _00082_);
  or _51296_ (_00084_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or _51297_ (_00085_, \oc8051_gm_cxrom_1.cell4.data [1], _00074_);
  nand _51298_ (_00086_, _00085_, _00084_);
  nand _51299_ (_00087_, _00086_, _43100_);
  or _51300_ (_00088_, \oc8051_gm_cxrom_1.cell4.data [1], _43100_);
  and _51301_ (_05322_, _00088_, _00087_);
  or _51302_ (_00089_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or _51303_ (_00090_, \oc8051_gm_cxrom_1.cell4.data [2], _00074_);
  nand _51304_ (_00091_, _00090_, _00089_);
  nand _51305_ (_00092_, _00091_, _43100_);
  or _51306_ (_00093_, \oc8051_gm_cxrom_1.cell4.data [2], _43100_);
  and _51307_ (_05326_, _00093_, _00092_);
  or _51308_ (_00094_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or _51309_ (_00095_, \oc8051_gm_cxrom_1.cell4.data [3], _00074_);
  nand _51310_ (_00096_, _00095_, _00094_);
  nand _51311_ (_00097_, _00096_, _43100_);
  or _51312_ (_00098_, \oc8051_gm_cxrom_1.cell4.data [3], _43100_);
  and _51313_ (_05329_, _00098_, _00097_);
  or _51314_ (_00099_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or _51315_ (_00100_, \oc8051_gm_cxrom_1.cell4.data [4], _00074_);
  nand _51316_ (_00101_, _00100_, _00099_);
  nand _51317_ (_00102_, _00101_, _43100_);
  or _51318_ (_00103_, \oc8051_gm_cxrom_1.cell4.data [4], _43100_);
  and _51319_ (_05333_, _00103_, _00102_);
  or _51320_ (_00104_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or _51321_ (_00105_, \oc8051_gm_cxrom_1.cell4.data [5], _00074_);
  nand _51322_ (_00106_, _00105_, _00104_);
  nand _51323_ (_00107_, _00106_, _43100_);
  or _51324_ (_00108_, \oc8051_gm_cxrom_1.cell4.data [5], _43100_);
  and _51325_ (_05337_, _00108_, _00107_);
  or _51326_ (_00109_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or _51327_ (_00110_, \oc8051_gm_cxrom_1.cell4.data [6], _00074_);
  nand _51328_ (_00111_, _00110_, _00109_);
  nand _51329_ (_00112_, _00111_, _43100_);
  or _51330_ (_00113_, \oc8051_gm_cxrom_1.cell4.data [6], _43100_);
  and _51331_ (_05341_, _00113_, _00112_);
  or _51332_ (_00114_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not _51333_ (_00115_, \oc8051_gm_cxrom_1.cell5.valid );
  or _51334_ (_00116_, _00115_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand _51335_ (_00117_, _00116_, _00114_);
  nand _51336_ (_00118_, _00117_, _43100_);
  or _51337_ (_00119_, \oc8051_gm_cxrom_1.cell5.data [7], _43100_);
  and _51338_ (_05363_, _00119_, _00118_);
  or _51339_ (_00120_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or _51340_ (_00121_, \oc8051_gm_cxrom_1.cell5.data [0], _00115_);
  nand _51341_ (_00122_, _00121_, _00120_);
  nand _51342_ (_00123_, _00122_, _43100_);
  or _51343_ (_00124_, \oc8051_gm_cxrom_1.cell5.data [0], _43100_);
  and _51344_ (_05369_, _00124_, _00123_);
  or _51345_ (_00125_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or _51346_ (_00126_, \oc8051_gm_cxrom_1.cell5.data [1], _00115_);
  nand _51347_ (_00127_, _00126_, _00125_);
  nand _51348_ (_00128_, _00127_, _43100_);
  or _51349_ (_00129_, \oc8051_gm_cxrom_1.cell5.data [1], _43100_);
  and _51350_ (_05373_, _00129_, _00128_);
  or _51351_ (_00130_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or _51352_ (_00132_, \oc8051_gm_cxrom_1.cell5.data [2], _00115_);
  nand _51353_ (_00134_, _00132_, _00130_);
  nand _51354_ (_00136_, _00134_, _43100_);
  or _51355_ (_00138_, \oc8051_gm_cxrom_1.cell5.data [2], _43100_);
  and _51356_ (_05377_, _00138_, _00136_);
  or _51357_ (_00141_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or _51358_ (_00143_, \oc8051_gm_cxrom_1.cell5.data [3], _00115_);
  nand _51359_ (_00145_, _00143_, _00141_);
  nand _51360_ (_00147_, _00145_, _43100_);
  or _51361_ (_00149_, \oc8051_gm_cxrom_1.cell5.data [3], _43100_);
  and _51362_ (_05381_, _00149_, _00147_);
  or _51363_ (_00152_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or _51364_ (_00154_, \oc8051_gm_cxrom_1.cell5.data [4], _00115_);
  nand _51365_ (_00156_, _00154_, _00152_);
  nand _51366_ (_00158_, _00156_, _43100_);
  or _51367_ (_00160_, \oc8051_gm_cxrom_1.cell5.data [4], _43100_);
  and _51368_ (_05385_, _00160_, _00158_);
  or _51369_ (_00163_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or _51370_ (_00165_, \oc8051_gm_cxrom_1.cell5.data [5], _00115_);
  nand _51371_ (_00167_, _00165_, _00163_);
  nand _51372_ (_00169_, _00167_, _43100_);
  or _51373_ (_00171_, \oc8051_gm_cxrom_1.cell5.data [5], _43100_);
  and _51374_ (_05389_, _00171_, _00169_);
  or _51375_ (_00174_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or _51376_ (_00176_, \oc8051_gm_cxrom_1.cell5.data [6], _00115_);
  nand _51377_ (_00178_, _00176_, _00174_);
  nand _51378_ (_00180_, _00178_, _43100_);
  or _51379_ (_00182_, \oc8051_gm_cxrom_1.cell5.data [6], _43100_);
  and _51380_ (_05393_, _00182_, _00180_);
  or _51381_ (_00185_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not _51382_ (_00187_, \oc8051_gm_cxrom_1.cell6.valid );
  or _51383_ (_00188_, _00187_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand _51384_ (_00189_, _00188_, _00185_);
  nand _51385_ (_00190_, _00189_, _43100_);
  or _51386_ (_00191_, \oc8051_gm_cxrom_1.cell6.data [7], _43100_);
  and _51387_ (_05414_, _00191_, _00190_);
  or _51388_ (_00192_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or _51389_ (_00193_, \oc8051_gm_cxrom_1.cell6.data [0], _00187_);
  nand _51390_ (_00194_, _00193_, _00192_);
  nand _51391_ (_00195_, _00194_, _43100_);
  or _51392_ (_00196_, \oc8051_gm_cxrom_1.cell6.data [0], _43100_);
  and _51393_ (_05421_, _00196_, _00195_);
  or _51394_ (_00197_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or _51395_ (_00198_, \oc8051_gm_cxrom_1.cell6.data [1], _00187_);
  nand _51396_ (_00199_, _00198_, _00197_);
  nand _51397_ (_00200_, _00199_, _43100_);
  or _51398_ (_00201_, \oc8051_gm_cxrom_1.cell6.data [1], _43100_);
  and _51399_ (_05425_, _00201_, _00200_);
  or _51400_ (_00202_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or _51401_ (_00203_, \oc8051_gm_cxrom_1.cell6.data [2], _00187_);
  nand _51402_ (_00204_, _00203_, _00202_);
  nand _51403_ (_00205_, _00204_, _43100_);
  or _51404_ (_00206_, \oc8051_gm_cxrom_1.cell6.data [2], _43100_);
  and _51405_ (_05429_, _00206_, _00205_);
  or _51406_ (_00207_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or _51407_ (_00208_, \oc8051_gm_cxrom_1.cell6.data [3], _00187_);
  nand _51408_ (_00209_, _00208_, _00207_);
  nand _51409_ (_00210_, _00209_, _43100_);
  or _51410_ (_00211_, \oc8051_gm_cxrom_1.cell6.data [3], _43100_);
  and _51411_ (_05433_, _00211_, _00210_);
  or _51412_ (_00212_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or _51413_ (_00213_, \oc8051_gm_cxrom_1.cell6.data [4], _00187_);
  nand _51414_ (_00214_, _00213_, _00212_);
  nand _51415_ (_00215_, _00214_, _43100_);
  or _51416_ (_00216_, \oc8051_gm_cxrom_1.cell6.data [4], _43100_);
  and _51417_ (_05437_, _00216_, _00215_);
  or _51418_ (_00217_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or _51419_ (_00218_, \oc8051_gm_cxrom_1.cell6.data [5], _00187_);
  nand _51420_ (_00219_, _00218_, _00217_);
  nand _51421_ (_00220_, _00219_, _43100_);
  or _51422_ (_00221_, \oc8051_gm_cxrom_1.cell6.data [5], _43100_);
  and _51423_ (_05441_, _00221_, _00220_);
  or _51424_ (_00222_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or _51425_ (_00223_, \oc8051_gm_cxrom_1.cell6.data [6], _00187_);
  nand _51426_ (_00224_, _00223_, _00222_);
  nand _51427_ (_00225_, _00224_, _43100_);
  or _51428_ (_00226_, \oc8051_gm_cxrom_1.cell6.data [6], _43100_);
  and _51429_ (_05445_, _00226_, _00225_);
  or _51430_ (_00227_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not _51431_ (_00228_, \oc8051_gm_cxrom_1.cell7.valid );
  or _51432_ (_00229_, _00228_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand _51433_ (_00230_, _00229_, _00227_);
  nand _51434_ (_00231_, _00230_, _43100_);
  or _51435_ (_00232_, \oc8051_gm_cxrom_1.cell7.data [7], _43100_);
  and _51436_ (_05467_, _00232_, _00231_);
  or _51437_ (_00233_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or _51438_ (_00234_, \oc8051_gm_cxrom_1.cell7.data [0], _00228_);
  nand _51439_ (_00235_, _00234_, _00233_);
  nand _51440_ (_00236_, _00235_, _43100_);
  or _51441_ (_00237_, \oc8051_gm_cxrom_1.cell7.data [0], _43100_);
  and _51442_ (_05474_, _00237_, _00236_);
  or _51443_ (_00238_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or _51444_ (_00239_, \oc8051_gm_cxrom_1.cell7.data [1], _00228_);
  nand _51445_ (_00240_, _00239_, _00238_);
  nand _51446_ (_00241_, _00240_, _43100_);
  or _51447_ (_00242_, \oc8051_gm_cxrom_1.cell7.data [1], _43100_);
  and _51448_ (_05478_, _00242_, _00241_);
  or _51449_ (_00243_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or _51450_ (_00244_, \oc8051_gm_cxrom_1.cell7.data [2], _00228_);
  nand _51451_ (_00245_, _00244_, _00243_);
  nand _51452_ (_00246_, _00245_, _43100_);
  or _51453_ (_00247_, \oc8051_gm_cxrom_1.cell7.data [2], _43100_);
  and _51454_ (_05482_, _00247_, _00246_);
  or _51455_ (_00248_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or _51456_ (_00249_, \oc8051_gm_cxrom_1.cell7.data [3], _00228_);
  nand _51457_ (_00250_, _00249_, _00248_);
  nand _51458_ (_00251_, _00250_, _43100_);
  or _51459_ (_00252_, \oc8051_gm_cxrom_1.cell7.data [3], _43100_);
  and _51460_ (_05486_, _00252_, _00251_);
  or _51461_ (_00253_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or _51462_ (_00254_, \oc8051_gm_cxrom_1.cell7.data [4], _00228_);
  nand _51463_ (_00255_, _00254_, _00253_);
  nand _51464_ (_00256_, _00255_, _43100_);
  or _51465_ (_00257_, \oc8051_gm_cxrom_1.cell7.data [4], _43100_);
  and _51466_ (_05490_, _00257_, _00256_);
  or _51467_ (_00258_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or _51468_ (_00259_, \oc8051_gm_cxrom_1.cell7.data [5], _00228_);
  nand _51469_ (_00260_, _00259_, _00258_);
  nand _51470_ (_00261_, _00260_, _43100_);
  or _51471_ (_00262_, \oc8051_gm_cxrom_1.cell7.data [5], _43100_);
  and _51472_ (_05494_, _00262_, _00261_);
  or _51473_ (_00263_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or _51474_ (_00264_, \oc8051_gm_cxrom_1.cell7.data [6], _00228_);
  nand _51475_ (_00265_, _00264_, _00263_);
  nand _51476_ (_00266_, _00265_, _43100_);
  or _51477_ (_00267_, \oc8051_gm_cxrom_1.cell7.data [6], _43100_);
  and _51478_ (_05498_, _00267_, _00266_);
  or _51479_ (_00268_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not _51480_ (_00269_, \oc8051_gm_cxrom_1.cell8.valid );
  or _51481_ (_00270_, _00269_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand _51482_ (_00271_, _00270_, _00268_);
  nand _51483_ (_00272_, _00271_, _43100_);
  or _51484_ (_00273_, \oc8051_gm_cxrom_1.cell8.data [7], _43100_);
  and _51485_ (_05520_, _00273_, _00272_);
  or _51486_ (_00274_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or _51487_ (_00275_, \oc8051_gm_cxrom_1.cell8.data [0], _00269_);
  nand _51488_ (_00276_, _00275_, _00274_);
  nand _51489_ (_00277_, _00276_, _43100_);
  or _51490_ (_00278_, \oc8051_gm_cxrom_1.cell8.data [0], _43100_);
  and _51491_ (_05527_, _00278_, _00277_);
  or _51492_ (_00279_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or _51493_ (_00280_, \oc8051_gm_cxrom_1.cell8.data [1], _00269_);
  nand _51494_ (_00281_, _00280_, _00279_);
  nand _51495_ (_00282_, _00281_, _43100_);
  or _51496_ (_00283_, \oc8051_gm_cxrom_1.cell8.data [1], _43100_);
  and _51497_ (_05531_, _00283_, _00282_);
  or _51498_ (_00284_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or _51499_ (_00285_, \oc8051_gm_cxrom_1.cell8.data [2], _00269_);
  nand _51500_ (_00286_, _00285_, _00284_);
  nand _51501_ (_00287_, _00286_, _43100_);
  or _51502_ (_00288_, \oc8051_gm_cxrom_1.cell8.data [2], _43100_);
  and _51503_ (_05535_, _00288_, _00287_);
  or _51504_ (_00289_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or _51505_ (_00290_, \oc8051_gm_cxrom_1.cell8.data [3], _00269_);
  nand _51506_ (_00291_, _00290_, _00289_);
  nand _51507_ (_00292_, _00291_, _43100_);
  or _51508_ (_00293_, \oc8051_gm_cxrom_1.cell8.data [3], _43100_);
  and _51509_ (_05539_, _00293_, _00292_);
  or _51510_ (_00294_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or _51511_ (_00295_, \oc8051_gm_cxrom_1.cell8.data [4], _00269_);
  nand _51512_ (_00296_, _00295_, _00294_);
  nand _51513_ (_00297_, _00296_, _43100_);
  or _51514_ (_00298_, \oc8051_gm_cxrom_1.cell8.data [4], _43100_);
  and _51515_ (_05543_, _00298_, _00297_);
  or _51516_ (_00299_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or _51517_ (_00300_, \oc8051_gm_cxrom_1.cell8.data [5], _00269_);
  nand _51518_ (_00301_, _00300_, _00299_);
  nand _51519_ (_00302_, _00301_, _43100_);
  or _51520_ (_00303_, \oc8051_gm_cxrom_1.cell8.data [5], _43100_);
  and _51521_ (_05547_, _00303_, _00302_);
  or _51522_ (_00304_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or _51523_ (_00305_, \oc8051_gm_cxrom_1.cell8.data [6], _00269_);
  nand _51524_ (_00306_, _00305_, _00304_);
  nand _51525_ (_00307_, _00306_, _43100_);
  or _51526_ (_00308_, \oc8051_gm_cxrom_1.cell8.data [6], _43100_);
  and _51527_ (_05551_, _00308_, _00307_);
  or _51528_ (_00309_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not _51529_ (_00310_, \oc8051_gm_cxrom_1.cell9.valid );
  or _51530_ (_00311_, _00310_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand _51531_ (_00312_, _00311_, _00309_);
  nand _51532_ (_00313_, _00312_, _43100_);
  or _51533_ (_00314_, \oc8051_gm_cxrom_1.cell9.data [7], _43100_);
  and _51534_ (_05573_, _00314_, _00313_);
  or _51535_ (_00315_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or _51536_ (_00316_, \oc8051_gm_cxrom_1.cell9.data [0], _00310_);
  nand _51537_ (_00317_, _00316_, _00315_);
  nand _51538_ (_00318_, _00317_, _43100_);
  or _51539_ (_00319_, \oc8051_gm_cxrom_1.cell9.data [0], _43100_);
  and _51540_ (_05580_, _00319_, _00318_);
  or _51541_ (_00320_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or _51542_ (_00321_, \oc8051_gm_cxrom_1.cell9.data [1], _00310_);
  nand _51543_ (_00322_, _00321_, _00320_);
  nand _51544_ (_00323_, _00322_, _43100_);
  or _51545_ (_00324_, \oc8051_gm_cxrom_1.cell9.data [1], _43100_);
  and _51546_ (_05584_, _00324_, _00323_);
  or _51547_ (_00325_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or _51548_ (_00326_, \oc8051_gm_cxrom_1.cell9.data [2], _00310_);
  nand _51549_ (_00327_, _00326_, _00325_);
  nand _51550_ (_00328_, _00327_, _43100_);
  or _51551_ (_00329_, \oc8051_gm_cxrom_1.cell9.data [2], _43100_);
  and _51552_ (_05588_, _00329_, _00328_);
  or _51553_ (_00330_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or _51554_ (_00331_, \oc8051_gm_cxrom_1.cell9.data [3], _00310_);
  nand _51555_ (_00332_, _00331_, _00330_);
  nand _51556_ (_00333_, _00332_, _43100_);
  or _51557_ (_00334_, \oc8051_gm_cxrom_1.cell9.data [3], _43100_);
  and _51558_ (_05592_, _00334_, _00333_);
  or _51559_ (_00335_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or _51560_ (_00336_, \oc8051_gm_cxrom_1.cell9.data [4], _00310_);
  nand _51561_ (_00337_, _00336_, _00335_);
  nand _51562_ (_00338_, _00337_, _43100_);
  or _51563_ (_00339_, \oc8051_gm_cxrom_1.cell9.data [4], _43100_);
  and _51564_ (_05596_, _00339_, _00338_);
  or _51565_ (_00340_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or _51566_ (_00341_, \oc8051_gm_cxrom_1.cell9.data [5], _00310_);
  nand _51567_ (_00342_, _00341_, _00340_);
  nand _51568_ (_00343_, _00342_, _43100_);
  or _51569_ (_00344_, \oc8051_gm_cxrom_1.cell9.data [5], _43100_);
  and _51570_ (_05600_, _00344_, _00343_);
  or _51571_ (_00345_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or _51572_ (_00346_, \oc8051_gm_cxrom_1.cell9.data [6], _00310_);
  nand _51573_ (_00347_, _00346_, _00345_);
  nand _51574_ (_00348_, _00347_, _43100_);
  or _51575_ (_00349_, \oc8051_gm_cxrom_1.cell9.data [6], _43100_);
  and _51576_ (_05604_, _00349_, _00348_);
  or _51577_ (_00350_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not _51578_ (_00351_, \oc8051_gm_cxrom_1.cell10.valid );
  or _51579_ (_00352_, _00351_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand _51580_ (_00353_, _00352_, _00350_);
  nand _51581_ (_00354_, _00353_, _43100_);
  or _51582_ (_00355_, \oc8051_gm_cxrom_1.cell10.data [7], _43100_);
  and _51583_ (_05626_, _00355_, _00354_);
  or _51584_ (_00356_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or _51585_ (_00357_, \oc8051_gm_cxrom_1.cell10.data [0], _00351_);
  nand _51586_ (_00358_, _00357_, _00356_);
  nand _51587_ (_00359_, _00358_, _43100_);
  or _51588_ (_00360_, \oc8051_gm_cxrom_1.cell10.data [0], _43100_);
  and _51589_ (_05633_, _00360_, _00359_);
  or _51590_ (_00361_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or _51591_ (_00362_, \oc8051_gm_cxrom_1.cell10.data [1], _00351_);
  nand _51592_ (_00363_, _00362_, _00361_);
  nand _51593_ (_00364_, _00363_, _43100_);
  or _51594_ (_00365_, \oc8051_gm_cxrom_1.cell10.data [1], _43100_);
  and _51595_ (_05637_, _00365_, _00364_);
  or _51596_ (_00366_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or _51597_ (_00367_, \oc8051_gm_cxrom_1.cell10.data [2], _00351_);
  nand _51598_ (_00368_, _00367_, _00366_);
  nand _51599_ (_00369_, _00368_, _43100_);
  or _51600_ (_00370_, \oc8051_gm_cxrom_1.cell10.data [2], _43100_);
  and _51601_ (_05641_, _00370_, _00369_);
  or _51602_ (_00371_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or _51603_ (_00372_, \oc8051_gm_cxrom_1.cell10.data [3], _00351_);
  nand _51604_ (_00373_, _00372_, _00371_);
  nand _51605_ (_00374_, _00373_, _43100_);
  or _51606_ (_00375_, \oc8051_gm_cxrom_1.cell10.data [3], _43100_);
  and _51607_ (_05645_, _00375_, _00374_);
  or _51608_ (_00376_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or _51609_ (_00377_, \oc8051_gm_cxrom_1.cell10.data [4], _00351_);
  nand _51610_ (_00378_, _00377_, _00376_);
  nand _51611_ (_00379_, _00378_, _43100_);
  or _51612_ (_00380_, \oc8051_gm_cxrom_1.cell10.data [4], _43100_);
  and _51613_ (_05649_, _00380_, _00379_);
  or _51614_ (_00381_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or _51615_ (_00382_, \oc8051_gm_cxrom_1.cell10.data [5], _00351_);
  nand _51616_ (_00383_, _00382_, _00381_);
  nand _51617_ (_00384_, _00383_, _43100_);
  or _51618_ (_00385_, \oc8051_gm_cxrom_1.cell10.data [5], _43100_);
  and _51619_ (_05653_, _00385_, _00384_);
  or _51620_ (_00386_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or _51621_ (_00387_, \oc8051_gm_cxrom_1.cell10.data [6], _00351_);
  nand _51622_ (_00388_, _00387_, _00386_);
  nand _51623_ (_00389_, _00388_, _43100_);
  or _51624_ (_00390_, \oc8051_gm_cxrom_1.cell10.data [6], _43100_);
  and _51625_ (_05657_, _00390_, _00389_);
  or _51626_ (_00391_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not _51627_ (_00392_, \oc8051_gm_cxrom_1.cell11.valid );
  or _51628_ (_00393_, _00392_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand _51629_ (_00394_, _00393_, _00391_);
  nand _51630_ (_00395_, _00394_, _43100_);
  or _51631_ (_00396_, \oc8051_gm_cxrom_1.cell11.data [7], _43100_);
  and _51632_ (_05679_, _00396_, _00395_);
  or _51633_ (_00397_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or _51634_ (_00398_, \oc8051_gm_cxrom_1.cell11.data [0], _00392_);
  nand _51635_ (_00399_, _00398_, _00397_);
  nand _51636_ (_00400_, _00399_, _43100_);
  or _51637_ (_00401_, \oc8051_gm_cxrom_1.cell11.data [0], _43100_);
  and _51638_ (_05686_, _00401_, _00400_);
  or _51639_ (_00402_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or _51640_ (_00403_, \oc8051_gm_cxrom_1.cell11.data [1], _00392_);
  nand _51641_ (_00404_, _00403_, _00402_);
  nand _51642_ (_00405_, _00404_, _43100_);
  or _51643_ (_00406_, \oc8051_gm_cxrom_1.cell11.data [1], _43100_);
  and _51644_ (_05690_, _00406_, _00405_);
  or _51645_ (_00407_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or _51646_ (_00408_, \oc8051_gm_cxrom_1.cell11.data [2], _00392_);
  nand _51647_ (_00409_, _00408_, _00407_);
  nand _51648_ (_00410_, _00409_, _43100_);
  or _51649_ (_00411_, \oc8051_gm_cxrom_1.cell11.data [2], _43100_);
  and _51650_ (_05694_, _00411_, _00410_);
  or _51651_ (_00412_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or _51652_ (_00413_, \oc8051_gm_cxrom_1.cell11.data [3], _00392_);
  nand _51653_ (_00414_, _00413_, _00412_);
  nand _51654_ (_00415_, _00414_, _43100_);
  or _51655_ (_00416_, \oc8051_gm_cxrom_1.cell11.data [3], _43100_);
  and _51656_ (_05698_, _00416_, _00415_);
  or _51657_ (_00417_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or _51658_ (_00418_, \oc8051_gm_cxrom_1.cell11.data [4], _00392_);
  nand _51659_ (_00419_, _00418_, _00417_);
  nand _51660_ (_00420_, _00419_, _43100_);
  or _51661_ (_00421_, \oc8051_gm_cxrom_1.cell11.data [4], _43100_);
  and _51662_ (_05702_, _00421_, _00420_);
  or _51663_ (_00422_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or _51664_ (_00423_, \oc8051_gm_cxrom_1.cell11.data [5], _00392_);
  nand _51665_ (_00424_, _00423_, _00422_);
  nand _51666_ (_00425_, _00424_, _43100_);
  or _51667_ (_00426_, \oc8051_gm_cxrom_1.cell11.data [5], _43100_);
  and _51668_ (_05706_, _00426_, _00425_);
  or _51669_ (_00427_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or _51670_ (_00428_, \oc8051_gm_cxrom_1.cell11.data [6], _00392_);
  nand _51671_ (_00429_, _00428_, _00427_);
  nand _51672_ (_00430_, _00429_, _43100_);
  or _51673_ (_00431_, \oc8051_gm_cxrom_1.cell11.data [6], _43100_);
  and _51674_ (_05710_, _00431_, _00430_);
  or _51675_ (_00432_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not _51676_ (_00433_, \oc8051_gm_cxrom_1.cell12.valid );
  or _51677_ (_00434_, _00433_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand _51678_ (_00435_, _00434_, _00432_);
  nand _51679_ (_00436_, _00435_, _43100_);
  or _51680_ (_00437_, \oc8051_gm_cxrom_1.cell12.data [7], _43100_);
  and _51681_ (_05732_, _00437_, _00436_);
  or _51682_ (_00438_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or _51683_ (_00439_, \oc8051_gm_cxrom_1.cell12.data [0], _00433_);
  nand _51684_ (_00440_, _00439_, _00438_);
  nand _51685_ (_00441_, _00440_, _43100_);
  or _51686_ (_00442_, \oc8051_gm_cxrom_1.cell12.data [0], _43100_);
  and _51687_ (_05739_, _00442_, _00441_);
  or _51688_ (_00443_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or _51689_ (_00444_, \oc8051_gm_cxrom_1.cell12.data [1], _00433_);
  nand _51690_ (_00445_, _00444_, _00443_);
  nand _51691_ (_00446_, _00445_, _43100_);
  or _51692_ (_00447_, \oc8051_gm_cxrom_1.cell12.data [1], _43100_);
  and _51693_ (_05743_, _00447_, _00446_);
  or _51694_ (_00448_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or _51695_ (_00449_, \oc8051_gm_cxrom_1.cell12.data [2], _00433_);
  nand _51696_ (_00450_, _00449_, _00448_);
  nand _51697_ (_00451_, _00450_, _43100_);
  or _51698_ (_00452_, \oc8051_gm_cxrom_1.cell12.data [2], _43100_);
  and _51699_ (_05747_, _00452_, _00451_);
  or _51700_ (_00453_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or _51701_ (_00454_, \oc8051_gm_cxrom_1.cell12.data [3], _00433_);
  nand _51702_ (_00455_, _00454_, _00453_);
  nand _51703_ (_00456_, _00455_, _43100_);
  or _51704_ (_00457_, \oc8051_gm_cxrom_1.cell12.data [3], _43100_);
  and _51705_ (_05751_, _00457_, _00456_);
  or _51706_ (_00458_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or _51707_ (_00459_, \oc8051_gm_cxrom_1.cell12.data [4], _00433_);
  nand _51708_ (_00460_, _00459_, _00458_);
  nand _51709_ (_00461_, _00460_, _43100_);
  or _51710_ (_00462_, \oc8051_gm_cxrom_1.cell12.data [4], _43100_);
  and _51711_ (_05755_, _00462_, _00461_);
  or _51712_ (_00463_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or _51713_ (_00464_, \oc8051_gm_cxrom_1.cell12.data [5], _00433_);
  nand _51714_ (_00465_, _00464_, _00463_);
  nand _51715_ (_00466_, _00465_, _43100_);
  or _51716_ (_00467_, \oc8051_gm_cxrom_1.cell12.data [5], _43100_);
  and _51717_ (_05759_, _00467_, _00466_);
  or _51718_ (_00468_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or _51719_ (_00469_, \oc8051_gm_cxrom_1.cell12.data [6], _00433_);
  nand _51720_ (_00470_, _00469_, _00468_);
  nand _51721_ (_00471_, _00470_, _43100_);
  or _51722_ (_00472_, \oc8051_gm_cxrom_1.cell12.data [6], _43100_);
  and _51723_ (_05763_, _00472_, _00471_);
  or _51724_ (_00473_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not _51725_ (_00474_, \oc8051_gm_cxrom_1.cell13.valid );
  or _51726_ (_00475_, _00474_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand _51727_ (_00476_, _00475_, _00473_);
  nand _51728_ (_00477_, _00476_, _43100_);
  or _51729_ (_00478_, \oc8051_gm_cxrom_1.cell13.data [7], _43100_);
  and _51730_ (_05785_, _00478_, _00477_);
  or _51731_ (_00479_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or _51732_ (_00480_, \oc8051_gm_cxrom_1.cell13.data [0], _00474_);
  nand _51733_ (_00481_, _00480_, _00479_);
  nand _51734_ (_00482_, _00481_, _43100_);
  or _51735_ (_00483_, \oc8051_gm_cxrom_1.cell13.data [0], _43100_);
  and _51736_ (_05792_, _00483_, _00482_);
  or _51737_ (_00484_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or _51738_ (_00485_, \oc8051_gm_cxrom_1.cell13.data [1], _00474_);
  nand _51739_ (_00486_, _00485_, _00484_);
  nand _51740_ (_00487_, _00486_, _43100_);
  or _51741_ (_00488_, \oc8051_gm_cxrom_1.cell13.data [1], _43100_);
  and _51742_ (_05796_, _00488_, _00487_);
  or _51743_ (_00489_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or _51744_ (_00490_, \oc8051_gm_cxrom_1.cell13.data [2], _00474_);
  nand _51745_ (_00491_, _00490_, _00489_);
  nand _51746_ (_00492_, _00491_, _43100_);
  or _51747_ (_00493_, \oc8051_gm_cxrom_1.cell13.data [2], _43100_);
  and _51748_ (_05800_, _00493_, _00492_);
  or _51749_ (_00494_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or _51750_ (_00495_, \oc8051_gm_cxrom_1.cell13.data [3], _00474_);
  nand _51751_ (_00496_, _00495_, _00494_);
  nand _51752_ (_00497_, _00496_, _43100_);
  or _51753_ (_00498_, \oc8051_gm_cxrom_1.cell13.data [3], _43100_);
  and _51754_ (_05804_, _00498_, _00497_);
  or _51755_ (_00499_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or _51756_ (_00500_, \oc8051_gm_cxrom_1.cell13.data [4], _00474_);
  nand _51757_ (_00501_, _00500_, _00499_);
  nand _51758_ (_00502_, _00501_, _43100_);
  or _51759_ (_00503_, \oc8051_gm_cxrom_1.cell13.data [4], _43100_);
  and _51760_ (_05808_, _00503_, _00502_);
  or _51761_ (_00504_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or _51762_ (_00505_, \oc8051_gm_cxrom_1.cell13.data [5], _00474_);
  nand _51763_ (_00506_, _00505_, _00504_);
  nand _51764_ (_00507_, _00506_, _43100_);
  or _51765_ (_00508_, \oc8051_gm_cxrom_1.cell13.data [5], _43100_);
  and _51766_ (_05812_, _00508_, _00507_);
  or _51767_ (_00509_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or _51768_ (_00510_, \oc8051_gm_cxrom_1.cell13.data [6], _00474_);
  nand _51769_ (_00511_, _00510_, _00509_);
  nand _51770_ (_00512_, _00511_, _43100_);
  or _51771_ (_00513_, \oc8051_gm_cxrom_1.cell13.data [6], _43100_);
  and _51772_ (_05816_, _00513_, _00512_);
  or _51773_ (_00514_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not _51774_ (_00515_, \oc8051_gm_cxrom_1.cell14.valid );
  or _51775_ (_00516_, _00515_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand _51776_ (_00517_, _00516_, _00514_);
  nand _51777_ (_00518_, _00517_, _43100_);
  or _51778_ (_00519_, \oc8051_gm_cxrom_1.cell14.data [7], _43100_);
  and _51779_ (_05838_, _00519_, _00518_);
  or _51780_ (_00520_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or _51781_ (_00521_, \oc8051_gm_cxrom_1.cell14.data [0], _00515_);
  nand _51782_ (_00522_, _00521_, _00520_);
  nand _51783_ (_00523_, _00522_, _43100_);
  or _51784_ (_00524_, \oc8051_gm_cxrom_1.cell14.data [0], _43100_);
  and _51785_ (_05845_, _00524_, _00523_);
  or _51786_ (_00525_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or _51787_ (_00526_, \oc8051_gm_cxrom_1.cell14.data [1], _00515_);
  nand _51788_ (_00527_, _00526_, _00525_);
  nand _51789_ (_00528_, _00527_, _43100_);
  or _51790_ (_00529_, \oc8051_gm_cxrom_1.cell14.data [1], _43100_);
  and _51791_ (_05849_, _00529_, _00528_);
  or _51792_ (_00530_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or _51793_ (_00531_, \oc8051_gm_cxrom_1.cell14.data [2], _00515_);
  nand _51794_ (_00532_, _00531_, _00530_);
  nand _51795_ (_00533_, _00532_, _43100_);
  or _51796_ (_00534_, \oc8051_gm_cxrom_1.cell14.data [2], _43100_);
  and _51797_ (_05853_, _00534_, _00533_);
  or _51798_ (_00535_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or _51799_ (_00536_, \oc8051_gm_cxrom_1.cell14.data [3], _00515_);
  nand _51800_ (_00537_, _00536_, _00535_);
  nand _51801_ (_00538_, _00537_, _43100_);
  or _51802_ (_00539_, \oc8051_gm_cxrom_1.cell14.data [3], _43100_);
  and _51803_ (_05857_, _00539_, _00538_);
  or _51804_ (_00540_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or _51805_ (_00541_, \oc8051_gm_cxrom_1.cell14.data [4], _00515_);
  nand _51806_ (_00542_, _00541_, _00540_);
  nand _51807_ (_00543_, _00542_, _43100_);
  or _51808_ (_00545_, \oc8051_gm_cxrom_1.cell14.data [4], _43100_);
  and _51809_ (_05861_, _00545_, _00543_);
  or _51810_ (_00547_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or _51811_ (_00548_, \oc8051_gm_cxrom_1.cell14.data [5], _00515_);
  nand _51812_ (_00550_, _00548_, _00547_);
  nand _51813_ (_00551_, _00550_, _43100_);
  or _51814_ (_00553_, \oc8051_gm_cxrom_1.cell14.data [5], _43100_);
  and _51815_ (_05865_, _00553_, _00551_);
  or _51816_ (_00555_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or _51817_ (_00556_, \oc8051_gm_cxrom_1.cell14.data [6], _00515_);
  nand _51818_ (_00558_, _00556_, _00555_);
  nand _51819_ (_00559_, _00558_, _43100_);
  or _51820_ (_00561_, \oc8051_gm_cxrom_1.cell14.data [6], _43100_);
  and _51821_ (_05869_, _00561_, _00559_);
  or _51822_ (_00563_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not _51823_ (_00564_, \oc8051_gm_cxrom_1.cell15.valid );
  or _51824_ (_00566_, _00564_, \oc8051_gm_cxrom_1.cell15.data [7]);
  and _51825_ (_00567_, _00566_, _00563_);
  or _51826_ (_00569_, _00567_, rst);
  or _51827_ (_00570_, \oc8051_gm_cxrom_1.cell15.data [7], _43100_);
  and _51828_ (_05891_, _00570_, _00569_);
  or _51829_ (_00572_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or _51830_ (_00574_, \oc8051_gm_cxrom_1.cell15.data [0], _00564_);
  and _51831_ (_00575_, _00574_, _00572_);
  or _51832_ (_00577_, _00575_, rst);
  or _51833_ (_00578_, \oc8051_gm_cxrom_1.cell15.data [0], _43100_);
  and _51834_ (_05898_, _00578_, _00577_);
  or _51835_ (_00580_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or _51836_ (_00582_, \oc8051_gm_cxrom_1.cell15.data [1], _00564_);
  and _51837_ (_00583_, _00582_, _00580_);
  or _51838_ (_00585_, _00583_, rst);
  or _51839_ (_00586_, \oc8051_gm_cxrom_1.cell15.data [1], _43100_);
  and _51840_ (_05902_, _00586_, _00585_);
  or _51841_ (_00588_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or _51842_ (_00590_, \oc8051_gm_cxrom_1.cell15.data [2], _00564_);
  and _51843_ (_00591_, _00590_, _00588_);
  or _51844_ (_00593_, _00591_, rst);
  or _51845_ (_00594_, \oc8051_gm_cxrom_1.cell15.data [2], _43100_);
  and _51846_ (_05906_, _00594_, _00593_);
  or _51847_ (_00595_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or _51848_ (_00596_, \oc8051_gm_cxrom_1.cell15.data [3], _00564_);
  and _51849_ (_00597_, _00596_, _00595_);
  or _51850_ (_00598_, _00597_, rst);
  or _51851_ (_00599_, \oc8051_gm_cxrom_1.cell15.data [3], _43100_);
  and _51852_ (_05910_, _00599_, _00598_);
  or _51853_ (_00600_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or _51854_ (_00601_, \oc8051_gm_cxrom_1.cell15.data [4], _00564_);
  and _51855_ (_00602_, _00601_, _00600_);
  or _51856_ (_00603_, _00602_, rst);
  or _51857_ (_00604_, \oc8051_gm_cxrom_1.cell15.data [4], _43100_);
  and _51858_ (_05914_, _00604_, _00603_);
  or _51859_ (_00605_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or _51860_ (_00606_, \oc8051_gm_cxrom_1.cell15.data [5], _00564_);
  and _51861_ (_00607_, _00606_, _00605_);
  or _51862_ (_00608_, _00607_, rst);
  or _51863_ (_00609_, \oc8051_gm_cxrom_1.cell15.data [5], _43100_);
  and _51864_ (_05918_, _00609_, _00608_);
  or _51865_ (_00610_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or _51866_ (_00611_, \oc8051_gm_cxrom_1.cell15.data [6], _00564_);
  and _51867_ (_00612_, _00611_, _00610_);
  or _51868_ (_00613_, _00612_, rst);
  or _51869_ (_00614_, \oc8051_gm_cxrom_1.cell15.data [6], _43100_);
  and _51870_ (_05922_, _00614_, _00613_);
  nor _51871_ (_09697_, _38475_, rst);
  and _51872_ (_00615_, _36509_, _43100_);
  nand _51873_ (_00616_, _00615_, _38483_);
  nor _51874_ (_00617_, _38467_, _38439_);
  or _51875_ (_09700_, _00617_, _00616_);
  not _51876_ (_00618_, _37164_);
  and _51877_ (_00619_, _37654_, _37426_);
  and _51878_ (_00620_, _00619_, _00618_);
  and _51879_ (_00621_, _38215_, _38410_);
  and _51880_ (_00622_, _00621_, _38432_);
  and _51881_ (_00623_, _00622_, _37951_);
  and _51882_ (_00624_, _00623_, _00620_);
  not _51883_ (_00625_, _37426_);
  and _51884_ (_00626_, _37654_, _00625_);
  not _51885_ (_00627_, _36890_);
  not _51886_ (_00628_, _38432_);
  nor _51887_ (_00629_, _00628_, _38410_);
  not _51888_ (_00630_, _37951_);
  nor _51889_ (_00631_, _00630_, _38215_);
  and _51890_ (_00632_, _00631_, _00629_);
  and _51891_ (_00633_, _00632_, _00627_);
  and _51892_ (_00634_, _00622_, _00630_);
  and _51893_ (_00635_, _00634_, _37164_);
  or _51894_ (_00636_, _00635_, _00633_);
  and _51895_ (_00637_, _00636_, _00626_);
  or _51896_ (_00638_, _00637_, _00624_);
  not _51897_ (_00639_, _38215_);
  and _51898_ (_00640_, _00629_, _00639_);
  and _51899_ (_00641_, _00640_, _00630_);
  and _51900_ (_00642_, _37164_, _36890_);
  nor _51901_ (_00643_, _37654_, _37426_);
  and _51902_ (_00644_, _00643_, _00642_);
  and _51903_ (_00645_, _00644_, _00641_);
  and _51904_ (_00646_, _00619_, _37164_);
  and _51905_ (_00647_, _00646_, _00623_);
  or _51906_ (_00648_, _00647_, _00645_);
  and _51907_ (_00649_, _37164_, _00627_);
  and _51908_ (_00650_, _00649_, _00626_);
  and _51909_ (_00651_, _38432_, _38410_);
  and _51910_ (_00652_, _00631_, _00651_);
  and _51911_ (_00653_, _00652_, _00650_);
  not _51912_ (_00654_, _00651_);
  nor _51913_ (_00655_, _37164_, _00627_);
  and _51914_ (_00656_, _00655_, _00626_);
  and _51915_ (_00657_, _00656_, _00654_);
  or _51916_ (_00658_, _00657_, _00653_);
  or _51917_ (_00659_, _00658_, _00648_);
  not _51918_ (_00660_, _00652_);
  nor _51919_ (_00661_, _37164_, _36890_);
  and _51920_ (_00662_, _00661_, _00619_);
  and _51921_ (_00663_, _00642_, _00619_);
  nor _51922_ (_00664_, _00663_, _00662_);
  nor _51923_ (_00665_, _00664_, _00660_);
  and _51924_ (_00666_, _00643_, _00618_);
  and _51925_ (_00667_, _00627_, _38432_);
  and _51926_ (_00668_, _00667_, _00621_);
  or _51927_ (_00669_, _00668_, _00652_);
  and _51928_ (_00670_, _00669_, _00666_);
  or _51929_ (_00671_, _00670_, _00665_);
  or _51930_ (_00672_, _00671_, _00659_);
  not _51931_ (_00673_, _37654_);
  and _51932_ (_00674_, _00673_, _37426_);
  and _51933_ (_00675_, _00674_, _00661_);
  nor _51934_ (_00676_, _00675_, _00630_);
  nor _51935_ (_00677_, _00654_, _38215_);
  not _51936_ (_00678_, _00677_);
  nor _51937_ (_00679_, _00678_, _00676_);
  not _51938_ (_00680_, _00679_);
  and _51939_ (_00681_, _00655_, _00619_);
  and _51940_ (_00682_, _00652_, _00681_);
  and _51941_ (_00683_, _00674_, _00649_);
  and _51942_ (_00684_, _00683_, _00652_);
  nor _51943_ (_00685_, _00684_, _00682_);
  and _51944_ (_00686_, _00685_, _00680_);
  and _51945_ (_00687_, _36890_, _38432_);
  and _51946_ (_00688_, _00687_, _00621_);
  and _51947_ (_00689_, _00688_, _00666_);
  and _51948_ (_00690_, _00644_, _00628_);
  or _51949_ (_00691_, _00690_, _00689_);
  and _51950_ (_00692_, _00674_, _00655_);
  and _51951_ (_00693_, _00692_, _00634_);
  and _51952_ (_00694_, _00674_, _36890_);
  and _51953_ (_00695_, _00694_, _00652_);
  or _51954_ (_00696_, _00695_, _00693_);
  nor _51955_ (_00697_, _00696_, _00691_);
  nand _51956_ (_00698_, _00697_, _00686_);
  or _51957_ (_00699_, _00698_, _00672_);
  or _51958_ (_00700_, _00699_, _00638_);
  and _51959_ (_00701_, _00700_, _36520_);
  not _51960_ (_00702_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _51961_ (_00703_, _36498_, _18201_);
  and _51962_ (_00704_, _00703_, _38464_);
  nor _51963_ (_00705_, _00704_, _00702_);
  or _51964_ (_00706_, _00705_, rst);
  or _51965_ (_09703_, _00706_, _00701_);
  nand _51966_ (_00707_, _37426_, _36444_);
  or _51967_ (_00708_, _36444_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _51968_ (_00709_, _00708_, _43100_);
  and _51969_ (_09706_, _00709_, _00707_);
  and _51970_ (_00710_, \oc8051_top_1.oc8051_sfr1.wait_data , _43100_);
  and _51971_ (_00711_, _00710_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _51972_ (_00712_, _38457_, _38484_);
  and _51973_ (_00713_, _38440_, _38448_);
  and _51974_ (_00714_, _00713_, _36967_);
  or _51975_ (_00715_, _00714_, _00712_);
  and _51976_ (_00716_, _38453_, _38467_);
  or _51977_ (_00717_, _00716_, _38468_);
  or _51978_ (_00718_, _00717_, _38543_);
  and _51979_ (_00719_, _38520_, _38439_);
  and _51980_ (_00720_, _38440_, _38517_);
  or _51981_ (_00721_, _00720_, _00719_);
  nor _51982_ (_00722_, _00721_, _00718_);
  nand _51983_ (_00723_, _00722_, _38561_);
  or _51984_ (_00724_, _00723_, _00715_);
  and _51985_ (_00725_, _00724_, _00615_);
  or _51986_ (_09709_, _00725_, _00711_);
  and _51987_ (_00726_, _36967_, _38437_);
  and _51988_ (_00727_, _00726_, _38516_);
  or _51989_ (_00728_, _00727_, _38599_);
  not _51990_ (_00729_, _38270_);
  and _51991_ (_00730_, _00729_, _38455_);
  and _51992_ (_00731_, _00730_, _38517_);
  or _51993_ (_00732_, _00731_, _00728_);
  and _51994_ (_00733_, _38467_, _38449_);
  or _51995_ (_00734_, _00733_, _38441_);
  or _51996_ (_00735_, _00734_, _00732_);
  and _51997_ (_00736_, _00735_, _36509_);
  and _51998_ (_00737_, _38570_, _00702_);
  not _51999_ (_00738_, _38460_);
  and _52000_ (_00739_, _00738_, _00737_);
  and _52001_ (_00740_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52002_ (_00741_, _00740_, _00739_);
  or _52003_ (_00742_, _00741_, _00736_);
  and _52004_ (_09712_, _00742_, _43100_);
  and _52005_ (_00743_, _00710_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _52006_ (_00744_, _38457_, _38508_);
  nor _52007_ (_00745_, _38520_, _38508_);
  nor _52008_ (_00746_, _00745_, _38490_);
  or _52009_ (_00747_, _00746_, _00744_);
  and _52010_ (_00748_, _00730_, _38530_);
  or _52011_ (_00749_, _00748_, _00747_);
  nor _52012_ (_00750_, _00745_, _38454_);
  and _52013_ (_00751_, _36956_, _38437_);
  and _52014_ (_00752_, _00751_, _38507_);
  nor _52015_ (_00753_, _00752_, _00750_);
  not _52016_ (_00754_, _00753_);
  and _52017_ (_00755_, _38457_, _36956_);
  and _52018_ (_00756_, _00755_, _37731_);
  and _52019_ (_00757_, _38491_, _38437_);
  or _52020_ (_00758_, _00757_, _38591_);
  or _52021_ (_00759_, _00758_, _00756_);
  or _52022_ (_00760_, _00759_, _00734_);
  or _52023_ (_00761_, _00760_, _00754_);
  or _52024_ (_00762_, _00761_, _00749_);
  and _52025_ (_00763_, _00762_, _00615_);
  or _52026_ (_09715_, _00763_, _00743_);
  and _52027_ (_00764_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _52028_ (_00765_, _38551_, _36509_);
  or _52029_ (_00766_, _00765_, _00764_);
  or _52030_ (_00767_, _00766_, _00739_);
  and _52031_ (_09718_, _00767_, _43100_);
  and _52032_ (_00768_, _38530_, _38504_);
  and _52033_ (_00769_, _38438_, _38480_);
  and _52034_ (_00770_, _00769_, _36956_);
  or _52035_ (_00771_, _00770_, _00768_);
  or _52036_ (_00772_, _00771_, _00714_);
  and _52037_ (_00773_, _00771_, _38466_);
  or _52038_ (_00774_, _00773_, _36455_);
  and _52039_ (_00775_, _00774_, _00772_);
  not _52040_ (_00776_, _38484_);
  nor _52041_ (_00777_, _00617_, _00776_);
  nor _52042_ (_00778_, _00777_, _00713_);
  not _52043_ (_00779_, _00778_);
  and _52044_ (_00780_, _00779_, _00737_);
  or _52045_ (_00781_, _00780_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52046_ (_00782_, _00781_, _00775_);
  or _52047_ (_00783_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18201_);
  and _52048_ (_00784_, _00783_, _43100_);
  and _52049_ (_09721_, _00784_, _00782_);
  and _52050_ (_00785_, _00710_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and _52051_ (_00786_, _00751_, _38516_);
  or _52052_ (_00787_, _00752_, _00786_);
  or _52053_ (_00788_, _38530_, _38517_);
  and _52054_ (_00789_, _00788_, _38487_);
  or _52055_ (_00790_, _00789_, _00787_);
  and _52056_ (_00791_, _38504_, _37742_);
  or _52057_ (_00792_, _00748_, _00719_);
  or _52058_ (_00793_, _00792_, _00791_);
  or _52059_ (_00794_, _00727_, _38518_);
  or _52060_ (_00795_, _38441_, _38536_);
  or _52061_ (_00796_, _00795_, _00794_);
  or _52062_ (_00797_, _00796_, _00793_);
  or _52063_ (_00798_, _00797_, _00790_);
  and _52064_ (_00799_, _00798_, _00615_);
  or _52065_ (_09724_, _00799_, _00785_);
  and _52066_ (_00800_, _00710_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _52067_ (_00801_, _00730_, _38514_);
  and _52068_ (_00802_, _38440_, _38496_);
  or _52069_ (_00803_, _00802_, _38532_);
  nor _52070_ (_00804_, _00803_, _00801_);
  nand _52071_ (_00805_, _00804_, _00753_);
  nor _52072_ (_00806_, _37219_, _37720_);
  and _52073_ (_00807_, _00806_, _38488_);
  or _52074_ (_00808_, _00807_, _38603_);
  and _52075_ (_00809_, _38520_, _38487_);
  or _52076_ (_00810_, _00809_, _00808_);
  or _52077_ (_00811_, _38535_, _38528_);
  and _52078_ (_00812_, _38457_, _38527_);
  or _52079_ (_00813_, _00812_, _00731_);
  or _52080_ (_00814_, _00813_, _00811_);
  or _52081_ (_00815_, _00814_, _00810_);
  or _52082_ (_00816_, _00815_, _00805_);
  and _52083_ (_00817_, _00726_, _00806_);
  and _52084_ (_00818_, _00726_, _38444_);
  or _52085_ (_00819_, _00818_, _00817_);
  nor _52086_ (_00820_, _38589_, _38563_);
  nand _52087_ (_00821_, _00820_, _38541_);
  or _52088_ (_00822_, _00821_, _00819_);
  or _52089_ (_00823_, _00822_, _00749_);
  or _52090_ (_00824_, _00823_, _00816_);
  and _52091_ (_00825_, _00824_, _00615_);
  or _52092_ (_09727_, _00825_, _00800_);
  and _52093_ (_00826_, _00730_, _38497_);
  or _52094_ (_00827_, _00826_, _38600_);
  and _52095_ (_00828_, _00751_, _38447_);
  and _52096_ (_00829_, _00828_, _37470_);
  or _52097_ (_00830_, _00829_, _38583_);
  and _52098_ (_00831_, _38497_, _38437_);
  or _52099_ (_00832_, _00831_, _00830_);
  or _52100_ (_00833_, _00832_, _00827_);
  and _52101_ (_00834_, _00730_, _38449_);
  or _52102_ (_00835_, _00834_, _00833_);
  and _52103_ (_00836_, _00835_, _36509_);
  nand _52104_ (_00837_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand _52105_ (_00838_, _00837_, _38472_);
  or _52106_ (_00839_, _00838_, _00836_);
  and _52107_ (_09730_, _00839_, _43100_);
  or _52108_ (_00840_, _38521_, _38518_);
  not _52109_ (_00841_, _38564_);
  or _52110_ (_00842_, _00746_, _00841_);
  or _52111_ (_00843_, _00842_, _00840_);
  and _52112_ (_00844_, _37219_, _37709_);
  and _52113_ (_00845_, _00844_, _36956_);
  and _52114_ (_00846_, _00845_, _38481_);
  or _52115_ (_00847_, _00846_, _38531_);
  or _52116_ (_00848_, _00847_, _38528_);
  or _52117_ (_00849_, _00848_, _00768_);
  nand _52118_ (_00850_, _38552_, _38544_);
  or _52119_ (_00851_, _00850_, _00849_);
  or _52120_ (_00852_, _00851_, _00843_);
  and _52121_ (_00853_, _00726_, _38448_);
  or _52122_ (_00854_, _00853_, _00770_);
  and _52123_ (_00855_, _00751_, _00844_);
  or _52124_ (_00856_, _00855_, _38510_);
  or _52125_ (_00857_, _00856_, _00728_);
  or _52126_ (_00858_, _00857_, _00854_);
  and _52127_ (_00859_, _00845_, _38487_);
  or _52128_ (_00860_, _00859_, _38589_);
  or _52129_ (_00861_, _00860_, _38489_);
  or _52130_ (_00862_, _38586_, _38548_);
  or _52131_ (_00863_, _00862_, _00861_);
  or _52132_ (_00864_, _00863_, _00858_);
  or _52133_ (_00865_, _00864_, _00754_);
  or _52134_ (_00866_, _00865_, _00852_);
  and _52135_ (_00867_, _00866_, _36509_);
  or _52136_ (_00868_, _00773_, _00739_);
  and _52137_ (_00869_, _38466_, _38559_);
  or _52138_ (_00870_, _00869_, _00868_);
  and _52139_ (_00871_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52140_ (_00872_, _00871_, _00870_);
  or _52141_ (_00873_, _00872_, _00867_);
  and _52142_ (_09733_, _00873_, _43100_);
  nor _52143_ (_09792_, _38612_, rst);
  nor _52144_ (_09794_, _38575_, rst);
  nand _52145_ (_09797_, _00779_, _00615_);
  nand _52146_ (_00874_, _00713_, _00615_);
  not _52147_ (_00875_, _38467_);
  or _52148_ (_00876_, _00616_, _00875_);
  and _52149_ (_09800_, _00876_, _00874_);
  or _52150_ (_00877_, _00638_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _52151_ (_00878_, _00877_, _00704_);
  nor _52152_ (_00879_, _00703_, _38464_);
  or _52153_ (_00880_, _00879_, rst);
  or _52154_ (_09803_, _00880_, _00878_);
  nand _52155_ (_00881_, _37951_, _36444_);
  or _52156_ (_00882_, _36444_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _52157_ (_00883_, _00882_, _43100_);
  and _52158_ (_09806_, _00883_, _00881_);
  not _52159_ (_00884_, _36444_);
  or _52160_ (_00885_, _38215_, _00884_);
  or _52161_ (_00886_, _36444_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _52162_ (_00887_, _00886_, _43100_);
  and _52163_ (_09809_, _00887_, _00885_);
  nand _52164_ (_00888_, _38410_, _36444_);
  or _52165_ (_00889_, _36444_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _52166_ (_00890_, _00889_, _43100_);
  and _52167_ (_09812_, _00890_, _00888_);
  nand _52168_ (_00891_, _38432_, _36444_);
  or _52169_ (_00892_, _36444_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _52170_ (_00893_, _00892_, _43100_);
  and _52171_ (_09815_, _00893_, _00891_);
  or _52172_ (_00894_, _36890_, _00884_);
  or _52173_ (_00895_, _36444_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _52174_ (_00896_, _00895_, _43100_);
  and _52175_ (_09818_, _00896_, _00894_);
  nand _52176_ (_00897_, _37164_, _36444_);
  or _52177_ (_00898_, _36444_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _52178_ (_00899_, _00898_, _43100_);
  and _52179_ (_09821_, _00899_, _00897_);
  nand _52180_ (_00900_, _37654_, _36444_);
  or _52181_ (_00901_, _36444_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _52182_ (_00902_, _00901_, _43100_);
  and _52183_ (_09824_, _00902_, _00900_);
  or _52184_ (_00903_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _18201_);
  and _52185_ (_00904_, _00903_, _43100_);
  and _52186_ (_00905_, _00904_, _00781_);
  and _52187_ (_00906_, _38449_, _38487_);
  or _52188_ (_00907_, _00826_, _00906_);
  and _52189_ (_00908_, _00726_, _38499_);
  or _52190_ (_00909_, _00834_, _00908_);
  or _52191_ (_00910_, _00909_, _00907_);
  or _52192_ (_00911_, _38441_, _38593_);
  or _52193_ (_00912_, _00911_, _00910_);
  and _52194_ (_00913_, _38499_, _38437_);
  and _52195_ (_00914_, _00913_, _36956_);
  or _52196_ (_00915_, _00914_, _00831_);
  or _52197_ (_00916_, _38520_, _38507_);
  and _52198_ (_00917_, _00916_, _38457_);
  or _52199_ (_00918_, _00917_, _00915_);
  or _52200_ (_00919_, _00918_, _00912_);
  and _52201_ (_00920_, _00730_, _38500_);
  or _52202_ (_00921_, _00920_, _00830_);
  and _52203_ (_00922_, _38457_, _38445_);
  and _52204_ (_00923_, _00730_, _38484_);
  or _52205_ (_00924_, _00923_, _00922_);
  or _52206_ (_00925_, _00924_, _00921_);
  or _52207_ (_00926_, _00802_, _38603_);
  or _52208_ (_00928_, _00818_, _00801_);
  or _52209_ (_00929_, _00928_, _00926_);
  or _52210_ (_00930_, _00929_, _00925_);
  or _52211_ (_00931_, _00733_, _38540_);
  or _52212_ (_00932_, _00931_, _00812_);
  and _52213_ (_00933_, _38500_, _38487_);
  and _52214_ (_00934_, _00726_, _38483_);
  and _52215_ (_00935_, _00755_, _38483_);
  or _52216_ (_00936_, _00935_, _00934_);
  or _52217_ (_00937_, _00936_, _00933_);
  or _52218_ (_00938_, _00937_, _00932_);
  or _52219_ (_00939_, _00938_, _00930_);
  or _52220_ (_00940_, _00939_, _00919_);
  and _52221_ (_00941_, _00940_, _00615_);
  or _52222_ (_09827_, _00941_, _00905_);
  and _52223_ (_00942_, _00710_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not _52224_ (_00943_, _38519_);
  or _52225_ (_00944_, _00819_, _00943_);
  or _52226_ (_00945_, _38527_, _38514_);
  and _52227_ (_00946_, _00945_, _38504_);
  not _52228_ (_00947_, _38457_);
  nor _52229_ (_00948_, _00947_, _38501_);
  or _52230_ (_00949_, _00948_, _00946_);
  or _52231_ (_00950_, _00949_, _00944_);
  or _52232_ (_00951_, _00932_, _00810_);
  and _52233_ (_00952_, _38457_, _38514_);
  and _52234_ (_00953_, _37219_, _37720_);
  and _52235_ (_00954_, _00751_, _00953_);
  and _52236_ (_00955_, _00954_, _37470_);
  nor _52237_ (_00956_, _00955_, _38588_);
  not _52238_ (_00958_, _00956_);
  or _52239_ (_00959_, _00958_, _00756_);
  or _52240_ (_00960_, _00959_, _00952_);
  or _52241_ (_00961_, _00960_, _00715_);
  or _52242_ (_00962_, _00961_, _00951_);
  or _52243_ (_00963_, _00962_, _00950_);
  and _52244_ (_00964_, _00963_, _00615_);
  or _52245_ (_34277_, _00964_, _00942_);
  or _52246_ (_00965_, _00862_, _00854_);
  or _52247_ (_00966_, _00965_, _00852_);
  and _52248_ (_00967_, _00966_, _36509_);
  and _52249_ (_00968_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52250_ (_00969_, _00968_, _00870_);
  or _52251_ (_00970_, _00969_, _00967_);
  and _52252_ (_34279_, _00970_, _43100_);
  and _52253_ (_00971_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52254_ (_00972_, _00971_, _00868_);
  and _52255_ (_00973_, _00972_, _43100_);
  and _52256_ (_00974_, _38562_, _36967_);
  or _52257_ (_00975_, _00974_, _38599_);
  or _52258_ (_00977_, _00975_, _00861_);
  or _52259_ (_00978_, _00977_, _00771_);
  and _52260_ (_00979_, _00978_, _00615_);
  or _52261_ (_34282_, _00979_, _00973_);
  or _52262_ (_00980_, _00713_, _38459_);
  and _52263_ (_00981_, _00826_, _36956_);
  or _52264_ (_00982_, _00981_, _00920_);
  or _52265_ (_00983_, _00982_, _00980_);
  or _52266_ (_00984_, _00830_, _38582_);
  or _52267_ (_00985_, _00915_, _00802_);
  or _52268_ (_00986_, _00985_, _00984_);
  or _52269_ (_00987_, _00986_, _00983_);
  and _52270_ (_00988_, _38457_, _38517_);
  or _52271_ (_00989_, _00935_, _38458_);
  or _52272_ (_00990_, _00989_, _00988_);
  and _52273_ (_00991_, _00730_, _38491_);
  or _52274_ (_00992_, _00991_, _00834_);
  or _52275_ (_00993_, _00992_, _00712_);
  or _52276_ (_00994_, _00993_, _00917_);
  or _52277_ (_00995_, _00994_, _00990_);
  or _52278_ (_00996_, _00855_, _00906_);
  or _52279_ (_00997_, _00996_, _00859_);
  or _52280_ (_00998_, _00812_, _38446_);
  or _52281_ (_00999_, _00922_, _00952_);
  or _52282_ (_01000_, _00999_, _00998_);
  or _52283_ (_01001_, _01000_, _00997_);
  and _52284_ (_01002_, _00826_, _36967_);
  and _52285_ (_01003_, _38504_, _38500_);
  and _52286_ (_01004_, _00846_, _37470_);
  or _52287_ (_01005_, _01004_, _01003_);
  or _52288_ (_01006_, _01005_, _01002_);
  or _52289_ (_01007_, _01006_, _00771_);
  or _52290_ (_01008_, _01007_, _01001_);
  or _52291_ (_01009_, _01008_, _00995_);
  or _52292_ (_01010_, _01009_, _00987_);
  and _52293_ (_01011_, _01010_, _36509_);
  and _52294_ (_01012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52295_ (_01013_, _00780_, _38473_);
  or _52296_ (_01014_, _01013_, _01012_);
  or _52297_ (_01015_, _01014_, _01011_);
  and _52298_ (_34284_, _01015_, _43100_);
  and _52299_ (_01016_, _00859_, _37470_);
  or _52300_ (_01017_, _38459_, _00906_);
  or _52301_ (_01018_, _01017_, _38548_);
  or _52302_ (_01019_, _01018_, _01016_);
  or _52303_ (_01020_, _01019_, _00984_);
  or _52304_ (_01021_, _01020_, _00985_);
  and _52305_ (_01022_, _00751_, _38483_);
  or _52306_ (_01023_, _00846_, _00733_);
  nor _52307_ (_01024_, _01023_, _01022_);
  nand _52308_ (_01025_, _01024_, _38451_);
  and _52309_ (_01026_, _00945_, _38440_);
  or _52310_ (_01027_, _01026_, _38502_);
  or _52311_ (_01028_, _01027_, _01025_);
  or _52312_ (_01029_, _01028_, _00995_);
  or _52313_ (_01030_, _01029_, _01021_);
  and _52314_ (_01031_, _01030_, _36509_);
  and _52315_ (_01032_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52316_ (_01033_, _01032_, _01013_);
  or _52317_ (_01034_, _01033_, _01031_);
  and _52318_ (_34286_, _01034_, _43100_);
  and _52319_ (_01035_, _00710_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not _52320_ (_01036_, _42525_);
  or _52321_ (_01037_, _00834_, _01036_);
  and _52322_ (_01038_, _38440_, _38520_);
  and _52323_ (_01039_, _38440_, _38507_);
  and _52324_ (_01040_, _01039_, _36956_);
  or _52325_ (_01041_, _01040_, _01038_);
  or _52326_ (_01042_, _01041_, _00790_);
  or _52327_ (_01043_, _01042_, _01037_);
  not _52328_ (_01044_, _42524_);
  or _52329_ (_01045_, _00795_, _01044_);
  and _52330_ (_01046_, _38457_, _38520_);
  or _52331_ (_01047_, _01046_, _00748_);
  or _52332_ (_01048_, _01047_, _00840_);
  or _52333_ (_01049_, _01048_, _01045_);
  or _52334_ (_01050_, _00829_, _00727_);
  and _52335_ (_01051_, _38581_, _38497_);
  and _52336_ (_01052_, _38440_, _38491_);
  or _52337_ (_01053_, _01052_, _01051_);
  or _52338_ (_01054_, _01053_, _01050_);
  and _52339_ (_01055_, _38554_, _38437_);
  or _52340_ (_01056_, _01055_, _00906_);
  or _52341_ (_01057_, _01056_, _38550_);
  and _52342_ (_01058_, _38440_, _38554_);
  or _52343_ (_01059_, _01058_, _00981_);
  or _52344_ (_01060_, _01059_, _01057_);
  or _52345_ (_01061_, _01060_, _01054_);
  or _52346_ (_01062_, _01061_, _01049_);
  or _52347_ (_01063_, _01062_, _01043_);
  and _52348_ (_01064_, _01063_, _00615_);
  or _52349_ (_34288_, _01064_, _01035_);
  or _52350_ (_01065_, _00809_, _00807_);
  or _52351_ (_01066_, _01065_, _01002_);
  or _52352_ (_01067_, _01066_, _00814_);
  or _52353_ (_01068_, _01067_, _00983_);
  or _52354_ (_01069_, _01058_, _01046_);
  or _52355_ (_01070_, _01040_, _00915_);
  or _52356_ (_01071_, _01070_, _01069_);
  nand _52357_ (_01072_, _38585_, _38549_);
  or _52358_ (_01073_, _00817_, _38441_);
  or _52359_ (_01074_, _38446_, _38540_);
  or _52360_ (_01075_, _01074_, _01073_);
  or _52361_ (_01076_, _01075_, _01072_);
  or _52362_ (_01077_, _01076_, _01071_);
  or _52363_ (_01078_, _01077_, _01068_);
  and _52364_ (_01079_, _01078_, _00615_);
  and _52365_ (_01080_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _52366_ (_01081_, _38459_, _36466_);
  or _52367_ (_01082_, _01081_, _01080_);
  and _52368_ (_01083_, _01082_, _43100_);
  or _52369_ (_34290_, _01083_, _01079_);
  or _52370_ (_01084_, _00933_, _00914_);
  nor _52371_ (_01085_, _00757_, _38539_);
  nand _52372_ (_01086_, _01085_, _38590_);
  or _52373_ (_01087_, _01086_, _00993_);
  or _52374_ (_01088_, _01087_, _01084_);
  nor _52375_ (_01089_, _00920_, _38548_);
  not _52376_ (_01090_, _01089_);
  nor _52377_ (_01091_, _01090_, _38547_);
  or _52378_ (_01092_, _00731_, _38602_);
  and _52379_ (_01093_, _38440_, _38497_);
  or _52380_ (_01094_, _01093_, _01050_);
  nor _52381_ (_01095_, _01094_, _01092_);
  nand _52382_ (_01096_, _01095_, _01091_);
  or _52383_ (_01097_, _01096_, _01088_);
  or _52384_ (_01098_, _00935_, _38542_);
  or _52385_ (_01099_, _01098_, _01052_);
  or _52386_ (_01100_, _01099_, _00754_);
  or _52387_ (_01101_, _01100_, _00749_);
  or _52388_ (_01102_, _01101_, _01097_);
  and _52389_ (_01103_, _01102_, _36509_);
  and _52390_ (_01104_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52391_ (_01105_, _01104_, _38470_);
  or _52392_ (_01106_, _01105_, _01103_);
  and _52393_ (_34292_, _01106_, _43100_);
  or _52394_ (_01107_, _01047_, _00794_);
  or _52395_ (_01108_, _01090_, _01084_);
  or _52396_ (_01109_, _01108_, _01107_);
  or _52397_ (_01110_, _38599_, _38589_);
  nor _52398_ (_01111_, _01110_, _01039_);
  nand _52399_ (_01112_, _01111_, _42525_);
  or _52400_ (_01113_, _01112_, _00747_);
  or _52401_ (_01114_, _01113_, _01109_);
  or _52402_ (_01115_, _01114_, _01100_);
  and _52403_ (_01116_, _01115_, _00615_);
  and _52404_ (_01117_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52405_ (_01118_, _01117_, _38471_);
  and _52406_ (_01119_, _01118_, _43100_);
  or _52407_ (_34294_, _01119_, _01116_);
  and _52408_ (_01120_, _00710_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor _52409_ (_01121_, _00720_, _38522_);
  nand _52410_ (_01122_, _01121_, _42524_);
  not _52411_ (_01123_, _38438_);
  or _52412_ (_01124_, _38440_, _01123_);
  and _52413_ (_01125_, _01124_, _38491_);
  or _52414_ (_01126_, _01125_, _01069_);
  or _52415_ (_01127_, _01126_, _01122_);
  or _52416_ (_01128_, _01041_, _00833_);
  or _52417_ (_01129_, _01128_, _01037_);
  or _52418_ (_01130_, _01129_, _01127_);
  and _52419_ (_01131_, _01130_, _00615_);
  or _52420_ (_34296_, _01131_, _01120_);
  nor _52421_ (_39173_, _37426_, rst);
  nor _52422_ (_39174_, _42516_, rst);
  and _52423_ (_01132_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _52424_ (_01133_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _52425_ (_01134_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _52426_ (_01135_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _52427_ (_01136_, _01135_, _01134_);
  and _52428_ (_01137_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _52429_ (_01138_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _52430_ (_01139_, _01138_, _01137_);
  and _52431_ (_01140_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _52432_ (_01141_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _52433_ (_01142_, _01141_, _01140_);
  and _52434_ (_01143_, _01142_, _01139_);
  and _52435_ (_01144_, _01143_, _01136_);
  nor _52436_ (_01145_, _01144_, _36694_);
  nor _52437_ (_01146_, _01145_, _01133_);
  nor _52438_ (_01147_, _01146_, _42500_);
  nor _52439_ (_01148_, _01147_, _01132_);
  nor _52440_ (_39176_, _01148_, rst);
  nor _52441_ (_39186_, _37951_, rst);
  and _52442_ (_39188_, _38215_, _43100_);
  nor _52443_ (_39189_, _38410_, rst);
  nor _52444_ (_39190_, _38432_, rst);
  and _52445_ (_39191_, _36890_, _43100_);
  nor _52446_ (_39192_, _37164_, rst);
  nor _52447_ (_39193_, _37654_, rst);
  nor _52448_ (_39194_, _42682_, rst);
  nor _52449_ (_39195_, _42611_, rst);
  nor _52450_ (_39197_, _42803_, rst);
  nor _52451_ (_39198_, _42646_, rst);
  nor _52452_ (_39199_, _42551_, rst);
  nor _52453_ (_39200_, _42777_, rst);
  nor _52454_ (_39201_, _42739_, rst);
  and _52455_ (_01149_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _52456_ (_01150_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _52457_ (_01151_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _52458_ (_01152_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _52459_ (_01153_, _01152_, _01151_);
  and _52460_ (_01154_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _52461_ (_01155_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _52462_ (_01156_, _01155_, _01154_);
  and _52463_ (_01157_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _52464_ (_01158_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _52465_ (_01159_, _01158_, _01157_);
  and _52466_ (_01160_, _01159_, _01156_);
  and _52467_ (_01161_, _01160_, _01153_);
  nor _52468_ (_01162_, _01161_, _36694_);
  nor _52469_ (_01163_, _01162_, _01150_);
  nor _52470_ (_01164_, _01163_, _42500_);
  nor _52471_ (_01165_, _01164_, _01149_);
  nor _52472_ (_39203_, _01165_, rst);
  and _52473_ (_01166_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _52474_ (_01167_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _52475_ (_01168_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _52476_ (_01169_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _52477_ (_01170_, _01169_, _01168_);
  and _52478_ (_01171_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _52479_ (_01172_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _52480_ (_01173_, _01172_, _01171_);
  and _52481_ (_01174_, _01173_, _01170_);
  and _52482_ (_01175_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _52483_ (_01176_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _52484_ (_01177_, _01176_, _01175_);
  and _52485_ (_01178_, _01177_, _01174_);
  nor _52486_ (_01179_, _01178_, _36694_);
  nor _52487_ (_01180_, _01179_, _01167_);
  nor _52488_ (_01181_, _01180_, _42500_);
  nor _52489_ (_01182_, _01181_, _01166_);
  nor _52490_ (_39204_, _01182_, rst);
  and _52491_ (_01183_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _52492_ (_01184_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _52493_ (_01185_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _52494_ (_01186_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _52495_ (_01187_, _01186_, _01185_);
  and _52496_ (_01188_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _52497_ (_01189_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _52498_ (_01190_, _01189_, _01188_);
  and _52499_ (_01191_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _52500_ (_01192_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _52501_ (_01193_, _01192_, _01191_);
  and _52502_ (_01194_, _01193_, _01190_);
  and _52503_ (_01195_, _01194_, _01187_);
  nor _52504_ (_01196_, _01195_, _36694_);
  nor _52505_ (_01197_, _01196_, _01184_);
  nor _52506_ (_01198_, _01197_, _42500_);
  nor _52507_ (_01199_, _01198_, _01183_);
  nor _52508_ (_39205_, _01199_, rst);
  and _52509_ (_01200_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _52510_ (_01201_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _52511_ (_01202_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _52512_ (_01203_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _52513_ (_01204_, _01203_, _01202_);
  and _52514_ (_01205_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _52515_ (_01206_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _52516_ (_01207_, _01206_, _01205_);
  and _52517_ (_01208_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _52518_ (_01209_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _52519_ (_01210_, _01209_, _01208_);
  and _52520_ (_01212_, _01210_, _01207_);
  and _52521_ (_01214_, _01212_, _01204_);
  nor _52522_ (_01216_, _01214_, _36694_);
  nor _52523_ (_01218_, _01216_, _01201_);
  nor _52524_ (_01220_, _01218_, _42500_);
  nor _52525_ (_01222_, _01220_, _01200_);
  nor _52526_ (_39206_, _01222_, rst);
  and _52527_ (_01225_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _52528_ (_01227_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _52529_ (_01229_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _52530_ (_01231_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _52531_ (_01233_, _01231_, _01229_);
  and _52532_ (_01235_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _52533_ (_01237_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _52534_ (_01239_, _01237_, _01235_);
  and _52535_ (_01241_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _52536_ (_01243_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _52537_ (_01245_, _01243_, _01241_);
  and _52538_ (_01247_, _01245_, _01239_);
  and _52539_ (_01249_, _01247_, _01233_);
  nor _52540_ (_01251_, _01249_, _36694_);
  nor _52541_ (_01253_, _01251_, _01227_);
  nor _52542_ (_01255_, _01253_, _42500_);
  nor _52543_ (_01257_, _01255_, _01225_);
  nor _52544_ (_39207_, _01257_, rst);
  and _52545_ (_01260_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _52546_ (_01262_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _52547_ (_01264_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _52548_ (_01266_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _52549_ (_01268_, _01266_, _01264_);
  and _52550_ (_01270_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _52551_ (_01272_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _52552_ (_01274_, _01272_, _01270_);
  and _52553_ (_01276_, _01274_, _01268_);
  and _52554_ (_01278_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _52555_ (_01280_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _52556_ (_01282_, _01280_, _01278_);
  and _52557_ (_01284_, _01282_, _01276_);
  nor _52558_ (_01286_, _01284_, _36694_);
  nor _52559_ (_01288_, _01286_, _01262_);
  nor _52560_ (_01290_, _01288_, _42500_);
  nor _52561_ (_01292_, _01290_, _01260_);
  nor _52562_ (_39209_, _01292_, rst);
  and _52563_ (_01295_, _42500_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _52564_ (_01297_, _36694_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _52565_ (_01299_, _36738_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _52566_ (_01301_, _36781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _52567_ (_01303_, _01301_, _01299_);
  and _52568_ (_01305_, _36575_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _52569_ (_01306_, _36607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _52570_ (_01307_, _01306_, _01305_);
  and _52571_ (_01308_, _36705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _52572_ (_01309_, _36651_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _52573_ (_01310_, _01309_, _01308_);
  and _52574_ (_01311_, _01310_, _01307_);
  and _52575_ (_01312_, _01311_, _01303_);
  nor _52576_ (_01313_, _01312_, _36694_);
  nor _52577_ (_01314_, _01313_, _01297_);
  nor _52578_ (_01315_, _01314_, _42500_);
  nor _52579_ (_01316_, _01315_, _01295_);
  nor _52580_ (_39210_, _01316_, rst);
  and _52581_ (_01317_, _36520_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _52582_ (_01318_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _52583_ (_01319_, _01317_, _38760_);
  and _52584_ (_01320_, _01319_, _43100_);
  and _52585_ (_39234_, _01320_, _01318_);
  not _52586_ (_01321_, _01317_);
  or _52587_ (_01322_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _52588_ (_01323_, _36520_, _43100_);
  and _52589_ (_00000_, _01323_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _52590_ (_01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _43100_);
  or _52591_ (_01325_, _01324_, _00000_);
  and _52592_ (_39235_, _01325_, _01322_);
  nor _52593_ (_39273_, _42521_, rst);
  and _52594_ (_39275_, _42559_, _43100_);
  and _52595_ (_39276_, _42495_, _43100_);
  nor _52596_ (_01326_, _38561_, _38570_);
  nor _52597_ (_01327_, _42665_, _27650_);
  and _52598_ (_01328_, _42665_, _27650_);
  nor _52599_ (_01329_, _01328_, _01327_);
  nor _52600_ (_01330_, _42579_, _27825_);
  and _52601_ (_01331_, _42579_, _27825_);
  nor _52602_ (_01332_, _01331_, _01330_);
  nor _52603_ (_01333_, _01332_, _01329_);
  nor _52604_ (_01334_, _42787_, _27343_);
  and _52605_ (_01335_, _42787_, _27343_);
  nor _52606_ (_01336_, _01335_, _01334_);
  nor _52607_ (_01337_, _42743_, _27211_);
  and _52608_ (_01338_, _42743_, _27211_);
  nor _52609_ (_01339_, _01338_, _01337_);
  nor _52610_ (_01340_, _01339_, _01336_);
  and _52611_ (_01341_, _01340_, _01333_);
  and _52612_ (_01342_, _01341_, _42858_);
  nor _52613_ (_01343_, _31308_, _40112_);
  and _52614_ (_01344_, _01343_, _01342_);
  and _52615_ (_01345_, _01344_, _01326_);
  not _52616_ (_01346_, _01345_);
  not _52617_ (_01347_, _00786_);
  nor _52618_ (_01348_, _00991_, _38536_);
  and _52619_ (_01349_, _01348_, _01347_);
  and _52620_ (_01350_, _01349_, _00956_);
  nor _52621_ (_01351_, _01326_, _38469_);
  or _52622_ (_01352_, _28571_, _28209_);
  nor _52623_ (_01353_, _01352_, _28538_);
  and _52624_ (_01354_, _01353_, _31460_);
  nand _52625_ (_01355_, _01354_, _33725_);
  nor _52626_ (_01356_, _01355_, _34573_);
  and _52627_ (_01357_, _01356_, _01351_);
  and _52628_ (_01358_, _01357_, _35748_);
  and _52629_ (_01359_, _01358_, _29196_);
  not _52630_ (_01360_, _01359_);
  and _52631_ (_01361_, _01326_, _28944_);
  not _52632_ (_01362_, _01361_);
  nor _52633_ (_01363_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _52634_ (_01364_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _52635_ (_01365_, _01364_, _01363_);
  nor _52636_ (_01366_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _52637_ (_01367_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _52638_ (_01368_, _01367_, _01366_);
  and _52639_ (_01369_, _01368_, _01365_);
  and _52640_ (_01370_, _01369_, _38610_);
  not _52641_ (_01371_, _38469_);
  nor _52642_ (_01372_, _01326_, _38498_);
  nor _52643_ (_01373_, _01372_, _01371_);
  and _52644_ (_01374_, _01373_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _52645_ (_01375_, _01374_, _01370_);
  and _52646_ (_01376_, _01375_, _01362_);
  and _52647_ (_01377_, _01376_, _01360_);
  not _52648_ (_01378_, _38500_);
  nor _52649_ (_01379_, _38554_, _38445_);
  and _52650_ (_01380_, _01379_, _01378_);
  nor _52651_ (_01381_, _01380_, _00875_);
  not _52652_ (_01382_, _01381_);
  and _52653_ (_01383_, _01382_, _01377_);
  and _52654_ (_01384_, _01383_, _01350_);
  and _52655_ (_01385_, _38468_, _36967_);
  or _52656_ (_01386_, _01385_, _38559_);
  or _52657_ (_01387_, _01386_, _01377_);
  nor _52658_ (_01388_, _01387_, _38558_);
  or _52659_ (_01389_, _01388_, _01384_);
  nor _52660_ (_01390_, _00729_, _38414_);
  and _52661_ (_01391_, _38006_, _38454_);
  and _52662_ (_01392_, _01391_, _01390_);
  and _52663_ (_01393_, _01392_, _38445_);
  nor _52664_ (_01394_, _01393_, _00716_);
  and _52665_ (_01395_, _01394_, _01389_);
  and _52666_ (_01396_, _01395_, _38506_);
  nor _52667_ (_01397_, _01396_, _42532_);
  and _52668_ (_01398_, _38507_, _38504_);
  nor _52669_ (_01399_, _01398_, _00769_);
  nor _52670_ (_01400_, _01399_, _36466_);
  nor _52671_ (_01401_, _01400_, _38572_);
  not _52672_ (_01402_, _01401_);
  nor _52673_ (_01403_, _01402_, _01397_);
  nor _52674_ (_01404_, _39115_, _39106_);
  and _52675_ (_01405_, _01404_, _39170_);
  not _52676_ (_01406_, _01405_);
  and _52677_ (_01407_, _01406_, _01373_);
  not _52678_ (_01408_, _39409_);
  and _52679_ (_01409_, _01408_, _38610_);
  nor _52680_ (_01410_, _01409_, _01407_);
  not _52681_ (_01411_, _01410_);
  nor _52682_ (_01412_, _01411_, _01403_);
  nor _52683_ (_01413_, _42617_, _26860_);
  and _52684_ (_01414_, _42617_, _26860_);
  nor _52685_ (_01415_, _01414_, _01413_);
  and _52686_ (_01416_, _42701_, _32582_);
  nor _52687_ (_01417_, _42701_, _32582_);
  or _52688_ (_01418_, _01417_, _01416_);
  nor _52689_ (_01419_, _01418_, _01415_);
  nor _52690_ (_01420_, _42823_, _26740_);
  and _52691_ (_01421_, _42823_, _26740_);
  nor _52692_ (_01422_, _01421_, _01420_);
  nor _52693_ (_01423_, _01422_, _39432_);
  and _52694_ (_01424_, _01423_, _01419_);
  and _52695_ (_01425_, _01424_, _01342_);
  nor _52696_ (_01426_, _27496_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _52697_ (_01427_, _01426_, _01425_);
  not _52698_ (_01428_, _01427_);
  and _52699_ (_01429_, _01428_, _01412_);
  and _52700_ (_01430_, _01429_, _01346_);
  nor _52701_ (_01431_, _38572_, rst);
  and _52702_ (_39280_, _01431_, _01430_);
  and _52703_ (_39281_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _43100_);
  and _52704_ (_39282_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _43100_);
  not _52705_ (_01432_, _38572_);
  nor _52706_ (_01433_, _01432_, _30574_);
  not _52707_ (_01434_, _38845_);
  and _52708_ (_01435_, _38446_, _38466_);
  and _52709_ (_01436_, _01435_, _01434_);
  not _52710_ (_01437_, _38468_);
  and _52711_ (_01438_, _00956_, _38561_);
  and _52712_ (_01439_, _01438_, _01437_);
  and _52713_ (_01440_, _01439_, _01394_);
  and _52714_ (_01441_, _01440_, _01349_);
  nor _52715_ (_01442_, _01441_, _42532_);
  nor _52716_ (_01443_, _01435_, _01400_);
  not _52717_ (_01444_, _01443_);
  and _52718_ (_01445_, _01438_, _01348_);
  nor _52719_ (_01446_, _01445_, _42532_);
  and _52720_ (_01447_, _01398_, _36455_);
  not _52721_ (_01448_, _01447_);
  and _52722_ (_01449_, _38467_, _38497_);
  and _52723_ (_01450_, _01449_, _36455_);
  nor _52724_ (_01451_, _01450_, _38572_);
  and _52725_ (_01452_, _01451_, _01448_);
  not _52726_ (_01453_, _01452_);
  nor _52727_ (_01454_, _01453_, _01446_);
  nand _52728_ (_01455_, _01454_, _01444_);
  nor _52729_ (_01456_, _01455_, _01442_);
  and _52730_ (_01457_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52731_ (_01458_, _01457_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _52732_ (_01459_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _52733_ (_01460_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _52734_ (_01461_, _01460_, _01459_);
  and _52735_ (_01462_, _01461_, _01458_);
  and _52736_ (_01463_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _52737_ (_01464_, _01463_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _52738_ (_01465_, _01464_, _01462_);
  and _52739_ (_01466_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _52740_ (_01467_, _01466_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52741_ (_01468_, _01467_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _52742_ (_01469_, _01468_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _52743_ (_01470_, _01469_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _52744_ (_01471_, _01469_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _52745_ (_01472_, _01471_, _01470_);
  and _52746_ (_01473_, _01472_, _01456_);
  and _52747_ (_01474_, _01447_, _42517_);
  or _52748_ (_01475_, _01474_, _01473_);
  nor _52749_ (_01476_, _01444_, _01442_);
  and _52750_ (_01477_, _01476_, _01454_);
  and _52751_ (_01478_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _52752_ (_01479_, _01478_, _01475_);
  nor _52753_ (_01480_, _01479_, _01436_);
  nand _52754_ (_01481_, _01480_, _01430_);
  or _52755_ (_01482_, _01481_, _01433_);
  and _52756_ (_01483_, _01454_, _42516_);
  not _52757_ (_01484_, _01148_);
  nor _52758_ (_01485_, _01454_, _01484_);
  nor _52759_ (_01486_, _01485_, _01483_);
  and _52760_ (_01487_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _52761_ (_01488_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _52762_ (_01489_, _01454_, _42739_);
  not _52763_ (_01490_, _01316_);
  nor _52764_ (_01491_, _01454_, _01490_);
  nor _52765_ (_01492_, _01491_, _01489_);
  and _52766_ (_01493_, _01492_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _52767_ (_01494_, _01492_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _52768_ (_01495_, _01494_, _01493_);
  and _52769_ (_01496_, _01454_, _42777_);
  not _52770_ (_01497_, _01292_);
  nor _52771_ (_01498_, _01454_, _01497_);
  nor _52772_ (_01499_, _01498_, _01496_);
  and _52773_ (_01500_, _01499_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _52774_ (_01501_, _01499_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _52775_ (_01502_, _01454_, _42551_);
  not _52776_ (_01503_, _01257_);
  nor _52777_ (_01504_, _01454_, _01503_);
  nor _52778_ (_01505_, _01504_, _01502_);
  nand _52779_ (_01506_, _01505_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52780_ (_01507_, _01454_, _42646_);
  not _52781_ (_01508_, _01222_);
  nor _52782_ (_01509_, _01454_, _01508_);
  nor _52783_ (_01510_, _01509_, _01507_);
  and _52784_ (_01511_, _01510_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _52785_ (_01512_, _01510_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _52786_ (_01513_, _01454_, _42803_);
  not _52787_ (_01514_, _01199_);
  nor _52788_ (_01515_, _01454_, _01514_);
  nor _52789_ (_01516_, _01515_, _01513_);
  and _52790_ (_01517_, _01516_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _52791_ (_01518_, _01454_, _42611_);
  not _52792_ (_01519_, _01182_);
  nor _52793_ (_01520_, _01454_, _01519_);
  nor _52794_ (_01521_, _01520_, _01518_);
  and _52795_ (_01522_, _01521_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _52796_ (_01523_, _01454_, _42682_);
  not _52797_ (_01524_, _01165_);
  nor _52798_ (_01525_, _01454_, _01524_);
  nor _52799_ (_01526_, _01525_, _01523_);
  and _52800_ (_01527_, _01526_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _52801_ (_01528_, _01521_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _52802_ (_01529_, _01528_, _01522_);
  and _52803_ (_01530_, _01529_, _01527_);
  nor _52804_ (_01531_, _01530_, _01522_);
  not _52805_ (_01532_, _01531_);
  nor _52806_ (_01533_, _01516_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _52807_ (_01534_, _01533_, _01517_);
  and _52808_ (_01535_, _01534_, _01532_);
  nor _52809_ (_01536_, _01535_, _01517_);
  nor _52810_ (_01537_, _01536_, _01512_);
  or _52811_ (_01538_, _01537_, _01511_);
  or _52812_ (_01539_, _01505_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52813_ (_01540_, _01539_, _01506_);
  nand _52814_ (_01541_, _01540_, _01538_);
  and _52815_ (_01542_, _01541_, _01506_);
  nor _52816_ (_01543_, _01542_, _01501_);
  or _52817_ (_01544_, _01543_, _01500_);
  and _52818_ (_01545_, _01544_, _01495_);
  nor _52819_ (_01546_, _01545_, _01493_);
  nor _52820_ (_01547_, _01546_, _01488_);
  or _52821_ (_01548_, _01547_, _01487_);
  and _52822_ (_01549_, _01548_, _01464_);
  and _52823_ (_01550_, _01549_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _52824_ (_01551_, _01550_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52825_ (_01552_, _01551_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _52826_ (_01553_, _01552_, _01486_);
  not _52827_ (_01554_, _01486_);
  nor _52828_ (_01555_, _01548_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _52829_ (_01556_, _01555_, _38782_);
  and _52830_ (_01557_, _01556_, _38787_);
  and _52831_ (_01558_, _01557_, _38772_);
  nor _52832_ (_01559_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52833_ (_01560_, _01559_, _01558_);
  nor _52834_ (_01561_, _01560_, _01554_);
  nor _52835_ (_01562_, _01561_, _01553_);
  or _52836_ (_01563_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _52837_ (_01564_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _52838_ (_01565_, _01564_, _01563_);
  and _52839_ (_01566_, _01565_, _01562_);
  or _52840_ (_01567_, _01566_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _52841_ (_01568_, _01566_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _52842_ (_01569_, _01568_, _01567_);
  and _52843_ (_01570_, _38497_, _36455_);
  and _52844_ (_01571_, _01570_, _38467_);
  or _52845_ (_01572_, _01571_, _01442_);
  and _52846_ (_01573_, _01572_, _01455_);
  and _52847_ (_01574_, _01573_, _01569_);
  or _52848_ (_01575_, _01574_, _01482_);
  and _52849_ (_01576_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _52850_ (_01577_, _36564_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _52851_ (_01578_, _01577_, _42500_);
  nor _52852_ (_01579_, _01578_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _52853_ (_01580_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _52854_ (_01581_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _52855_ (_01582_, _01581_, _01580_);
  not _52856_ (_01583_, _01582_);
  nor _52857_ (_01584_, _01583_, _01579_);
  and _52858_ (_01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _52859_ (_01586_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _52860_ (_01587_, _01586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _52861_ (_01588_, _01587_, _01584_);
  and _52862_ (_01589_, _01588_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _52863_ (_01590_, _01589_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _52864_ (_01591_, _01590_, _01576_);
  and _52865_ (_01592_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _52866_ (_01593_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _52867_ (_01594_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _52868_ (_01595_, _01594_, _01593_);
  or _52869_ (_01596_, _01595_, _01430_);
  and _52870_ (_01597_, _01596_, _43100_);
  and _52871_ (_39283_, _01597_, _01575_);
  and _52872_ (_01598_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _43100_);
  and _52873_ (_01599_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _52874_ (_01600_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _52875_ (_01601_, _36509_, _01600_);
  not _52876_ (_01602_, _01601_);
  not _52877_ (_01603_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _52878_ (_01604_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _52879_ (_01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _52880_ (_01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _52881_ (_01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _52882_ (_01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _52883_ (_01609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _52884_ (_01610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _52885_ (_01611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _52886_ (_01612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _52887_ (_01613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _52888_ (_01614_, _01613_, _01612_);
  and _52889_ (_01615_, _01614_, _01611_);
  and _52890_ (_01616_, _01615_, _01610_);
  and _52891_ (_01617_, _01616_, _01609_);
  and _52892_ (_01618_, _01617_, _01608_);
  and _52893_ (_01619_, _01618_, _01607_);
  and _52894_ (_01620_, _01619_, _01606_);
  and _52895_ (_01621_, _01620_, _01605_);
  and _52896_ (_01622_, _01621_, _01604_);
  nor _52897_ (_01623_, _01622_, _01603_);
  and _52898_ (_01624_, _01622_, _01603_);
  nor _52899_ (_01625_, _01624_, _01623_);
  nor _52900_ (_01626_, _01621_, _01604_);
  nor _52901_ (_01627_, _01626_, _01622_);
  and _52902_ (_01628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _52903_ (_01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _52904_ (_01631_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _52905_ (_01632_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _52906_ (_01634_, _01632_, _01629_);
  and _52907_ (_01635_, _01634_, _01631_);
  nor _52908_ (_01637_, _01635_, _01629_);
  nor _52909_ (_01638_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _52910_ (_01640_, _01638_, _01628_);
  not _52911_ (_01641_, _01640_);
  nor _52912_ (_01643_, _01641_, _01637_);
  nor _52913_ (_01644_, _01643_, _01628_);
  not _52914_ (_01646_, _01644_);
  and _52915_ (_01647_, _01646_, _01619_);
  and _52916_ (_01649_, _01647_, _01606_);
  and _52917_ (_01650_, _01649_, _01605_);
  not _52918_ (_01652_, _01650_);
  nor _52919_ (_01653_, _01652_, _01627_);
  and _52920_ (_01655_, _01652_, _01627_);
  or _52921_ (_01656_, _01655_, _01653_);
  not _52922_ (_01658_, _01656_);
  and _52923_ (_01659_, _01644_, _01621_);
  and _52924_ (_01661_, _01644_, _01620_);
  nor _52925_ (_01662_, _01661_, _01605_);
  nor _52926_ (_01663_, _01662_, _01659_);
  not _52927_ (_01664_, _01663_);
  and _52928_ (_01665_, _01644_, _01619_);
  nor _52929_ (_01666_, _01665_, _01606_);
  nor _52930_ (_01667_, _01666_, _01661_);
  not _52931_ (_01668_, _01667_);
  and _52932_ (_01669_, _01644_, _01617_);
  and _52933_ (_01670_, _01669_, _01608_);
  nor _52934_ (_01671_, _01670_, _01607_);
  nor _52935_ (_01672_, _01671_, _01665_);
  not _52936_ (_01673_, _01672_);
  nor _52937_ (_01674_, _01669_, _01608_);
  nor _52938_ (_01675_, _01674_, _01670_);
  not _52939_ (_01676_, _01675_);
  not _52940_ (_01677_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _52941_ (_01678_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _52942_ (_01679_, _01644_, _01616_);
  and _52943_ (_01680_, _01679_, _01678_);
  nor _52944_ (_01681_, _01680_, _01677_);
  nor _52945_ (_01682_, _01681_, _01669_);
  not _52946_ (_01683_, _01682_);
  and _52947_ (_01684_, _01644_, _01614_);
  and _52948_ (_01685_, _01684_, _01611_);
  nor _52949_ (_01686_, _01685_, _01610_);
  nor _52950_ (_01687_, _01686_, _01679_);
  not _52951_ (_01688_, _01687_);
  nor _52952_ (_01689_, _01684_, _01611_);
  nor _52953_ (_01690_, _01689_, _01685_);
  not _52954_ (_01691_, _01690_);
  and _52955_ (_01692_, _01644_, _01613_);
  nor _52956_ (_01693_, _01692_, _01612_);
  nor _52957_ (_01694_, _01693_, _01684_);
  not _52958_ (_01695_, _01694_);
  not _52959_ (_01696_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _52960_ (_01697_, _01644_, _01696_);
  nor _52961_ (_01698_, _01644_, _01696_);
  nor _52962_ (_01699_, _01698_, _01697_);
  not _52963_ (_01700_, _01699_);
  nor _52964_ (_01701_, _00695_, _00653_);
  not _52965_ (_01702_, _00690_);
  and _52966_ (_01703_, _01702_, _00686_);
  and _52967_ (_01704_, _01703_, _01701_);
  nand _52968_ (_01705_, _00646_, _00641_);
  and _52969_ (_01706_, _00656_, _00641_);
  and _52970_ (_01707_, _00674_, _00642_);
  and _52971_ (_01708_, _01707_, _00634_);
  nor _52972_ (_01709_, _01708_, _01706_);
  and _52973_ (_01710_, _01709_, _01705_);
  and _52974_ (_01711_, _00661_, _00626_);
  and _52975_ (_01712_, _00642_, _00626_);
  or _52976_ (_01713_, _01712_, _01711_);
  and _52977_ (_01714_, _01713_, _00623_);
  not _52978_ (_01715_, _00641_);
  nor _52979_ (_01716_, _00692_, _00650_);
  nor _52980_ (_01717_, _01716_, _01715_);
  nor _52981_ (_01718_, _01717_, _01714_);
  and _52982_ (_01719_, _01718_, _01710_);
  not _52983_ (_01720_, _00623_);
  and _52984_ (_01721_, _00643_, _00649_);
  nor _52985_ (_01722_, _01721_, _00656_);
  or _52986_ (_01723_, _01722_, _01720_);
  nand _52987_ (_01724_, _00641_, _00620_);
  and _52988_ (_01725_, _01724_, _01723_);
  and _52989_ (_01726_, _00643_, _00655_);
  nor _52990_ (_01727_, _01726_, _00683_);
  nor _52991_ (_01728_, _01727_, _01715_);
  nor _52992_ (_01729_, _01728_, _00647_);
  and _52993_ (_01730_, _01729_, _01725_);
  and _52994_ (_01731_, _01730_, _01719_);
  and _52995_ (_01732_, _01731_, _01704_);
  not _52996_ (_01733_, _00665_);
  and _52997_ (_01734_, _00656_, _00632_);
  nor _52998_ (_01735_, _01734_, _00645_);
  and _52999_ (_01736_, _01735_, _01733_);
  not _53000_ (_01737_, _01707_);
  nor _53001_ (_01738_, _00640_, _00623_);
  nor _53002_ (_01739_, _01738_, _01737_);
  and _53003_ (_01740_, _00643_, _37164_);
  nor _53004_ (_01741_, _01740_, _01711_);
  nor _53005_ (_01742_, _01741_, _00660_);
  nor _53006_ (_01743_, _01742_, _01739_);
  and _53007_ (_01744_, _01743_, _01736_);
  nand _53008_ (_01745_, _00633_, _00620_);
  and _53009_ (_01746_, _00674_, _00618_);
  nor _53010_ (_01747_, _00639_, _38410_);
  and _53011_ (_01748_, _01747_, _00687_);
  and _53012_ (_01749_, _01748_, _01746_);
  and _53013_ (_01750_, _00650_, _00623_);
  and _53014_ (_01751_, _00681_, _00632_);
  or _53015_ (_01752_, _01751_, _01750_);
  nor _53016_ (_01753_, _01752_, _01749_);
  and _53017_ (_01754_, _01753_, _01745_);
  and _53018_ (_01755_, _00643_, _00661_);
  nand _53019_ (_01756_, _01755_, _00641_);
  and _53020_ (_01757_, _00652_, _01712_);
  and _53021_ (_01758_, _00692_, _00632_);
  nor _53022_ (_01759_, _01758_, _01757_);
  and _53023_ (_01760_, _01759_, _01756_);
  and _53024_ (_01761_, _01721_, _00641_);
  and _53025_ (_01762_, _00656_, _00652_);
  nor _53026_ (_01763_, _01762_, _01761_);
  nor _53027_ (_01764_, _01747_, _00628_);
  not _53028_ (_01765_, _01764_);
  and _53029_ (_01766_, _01765_, _00656_);
  and _53030_ (_01767_, _00683_, _00634_);
  nor _53031_ (_01768_, _01767_, _01766_);
  and _53032_ (_01769_, _01768_, _01763_);
  and _53033_ (_01770_, _01769_, _01760_);
  and _53034_ (_01771_, _01770_, _01754_);
  and _53035_ (_01772_, _01771_, _01744_);
  and _53036_ (_01773_, _01772_, _01732_);
  and _53037_ (_01774_, _00650_, _00628_);
  and _53038_ (_01775_, _01747_, _00626_);
  and _53039_ (_01776_, _01775_, _00667_);
  nor _53040_ (_01777_, _00692_, _01711_);
  nor _53041_ (_01778_, _01777_, _38432_);
  or _53042_ (_01779_, _01778_, _01776_);
  nor _53043_ (_01780_, _01779_, _01774_);
  nor _53044_ (_01781_, _00675_, _01712_);
  not _53045_ (_01782_, _01781_);
  and _53046_ (_01783_, _01782_, _00640_);
  and _53047_ (_01784_, _00683_, _00632_);
  nor _53048_ (_01785_, _01784_, _00623_);
  not _53049_ (_01786_, _00683_);
  nor _53050_ (_01787_, _00692_, _00644_);
  and _53051_ (_01788_, _01787_, _01786_);
  nor _53052_ (_01789_, _01788_, _01785_);
  and _53053_ (_01790_, _00675_, _00622_);
  or _53054_ (_01791_, _01790_, _01789_);
  nor _53055_ (_01792_, _01791_, _01783_);
  and _53056_ (_01793_, _01792_, _01780_);
  and _53057_ (_01794_, _01793_, _01773_);
  nor _53058_ (_01795_, _01634_, _01631_);
  nor _53059_ (_01796_, _01795_, _01635_);
  not _53060_ (_01797_, _01796_);
  nor _53061_ (_01798_, _01797_, _01794_);
  and _53062_ (_01799_, _00675_, _00634_);
  nor _53063_ (_01800_, _01767_, _01799_);
  nor _53064_ (_01801_, _00682_, _00647_);
  nor _53065_ (_01802_, _01717_, _01757_);
  and _53066_ (_01803_, _01802_, _01801_);
  and _53067_ (_01804_, _01803_, _01800_);
  not _53068_ (_01805_, _01766_);
  and _53069_ (_01806_, _01709_, _01736_);
  and _53070_ (_01807_, _01806_, _01805_);
  and _53071_ (_01808_, _01807_, _01804_);
  not _53072_ (_01809_, _01808_);
  nor _53073_ (_01810_, _01809_, _01794_);
  not _53074_ (_01811_, _01810_);
  nor _53075_ (_01812_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _53076_ (_01813_, _01812_, _01631_);
  and _53077_ (_01814_, _01813_, _01811_);
  and _53078_ (_01815_, _01797_, _01794_);
  nor _53079_ (_01816_, _01815_, _01798_);
  and _53080_ (_01817_, _01816_, _01814_);
  nor _53081_ (_01818_, _01817_, _01798_);
  not _53082_ (_01819_, _01818_);
  and _53083_ (_01820_, _01641_, _01637_);
  nor _53084_ (_01821_, _01820_, _01643_);
  and _53085_ (_01822_, _01821_, _01819_);
  and _53086_ (_01823_, _01822_, _01700_);
  not _53087_ (_01824_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53088_ (_01825_, _01697_, _01824_);
  or _53089_ (_01826_, _01825_, _01692_);
  and _53090_ (_01827_, _01826_, _01823_);
  and _53091_ (_01828_, _01827_, _01695_);
  and _53092_ (_01829_, _01828_, _01691_);
  and _53093_ (_01830_, _01829_, _01688_);
  nor _53094_ (_01831_, _01679_, _01678_);
  or _53095_ (_01832_, _01831_, _01680_);
  and _53096_ (_01833_, _01832_, _01830_);
  and _53097_ (_01834_, _01833_, _01683_);
  and _53098_ (_01835_, _01834_, _01676_);
  and _53099_ (_01836_, _01835_, _01673_);
  and _53100_ (_01837_, _01836_, _01668_);
  and _53101_ (_01838_, _01837_, _01664_);
  and _53102_ (_01839_, _01838_, _01658_);
  nor _53103_ (_01840_, _01839_, _01653_);
  not _53104_ (_01841_, _01840_);
  nor _53105_ (_01842_, _01841_, _01625_);
  and _53106_ (_01843_, _01841_, _01625_);
  or _53107_ (_01844_, _01843_, _01842_);
  or _53108_ (_01845_, _01844_, _01602_);
  or _53109_ (_01846_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _53110_ (_01847_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _53111_ (_01848_, _01847_, _01846_);
  and _53112_ (_01849_, _01848_, _01845_);
  or _53113_ (_39285_, _01849_, _01599_);
  nor _53114_ (_01850_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _53115_ (_39286_, _01850_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _53116_ (_39287_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _43100_);
  not _53117_ (_01851_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor _53118_ (_01852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _53119_ (_01853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _53120_ (_01854_, _01853_, _01852_);
  not _53121_ (_01855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _53122_ (_01856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _53123_ (_01857_, _01856_, _01855_);
  and _53124_ (_01858_, _01857_, _01854_);
  and _53125_ (_01859_, _01858_, _01851_);
  and _53126_ (_01860_, \oc8051_top_1.oc8051_rom1.ea_int , _36477_);
  nand _53127_ (_01861_, _01860_, _36509_);
  nand _53128_ (_01862_, _01861_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _53129_ (_01863_, _01862_, _01859_);
  and _53130_ (_39288_, _01863_, _43100_);
  and _53131_ (_01864_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _53132_ (_01865_, _01864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _53133_ (_39290_, _01865_, _43100_);
  nor _53134_ (_01866_, _01579_, _42500_);
  nor _53135_ (_01867_, _01794_, _36760_);
  nor _53136_ (_01868_, _01810_, _36629_);
  and _53137_ (_01869_, _01794_, _36760_);
  nor _53138_ (_01870_, _01869_, _01867_);
  and _53139_ (_01871_, _01870_, _01868_);
  nor _53140_ (_01872_, _01871_, _01867_);
  nor _53141_ (_01873_, _01872_, _42500_);
  and _53142_ (_01874_, _01873_, _36553_);
  nor _53143_ (_01875_, _01873_, _36553_);
  nor _53144_ (_01876_, _01875_, _01874_);
  nor _53145_ (_01877_, _01876_, _01866_);
  and _53146_ (_01878_, _36770_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _53147_ (_01879_, _01878_, _01866_);
  nor _53148_ (_01880_, _01879_, _01808_);
  or _53149_ (_01881_, _01880_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _53150_ (_01882_, _01881_, _01877_);
  and _53151_ (_39291_, _01882_, _43100_);
  nor _53152_ (_01883_, _36825_, _38149_);
  and _53153_ (_01884_, _37612_, _37382_);
  and _53154_ (_01885_, _01884_, _01883_);
  nand _53155_ (_01886_, _01323_, _38406_);
  nor _53156_ (_01887_, _01886_, _37907_);
  not _53157_ (_01888_, _38428_);
  and _53158_ (_01889_, _37121_, _01888_);
  and _53159_ (_01890_, _01889_, _01887_);
  and _53160_ (_39294_, _01890_, _01885_);
  nor _53161_ (_01891_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _53162_ (_01892_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _53163_ (_01893_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _53164_ (_39297_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _43100_);
  and _53165_ (_01894_, _39297_, _01893_);
  or _53166_ (_39295_, _01894_, _01892_);
  not _53167_ (_01895_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _53168_ (_01896_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _53169_ (_01897_, _01896_, _01895_);
  and _53170_ (_01898_, _01896_, _01895_);
  nor _53171_ (_01899_, _01898_, _01897_);
  not _53172_ (_01900_, _01899_);
  and _53173_ (_01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _53174_ (_01902_, _01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _53175_ (_01903_, _01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _53176_ (_01904_, _01903_, _01902_);
  or _53177_ (_01905_, _01904_, _01896_);
  and _53178_ (_01906_, _01905_, _01900_);
  nor _53179_ (_01907_, _01897_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _53180_ (_01908_, _01897_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _53181_ (_01909_, _01908_, _01907_);
  or _53182_ (_01910_, _01902_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _53183_ (_39299_, _01910_, _43100_);
  and _53184_ (_01911_, _39299_, _01909_);
  and _53185_ (_39298_, _01911_, _01906_);
  not _53186_ (_01912_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _53187_ (_01913_, _01579_, _01912_);
  and _53188_ (_01914_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _53189_ (_01915_, _01913_);
  and _53190_ (_01916_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _53191_ (_01917_, _01916_, _01914_);
  and _53192_ (_39300_, _01917_, _43100_);
  and _53193_ (_01918_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _53194_ (_01919_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _53195_ (_01920_, _01919_, _01918_);
  and _53196_ (_39301_, _01920_, _43100_);
  and _53197_ (_01921_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _53198_ (_01922_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53199_ (_01923_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _01922_);
  and _53200_ (_01924_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _53201_ (_01925_, _01924_, _01921_);
  and _53202_ (_39302_, _01925_, _43100_);
  and _53203_ (_01926_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53204_ (_01927_, _01926_, _01923_);
  and _53205_ (_39303_, _01927_, _43100_);
  or _53206_ (_01928_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _53207_ (_39305_, _01928_, _43100_);
  not _53208_ (_01929_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _53209_ (_01930_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _53210_ (_01931_, _01930_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53211_ (_01932_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _53212_ (_01933_, _01932_, _43100_);
  and _53213_ (_39306_, _01933_, _01931_);
  or _53214_ (_01934_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _53215_ (_39307_, _01934_, _43100_);
  nor _53216_ (_01935_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _53217_ (_01936_, _01935_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53218_ (_01937_, _01936_, _43100_);
  and _53219_ (_01938_, _39297_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _53220_ (_39308_, _01938_, _01937_);
  and _53221_ (_01939_, _01912_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _53222_ (_01940_, _01939_, _01936_);
  and _53223_ (_39309_, _01940_, _43100_);
  nand _53224_ (_01941_, _01936_, _38845_);
  or _53225_ (_01942_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _53226_ (_01943_, _01942_, _43100_);
  and _53227_ (_39310_, _01943_, _01941_);
  nand _53228_ (_01944_, _38477_, _43100_);
  nor _53229_ (_39311_, _01944_, _38614_);
  or _53230_ (_01945_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _53231_ (_01946_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand _53232_ (_01947_, _01317_, _01946_);
  and _53233_ (_01948_, _01947_, _43100_);
  and _53234_ (_39347_, _01948_, _01945_);
  or _53235_ (_01949_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _53236_ (_01950_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _53237_ (_01951_, _01317_, _01950_);
  and _53238_ (_01952_, _01951_, _43100_);
  and _53239_ (_39348_, _01952_, _01949_);
  or _53240_ (_01953_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _53241_ (_01954_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _53242_ (_01955_, _01317_, _01954_);
  and _53243_ (_01956_, _01955_, _43100_);
  and _53244_ (_39349_, _01956_, _01953_);
  or _53245_ (_01957_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _53246_ (_01958_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _53247_ (_01959_, _01317_, _01958_);
  and _53248_ (_01960_, _01959_, _43100_);
  and _53249_ (_39350_, _01960_, _01957_);
  or _53250_ (_01961_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not _53251_ (_01962_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand _53252_ (_01963_, _01317_, _01962_);
  and _53253_ (_01964_, _01963_, _43100_);
  and _53254_ (_39351_, _01964_, _01961_);
  or _53255_ (_01965_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not _53256_ (_01966_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand _53257_ (_01967_, _01317_, _01966_);
  and _53258_ (_01968_, _01967_, _43100_);
  and _53259_ (_39353_, _01968_, _01965_);
  or _53260_ (_01969_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or _53261_ (_01970_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _53262_ (_01971_, _01970_, _43100_);
  and _53263_ (_39354_, _01971_, _01969_);
  or _53264_ (_01972_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _53265_ (_01973_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand _53266_ (_01974_, _01317_, _01973_);
  and _53267_ (_01975_, _01974_, _43100_);
  and _53268_ (_39355_, _01975_, _01972_);
  or _53269_ (_01976_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _53270_ (_01977_, _01317_, _38776_);
  and _53271_ (_01978_, _01977_, _43100_);
  and _53272_ (_39356_, _01978_, _01976_);
  or _53273_ (_01979_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _53274_ (_01980_, _01317_, _38782_);
  and _53275_ (_01981_, _01980_, _43100_);
  and _53276_ (_39357_, _01981_, _01979_);
  or _53277_ (_01982_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _53278_ (_01983_, _01317_, _38787_);
  and _53279_ (_01984_, _01983_, _43100_);
  and _53280_ (_39358_, _01984_, _01982_);
  or _53281_ (_01985_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _53282_ (_01986_, _01317_, _38772_);
  and _53283_ (_01987_, _01986_, _43100_);
  and _53284_ (_39359_, _01987_, _01985_);
  or _53285_ (_01988_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _53286_ (_01989_, _01317_, _38793_);
  and _53287_ (_01990_, _01989_, _43100_);
  and _53288_ (_39360_, _01990_, _01988_);
  or _53289_ (_01991_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _53290_ (_01992_, _01317_, _38768_);
  and _53291_ (_01993_, _01992_, _43100_);
  and _53292_ (_39361_, _01993_, _01991_);
  or _53293_ (_01994_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _53294_ (_01995_, _01317_, _38764_);
  and _53295_ (_01996_, _01995_, _43100_);
  and _53296_ (_39362_, _01996_, _01994_);
  and _53297_ (_01997_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _53298_ (_01998_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _53299_ (_01999_, _01998_, _01997_);
  and _53300_ (_39367_, _01999_, _43100_);
  and _53301_ (_02000_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53302_ (_02001_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _53303_ (_02002_, _02001_, _02000_);
  and _53304_ (_39368_, _02002_, _43100_);
  and _53305_ (_02003_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _53306_ (_02004_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _53307_ (_02005_, _02004_, _02003_);
  and _53308_ (_39369_, _02005_, _43100_);
  and _53309_ (_02006_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53310_ (_02007_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _53311_ (_02008_, _02007_, _02006_);
  and _53312_ (_39370_, _02008_, _43100_);
  and _53313_ (_02009_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _53314_ (_02010_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or _53315_ (_02011_, _02010_, _02009_);
  and _53316_ (_39371_, _02011_, _43100_);
  and _53317_ (_02012_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _53318_ (_02013_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or _53319_ (_02014_, _02013_, _02012_);
  and _53320_ (_39372_, _02014_, _43100_);
  and _53321_ (_02015_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _53322_ (_02016_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or _53323_ (_02017_, _02016_, _02015_);
  and _53324_ (_39373_, _02017_, _43100_);
  and _53325_ (_02018_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _53326_ (_02019_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or _53327_ (_02020_, _02019_, _02018_);
  and _53328_ (_39374_, _02020_, _43100_);
  and _53329_ (_02021_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _53330_ (_02022_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or _53331_ (_02023_, _02022_, _02021_);
  and _53332_ (_39375_, _02023_, _43100_);
  and _53333_ (_02024_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _53334_ (_02025_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or _53335_ (_02026_, _02025_, _02024_);
  and _53336_ (_39376_, _02026_, _43100_);
  and _53337_ (_02027_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _53338_ (_02028_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or _53339_ (_02029_, _02028_, _02027_);
  and _53340_ (_39378_, _02029_, _43100_);
  and _53341_ (_02030_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _53342_ (_02031_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or _53343_ (_02032_, _02031_, _02030_);
  and _53344_ (_39379_, _02032_, _43100_);
  and _53345_ (_02033_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _53346_ (_02034_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or _53347_ (_02035_, _02034_, _02033_);
  and _53348_ (_39380_, _02035_, _43100_);
  and _53349_ (_02036_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _53350_ (_02037_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or _53351_ (_02038_, _02037_, _02036_);
  and _53352_ (_39381_, _02038_, _43100_);
  and _53353_ (_02039_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _53354_ (_02040_, _01321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or _53355_ (_02041_, _02040_, _02039_);
  and _53356_ (_39382_, _02041_, _43100_);
  and _53357_ (_39558_, _38006_, _43100_);
  and _53358_ (_39559_, _38270_, _43100_);
  and _53359_ (_39560_, _38414_, _43100_);
  nor _53360_ (_39561_, _42476_, rst);
  and _53361_ (_02042_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _53362_ (_02043_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or _53363_ (_02044_, _02043_, _02042_);
  and _53364_ (_39562_, _02044_, _43100_);
  and _53365_ (_02045_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _53366_ (_02046_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _53367_ (_02047_, _02046_, _02045_);
  and _53368_ (_39563_, _02047_, _43100_);
  and _53369_ (_02048_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _53370_ (_02049_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _53371_ (_02050_, _02049_, _02048_);
  and _53372_ (_39564_, _02050_, _43100_);
  and _53373_ (_02051_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _53374_ (_02052_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or _53375_ (_02053_, _02052_, _02051_);
  and _53376_ (_39565_, _02053_, _43100_);
  and _53377_ (_02054_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _53378_ (_02055_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _53379_ (_02056_, _02055_, _02054_);
  and _53380_ (_39567_, _02056_, _43100_);
  and _53381_ (_02057_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _53382_ (_02058_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or _53383_ (_02059_, _02058_, _02057_);
  and _53384_ (_39568_, _02059_, _43100_);
  and _53385_ (_02060_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _53386_ (_02061_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or _53387_ (_02062_, _02061_, _02060_);
  and _53388_ (_39569_, _02062_, _43100_);
  and _53389_ (_02063_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _53390_ (_02064_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or _53391_ (_02065_, _02064_, _02063_);
  and _53392_ (_39570_, _02065_, _43100_);
  and _53393_ (_02066_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and _53394_ (_02067_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _53395_ (_02068_, _02067_, _02066_);
  and _53396_ (_39571_, _02068_, _43100_);
  and _53397_ (_02069_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and _53398_ (_02070_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _53399_ (_02071_, _02070_, _02069_);
  and _53400_ (_39572_, _02071_, _43100_);
  and _53401_ (_02072_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and _53402_ (_02073_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _53403_ (_02074_, _02073_, _02072_);
  and _53404_ (_39573_, _02074_, _43100_);
  and _53405_ (_02075_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and _53406_ (_02076_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _53407_ (_02077_, _02076_, _02075_);
  and _53408_ (_39574_, _02077_, _43100_);
  and _53409_ (_02078_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and _53410_ (_02079_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _53411_ (_02080_, _02079_, _02078_);
  and _53412_ (_39575_, _02080_, _43100_);
  and _53413_ (_02081_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and _53414_ (_02082_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _53415_ (_02083_, _02082_, _02081_);
  and _53416_ (_39576_, _02083_, _43100_);
  and _53417_ (_02084_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and _53418_ (_02085_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _53419_ (_02086_, _02085_, _02084_);
  and _53420_ (_39578_, _02086_, _43100_);
  and _53421_ (_02087_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and _53422_ (_02088_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _53423_ (_02089_, _02088_, _02087_);
  and _53424_ (_39579_, _02089_, _43100_);
  and _53425_ (_02090_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _53426_ (_02091_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _53427_ (_02092_, _02091_, _02090_);
  and _53428_ (_39580_, _02092_, _43100_);
  and _53429_ (_02093_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _53430_ (_02094_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _53431_ (_02095_, _02094_, _02093_);
  and _53432_ (_39581_, _02095_, _43100_);
  and _53433_ (_02096_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _53434_ (_02097_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _53435_ (_02098_, _02097_, _02096_);
  and _53436_ (_39582_, _02098_, _43100_);
  and _53437_ (_02099_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _53438_ (_02100_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _53439_ (_02101_, _02100_, _02099_);
  and _53440_ (_39583_, _02101_, _43100_);
  and _53441_ (_02102_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _53442_ (_02103_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _53443_ (_02104_, _02103_, _02102_);
  and _53444_ (_39584_, _02104_, _43100_);
  and _53445_ (_02105_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _53446_ (_02106_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _53447_ (_02107_, _02106_, _02105_);
  and _53448_ (_39585_, _02107_, _43100_);
  and _53449_ (_02108_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _53450_ (_02109_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _53451_ (_02110_, _02109_, _02108_);
  and _53452_ (_39586_, _02110_, _43100_);
  and _53453_ (_02111_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _53454_ (_02113_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _53455_ (_02115_, _02113_, _02111_);
  and _53456_ (_39587_, _02115_, _43100_);
  and _53457_ (_02118_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _53458_ (_02120_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _53459_ (_02122_, _02120_, _02118_);
  and _53460_ (_39589_, _02122_, _43100_);
  and _53461_ (_02125_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _53462_ (_02127_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _53463_ (_02129_, _02127_, _02125_);
  and _53464_ (_39590_, _02129_, _43100_);
  and _53465_ (_02132_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _53466_ (_02134_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _53467_ (_02136_, _02134_, _02132_);
  and _53468_ (_39591_, _02136_, _43100_);
  and _53469_ (_02139_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _53470_ (_02141_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _53471_ (_02143_, _02141_, _02139_);
  and _53472_ (_39592_, _02143_, _43100_);
  and _53473_ (_02146_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _53474_ (_02148_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _53475_ (_02150_, _02148_, _02146_);
  and _53476_ (_39593_, _02150_, _43100_);
  and _53477_ (_02153_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _53478_ (_02155_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _53479_ (_02157_, _02155_, _02153_);
  and _53480_ (_39594_, _02157_, _43100_);
  and _53481_ (_02160_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _53482_ (_02162_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _53483_ (_02164_, _02162_, _02160_);
  and _53484_ (_39595_, _02164_, _43100_);
  nor _53485_ (_39596_, _42697_, rst);
  nor _53486_ (_39598_, _42591_, rst);
  nor _53487_ (_39599_, _42815_, rst);
  nor _53488_ (_39600_, _42661_, rst);
  nor _53489_ (_39601_, _42575_, rst);
  and _53490_ (_39602_, _42762_, _43100_);
  nor _53491_ (_39604_, _42720_, rst);
  and _53492_ (_39620_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _43100_);
  and _53493_ (_39621_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _43100_);
  and _53494_ (_39622_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _43100_);
  and _53495_ (_39623_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _43100_);
  and _53496_ (_39624_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _43100_);
  and _53497_ (_39626_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _43100_);
  and _53498_ (_39627_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _43100_);
  or _53499_ (_02170_, _01477_, _01435_);
  and _53500_ (_02171_, _02170_, _31809_);
  or _53501_ (_02172_, _01526_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _53502_ (_02173_, _01527_);
  nor _53503_ (_02174_, _01450_, _01442_);
  not _53504_ (_02175_, _02174_);
  and _53505_ (_02176_, _02175_, _01455_);
  and _53506_ (_02177_, _02176_, _02173_);
  and _53507_ (_02178_, _02177_, _02172_);
  and _53508_ (_02179_, _01456_, _42683_);
  and _53509_ (_02180_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _53510_ (_02181_, _02180_, _02179_);
  and _53511_ (_02182_, _01447_, _01524_);
  or _53512_ (_02183_, _02182_, _02181_);
  nor _53513_ (_02184_, _02183_, _02178_);
  nand _53514_ (_02185_, _02184_, _01430_);
  or _53515_ (_02186_, _02185_, _02171_);
  or _53516_ (_02187_, _01430_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _53517_ (_02188_, _02187_, _43100_);
  and _53518_ (_39628_, _02188_, _02186_);
  and _53519_ (_02189_, _02170_, _32506_);
  or _53520_ (_02190_, _01529_, _01527_);
  not _53521_ (_02191_, _01530_);
  and _53522_ (_02192_, _02176_, _02191_);
  and _53523_ (_02193_, _02192_, _02190_);
  and _53524_ (_02194_, _01456_, _42612_);
  and _53525_ (_02195_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _53526_ (_02196_, _02195_, _02194_);
  and _53527_ (_02197_, _01447_, _01519_);
  or _53528_ (_02198_, _02197_, _02196_);
  nor _53529_ (_02199_, _02198_, _02193_);
  nand _53530_ (_02200_, _02199_, _01430_);
  or _53531_ (_02201_, _02200_, _02189_);
  or _53532_ (_02202_, _01430_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _53533_ (_02203_, _02202_, _43100_);
  and _53534_ (_39629_, _02203_, _02201_);
  and _53535_ (_02204_, _02170_, _33213_);
  or _53536_ (_02205_, _01534_, _01532_);
  not _53537_ (_02206_, _01535_);
  and _53538_ (_02207_, _02176_, _02206_);
  and _53539_ (_02208_, _02207_, _02205_);
  and _53540_ (_02209_, _01456_, _42804_);
  and _53541_ (_02210_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _53542_ (_02211_, _02210_, _02209_);
  and _53543_ (_02212_, _01447_, _01514_);
  or _53544_ (_02213_, _02212_, _02211_);
  nor _53545_ (_02214_, _02213_, _02208_);
  nand _53546_ (_02215_, _02214_, _01430_);
  or _53547_ (_02216_, _02215_, _02204_);
  not _53548_ (_02217_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _53549_ (_02218_, _01579_, _02217_);
  and _53550_ (_02219_, _01579_, _02217_);
  nor _53551_ (_02220_, _02219_, _02218_);
  or _53552_ (_02221_, _02220_, _01430_);
  and _53553_ (_02222_, _02221_, _43100_);
  and _53554_ (_39630_, _02222_, _02216_);
  and _53555_ (_02223_, _02170_, _33964_);
  or _53556_ (_02224_, _01512_, _01511_);
  or _53557_ (_02225_, _02224_, _01536_);
  nand _53558_ (_02226_, _02224_, _01536_);
  and _53559_ (_02227_, _02226_, _02176_);
  and _53560_ (_02228_, _02227_, _02225_);
  and _53561_ (_02229_, _01456_, _42647_);
  and _53562_ (_02230_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _53563_ (_02231_, _02230_, _02229_);
  and _53564_ (_02232_, _01447_, _01508_);
  or _53565_ (_02233_, _02232_, _02231_);
  nor _53566_ (_02234_, _02233_, _02228_);
  nand _53567_ (_02235_, _02234_, _01430_);
  or _53568_ (_02236_, _02235_, _02223_);
  and _53569_ (_02237_, _02218_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53570_ (_02238_, _02218_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53571_ (_02239_, _02238_, _02237_);
  or _53572_ (_02240_, _02239_, _01430_);
  and _53573_ (_02241_, _02240_, _43100_);
  and _53574_ (_39631_, _02241_, _02236_);
  and _53575_ (_02242_, _02170_, _34704_);
  or _53576_ (_02243_, _01540_, _01538_);
  and _53577_ (_02244_, _02176_, _01541_);
  and _53578_ (_02245_, _02244_, _02243_);
  and _53579_ (_02246_, _01456_, _42552_);
  and _53580_ (_02247_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _53581_ (_02248_, _02247_, _02246_);
  and _53582_ (_02249_, _01447_, _01503_);
  or _53583_ (_02250_, _02249_, _02248_);
  nor _53584_ (_02251_, _02250_, _02245_);
  nand _53585_ (_02252_, _02251_, _01430_);
  or _53586_ (_02253_, _02252_, _02242_);
  and _53587_ (_02254_, _02237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53588_ (_02255_, _02237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53589_ (_02256_, _02255_, _02254_);
  or _53590_ (_02257_, _02256_, _01430_);
  and _53591_ (_02258_, _02257_, _43100_);
  and _53592_ (_39632_, _02258_, _02253_);
  and _53593_ (_02259_, _02170_, _35531_);
  and _53594_ (_02260_, _01456_, _42778_);
  and _53595_ (_02261_, _01447_, _01497_);
  and _53596_ (_02262_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _53597_ (_02263_, _02262_, _02261_);
  or _53598_ (_02264_, _02263_, _02260_);
  or _53599_ (_02265_, _01501_, _01500_);
  or _53600_ (_02266_, _02265_, _01542_);
  nand _53601_ (_02267_, _02265_, _01542_);
  and _53602_ (_02268_, _02267_, _02176_);
  and _53603_ (_02269_, _02268_, _02266_);
  nor _53604_ (_02270_, _02269_, _02264_);
  nand _53605_ (_02271_, _02270_, _01430_);
  or _53606_ (_02272_, _02271_, _02259_);
  nor _53607_ (_02273_, _02254_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _53608_ (_02274_, _02273_, _01584_);
  or _53609_ (_02275_, _02274_, _01430_);
  and _53610_ (_02276_, _02275_, _43100_);
  and _53611_ (_39633_, _02276_, _02272_);
  nor _53612_ (_02277_, _01584_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _53613_ (_02278_, _01584_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _53614_ (_02279_, _02278_, _02277_);
  or _53615_ (_02280_, _02279_, _01430_);
  and _53616_ (_02281_, _02280_, _43100_);
  and _53617_ (_02282_, _02170_, _36249_);
  or _53618_ (_02283_, _01544_, _01495_);
  not _53619_ (_02284_, _01545_);
  and _53620_ (_02285_, _02176_, _02284_);
  and _53621_ (_02286_, _02285_, _02283_);
  and _53622_ (_02287_, _01456_, _42740_);
  and _53623_ (_02288_, _01447_, _01490_);
  and _53624_ (_02289_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _53625_ (_02290_, _02289_, _02288_);
  or _53626_ (_02291_, _02290_, _02287_);
  nor _53627_ (_02292_, _02291_, _02286_);
  nand _53628_ (_02293_, _02292_, _01430_);
  or _53629_ (_02294_, _02293_, _02282_);
  and _53630_ (_39634_, _02294_, _02281_);
  and _53631_ (_02295_, _02170_, _30585_);
  or _53632_ (_02296_, _01487_, _01488_);
  or _53633_ (_02297_, _02296_, _01546_);
  nand _53634_ (_02298_, _02296_, _01546_);
  and _53635_ (_02299_, _02298_, _02176_);
  and _53636_ (_02300_, _02299_, _02297_);
  and _53637_ (_02301_, _01456_, _42517_);
  and _53638_ (_02302_, _01447_, _01484_);
  and _53639_ (_02303_, _38572_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _53640_ (_02304_, _02303_, _02302_);
  nor _53641_ (_02305_, _02304_, _02301_);
  nand _53642_ (_02306_, _02305_, _01430_);
  or _53643_ (_02307_, _02306_, _02300_);
  or _53644_ (_02308_, _02307_, _02295_);
  nor _53645_ (_02309_, _02278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _53646_ (_02310_, _02278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _53647_ (_02311_, _02310_, _02309_);
  or _53648_ (_02312_, _02311_, _01430_);
  and _53649_ (_02313_, _02312_, _43100_);
  and _53650_ (_39635_, _02313_, _02308_);
  nor _53651_ (_02314_, _01432_, _31808_);
  not _53652_ (_02315_, _38882_);
  and _53653_ (_02316_, _01435_, _02315_);
  and _53654_ (_02317_, _01548_, _38776_);
  nor _53655_ (_02318_, _01548_, _38776_);
  nor _53656_ (_02319_, _02318_, _02317_);
  nor _53657_ (_02320_, _02319_, _01486_);
  and _53658_ (_02321_, _02319_, _01486_);
  or _53659_ (_02322_, _02321_, _02320_);
  and _53660_ (_02323_, _02322_, _02176_);
  nand _53661_ (_02324_, _01447_, _42683_);
  and _53662_ (_02325_, _01456_, _00618_);
  and _53663_ (_02326_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _53664_ (_02327_, _02326_, _02325_);
  and _53665_ (_02328_, _02327_, _02324_);
  nand _53666_ (_02329_, _02328_, _01430_);
  or _53667_ (_02330_, _02329_, _02323_);
  or _53668_ (_02331_, _02330_, _02316_);
  or _53669_ (_02332_, _02331_, _02314_);
  or _53670_ (_02333_, _02310_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand _53671_ (_02334_, _01586_, _01584_);
  and _53672_ (_02335_, _02334_, _02333_);
  or _53673_ (_02336_, _02335_, _01430_);
  and _53674_ (_02337_, _02336_, _43100_);
  and _53675_ (_39636_, _02337_, _02332_);
  nor _53676_ (_02338_, _01432_, _32495_);
  and _53677_ (_02339_, _01548_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _53678_ (_02340_, _02339_, _01554_);
  and _53679_ (_02341_, _01555_, _01486_);
  nor _53680_ (_02342_, _02341_, _02340_);
  nand _53681_ (_02343_, _02342_, _38782_);
  or _53682_ (_02344_, _02342_, _38782_);
  and _53683_ (_02345_, _02344_, _02176_);
  and _53684_ (_02346_, _02345_, _02343_);
  not _53685_ (_02347_, _38916_);
  and _53686_ (_02348_, _01435_, _02347_);
  and _53687_ (_02349_, _01456_, _00673_);
  and _53688_ (_02350_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _53689_ (_02351_, _01447_, _42612_);
  or _53690_ (_02352_, _02351_, _02350_);
  or _53691_ (_02353_, _02352_, _02349_);
  nor _53692_ (_02354_, _02353_, _02348_);
  nand _53693_ (_02355_, _02354_, _01430_);
  or _53694_ (_02356_, _02355_, _02346_);
  or _53695_ (_02357_, _02356_, _02338_);
  nand _53696_ (_02358_, _02334_, _01677_);
  or _53697_ (_02360_, _02334_, _01677_);
  and _53698_ (_02361_, _02360_, _02358_);
  or _53699_ (_02362_, _02361_, _01430_);
  and _53700_ (_02363_, _02362_, _43100_);
  and _53701_ (_39637_, _02363_, _02357_);
  nor _53702_ (_02364_, _01432_, _33202_);
  and _53703_ (_02365_, _01556_, _01486_);
  and _53704_ (_02366_, _02340_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _53705_ (_02367_, _02366_, _02365_);
  nor _53706_ (_02368_, _02367_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _53707_ (_02369_, _02367_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _53708_ (_02370_, _02369_, _02368_);
  and _53709_ (_02371_, _02370_, _02176_);
  not _53710_ (_02372_, _38947_);
  and _53711_ (_02373_, _01435_, _02372_);
  and _53712_ (_02374_, _01456_, _00625_);
  and _53713_ (_02375_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _53714_ (_02376_, _01447_, _42804_);
  or _53715_ (_02377_, _02376_, _02375_);
  or _53716_ (_02378_, _02377_, _02374_);
  nor _53717_ (_02379_, _02378_, _02373_);
  nand _53718_ (_02380_, _02379_, _01430_);
  or _53719_ (_02381_, _02380_, _02371_);
  or _53720_ (_02382_, _02381_, _02364_);
  nor _53721_ (_02383_, _01588_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _53722_ (_02384_, _02383_, _01589_);
  or _53723_ (_02385_, _02384_, _01430_);
  and _53724_ (_02386_, _02385_, _43100_);
  and _53725_ (_39638_, _02386_, _02382_);
  nor _53726_ (_02387_, _01432_, _33953_);
  and _53727_ (_02388_, _01549_, _01554_);
  and _53728_ (_02389_, _01557_, _01486_);
  nor _53729_ (_02390_, _02389_, _02388_);
  nand _53730_ (_02391_, _02390_, _38772_);
  or _53731_ (_02392_, _02390_, _38772_);
  and _53732_ (_02393_, _02392_, _02176_);
  and _53733_ (_02394_, _02393_, _02391_);
  not _53734_ (_02395_, _38976_);
  and _53735_ (_02396_, _01435_, _02395_);
  and _53736_ (_02397_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _53737_ (_02398_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _53738_ (_02399_, _02398_, _01466_);
  and _53739_ (_02400_, _02399_, _01456_);
  and _53740_ (_02401_, _01447_, _42647_);
  or _53741_ (_02402_, _02401_, _02400_);
  or _53742_ (_02403_, _02402_, _02397_);
  nor _53743_ (_02404_, _02403_, _02396_);
  nand _53744_ (_02405_, _02404_, _01430_);
  or _53745_ (_02406_, _02405_, _02394_);
  or _53746_ (_02407_, _02406_, _02387_);
  nor _53747_ (_02408_, _01589_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _53748_ (_02409_, _02408_, _01590_);
  or _53749_ (_02410_, _02409_, _01430_);
  and _53750_ (_02411_, _02410_, _43100_);
  and _53751_ (_39639_, _02411_, _02407_);
  nor _53752_ (_02412_, _01432_, _34693_);
  and _53753_ (_02413_, _01550_, _01554_);
  and _53754_ (_02414_, _01558_, _01486_);
  nor _53755_ (_02415_, _02414_, _02413_);
  nand _53756_ (_02416_, _02415_, _38793_);
  or _53757_ (_02417_, _02415_, _38793_);
  and _53758_ (_02418_, _02417_, _02176_);
  and _53759_ (_02419_, _02418_, _02416_);
  not _53760_ (_02420_, _39007_);
  nand _53761_ (_02421_, _01435_, _02420_);
  nor _53762_ (_02422_, _01466_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _53763_ (_02423_, _02422_, _01467_);
  and _53764_ (_02424_, _02423_, _01456_);
  and _53765_ (_02425_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _53766_ (_02426_, _01447_, _42552_);
  or _53767_ (_02427_, _02426_, _02425_);
  nor _53768_ (_02428_, _02427_, _02424_);
  and _53769_ (_02429_, _02428_, _02421_);
  nand _53770_ (_02430_, _02429_, _01430_);
  or _53771_ (_02431_, _02430_, _02419_);
  or _53772_ (_02432_, _02431_, _02412_);
  nor _53773_ (_02433_, _01590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _53774_ (_02434_, _01590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _53775_ (_02435_, _02434_, _02433_);
  or _53776_ (_02436_, _02435_, _01430_);
  and _53777_ (_02437_, _02436_, _43100_);
  and _53778_ (_39640_, _02437_, _02432_);
  nor _53779_ (_02438_, _01432_, _35520_);
  and _53780_ (_02439_, _01551_, _01554_);
  and _53781_ (_02440_, _02414_, _38793_);
  nor _53782_ (_02441_, _02440_, _02439_);
  nand _53783_ (_02442_, _02441_, _38768_);
  or _53784_ (_02443_, _02441_, _38768_);
  and _53785_ (_02444_, _02443_, _02176_);
  and _53786_ (_02445_, _02444_, _02442_);
  not _53787_ (_02446_, _39041_);
  nand _53788_ (_02447_, _01435_, _02446_);
  nor _53789_ (_02448_, _01467_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _53790_ (_02449_, _02448_, _01468_);
  and _53791_ (_02450_, _02449_, _01456_);
  and _53792_ (_02451_, _01447_, _42778_);
  or _53793_ (_02452_, _02451_, _02450_);
  and _53794_ (_02453_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _53795_ (_02454_, _02453_, _02452_);
  and _53796_ (_02455_, _02454_, _02447_);
  nand _53797_ (_02456_, _02455_, _01430_);
  or _53798_ (_02457_, _02456_, _02445_);
  or _53799_ (_02458_, _02457_, _02438_);
  or _53800_ (_02459_, _02434_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand _53801_ (_02460_, _02434_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _53802_ (_02461_, _02460_, _02459_);
  or _53803_ (_02462_, _02461_, _01430_);
  and _53804_ (_02463_, _02462_, _43100_);
  and _53805_ (_39641_, _02463_, _02458_);
  nor _53806_ (_02464_, _01432_, _36239_);
  nor _53807_ (_02465_, _01562_, _38764_);
  and _53808_ (_02466_, _01562_, _38764_);
  or _53809_ (_02467_, _02466_, _02465_);
  and _53810_ (_02468_, _02467_, _02176_);
  not _53811_ (_02469_, _39071_);
  nand _53812_ (_02470_, _01435_, _02469_);
  nor _53813_ (_02471_, _01468_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _53814_ (_02472_, _02471_, _01469_);
  and _53815_ (_02473_, _02472_, _01456_);
  and _53816_ (_02474_, _01447_, _42740_);
  or _53817_ (_02475_, _02474_, _02473_);
  and _53818_ (_02476_, _01477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _53819_ (_02477_, _02476_, _02475_);
  and _53820_ (_02478_, _02477_, _02470_);
  nand _53821_ (_02479_, _02478_, _01430_);
  or _53822_ (_02480_, _02479_, _02468_);
  or _53823_ (_02481_, _02480_, _02464_);
  nor _53824_ (_02482_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _53825_ (_02483_, _02482_, _01592_);
  or _53826_ (_02484_, _02483_, _01430_);
  and _53827_ (_02485_, _02484_, _43100_);
  and _53828_ (_39642_, _02485_, _02481_);
  and _53829_ (_02486_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _53830_ (_02487_, _01813_, _01811_);
  nor _53831_ (_02488_, _02487_, _01814_);
  or _53832_ (_02489_, _02488_, _01602_);
  or _53833_ (_02490_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _53834_ (_02491_, _02490_, _01847_);
  and _53835_ (_02492_, _02491_, _02489_);
  or _53836_ (_39643_, _02492_, _02486_);
  nor _53837_ (_02493_, _01816_, _01814_);
  nor _53838_ (_02494_, _02493_, _01817_);
  or _53839_ (_02495_, _02494_, _01602_);
  or _53840_ (_02496_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _53841_ (_02497_, _02496_, _01847_);
  and _53842_ (_02498_, _02497_, _02495_);
  and _53843_ (_02499_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _53844_ (_39644_, _02499_, _02498_);
  or _53845_ (_02500_, _01821_, _01819_);
  nor _53846_ (_02501_, _01602_, _01822_);
  and _53847_ (_02502_, _02501_, _02500_);
  nor _53848_ (_02503_, _01601_, _01954_);
  or _53849_ (_02504_, _02503_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _53850_ (_02505_, _02504_, _02502_);
  or _53851_ (_02506_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _36477_);
  and _53852_ (_02507_, _02506_, _43100_);
  and _53853_ (_39645_, _02507_, _02505_);
  and _53854_ (_02508_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53855_ (_02509_, _01822_, _01700_);
  nor _53856_ (_02510_, _02509_, _01823_);
  or _53857_ (_02511_, _02510_, _01602_);
  or _53858_ (_02512_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _53859_ (_02513_, _02512_, _01847_);
  and _53860_ (_02514_, _02513_, _02511_);
  or _53861_ (_39647_, _02514_, _02508_);
  and _53862_ (_02515_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53863_ (_02516_, _01826_, _01823_);
  nor _53864_ (_02517_, _02516_, _01827_);
  or _53865_ (_02518_, _02517_, _01602_);
  or _53866_ (_02519_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _53867_ (_02520_, _02519_, _01847_);
  and _53868_ (_02521_, _02520_, _02518_);
  or _53869_ (_39648_, _02521_, _02515_);
  and _53870_ (_02522_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _53871_ (_02523_, _01827_, _01695_);
  nor _53872_ (_02524_, _02523_, _01828_);
  or _53873_ (_02525_, _02524_, _01602_);
  or _53874_ (_02526_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _53875_ (_02527_, _02526_, _01847_);
  and _53876_ (_02528_, _02527_, _02525_);
  or _53877_ (_39649_, _02528_, _02522_);
  nor _53878_ (_02529_, _01828_, _01691_);
  nor _53879_ (_02530_, _02529_, _01829_);
  or _53880_ (_02531_, _02530_, _01602_);
  or _53881_ (_02532_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _53882_ (_02533_, _02532_, _01847_);
  and _53883_ (_02534_, _02533_, _02531_);
  and _53884_ (_02535_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _53885_ (_39650_, _02535_, _02534_);
  nor _53886_ (_02536_, _01829_, _01688_);
  nor _53887_ (_02537_, _02536_, _01830_);
  or _53888_ (_02538_, _02537_, _01602_);
  or _53889_ (_02539_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _53890_ (_02540_, _02539_, _01847_);
  and _53891_ (_02541_, _02540_, _02538_);
  and _53892_ (_02542_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _53893_ (_39651_, _02542_, _02541_);
  and _53894_ (_02543_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _53895_ (_02544_, _01832_, _01830_);
  nor _53896_ (_02545_, _02544_, _01833_);
  or _53897_ (_02547_, _02545_, _01602_);
  or _53898_ (_02548_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _53899_ (_02549_, _02548_, _01847_);
  and _53900_ (_02550_, _02549_, _02547_);
  or _53901_ (_39652_, _02550_, _02543_);
  nor _53902_ (_02551_, _01833_, _01683_);
  nor _53903_ (_02552_, _02551_, _01834_);
  or _53904_ (_02553_, _02552_, _01602_);
  or _53905_ (_02554_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _53906_ (_02555_, _02554_, _01847_);
  and _53907_ (_02556_, _02555_, _02553_);
  and _53908_ (_02557_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _53909_ (_39653_, _02557_, _02556_);
  or _53910_ (_02558_, _01834_, _01676_);
  nor _53911_ (_02559_, _01602_, _01835_);
  and _53912_ (_02560_, _02559_, _02558_);
  nor _53913_ (_02561_, _01601_, _38787_);
  or _53914_ (_02562_, _02561_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _53915_ (_02563_, _02562_, _02560_);
  or _53916_ (_02564_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _36477_);
  and _53917_ (_02565_, _02564_, _43100_);
  and _53918_ (_39654_, _02565_, _02563_);
  nor _53919_ (_02566_, _01835_, _01673_);
  nor _53920_ (_02568_, _02566_, _01836_);
  or _53921_ (_02569_, _02568_, _01602_);
  or _53922_ (_02570_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _53923_ (_02571_, _02570_, _01847_);
  and _53924_ (_02572_, _02571_, _02569_);
  and _53925_ (_02573_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _53926_ (_39655_, _02573_, _02572_);
  and _53927_ (_02574_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _53928_ (_02575_, _01836_, _01668_);
  nor _53929_ (_02576_, _02575_, _01837_);
  or _53930_ (_02577_, _02576_, _01602_);
  or _53931_ (_02579_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _53932_ (_02580_, _02579_, _01847_);
  and _53933_ (_02581_, _02580_, _02577_);
  or _53934_ (_39656_, _02581_, _02574_);
  nor _53935_ (_02582_, _01837_, _01664_);
  nor _53936_ (_02583_, _02582_, _01838_);
  or _53937_ (_02584_, _02583_, _01602_);
  or _53938_ (_02585_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _53939_ (_02586_, _02585_, _01847_);
  and _53940_ (_02587_, _02586_, _02584_);
  and _53941_ (_02588_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _53942_ (_39658_, _02588_, _02587_);
  nor _53943_ (_02589_, _01838_, _01658_);
  nor _53944_ (_02590_, _02589_, _01839_);
  or _53945_ (_02591_, _02590_, _01602_);
  or _53946_ (_02592_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _53947_ (_02593_, _02592_, _01847_);
  and _53948_ (_02594_, _02593_, _02591_);
  and _53949_ (_02595_, _01598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _53950_ (_39659_, _02595_, _02594_);
  and _53951_ (_02596_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _53952_ (_02597_, _02596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _53953_ (_39660_, _02597_, _43100_);
  and _53954_ (_02598_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _53955_ (_02599_, _02598_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _53956_ (_39661_, _02599_, _43100_);
  and _53957_ (_02600_, _01858_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _53958_ (_02601_, _02600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _53959_ (_39662_, _02601_, _43100_);
  and _53960_ (_02602_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _53961_ (_02603_, _02602_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _53962_ (_39663_, _02603_, _43100_);
  and _53963_ (_02604_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _53964_ (_02605_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _53965_ (_39664_, _02605_, _43100_);
  and _53966_ (_02606_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _53967_ (_02607_, _02606_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _53968_ (_39665_, _02607_, _43100_);
  and _53969_ (_02608_, _01859_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _53970_ (_02609_, _02608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _53971_ (_39666_, _02609_, _43100_);
  nor _53972_ (_02610_, _01810_, _42500_);
  nand _53973_ (_02611_, _02610_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _53974_ (_02612_, _02610_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _53975_ (_02613_, _02612_, _01847_);
  and _53976_ (_39667_, _02613_, _02611_);
  nor _53977_ (_02614_, _01870_, _01868_);
  nor _53978_ (_02615_, _02614_, _01871_);
  or _53979_ (_02616_, _02615_, _42500_);
  or _53980_ (_02617_, _36509_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _53981_ (_02618_, _02617_, _01847_);
  and _53982_ (_39669_, _02618_, _02616_);
  and _53983_ (_02619_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _53984_ (_02620_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _53985_ (_02621_, _02620_, _39297_);
  or _53986_ (_39685_, _02621_, _02619_);
  and _53987_ (_02622_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _53988_ (_02623_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _53989_ (_02624_, _02623_, _39297_);
  or _53990_ (_39686_, _02624_, _02622_);
  and _53991_ (_02625_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _53992_ (_02626_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _53993_ (_02627_, _02626_, _39297_);
  or _53994_ (_39687_, _02627_, _02625_);
  and _53995_ (_02628_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _53996_ (_02629_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _53997_ (_02630_, _02629_, _39297_);
  or _53998_ (_39688_, _02630_, _02628_);
  and _53999_ (_02631_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _54000_ (_02632_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _54001_ (_02633_, _02632_, _39297_);
  or _54002_ (_39689_, _02633_, _02631_);
  and _54003_ (_02634_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _54004_ (_02635_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _54005_ (_02636_, _02635_, _39297_);
  or _54006_ (_39691_, _02636_, _02634_);
  and _54007_ (_02637_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _54008_ (_02638_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _54009_ (_02639_, _02638_, _39297_);
  or _54010_ (_39692_, _02639_, _02637_);
  and _54011_ (_39693_, _01899_, _43100_);
  nor _54012_ (_39694_, _01909_, rst);
  and _54013_ (_39695_, _01905_, _43100_);
  and _54014_ (_02640_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _54015_ (_02641_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or _54016_ (_02642_, _02641_, _02640_);
  and _54017_ (_39696_, _02642_, _43100_);
  and _54018_ (_02643_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _54019_ (_02644_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or _54020_ (_02645_, _02644_, _02643_);
  and _54021_ (_39697_, _02645_, _43100_);
  and _54022_ (_02646_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _54023_ (_02647_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or _54024_ (_02648_, _02647_, _02646_);
  and _54025_ (_39698_, _02648_, _43100_);
  and _54026_ (_02649_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _54027_ (_02650_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or _54028_ (_02651_, _02650_, _02649_);
  and _54029_ (_39699_, _02651_, _43100_);
  and _54030_ (_02652_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _54031_ (_02653_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or _54032_ (_02654_, _02653_, _02652_);
  and _54033_ (_39700_, _02654_, _43100_);
  and _54034_ (_02655_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _54035_ (_02656_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or _54036_ (_02657_, _02656_, _02655_);
  and _54037_ (_39702_, _02657_, _43100_);
  and _54038_ (_02658_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _54039_ (_02659_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or _54040_ (_02660_, _02659_, _02658_);
  and _54041_ (_39703_, _02660_, _43100_);
  and _54042_ (_02661_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _54043_ (_02662_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or _54044_ (_02663_, _02662_, _02661_);
  and _54045_ (_39704_, _02663_, _43100_);
  and _54046_ (_02664_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _54047_ (_02665_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or _54048_ (_02666_, _02665_, _02664_);
  and _54049_ (_39705_, _02666_, _43100_);
  and _54050_ (_02667_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _54051_ (_02668_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _54052_ (_02669_, _02668_, _02667_);
  and _54053_ (_39706_, _02669_, _43100_);
  and _54054_ (_02670_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _54055_ (_02671_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _54056_ (_02672_, _02671_, _02670_);
  and _54057_ (_39707_, _02672_, _43100_);
  and _54058_ (_02673_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _54059_ (_02674_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _54060_ (_02675_, _02674_, _02673_);
  and _54061_ (_39708_, _02675_, _43100_);
  and _54062_ (_02676_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _54063_ (_02677_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _54064_ (_02678_, _02677_, _02676_);
  and _54065_ (_39709_, _02678_, _43100_);
  and _54066_ (_02679_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _54067_ (_02680_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _54068_ (_02681_, _02680_, _02679_);
  and _54069_ (_39710_, _02681_, _43100_);
  and _54070_ (_02682_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _54071_ (_02683_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _54072_ (_02684_, _02683_, _02682_);
  and _54073_ (_39711_, _02684_, _43100_);
  and _54074_ (_02685_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _54075_ (_02686_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _54076_ (_02687_, _02686_, _02685_);
  and _54077_ (_39713_, _02687_, _43100_);
  and _54078_ (_02688_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _54079_ (_02689_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _54080_ (_02690_, _02689_, _02688_);
  and _54081_ (_39714_, _02690_, _43100_);
  and _54082_ (_02691_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _54083_ (_02692_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _54084_ (_02693_, _02692_, _02691_);
  and _54085_ (_39715_, _02693_, _43100_);
  and _54086_ (_02694_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _54087_ (_02695_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _54088_ (_02696_, _02695_, _02694_);
  and _54089_ (_39716_, _02696_, _43100_);
  and _54090_ (_02697_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _54091_ (_02698_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _54092_ (_02699_, _02698_, _02697_);
  and _54093_ (_39717_, _02699_, _43100_);
  and _54094_ (_02700_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _54095_ (_02701_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _54096_ (_02702_, _02701_, _02700_);
  and _54097_ (_39718_, _02702_, _43100_);
  and _54098_ (_02704_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _54099_ (_02705_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _54100_ (_02706_, _02705_, _02704_);
  and _54101_ (_39719_, _02706_, _43100_);
  and _54102_ (_02707_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _54103_ (_02708_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _54104_ (_02709_, _02708_, _02707_);
  and _54105_ (_39720_, _02709_, _43100_);
  and _54106_ (_02710_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _54107_ (_02711_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _54108_ (_02712_, _02711_, _02710_);
  and _54109_ (_39721_, _02712_, _43100_);
  and _54110_ (_02713_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _54111_ (_02714_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _54112_ (_02715_, _02714_, _02713_);
  and _54113_ (_39722_, _02715_, _43100_);
  and _54114_ (_02716_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _54115_ (_02717_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _54116_ (_02718_, _02717_, _02716_);
  and _54117_ (_39724_, _02718_, _43100_);
  and _54118_ (_02719_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _54119_ (_02720_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _54120_ (_02721_, _02720_, _02719_);
  and _54121_ (_39725_, _02721_, _43100_);
  and _54122_ (_02722_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _54123_ (_02723_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _54124_ (_02724_, _02723_, _02722_);
  and _54125_ (_39726_, _02724_, _43100_);
  and _54126_ (_02725_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _54127_ (_02726_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _54128_ (_02727_, _02726_, _02725_);
  and _54129_ (_39727_, _02727_, _43100_);
  and _54130_ (_02728_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _54131_ (_02729_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _54132_ (_02730_, _02729_, _02728_);
  and _54133_ (_39728_, _02730_, _43100_);
  and _54134_ (_02731_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _54135_ (_02732_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _54136_ (_02733_, _02732_, _02731_);
  and _54137_ (_39729_, _02733_, _43100_);
  and _54138_ (_02734_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54139_ (_02735_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _54140_ (_02736_, _02735_, _02734_);
  and _54141_ (_39730_, _02736_, _43100_);
  and _54142_ (_02737_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54143_ (_02738_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _54144_ (_02739_, _02738_, _02737_);
  and _54145_ (_39731_, _02739_, _43100_);
  and _54146_ (_02740_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54147_ (_02741_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _54148_ (_02742_, _02741_, _02740_);
  and _54149_ (_39732_, _02742_, _43100_);
  and _54150_ (_02743_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54151_ (_02744_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _54152_ (_02745_, _02744_, _02743_);
  and _54153_ (_39733_, _02745_, _43100_);
  and _54154_ (_02746_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54155_ (_02747_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _54156_ (_02748_, _02747_, _02746_);
  and _54157_ (_39735_, _02748_, _43100_);
  and _54158_ (_02749_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54159_ (_02750_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _54160_ (_02751_, _02750_, _02749_);
  and _54161_ (_39736_, _02751_, _43100_);
  and _54162_ (_02752_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54163_ (_02753_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _54164_ (_02754_, _02753_, _02752_);
  and _54165_ (_39737_, _02754_, _43100_);
  and _54166_ (_02755_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54167_ (_02756_, _42697_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54168_ (_02757_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _54169_ (_02758_, _02757_, _01922_);
  and _54170_ (_02759_, _02758_, _02756_);
  or _54171_ (_02760_, _02759_, _02755_);
  and _54172_ (_39738_, _02760_, _43100_);
  and _54173_ (_02761_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54174_ (_02762_, _42591_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54175_ (_02763_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _54176_ (_02764_, _02763_, _01922_);
  and _54177_ (_02765_, _02764_, _02762_);
  or _54178_ (_02766_, _02765_, _02761_);
  and _54179_ (_39739_, _02766_, _43100_);
  and _54180_ (_02767_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54181_ (_02768_, _42815_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54182_ (_02769_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _54183_ (_02770_, _02769_, _01922_);
  and _54184_ (_02771_, _02770_, _02768_);
  or _54185_ (_02772_, _02771_, _02767_);
  and _54186_ (_39740_, _02772_, _43100_);
  and _54187_ (_02773_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54188_ (_02774_, _42661_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54189_ (_02775_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _54190_ (_02776_, _02775_, _01922_);
  and _54191_ (_02777_, _02776_, _02774_);
  or _54192_ (_02778_, _02777_, _02773_);
  and _54193_ (_39741_, _02778_, _43100_);
  and _54194_ (_02779_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54195_ (_02780_, _42575_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54196_ (_02781_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _54197_ (_02782_, _02781_, _01922_);
  and _54198_ (_02783_, _02782_, _02780_);
  or _54199_ (_02784_, _02783_, _02779_);
  and _54200_ (_39742_, _02784_, _43100_);
  and _54201_ (_02785_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54202_ (_02786_, _42762_, _01929_);
  or _54203_ (_02787_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _54204_ (_02788_, _02787_, _01922_);
  and _54205_ (_02789_, _02788_, _02786_);
  or _54206_ (_02790_, _02789_, _02785_);
  and _54207_ (_39743_, _02790_, _43100_);
  and _54208_ (_02791_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54209_ (_02792_, _42720_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54210_ (_02793_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _54211_ (_02794_, _02793_, _01922_);
  and _54212_ (_02795_, _02794_, _02792_);
  or _54213_ (_02796_, _02795_, _02791_);
  and _54214_ (_39744_, _02796_, _43100_);
  and _54215_ (_02797_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54216_ (_02798_, _42495_, _01929_);
  or _54217_ (_02799_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _54218_ (_02800_, _02799_, _01922_);
  and _54219_ (_02801_, _02800_, _02798_);
  or _54220_ (_02803_, _02801_, _02797_);
  and _54221_ (_39746_, _02803_, _43100_);
  and _54222_ (_02804_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _54223_ (_02805_, _02804_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54224_ (_02806_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _01922_);
  and _54225_ (_02808_, _02806_, _43100_);
  and _54226_ (_39747_, _02808_, _02805_);
  and _54227_ (_02809_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _54228_ (_02810_, _02809_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54229_ (_02811_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _01922_);
  and _54230_ (_02813_, _02811_, _43100_);
  and _54231_ (_39748_, _02813_, _02810_);
  and _54232_ (_02814_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _54233_ (_02815_, _02814_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54234_ (_02816_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _01922_);
  and _54235_ (_02818_, _02816_, _43100_);
  and _54236_ (_39749_, _02818_, _02815_);
  and _54237_ (_02819_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _54238_ (_02820_, _02819_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54239_ (_02821_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _01922_);
  and _54240_ (_02823_, _02821_, _43100_);
  and _54241_ (_39750_, _02823_, _02820_);
  and _54242_ (_02824_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _54243_ (_02825_, _02824_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54244_ (_02826_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _01922_);
  and _54245_ (_02828_, _02826_, _43100_);
  and _54246_ (_39751_, _02828_, _02825_);
  and _54247_ (_02829_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _54248_ (_02830_, _02829_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54249_ (_02831_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _01922_);
  and _54250_ (_02833_, _02831_, _43100_);
  and _54251_ (_39752_, _02833_, _02830_);
  and _54252_ (_02835_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _54253_ (_02836_, _02835_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54254_ (_02837_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _01922_);
  and _54255_ (_02838_, _02837_, _43100_);
  and _54256_ (_39753_, _02838_, _02836_);
  nand _54257_ (_02840_, _01936_, _31808_);
  or _54258_ (_02841_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _54259_ (_02843_, _02841_, _43100_);
  and _54260_ (_39754_, _02843_, _02840_);
  nand _54261_ (_02844_, _01936_, _32495_);
  or _54262_ (_02846_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _54263_ (_02847_, _02846_, _43100_);
  and _54264_ (_39755_, _02847_, _02844_);
  nand _54265_ (_02849_, _01936_, _33202_);
  or _54266_ (_02850_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _54267_ (_02852_, _02850_, _43100_);
  and _54268_ (_39757_, _02852_, _02849_);
  nand _54269_ (_02854_, _01936_, _33953_);
  or _54270_ (_02855_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _54271_ (_02857_, _02855_, _43100_);
  and _54272_ (_39758_, _02857_, _02854_);
  nand _54273_ (_02858_, _01936_, _34693_);
  or _54274_ (_02860_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _54275_ (_02861_, _02860_, _43100_);
  and _54276_ (_39759_, _02861_, _02858_);
  nand _54277_ (_02863_, _01936_, _35520_);
  or _54278_ (_02864_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _54279_ (_02866_, _02864_, _43100_);
  and _54280_ (_39760_, _02866_, _02863_);
  nand _54281_ (_02867_, _01936_, _36239_);
  or _54282_ (_02868_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _54283_ (_02869_, _02868_, _43100_);
  and _54284_ (_39761_, _02869_, _02867_);
  nand _54285_ (_02870_, _01936_, _30574_);
  or _54286_ (_02872_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _54287_ (_02874_, _02872_, _43100_);
  and _54288_ (_39762_, _02874_, _02870_);
  nand _54289_ (_02876_, _01936_, _38882_);
  or _54290_ (_02877_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _54291_ (_02878_, _02877_, _43100_);
  and _54292_ (_39763_, _02878_, _02876_);
  nand _54293_ (_02880_, _01936_, _38916_);
  or _54294_ (_02881_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _54295_ (_02883_, _02881_, _43100_);
  and _54296_ (_39764_, _02883_, _02880_);
  nand _54297_ (_02885_, _01936_, _38947_);
  or _54298_ (_02887_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _54299_ (_02888_, _02887_, _43100_);
  and _54300_ (_39765_, _02888_, _02885_);
  nand _54301_ (_02890_, _01936_, _38976_);
  or _54302_ (_02891_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _54303_ (_02892_, _02891_, _43100_);
  and _54304_ (_39766_, _02892_, _02890_);
  nand _54305_ (_02894_, _01936_, _39007_);
  or _54306_ (_02896_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _54307_ (_02898_, _02896_, _43100_);
  and _54308_ (_39768_, _02898_, _02894_);
  nand _54309_ (_02899_, _01936_, _39041_);
  or _54310_ (_02900_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _54311_ (_02902_, _02900_, _43100_);
  and _54312_ (_39769_, _02902_, _02899_);
  nand _54313_ (_02903_, _01936_, _39071_);
  or _54314_ (_02905_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _54315_ (_02906_, _02905_, _43100_);
  and _54316_ (_39770_, _02906_, _02903_);
  nor _54317_ (_39980_, _42534_, rst);
  and _54318_ (_02908_, _39237_, _27496_);
  and _54319_ (_02909_, _02908_, _42467_);
  nand _54320_ (_02911_, _02909_, _38704_);
  or _54321_ (_02912_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _54322_ (_02913_, _02912_, _43100_);
  and _54323_ (_39981_, _02913_, _02911_);
  and _54324_ (_02915_, _39497_, _27496_);
  not _54325_ (_02916_, _02915_);
  nor _54326_ (_02918_, _02916_, _38704_);
  not _54327_ (_02920_, _42467_);
  and _54328_ (_02921_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _54329_ (_02923_, _02921_, _02920_);
  or _54330_ (_02924_, _02923_, _02918_);
  or _54331_ (_02926_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _54332_ (_02927_, _02926_, _43100_);
  and _54333_ (_39982_, _02927_, _02924_);
  and _54334_ (_02928_, _27003_, _27661_);
  and _54335_ (_02929_, _02928_, _27496_);
  not _54336_ (_02930_, _02929_);
  nor _54337_ (_02932_, _02930_, _38704_);
  and _54338_ (_02934_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or _54339_ (_02935_, _02934_, _02920_);
  or _54340_ (_02936_, _02935_, _02932_);
  or _54341_ (_02938_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _54342_ (_02939_, _02938_, _43100_);
  and _54343_ (_39983_, _02939_, _02936_);
  and _54344_ (_02941_, _41582_, _27496_);
  not _54345_ (_02942_, _02941_);
  nor _54346_ (_02943_, _02942_, _38704_);
  and _54347_ (_02946_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _54348_ (_02947_, _02946_, _02920_);
  or _54349_ (_02948_, _02947_, _02943_);
  or _54350_ (_02950_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _54351_ (_02951_, _02950_, _43100_);
  and _54352_ (_39985_, _02951_, _02948_);
  nand _54353_ (_02953_, _02909_, _38682_);
  or _54354_ (_02954_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _54355_ (_02955_, _02954_, _43100_);
  and _54356_ (_40013_, _02955_, _02953_);
  nand _54357_ (_02958_, _02909_, _38672_);
  or _54358_ (_02960_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _54359_ (_02961_, _02960_, _43100_);
  and _54360_ (_40014_, _02961_, _02958_);
  nand _54361_ (_02962_, _02909_, _38665_);
  or _54362_ (_02964_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _54363_ (_02965_, _02964_, _43100_);
  and _54364_ (_40015_, _02965_, _02962_);
  nand _54365_ (_02967_, _02909_, _38658_);
  or _54366_ (_02968_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _54367_ (_02970_, _02968_, _43100_);
  and _54368_ (_40016_, _02970_, _02967_);
  nand _54369_ (_02972_, _02909_, _38650_);
  or _54370_ (_02973_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _54371_ (_02975_, _02973_, _43100_);
  and _54372_ (_40017_, _02975_, _02972_);
  nand _54373_ (_02976_, _02909_, _38642_);
  or _54374_ (_02978_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _54375_ (_02979_, _02978_, _43100_);
  and _54376_ (_40018_, _02979_, _02976_);
  nand _54377_ (_02982_, _02909_, _38635_);
  or _54378_ (_02983_, _02909_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _54379_ (_02984_, _02983_, _43100_);
  and _54380_ (_40019_, _02984_, _02982_);
  nor _54381_ (_02986_, _02916_, _38682_);
  and _54382_ (_02988_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or _54383_ (_02989_, _02988_, _02920_);
  or _54384_ (_02990_, _02989_, _02986_);
  or _54385_ (_02991_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _54386_ (_02993_, _02991_, _43100_);
  and _54387_ (_40021_, _02993_, _02990_);
  nor _54388_ (_02995_, _02916_, _38672_);
  and _54389_ (_02997_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _54390_ (_02998_, _02997_, _02920_);
  or _54391_ (_02999_, _02998_, _02995_);
  or _54392_ (_03001_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _54393_ (_03002_, _03001_, _43100_);
  and _54394_ (_40022_, _03002_, _02999_);
  nor _54395_ (_03004_, _02916_, _38665_);
  and _54396_ (_03005_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _54397_ (_03007_, _03005_, _02920_);
  or _54398_ (_03009_, _03007_, _03004_);
  or _54399_ (_03010_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _54400_ (_03011_, _03010_, _43100_);
  and _54401_ (_40023_, _03011_, _03009_);
  nor _54402_ (_03013_, _02916_, _38658_);
  and _54403_ (_03014_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _54404_ (_03016_, _03014_, _02920_);
  or _54405_ (_03017_, _03016_, _03013_);
  or _54406_ (_03019_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _54407_ (_03021_, _03019_, _43100_);
  and _54408_ (_40024_, _03021_, _03017_);
  nor _54409_ (_03022_, _02916_, _38650_);
  and _54410_ (_03024_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _54411_ (_03025_, _03024_, _02920_);
  or _54412_ (_03026_, _03025_, _03022_);
  or _54413_ (_03028_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _54414_ (_03029_, _03028_, _43100_);
  and _54415_ (_40025_, _03029_, _03026_);
  nor _54416_ (_03031_, _02916_, _38642_);
  and _54417_ (_03032_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _54418_ (_03033_, _03032_, _02920_);
  or _54419_ (_03035_, _03033_, _03031_);
  or _54420_ (_03036_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _54421_ (_03037_, _03036_, _43100_);
  and _54422_ (_40026_, _03037_, _03035_);
  nor _54423_ (_03039_, _02916_, _38635_);
  and _54424_ (_03040_, _02916_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _54425_ (_03042_, _03040_, _02920_);
  or _54426_ (_03043_, _03042_, _03039_);
  or _54427_ (_03044_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _54428_ (_03046_, _03044_, _43100_);
  and _54429_ (_40027_, _03046_, _03043_);
  or _54430_ (_03048_, _02929_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand _54431_ (_03049_, _02929_, _38682_);
  and _54432_ (_03050_, _03049_, _03048_);
  or _54433_ (_03051_, _03050_, _02920_);
  or _54434_ (_03052_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _54435_ (_03053_, _03052_, _43100_);
  and _54436_ (_40028_, _03053_, _03051_);
  nor _54437_ (_03055_, _02930_, _38672_);
  and _54438_ (_03056_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or _54439_ (_03057_, _03056_, _02920_);
  or _54440_ (_03059_, _03057_, _03055_);
  or _54441_ (_03060_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _54442_ (_03061_, _03060_, _43100_);
  and _54443_ (_40029_, _03061_, _03059_);
  nor _54444_ (_03063_, _02930_, _38665_);
  and _54445_ (_03064_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or _54446_ (_03066_, _03064_, _02920_);
  or _54447_ (_03067_, _03066_, _03063_);
  or _54448_ (_03068_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _54449_ (_03070_, _03068_, _43100_);
  and _54450_ (_40030_, _03070_, _03067_);
  not _54451_ (_03071_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _54452_ (_03073_, _02929_, _42467_);
  nor _54453_ (_03074_, _03073_, _03071_);
  and _54454_ (_03075_, _03073_, _40346_);
  or _54455_ (_03077_, _03075_, _03074_);
  and _54456_ (_40032_, _03077_, _43100_);
  nor _54457_ (_03079_, _02930_, _38650_);
  and _54458_ (_03080_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or _54459_ (_03081_, _03080_, _02920_);
  or _54460_ (_03082_, _03081_, _03079_);
  or _54461_ (_03084_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _54462_ (_03085_, _03084_, _43100_);
  and _54463_ (_40033_, _03085_, _03082_);
  nor _54464_ (_03087_, _02930_, _38642_);
  and _54465_ (_03088_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _54466_ (_03089_, _03088_, _02920_);
  or _54467_ (_03091_, _03089_, _03087_);
  or _54468_ (_03092_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _54469_ (_03093_, _03092_, _43100_);
  and _54470_ (_40034_, _03093_, _03091_);
  nor _54471_ (_03095_, _02930_, _38635_);
  and _54472_ (_03096_, _02930_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _54473_ (_03098_, _03096_, _02920_);
  or _54474_ (_03099_, _03098_, _03095_);
  or _54475_ (_03100_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _54476_ (_03102_, _03100_, _43100_);
  and _54477_ (_40035_, _03102_, _03099_);
  and _54478_ (_03103_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _54479_ (_03105_, _02942_, _38682_);
  or _54480_ (_03106_, _03105_, _02920_);
  or _54481_ (_03108_, _03106_, _03103_);
  or _54482_ (_03109_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _54483_ (_03110_, _03109_, _43100_);
  and _54484_ (_40036_, _03110_, _03108_);
  nor _54485_ (_03112_, _02942_, _38672_);
  and _54486_ (_03113_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _54487_ (_03114_, _03113_, _02920_);
  or _54488_ (_03116_, _03114_, _03112_);
  or _54489_ (_03117_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _54490_ (_03118_, _03117_, _43100_);
  and _54491_ (_40037_, _03118_, _03116_);
  nor _54492_ (_03120_, _02942_, _38665_);
  and _54493_ (_03121_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or _54494_ (_03123_, _03121_, _02920_);
  or _54495_ (_03124_, _03123_, _03120_);
  or _54496_ (_03125_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _54497_ (_03128_, _03125_, _43100_);
  and _54498_ (_40038_, _03128_, _03124_);
  nor _54499_ (_03129_, _02942_, _38658_);
  and _54500_ (_03131_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _54501_ (_03132_, _03131_, _02920_);
  or _54502_ (_03133_, _03132_, _03129_);
  or _54503_ (_03135_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _54504_ (_03136_, _03135_, _43100_);
  and _54505_ (_40039_, _03136_, _03133_);
  nor _54506_ (_03138_, _02942_, _38650_);
  and _54507_ (_03139_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or _54508_ (_03140_, _03139_, _02920_);
  or _54509_ (_03142_, _03140_, _03138_);
  or _54510_ (_03143_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _54511_ (_03144_, _03143_, _43100_);
  and _54512_ (_40040_, _03144_, _03142_);
  nor _54513_ (_03146_, _02942_, _38642_);
  and _54514_ (_03147_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or _54515_ (_03149_, _03147_, _02920_);
  or _54516_ (_03150_, _03149_, _03146_);
  or _54517_ (_03151_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _54518_ (_03153_, _03151_, _43100_);
  and _54519_ (_40041_, _03153_, _03150_);
  nor _54520_ (_03154_, _02942_, _38635_);
  and _54521_ (_03156_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _54522_ (_03157_, _03156_, _02920_);
  or _54523_ (_03158_, _03157_, _03154_);
  or _54524_ (_03160_, _42467_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _54525_ (_03161_, _03160_, _43100_);
  and _54526_ (_40043_, _03161_, _03158_);
  not _54527_ (_03163_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _54528_ (_03164_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _54529_ (_03166_, _03164_, _03163_);
  and _54530_ (_03167_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _43100_);
  and _54531_ (_40070_, _03167_, _03166_);
  nor _54532_ (_03168_, _03166_, rst);
  nand _54533_ (_03169_, _03164_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _54534_ (_03171_, _03164_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _54535_ (_03172_, _03171_, _03169_);
  and _54536_ (_40072_, _03172_, _03168_);
  nor _54537_ (_03174_, _42743_, _42787_);
  not _54538_ (_03175_, _42521_);
  and _54539_ (_03176_, _42579_, _03175_);
  and _54540_ (_03178_, _03176_, _03174_);
  and _54541_ (_03179_, _03178_, _42665_);
  and _54542_ (_03180_, _03179_, _39236_);
  nor _54543_ (_03182_, _03180_, _01344_);
  nor _54544_ (_03183_, _42743_, _42788_);
  nor _54545_ (_03184_, _42666_, _42579_);
  and _54546_ (_03186_, _03184_, _03175_);
  and _54547_ (_03187_, _03186_, _03183_);
  not _54548_ (_03188_, _42823_);
  nor _54549_ (_03190_, _39326_, _39314_);
  and _54550_ (_03191_, _39326_, _39314_);
  nor _54551_ (_03192_, _03191_, _03190_);
  nor _54552_ (_03194_, _39383_, _39338_);
  and _54553_ (_03195_, _39383_, _39338_);
  nor _54554_ (_03197_, _03195_, _03194_);
  nor _54555_ (_03198_, _03197_, _03192_);
  and _54556_ (_03199_, _03197_, _03192_);
  or _54557_ (_03200_, _03199_, _03198_);
  and _54558_ (_03202_, _39407_, _39395_);
  nor _54559_ (_03203_, _39407_, _39395_);
  nor _54560_ (_03204_, _03203_, _03202_);
  nor _54561_ (_03206_, _39419_, _39260_);
  and _54562_ (_03207_, _39419_, _39260_);
  nor _54563_ (_03208_, _03207_, _03206_);
  or _54564_ (_03210_, _03208_, _03204_);
  nand _54565_ (_03211_, _03208_, _03204_);
  and _54566_ (_03212_, _03211_, _03210_);
  nor _54567_ (_03214_, _03212_, _03200_);
  and _54568_ (_03215_, _03212_, _03200_);
  nor _54569_ (_03216_, _03215_, _03214_);
  or _54570_ (_03218_, _03216_, _03188_);
  and _54571_ (_03219_, _42701_, _42617_);
  or _54572_ (_03220_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _54573_ (_03222_, _03220_, _03219_);
  and _54574_ (_03223_, _03222_, _03218_);
  nor _54575_ (_03224_, _42701_, _42617_);
  and _54576_ (_03226_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not _54577_ (_03227_, _42701_);
  and _54578_ (_03229_, _03227_, _42617_);
  and _54579_ (_03230_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _54580_ (_03231_, _03230_, _03226_);
  and _54581_ (_03232_, _03231_, _03188_);
  or _54582_ (_03234_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _54583_ (_03235_, _03227_, _42617_);
  or _54584_ (_03236_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _54585_ (_03238_, _03236_, _03235_);
  and _54586_ (_03239_, _03238_, _03234_);
  and _54587_ (_03240_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _54588_ (_03242_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _54589_ (_03243_, _03242_, _03240_);
  and _54590_ (_03244_, _03243_, _42823_);
  or _54591_ (_03246_, _03244_, _03239_);
  or _54592_ (_03247_, _03246_, _03232_);
  or _54593_ (_03248_, _03247_, _03223_);
  and _54594_ (_03250_, _03248_, _03187_);
  nor _54595_ (_03251_, _03187_, _28636_);
  and _54596_ (_03252_, _42743_, _03175_);
  nand _54597_ (_03254_, _03252_, _42666_);
  not _54598_ (_03255_, _03183_);
  nand _54599_ (_03256_, _03186_, _03255_);
  and _54600_ (_03258_, _03256_, _03254_);
  and _54601_ (_03259_, _03258_, _03251_);
  and _54602_ (_03261_, _03176_, _42666_);
  and _54603_ (_03262_, _03261_, _03183_);
  nor _54604_ (_03263_, _03262_, _03179_);
  and _54605_ (_03264_, _42743_, _42787_);
  and _54606_ (_03266_, _03264_, _03176_);
  and _54607_ (_03267_, _03266_, _42665_);
  and _54608_ (_03268_, _42743_, _42788_);
  and _54609_ (_03270_, _03268_, _03176_);
  and _54610_ (_03271_, _03270_, _42665_);
  nor _54611_ (_03272_, _03271_, _03267_);
  and _54612_ (_03274_, _03272_, _03263_);
  and _54613_ (_03275_, _03274_, _03259_);
  and _54614_ (_03276_, _01425_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  nor _54615_ (_03278_, _00818_, _38521_);
  and _54616_ (_03279_, _38443_, _38488_);
  nor _54617_ (_03280_, _03279_, _00933_);
  and _54618_ (_03282_, _03280_, _03278_);
  not _54619_ (_03283_, _38515_);
  nor _54620_ (_03284_, _00913_, _38509_);
  and _54621_ (_03286_, _03284_, _03283_);
  and _54622_ (_03287_, _03286_, _00820_);
  and _54623_ (_03288_, _03287_, _03282_);
  and _54624_ (_03290_, _01091_, _00753_);
  and _54625_ (_03291_, _03290_, _03288_);
  and _54626_ (_03292_, _03291_, _38546_);
  nor _54627_ (_03293_, _03292_, _36466_);
  or _54628_ (_03294_, _03293_, p2_in[5]);
  not _54629_ (_03295_, _03293_);
  or _54630_ (_03296_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _54631_ (_03297_, _03296_, _03294_);
  and _54632_ (_03298_, _03297_, _03188_);
  or _54633_ (_03299_, _03293_, p2_in[1]);
  or _54634_ (_03300_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _54635_ (_03301_, _03300_, _03299_);
  and _54636_ (_03302_, _03301_, _42823_);
  or _54637_ (_03303_, _03302_, _03298_);
  and _54638_ (_03304_, _03303_, _03229_);
  or _54639_ (_03305_, _03293_, p2_in[2]);
  or _54640_ (_03306_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _54641_ (_03307_, _03306_, _03305_);
  or _54642_ (_03308_, _03307_, _03188_);
  or _54643_ (_03309_, _03293_, p2_in[6]);
  or _54644_ (_03310_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _54645_ (_03311_, _03310_, _03309_);
  or _54646_ (_03312_, _03311_, _42823_);
  and _54647_ (_03313_, _03312_, _03235_);
  and _54648_ (_03314_, _03313_, _03308_);
  or _54649_ (_03315_, _03293_, p2_in[4]);
  or _54650_ (_03316_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _54651_ (_03317_, _03316_, _03315_);
  and _54652_ (_03318_, _03317_, _03188_);
  nor _54653_ (_03319_, _03293_, p2_in[0]);
  and _54654_ (_03320_, _03293_, _39860_);
  nor _54655_ (_03321_, _03320_, _03319_);
  and _54656_ (_03322_, _03321_, _42823_);
  or _54657_ (_03323_, _03322_, _03318_);
  and _54658_ (_03324_, _03323_, _03219_);
  or _54659_ (_03325_, _03293_, p2_in[3]);
  or _54660_ (_03326_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _54661_ (_03327_, _03326_, _03325_);
  or _54662_ (_03328_, _03327_, _03188_);
  or _54663_ (_03329_, _03293_, p2_in[7]);
  or _54664_ (_03330_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _54665_ (_03331_, _03330_, _03329_);
  or _54666_ (_03332_, _03331_, _42823_);
  and _54667_ (_03333_, _03332_, _03224_);
  and _54668_ (_03334_, _03333_, _03328_);
  or _54669_ (_03335_, _03334_, _03324_);
  or _54670_ (_03336_, _03335_, _03314_);
  or _54671_ (_03337_, _03336_, _03304_);
  and _54672_ (_03338_, _03337_, _03271_);
  and _54673_ (_03339_, _03219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _54674_ (_03340_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _54675_ (_03341_, _03340_, _03339_);
  and _54676_ (_03342_, _03235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _54677_ (_03343_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _54678_ (_03344_, _03343_, _03342_);
  or _54679_ (_03345_, _03344_, _03341_);
  and _54680_ (_03346_, _03345_, _03188_);
  and _54681_ (_03347_, _03219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _54682_ (_03348_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _54683_ (_03349_, _03348_, _03347_);
  and _54684_ (_03350_, _03235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _54685_ (_03351_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _54686_ (_03352_, _03351_, _03350_);
  or _54687_ (_03353_, _03352_, _03349_);
  and _54688_ (_03354_, _03353_, _42823_);
  or _54689_ (_03355_, _03354_, _03346_);
  and _54690_ (_03356_, _03355_, _03262_);
  or _54691_ (_03357_, _03356_, _03338_);
  or _54692_ (_03358_, _03357_, _03276_);
  or _54693_ (_03359_, _03358_, _03275_);
  nor _54694_ (_03360_, _42823_, _40899_);
  and _54695_ (_03361_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _54696_ (_03362_, _03361_, _03360_);
  and _54697_ (_03364_, _03362_, _03219_);
  or _54698_ (_03365_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _54699_ (_03366_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _54700_ (_03367_, _03366_, _03224_);
  and _54701_ (_03368_, _03367_, _03365_);
  or _54702_ (_03369_, _03368_, _03364_);
  and _54703_ (_03370_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _54704_ (_03371_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _54705_ (_03372_, _03371_, _03370_);
  and _54706_ (_03373_, _03372_, _03235_);
  or _54707_ (_03374_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _54708_ (_03375_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _54709_ (_03376_, _03375_, _03229_);
  and _54710_ (_03377_, _03376_, _03374_);
  or _54711_ (_03378_, _03377_, _03373_);
  or _54712_ (_03379_, _03378_, _03369_);
  and _54713_ (_03380_, _03379_, _03268_);
  and _54714_ (_03381_, _03219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _54715_ (_03382_, _03235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _54716_ (_03383_, _03382_, _03381_);
  and _54717_ (_03384_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _54718_ (_03385_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _54719_ (_03386_, _03385_, _03384_);
  or _54720_ (_03387_, _03386_, _03383_);
  and _54721_ (_03388_, _03387_, _42823_);
  and _54722_ (_03389_, _03219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _54723_ (_03390_, _03235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _54724_ (_03391_, _03390_, _03389_);
  and _54725_ (_03392_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _54726_ (_03393_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _54727_ (_03394_, _03393_, _03392_);
  or _54728_ (_03395_, _03394_, _03391_);
  and _54729_ (_03396_, _03395_, _03188_);
  or _54730_ (_03397_, _03396_, _03388_);
  and _54731_ (_03398_, _03397_, _03264_);
  or _54732_ (_03399_, _03398_, _03380_);
  and _54733_ (_03400_, _03399_, _03261_);
  and _54734_ (_03401_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _54735_ (_03402_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _54736_ (_03403_, _03402_, _03401_);
  and _54737_ (_03404_, _03403_, _03188_);
  and _54738_ (_03405_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _54739_ (_03406_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _54740_ (_03407_, _03406_, _03405_);
  and _54741_ (_03408_, _03407_, _03219_);
  and _54742_ (_03409_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _54743_ (_03410_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _54744_ (_03411_, _03410_, _03409_);
  and _54745_ (_03412_, _03411_, _03235_);
  or _54746_ (_03413_, _03412_, _03408_);
  and _54747_ (_03414_, _03224_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _54748_ (_03415_, _03229_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _54749_ (_03416_, _03415_, _03414_);
  and _54750_ (_03417_, _03416_, _42823_);
  or _54751_ (_03418_, _03417_, _03413_);
  or _54752_ (_03419_, _03418_, _03404_);
  and _54753_ (_03420_, _03419_, _03179_);
  or _54754_ (_03421_, _42665_, _42521_);
  nor _54755_ (_03422_, _03421_, _42579_);
  and _54756_ (_03423_, _03422_, _03264_);
  nor _54757_ (_03424_, _42823_, _41473_);
  and _54758_ (_03425_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _54759_ (_03426_, _03425_, _03424_);
  and _54760_ (_03427_, _03426_, _03224_);
  or _54761_ (_03428_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand _54762_ (_03429_, _42823_, _41490_);
  and _54763_ (_03430_, _03429_, _03219_);
  and _54764_ (_03431_, _03430_, _03428_);
  or _54765_ (_03432_, _03431_, _03427_);
  nor _54766_ (_03433_, _42823_, _41899_);
  and _54767_ (_03434_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _54768_ (_03435_, _03434_, _03433_);
  and _54769_ (_03436_, _03435_, _03229_);
  nand _54770_ (_03437_, _42823_, _41924_);
  or _54771_ (_03438_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _54772_ (_03439_, _03438_, _03235_);
  and _54773_ (_03440_, _03439_, _03437_);
  or _54774_ (_03441_, _03440_, _03436_);
  or _54775_ (_03442_, _03441_, _03432_);
  and _54776_ (_03443_, _03442_, _03423_);
  or _54777_ (_03444_, _03293_, p0_in[5]);
  or _54778_ (_03445_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _54779_ (_03446_, _03445_, _03444_);
  and _54780_ (_03447_, _03446_, _03188_);
  or _54781_ (_03448_, _03293_, p0_in[1]);
  or _54782_ (_03449_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _54783_ (_03450_, _03449_, _03448_);
  and _54784_ (_03451_, _03450_, _42823_);
  or _54785_ (_03452_, _03451_, _03447_);
  and _54786_ (_03453_, _03452_, _03229_);
  or _54787_ (_03454_, _03293_, p0_in[2]);
  nand _54788_ (_03455_, _03293_, _39510_);
  and _54789_ (_03456_, _03455_, _03454_);
  or _54790_ (_03457_, _03456_, _03188_);
  or _54791_ (_03458_, _03293_, p0_in[6]);
  or _54792_ (_03459_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _54793_ (_03460_, _03459_, _03458_);
  or _54794_ (_03461_, _03460_, _42823_);
  and _54795_ (_03462_, _03461_, _03235_);
  and _54796_ (_03463_, _03462_, _03457_);
  or _54797_ (_03464_, _03293_, p0_in[4]);
  or _54798_ (_03465_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _54799_ (_03466_, _03465_, _03464_);
  and _54800_ (_03467_, _03466_, _03188_);
  nor _54801_ (_03468_, _03293_, p0_in[0]);
  and _54802_ (_03469_, _03293_, _39493_);
  nor _54803_ (_03470_, _03469_, _03468_);
  and _54804_ (_03471_, _03470_, _42823_);
  or _54805_ (_03472_, _03471_, _03467_);
  and _54806_ (_03473_, _03472_, _03219_);
  or _54807_ (_03474_, _03293_, p0_in[3]);
  or _54808_ (_03475_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _54809_ (_03476_, _03475_, _03474_);
  or _54810_ (_03477_, _03476_, _03188_);
  or _54811_ (_03478_, _03293_, p0_in[7]);
  or _54812_ (_03479_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _54813_ (_03480_, _03479_, _03478_);
  or _54814_ (_03481_, _03480_, _42823_);
  and _54815_ (_03482_, _03481_, _03224_);
  and _54816_ (_03483_, _03482_, _03477_);
  or _54817_ (_03484_, _03483_, _03473_);
  or _54818_ (_03485_, _03484_, _03463_);
  or _54819_ (_03486_, _03485_, _03453_);
  and _54820_ (_03487_, _03486_, _03267_);
  or _54821_ (_03488_, _03487_, _03443_);
  or _54822_ (_03489_, _03488_, _03420_);
  or _54823_ (_03490_, _03489_, _03400_);
  and _54824_ (_03491_, _03188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _54825_ (_03492_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _54826_ (_03493_, _03492_, _03491_);
  and _54827_ (_03494_, _03493_, _03224_);
  or _54828_ (_03495_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nand _54829_ (_03496_, _42823_, _40918_);
  and _54830_ (_03497_, _03496_, _03219_);
  and _54831_ (_03498_, _03497_, _03495_);
  or _54832_ (_03499_, _03498_, _03494_);
  nor _54833_ (_03500_, _42823_, _40930_);
  and _54834_ (_03501_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _54835_ (_03502_, _03501_, _03500_);
  and _54836_ (_03503_, _03502_, _03229_);
  nand _54837_ (_03504_, _42823_, _40923_);
  or _54838_ (_03505_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _54839_ (_03506_, _03505_, _03235_);
  and _54840_ (_03507_, _03506_, _03504_);
  or _54841_ (_03508_, _03507_, _03503_);
  or _54842_ (_03509_, _03508_, _03499_);
  and _54843_ (_03510_, _03509_, _03422_);
  or _54844_ (_03511_, _03293_, p3_in[7]);
  or _54845_ (_03512_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _54846_ (_03513_, _03512_, _03511_);
  and _54847_ (_03514_, _03513_, _03188_);
  or _54848_ (_03515_, _03293_, p3_in[3]);
  or _54849_ (_03516_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _54850_ (_03517_, _03516_, _03515_);
  and _54851_ (_03518_, _03517_, _42823_);
  or _54852_ (_03519_, _03518_, _03514_);
  and _54853_ (_03520_, _03519_, _03224_);
  nor _54854_ (_03521_, _03293_, p3_in[0]);
  and _54855_ (_03522_, _03293_, _39947_);
  nor _54856_ (_03523_, _03522_, _03521_);
  or _54857_ (_03524_, _03523_, _03188_);
  or _54858_ (_03525_, _03293_, p3_in[4]);
  or _54859_ (_03526_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _54860_ (_03527_, _03526_, _03525_);
  or _54861_ (_03528_, _03527_, _42823_);
  and _54862_ (_03529_, _03528_, _03219_);
  and _54863_ (_03530_, _03529_, _03524_);
  or _54864_ (_03531_, _03530_, _03520_);
  or _54865_ (_03532_, _03293_, p3_in[6]);
  or _54866_ (_03533_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _54867_ (_03534_, _03533_, _03532_);
  and _54868_ (_03535_, _03534_, _03188_);
  or _54869_ (_03536_, _03293_, p3_in[2]);
  or _54870_ (_03537_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _54871_ (_03538_, _03537_, _03536_);
  and _54872_ (_03539_, _03538_, _42823_);
  or _54873_ (_03540_, _03539_, _03535_);
  and _54874_ (_03541_, _03540_, _03235_);
  or _54875_ (_03542_, _03293_, p3_in[1]);
  or _54876_ (_03543_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _54877_ (_03544_, _03543_, _03542_);
  or _54878_ (_03545_, _03544_, _03188_);
  or _54879_ (_03546_, _03293_, p3_in[5]);
  or _54880_ (_03547_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _54881_ (_03548_, _03547_, _03546_);
  or _54882_ (_03549_, _03548_, _42823_);
  and _54883_ (_03550_, _03549_, _03229_);
  and _54884_ (_03551_, _03550_, _03545_);
  or _54885_ (_03552_, _03551_, _03541_);
  or _54886_ (_03553_, _03552_, _03531_);
  and _54887_ (_03554_, _03553_, _03186_);
  or _54888_ (_03555_, _03554_, _03510_);
  and _54889_ (_03556_, _03555_, _03268_);
  nor _54890_ (_03557_, _42823_, _30661_);
  and _54891_ (_03558_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _54892_ (_03559_, _03558_, _03557_);
  and _54893_ (_03560_, _03559_, _03224_);
  or _54894_ (_03561_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _54895_ (_03562_, _42823_, _31831_);
  and _54896_ (_03563_, _03562_, _03219_);
  and _54897_ (_03565_, _03563_, _03561_);
  or _54898_ (_03566_, _03565_, _03560_);
  nor _54899_ (_03567_, _42823_, _35553_);
  and _54900_ (_03568_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _54901_ (_03569_, _03568_, _03567_);
  and _54902_ (_03570_, _03569_, _03229_);
  nand _54903_ (_03571_, _42823_, _33235_);
  or _54904_ (_03572_, _42823_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _54905_ (_03573_, _03572_, _03235_);
  and _54906_ (_03574_, _03573_, _03571_);
  or _54907_ (_03575_, _03574_, _03570_);
  or _54908_ (_03576_, _03575_, _03566_);
  and _54909_ (_03577_, _03576_, _03174_);
  or _54910_ (_03578_, _03293_, p1_in[5]);
  or _54911_ (_03579_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _54912_ (_03580_, _03579_, _03578_);
  and _54913_ (_03581_, _03580_, _03188_);
  or _54914_ (_03582_, _03293_, p1_in[1]);
  or _54915_ (_03583_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _54916_ (_03584_, _03583_, _03582_);
  and _54917_ (_03585_, _03584_, _42823_);
  or _54918_ (_03586_, _03585_, _03581_);
  and _54919_ (_03587_, _03586_, _03229_);
  or _54920_ (_03588_, _03293_, p1_in[2]);
  or _54921_ (_03589_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _54922_ (_03590_, _03589_, _03588_);
  or _54923_ (_03591_, _03590_, _03188_);
  or _54924_ (_03592_, _03293_, p1_in[6]);
  or _54925_ (_03593_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _54926_ (_03594_, _03593_, _03592_);
  or _54927_ (_03595_, _03594_, _42823_);
  and _54928_ (_03596_, _03595_, _03235_);
  and _54929_ (_03597_, _03596_, _03591_);
  or _54930_ (_03598_, _03293_, p1_in[4]);
  or _54931_ (_03599_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _54932_ (_03600_, _03599_, _03598_);
  and _54933_ (_03601_, _03600_, _03188_);
  nor _54934_ (_03602_, _03293_, p1_in[0]);
  and _54935_ (_03603_, _03293_, _39779_);
  nor _54936_ (_03604_, _03603_, _03602_);
  and _54937_ (_03605_, _03604_, _42823_);
  or _54938_ (_03606_, _03605_, _03601_);
  and _54939_ (_03607_, _03606_, _03219_);
  or _54940_ (_03608_, _03293_, p1_in[3]);
  or _54941_ (_03609_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _54942_ (_03610_, _03609_, _03608_);
  or _54943_ (_03611_, _03610_, _03188_);
  or _54944_ (_03612_, _03293_, p1_in[7]);
  or _54945_ (_03613_, _03295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _54946_ (_03614_, _03613_, _03612_);
  or _54947_ (_03615_, _03614_, _42823_);
  and _54948_ (_03616_, _03615_, _03224_);
  and _54949_ (_03617_, _03616_, _03611_);
  or _54950_ (_03618_, _03617_, _03607_);
  or _54951_ (_03619_, _03618_, _03597_);
  or _54952_ (_03620_, _03619_, _03587_);
  and _54953_ (_03621_, _03620_, _03264_);
  or _54954_ (_03622_, _03621_, _03577_);
  and _54955_ (_03623_, _03622_, _03186_);
  or _54956_ (_03624_, _03623_, _03556_);
  or _54957_ (_03625_, _03624_, _03490_);
  or _54958_ (_03626_, _03625_, _03359_);
  or _54959_ (_03627_, _03626_, _03250_);
  nand _54960_ (_03628_, _03276_, _31265_);
  nand _54961_ (_03629_, _03628_, _03627_);
  nand _54962_ (_03630_, _03629_, _03182_);
  and _54963_ (_03631_, _03219_, _38683_);
  or _54964_ (_03632_, _03631_, _03188_);
  and _54965_ (_03633_, _03224_, _40346_);
  and _54966_ (_03634_, _03229_, _41428_);
  and _54967_ (_03635_, _03235_, _40334_);
  or _54968_ (_03636_, _03635_, _03634_);
  or _54969_ (_03637_, _03636_, _03633_);
  or _54970_ (_03638_, _03637_, _03632_);
  and _54971_ (_03639_, _03219_, _40357_);
  or _54972_ (_03640_, _03639_, _42823_);
  and _54973_ (_03641_, _03224_, _40145_);
  and _54974_ (_03642_, _03229_, _40370_);
  and _54975_ (_03643_, _03235_, _40383_);
  or _54976_ (_03644_, _03643_, _03642_);
  or _54977_ (_03645_, _03644_, _03641_);
  or _54978_ (_03646_, _03645_, _03640_);
  and _54979_ (_03647_, _03646_, _03638_);
  or _54980_ (_03648_, _03647_, _03182_);
  and _54981_ (_03649_, _03648_, _43100_);
  and _54982_ (_40073_, _03649_, _03630_);
  and _54983_ (_03650_, _42665_, _42823_);
  and _54984_ (_03651_, _03650_, _03219_);
  and _54985_ (_03652_, _03651_, _03178_);
  and _54986_ (_03653_, _03652_, _39231_);
  nor _54987_ (_03654_, _42788_, _42579_);
  nor _54988_ (_03655_, _42743_, _42521_);
  and _54989_ (_03656_, _03651_, _03655_);
  and _54990_ (_03657_, _03656_, _03654_);
  and _54991_ (_03658_, _03657_, _39106_);
  nor _54992_ (_03659_, _03658_, _03653_);
  and _54993_ (_03660_, _03650_, _03224_);
  and _54994_ (_03661_, _03660_, _03266_);
  nand _54995_ (_03662_, _03661_, _38755_);
  and _54996_ (_03663_, _03662_, _03659_);
  nor _54997_ (_03664_, _03663_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _54998_ (_03665_, _03664_);
  and _54999_ (_03666_, _03652_, _39236_);
  not _55000_ (_03667_, _39247_);
  and _55001_ (_03668_, _03224_, _03188_);
  nor _55002_ (_03669_, _03668_, _03667_);
  and _55003_ (_03670_, _03669_, _01342_);
  nor _55004_ (_03671_, _03670_, _03666_);
  and _55005_ (_03672_, _03671_, _01428_);
  and _55006_ (_03673_, _03672_, _03665_);
  and _55007_ (_03674_, _03266_, _03235_);
  and _55008_ (_03675_, _03674_, _03650_);
  and _55009_ (_03676_, _03675_, _38755_);
  or _55010_ (_03677_, _03676_, rst);
  nor _55011_ (_40074_, _03677_, _03673_);
  nand _55012_ (_03678_, _03676_, _30574_);
  and _55013_ (_03679_, _03183_, _03176_);
  nor _55014_ (_03680_, _42665_, _42823_);
  and _55015_ (_03681_, _03680_, _03219_);
  and _55016_ (_03682_, _03681_, _03679_);
  and _55017_ (_03683_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _55018_ (_03684_, _42666_, _42823_);
  and _55019_ (_03685_, _03684_, _03219_);
  and _55020_ (_03686_, _03685_, _03679_);
  and _55021_ (_03687_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _55022_ (_03688_, _03687_, _03683_);
  and _55023_ (_03689_, _03684_, _03235_);
  and _55024_ (_03690_, _03689_, _03679_);
  and _55025_ (_03691_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _55026_ (_03692_, _03680_, _03229_);
  and _55027_ (_03693_, _03692_, _03679_);
  and _55028_ (_03694_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _55029_ (_03695_, _03694_, _03691_);
  or _55030_ (_03696_, _03695_, _03688_);
  and _55031_ (_03697_, _03684_, _03224_);
  and _55032_ (_03698_, _03697_, _03679_);
  and _55033_ (_03699_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _55034_ (_03700_, _03685_, _03266_);
  and _55035_ (_03701_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _55036_ (_03702_, _03701_, _03699_);
  and _55037_ (_03703_, _03685_, _03270_);
  and _55038_ (_03704_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _55039_ (_03705_, _03668_, _42665_);
  nor _55040_ (_03706_, _42787_, _42579_);
  and _55041_ (_03707_, _03706_, _03252_);
  and _55042_ (_03708_, _03707_, _03705_);
  and _55043_ (_03709_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _55044_ (_03710_, _03709_, _03704_);
  or _55045_ (_03711_, _03710_, _03702_);
  or _55046_ (_03712_, _03711_, _03696_);
  and _55047_ (_03713_, _03684_, _03229_);
  and _55048_ (_03714_, _03713_, _03266_);
  and _55049_ (_03715_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _55050_ (_03716_, _03697_, _03266_);
  and _55051_ (_03717_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or _55052_ (_03718_, _03717_, _03715_);
  and _55053_ (_03719_, _03692_, _03266_);
  and _55054_ (_03720_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _55055_ (_03721_, _03689_, _03266_);
  and _55056_ (_03722_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _55057_ (_03723_, _03722_, _03720_);
  or _55058_ (_03724_, _03723_, _03718_);
  and _55059_ (_03725_, _03654_, _03252_);
  and _55060_ (_03726_, _03725_, _03713_);
  and _55061_ (_03727_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _55062_ (_03728_, _03725_, _03685_);
  and _55063_ (_03729_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _55064_ (_03730_, _03729_, _03727_);
  and _55065_ (_03731_, _03681_, _03266_);
  and _55066_ (_03732_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _55067_ (_03733_, _03668_, _03267_);
  and _55068_ (_03734_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _55069_ (_03735_, _03734_, _03732_);
  or _55070_ (_03736_, _03735_, _03730_);
  or _55071_ (_03737_, _03736_, _03724_);
  or _55072_ (_03738_, _03737_, _03712_);
  and _55073_ (_03739_, _03266_, _03229_);
  and _55074_ (_03740_, _03739_, _03650_);
  and _55075_ (_03741_, _03740_, _38706_);
  and _55076_ (_03742_, _03706_, _03656_);
  and _55077_ (_03743_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _55078_ (_03744_, _03743_, _03741_);
  and _55079_ (_03745_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _55080_ (_03746_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _55081_ (_03747_, _03746_, _03745_);
  or _55082_ (_03748_, _03747_, _03744_);
  and _55083_ (_03749_, _03651_, _03270_);
  and _55084_ (_03750_, _03749_, _03331_);
  and _55085_ (_03751_, _03707_, _03651_);
  and _55086_ (_03752_, _03751_, _03513_);
  or _55087_ (_03753_, _03752_, _03750_);
  and _55088_ (_03754_, _03651_, _03266_);
  and _55089_ (_03755_, _03754_, _03480_);
  and _55090_ (_03756_, _03725_, _03651_);
  and _55091_ (_03757_, _03756_, _03614_);
  or _55092_ (_03758_, _03757_, _03755_);
  or _55093_ (_03759_, _03758_, _03753_);
  or _55094_ (_03760_, _03759_, _03748_);
  and _55095_ (_03761_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _55096_ (_03762_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _55097_ (_03764_, _03762_, _03761_);
  or _55098_ (_03765_, _03764_, _03760_);
  or _55099_ (_03766_, _03765_, _03738_);
  and _55100_ (_03767_, _03651_, _03252_);
  or _55101_ (_03768_, _03742_, _03767_);
  or _55102_ (_03769_, _03768_, _03740_);
  and _55103_ (_03770_, _03266_, _03224_);
  nand _55104_ (_03771_, _03684_, _03770_);
  nor _55105_ (_03772_, _03726_, _03731_);
  nor _55106_ (_03773_, _03719_, _03728_);
  and _55107_ (_03774_, _03773_, _03772_);
  nand _55108_ (_03775_, _03774_, _03771_);
  or _55109_ (_03776_, _03775_, _03769_);
  or _55110_ (_03777_, _03708_, _03652_);
  or _55111_ (_03778_, _03733_, _03657_);
  or _55112_ (_03779_, _03778_, _03777_);
  and _55113_ (_03780_, _03770_, _03650_);
  or _55114_ (_03781_, _03698_, _03690_);
  or _55115_ (_03782_, _03693_, _03700_);
  or _55116_ (_03783_, _03782_, _03781_);
  or _55117_ (_03784_, _03783_, _03780_);
  or _55118_ (_03785_, _03784_, _03779_);
  nand _55119_ (_03786_, _03684_, _03674_);
  nor _55120_ (_03787_, _03703_, _03714_);
  nand _55121_ (_03788_, _03787_, _03786_);
  and _55122_ (_03789_, _03262_, _03219_);
  or _55123_ (_03790_, _03789_, _03675_);
  or _55124_ (_03791_, _03790_, _03788_);
  or _55125_ (_03792_, _03791_, _03785_);
  or _55126_ (_03793_, _03792_, _03776_);
  nand _55127_ (_03794_, _03793_, _03673_);
  and _55128_ (_03795_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _55129_ (_03796_, _03795_, _03766_);
  or _55130_ (_03797_, _03673_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _55131_ (_03798_, _03797_, _03796_);
  or _55132_ (_03799_, _03798_, _03676_);
  and _55133_ (_03800_, _03799_, _43100_);
  and _55134_ (_40075_, _03800_, _03678_);
  nor _55135_ (_40156_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _55136_ (_03801_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _55137_ (_03802_, _03164_, rst);
  and _55138_ (_40157_, _03802_, _03801_);
  nor _55139_ (_03803_, _03164_, _03163_);
  or _55140_ (_03804_, _03803_, _03166_);
  and _55141_ (_03805_, _03169_, _43100_);
  and _55142_ (_40158_, _03805_, _03804_);
  not _55143_ (_03806_, _03673_);
  nand _55144_ (_03807_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _55145_ (_03808_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _55146_ (_03809_, _03808_, _03807_);
  nand _55147_ (_03810_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _55148_ (_03811_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _55149_ (_03812_, _03811_, _03810_);
  and _55150_ (_03813_, _03812_, _03809_);
  nand _55151_ (_03814_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand _55152_ (_03815_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _55153_ (_03816_, _03815_, _03814_);
  nand _55154_ (_03817_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _55155_ (_03818_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _55156_ (_03819_, _03818_, _03817_);
  and _55157_ (_03820_, _03819_, _03816_);
  and _55158_ (_03821_, _03820_, _03813_);
  nand _55159_ (_03822_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _55160_ (_03823_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _55161_ (_03824_, _03823_, _03822_);
  nand _55162_ (_03825_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _55163_ (_03826_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _55164_ (_03827_, _03826_, _03825_);
  and _55165_ (_03828_, _03827_, _03824_);
  nand _55166_ (_03829_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand _55167_ (_03830_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _55168_ (_03831_, _03830_, _03829_);
  nand _55169_ (_03832_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _55170_ (_03833_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _55171_ (_03834_, _03833_, _03832_);
  and _55172_ (_03835_, _03834_, _03831_);
  and _55173_ (_03836_, _03835_, _03828_);
  and _55174_ (_03837_, _03836_, _03821_);
  nand _55175_ (_03838_, _03740_, _42686_);
  nand _55176_ (_03839_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _55177_ (_03840_, _03839_, _03838_);
  nand _55178_ (_03841_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _55179_ (_03842_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _55180_ (_03843_, _03842_, _03841_);
  and _55181_ (_03844_, _03843_, _03840_);
  nand _55182_ (_03845_, _03749_, _03321_);
  nand _55183_ (_03846_, _03751_, _03523_);
  and _55184_ (_03847_, _03846_, _03845_);
  nand _55185_ (_03848_, _03756_, _03604_);
  nand _55186_ (_03849_, _03754_, _03470_);
  and _55187_ (_03850_, _03849_, _03848_);
  and _55188_ (_03851_, _03850_, _03847_);
  and _55189_ (_03852_, _03851_, _03844_);
  nand _55190_ (_03853_, _03657_, _03216_);
  nand _55191_ (_03854_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _55192_ (_03855_, _03854_, _03853_);
  and _55193_ (_03856_, _03855_, _03852_);
  and _55194_ (_03857_, _03856_, _03837_);
  nor _55195_ (_03858_, _03857_, _03806_);
  and _55196_ (_03859_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or _55197_ (_03860_, _03859_, _03676_);
  or _55198_ (_03861_, _03860_, _03858_);
  nand _55199_ (_03862_, _03676_, _31808_);
  and _55200_ (_03863_, _03862_, _43100_);
  and _55201_ (_40159_, _03863_, _03861_);
  nand _55202_ (_03864_, _03676_, _32495_);
  and _55203_ (_03865_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _55204_ (_03866_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _55205_ (_03867_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _55206_ (_03868_, _03867_, _03866_);
  and _55207_ (_03869_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _55208_ (_03870_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _55209_ (_03871_, _03870_, _03869_);
  or _55210_ (_03872_, _03871_, _03868_);
  and _55211_ (_03873_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _55212_ (_03874_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _55213_ (_03875_, _03874_, _03873_);
  and _55214_ (_03876_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _55215_ (_03877_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _55216_ (_03878_, _03877_, _03876_);
  or _55217_ (_03879_, _03878_, _03875_);
  or _55218_ (_03880_, _03879_, _03872_);
  and _55219_ (_03881_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _55220_ (_03882_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _55221_ (_03883_, _03882_, _03881_);
  and _55222_ (_03884_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _55223_ (_03885_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _55224_ (_03886_, _03885_, _03884_);
  or _55225_ (_03887_, _03886_, _03883_);
  and _55226_ (_03888_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _55227_ (_03889_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _55228_ (_03890_, _03889_, _03888_);
  and _55229_ (_03891_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _55230_ (_03892_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _55231_ (_03893_, _03892_, _03891_);
  or _55232_ (_03894_, _03893_, _03890_);
  or _55233_ (_03895_, _03894_, _03887_);
  or _55234_ (_03896_, _03895_, _03880_);
  and _55235_ (_03897_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _55236_ (_03898_, _03740_, _42595_);
  or _55237_ (_03899_, _03898_, _03897_);
  and _55238_ (_03900_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _55239_ (_03901_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _55240_ (_03902_, _03901_, _03900_);
  or _55241_ (_03903_, _03902_, _03899_);
  and _55242_ (_03904_, _03749_, _03301_);
  and _55243_ (_03905_, _03751_, _03544_);
  or _55244_ (_03906_, _03905_, _03904_);
  and _55245_ (_03907_, _03756_, _03584_);
  and _55246_ (_03908_, _03754_, _03450_);
  or _55247_ (_03909_, _03908_, _03907_);
  or _55248_ (_03910_, _03909_, _03906_);
  or _55249_ (_03911_, _03910_, _03903_);
  and _55250_ (_03912_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _55251_ (_03913_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _55252_ (_03914_, _03913_, _03912_);
  or _55253_ (_03915_, _03914_, _03911_);
  or _55254_ (_03916_, _03915_, _03896_);
  and _55255_ (_03917_, _03916_, _03673_);
  or _55256_ (_03918_, _03917_, _03865_);
  or _55257_ (_03919_, _03918_, _03676_);
  and _55258_ (_03920_, _03919_, _43100_);
  and _55259_ (_40161_, _03920_, _03864_);
  nand _55260_ (_03921_, _03676_, _33202_);
  and _55261_ (_03922_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _55262_ (_03923_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _55263_ (_03924_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _55264_ (_03925_, _03924_, _03923_);
  and _55265_ (_03926_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _55266_ (_03927_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _55267_ (_03928_, _03927_, _03926_);
  or _55268_ (_03929_, _03928_, _03925_);
  and _55269_ (_03930_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _55270_ (_03931_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _55271_ (_03932_, _03931_, _03930_);
  and _55272_ (_03933_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _55273_ (_03934_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _55274_ (_03935_, _03934_, _03933_);
  or _55275_ (_03936_, _03935_, _03932_);
  or _55276_ (_03937_, _03936_, _03929_);
  and _55277_ (_03938_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _55278_ (_03939_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _55279_ (_03940_, _03939_, _03938_);
  and _55280_ (_03941_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _55281_ (_03942_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _55282_ (_03943_, _03942_, _03941_);
  or _55283_ (_03944_, _03943_, _03940_);
  and _55284_ (_03945_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _55285_ (_03946_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _55286_ (_03947_, _03946_, _03945_);
  and _55287_ (_03948_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _55288_ (_03949_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _55289_ (_03950_, _03949_, _03948_);
  or _55290_ (_03951_, _03950_, _03947_);
  or _55291_ (_03952_, _03951_, _03944_);
  or _55292_ (_03953_, _03952_, _03937_);
  and _55293_ (_03954_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _55294_ (_03955_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _55295_ (_03956_, _03955_, _03954_);
  and _55296_ (_03957_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _55297_ (_03959_, _03740_, _42819_);
  or _55298_ (_03960_, _03959_, _03957_);
  and _55299_ (_03961_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _55300_ (_03962_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _55301_ (_03963_, _03962_, _03961_);
  or _55302_ (_03964_, _03963_, _03960_);
  and _55303_ (_03965_, _03749_, _03307_);
  and _55304_ (_03966_, _03751_, _03538_);
  or _55305_ (_03967_, _03966_, _03965_);
  and _55306_ (_03968_, _03754_, _03456_);
  and _55307_ (_03969_, _03756_, _03590_);
  or _55308_ (_03970_, _03969_, _03968_);
  or _55309_ (_03971_, _03970_, _03967_);
  or _55310_ (_03972_, _03971_, _03964_);
  or _55311_ (_03973_, _03972_, _03956_);
  or _55312_ (_03974_, _03973_, _03953_);
  and _55313_ (_03975_, _03974_, _03673_);
  or _55314_ (_03976_, _03975_, _03922_);
  or _55315_ (_03977_, _03976_, _03676_);
  and _55316_ (_03978_, _03977_, _43100_);
  and _55317_ (_40162_, _03978_, _03921_);
  nand _55318_ (_03979_, _03676_, _33953_);
  and _55319_ (_03980_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _55320_ (_03981_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _55321_ (_03982_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _55322_ (_03983_, _03982_, _03981_);
  and _55323_ (_03984_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _55324_ (_03985_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _55325_ (_03986_, _03985_, _03984_);
  or _55326_ (_03987_, _03986_, _03983_);
  and _55327_ (_03988_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _55328_ (_03989_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _55329_ (_03990_, _03989_, _03988_);
  and _55330_ (_03991_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _55331_ (_03992_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _55332_ (_03993_, _03992_, _03991_);
  or _55333_ (_03994_, _03993_, _03990_);
  or _55334_ (_03995_, _03994_, _03987_);
  and _55335_ (_03996_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _55336_ (_03997_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _55337_ (_03998_, _03997_, _03996_);
  and _55338_ (_03999_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _55339_ (_04000_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _55340_ (_04001_, _04000_, _03999_);
  or _55341_ (_04002_, _04001_, _03998_);
  and _55342_ (_04003_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _55343_ (_04004_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _55344_ (_04005_, _04004_, _04003_);
  and _55345_ (_04006_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _55346_ (_04007_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _55347_ (_04008_, _04007_, _04006_);
  or _55348_ (_04009_, _04008_, _04005_);
  or _55349_ (_04010_, _04009_, _04002_);
  or _55350_ (_04011_, _04010_, _03995_);
  and _55351_ (_04012_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _55352_ (_04013_, _03740_, _42650_);
  or _55353_ (_04014_, _04013_, _04012_);
  and _55354_ (_04015_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _55355_ (_04016_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _55356_ (_04017_, _04016_, _04015_);
  or _55357_ (_04018_, _04017_, _04014_);
  and _55358_ (_04019_, _03749_, _03327_);
  and _55359_ (_04020_, _03751_, _03517_);
  or _55360_ (_04021_, _04020_, _04019_);
  and _55361_ (_04022_, _03756_, _03610_);
  and _55362_ (_04023_, _03754_, _03476_);
  or _55363_ (_04024_, _04023_, _04022_);
  or _55364_ (_04025_, _04024_, _04021_);
  or _55365_ (_04026_, _04025_, _04018_);
  and _55366_ (_04027_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _55367_ (_04028_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _55368_ (_04029_, _04028_, _04027_);
  or _55369_ (_04030_, _04029_, _04026_);
  or _55370_ (_04031_, _04030_, _04011_);
  and _55371_ (_04032_, _04031_, _03673_);
  or _55372_ (_04033_, _04032_, _03980_);
  or _55373_ (_04034_, _04033_, _03676_);
  and _55374_ (_04035_, _04034_, _43100_);
  and _55375_ (_40163_, _04035_, _03979_);
  nand _55376_ (_04036_, _03676_, _34693_);
  and _55377_ (_04037_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _55378_ (_04038_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _55379_ (_04039_, _04038_, _04037_);
  and _55380_ (_04040_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _55381_ (_04041_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _55382_ (_04042_, _04041_, _04040_);
  or _55383_ (_04043_, _04042_, _04039_);
  and _55384_ (_04044_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _55385_ (_04045_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _55386_ (_04046_, _04045_, _04044_);
  and _55387_ (_04047_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _55388_ (_04048_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _55389_ (_04049_, _04048_, _04047_);
  or _55390_ (_04050_, _04049_, _04046_);
  or _55391_ (_04051_, _04050_, _04043_);
  and _55392_ (_04052_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _55393_ (_04053_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _55394_ (_04054_, _04053_, _04052_);
  and _55395_ (_04055_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _55396_ (_04056_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _55397_ (_04058_, _04056_, _04055_);
  or _55398_ (_04059_, _04058_, _04054_);
  and _55399_ (_04060_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and _55400_ (_04061_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _55401_ (_04062_, _04061_, _04060_);
  and _55402_ (_04063_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _55403_ (_04064_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _55404_ (_04065_, _04064_, _04063_);
  or _55405_ (_04066_, _04065_, _04062_);
  or _55406_ (_04067_, _04066_, _04059_);
  or _55407_ (_04068_, _04067_, _04051_);
  and _55408_ (_04069_, _03740_, _42563_);
  and _55409_ (_04070_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _55410_ (_04071_, _04070_, _04069_);
  and _55411_ (_04072_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _55412_ (_04073_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _55413_ (_04074_, _04073_, _04072_);
  or _55414_ (_04075_, _04074_, _04071_);
  and _55415_ (_04076_, _03749_, _03317_);
  and _55416_ (_04077_, _03751_, _03527_);
  or _55417_ (_04078_, _04077_, _04076_);
  and _55418_ (_04079_, _03756_, _03600_);
  and _55419_ (_04080_, _03754_, _03466_);
  or _55420_ (_04081_, _04080_, _04079_);
  or _55421_ (_04082_, _04081_, _04078_);
  or _55422_ (_04083_, _04082_, _04075_);
  and _55423_ (_04084_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _55424_ (_04085_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _55425_ (_04086_, _04085_, _04084_);
  or _55426_ (_04087_, _04086_, _04083_);
  or _55427_ (_04088_, _04087_, _04068_);
  and _55428_ (_04089_, _04088_, _03673_);
  and _55429_ (_04090_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or _55430_ (_04091_, _04090_, _03676_);
  or _55431_ (_04092_, _04091_, _04089_);
  and _55432_ (_04093_, _04092_, _43100_);
  and _55433_ (_40164_, _04093_, _04036_);
  nand _55434_ (_04094_, _03676_, _35520_);
  and _55435_ (_04095_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _55436_ (_04096_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _55437_ (_04097_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _55438_ (_04098_, _04097_, _04096_);
  and _55439_ (_04099_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _55440_ (_04100_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _55441_ (_04101_, _04100_, _04099_);
  or _55442_ (_04102_, _04101_, _04098_);
  and _55443_ (_04103_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _55444_ (_04104_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _55445_ (_04105_, _04104_, _04103_);
  and _55446_ (_04106_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _55447_ (_04107_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _55448_ (_04108_, _04107_, _04106_);
  or _55449_ (_04109_, _04108_, _04105_);
  or _55450_ (_04110_, _04109_, _04102_);
  and _55451_ (_04111_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _55452_ (_04112_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _55453_ (_04113_, _04112_, _04111_);
  and _55454_ (_04114_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _55455_ (_04115_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _55456_ (_04116_, _04115_, _04114_);
  or _55457_ (_04117_, _04116_, _04113_);
  and _55458_ (_04118_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _55459_ (_04119_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _55460_ (_04120_, _04119_, _04118_);
  and _55461_ (_04121_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _55462_ (_04122_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _55463_ (_04123_, _04122_, _04121_);
  or _55464_ (_04124_, _04123_, _04120_);
  or _55465_ (_04125_, _04124_, _04117_);
  or _55466_ (_04126_, _04125_, _04110_);
  and _55467_ (_04127_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not _55468_ (_04128_, _38744_);
  and _55469_ (_04129_, _03740_, _04128_);
  or _55470_ (_04130_, _04129_, _04127_);
  and _55471_ (_04131_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _55472_ (_04132_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _55473_ (_04133_, _04132_, _04131_);
  or _55474_ (_04134_, _04133_, _04130_);
  and _55475_ (_04135_, _03749_, _03297_);
  and _55476_ (_04136_, _03751_, _03548_);
  or _55477_ (_04137_, _04136_, _04135_);
  and _55478_ (_04138_, _03756_, _03580_);
  and _55479_ (_04139_, _03754_, _03446_);
  or _55480_ (_04140_, _04139_, _04138_);
  or _55481_ (_04141_, _04140_, _04137_);
  or _55482_ (_04142_, _04141_, _04134_);
  and _55483_ (_04143_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _55484_ (_04144_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _55485_ (_04145_, _04144_, _04143_);
  or _55486_ (_04146_, _04145_, _04142_);
  or _55487_ (_04147_, _04146_, _04126_);
  and _55488_ (_04148_, _04147_, _03673_);
  or _55489_ (_04149_, _04148_, _04095_);
  or _55490_ (_04150_, _04149_, _03676_);
  and _55491_ (_04151_, _04150_, _43100_);
  and _55492_ (_40165_, _04151_, _04094_);
  nand _55493_ (_04152_, _03676_, _36239_);
  and _55494_ (_04153_, _03682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _55495_ (_04154_, _03686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _55496_ (_04155_, _04154_, _04153_);
  and _55497_ (_04157_, _03690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _55498_ (_04158_, _03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _55499_ (_04159_, _04158_, _04157_);
  or _55500_ (_04160_, _04159_, _04155_);
  and _55501_ (_04161_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _55502_ (_04162_, _03698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _55503_ (_04163_, _04162_, _04161_);
  and _55504_ (_04164_, _03703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _55505_ (_04165_, _03708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _55506_ (_04166_, _04165_, _04164_);
  or _55507_ (_04167_, _04166_, _04163_);
  or _55508_ (_04168_, _04167_, _04160_);
  and _55509_ (_04169_, _03714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _55510_ (_04170_, _03716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _55511_ (_04171_, _04170_, _04169_);
  and _55512_ (_04172_, _03719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _55513_ (_04173_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _55514_ (_04174_, _04173_, _04172_);
  or _55515_ (_04175_, _04174_, _04171_);
  and _55516_ (_04176_, _03728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _55517_ (_04177_, _03726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or _55518_ (_04178_, _04177_, _04176_);
  and _55519_ (_04179_, _03733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _55520_ (_04180_, _03731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _55521_ (_04181_, _04180_, _04179_);
  or _55522_ (_04182_, _04181_, _04178_);
  or _55523_ (_04183_, _04182_, _04175_);
  or _55524_ (_04184_, _04183_, _04168_);
  and _55525_ (_04185_, _03740_, _42724_);
  and _55526_ (_04186_, _03742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _55527_ (_04187_, _04186_, _04185_);
  and _55528_ (_04188_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _55529_ (_04189_, _03661_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _55530_ (_04190_, _04189_, _04188_);
  or _55531_ (_04191_, _04190_, _04187_);
  and _55532_ (_04192_, _03749_, _03311_);
  and _55533_ (_04193_, _03751_, _03534_);
  or _55534_ (_04194_, _04193_, _04192_);
  and _55535_ (_04195_, _03756_, _03594_);
  and _55536_ (_04196_, _03754_, _03460_);
  or _55537_ (_04197_, _04196_, _04195_);
  or _55538_ (_04198_, _04197_, _04194_);
  or _55539_ (_04199_, _04198_, _04191_);
  and _55540_ (_04200_, _03657_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _55541_ (_04201_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _55542_ (_04202_, _04201_, _04200_);
  or _55543_ (_04203_, _04202_, _04199_);
  or _55544_ (_04204_, _04203_, _04184_);
  and _55545_ (_04205_, _04204_, _03673_);
  and _55546_ (_04206_, _03794_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or _55547_ (_04207_, _04206_, _03676_);
  or _55548_ (_04208_, _04207_, _04205_);
  and _55549_ (_04209_, _04208_, _43100_);
  and _55550_ (_40166_, _04209_, _04152_);
  and _55551_ (_40237_, _42861_, _43100_);
  nor _55552_ (_40241_, _42823_, rst);
  and _55553_ (_40262_, _43005_, _43100_);
  nor _55554_ (_40265_, _42701_, rst);
  nor _55555_ (_40266_, _42617_, rst);
  not _55556_ (_04210_, _00394_);
  nor _55557_ (_04211_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _55558_ (_04212_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55559_ (_04213_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04212_);
  nor _55560_ (_04214_, _04213_, _04211_);
  nor _55561_ (_04215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55562_ (_04216_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04212_);
  nor _55563_ (_04217_, _04216_, _04215_);
  not _55564_ (_04218_, _04217_);
  nor _55565_ (_04219_, _04218_, _04214_);
  and _55566_ (_04220_, _04217_, _04214_);
  nor _55567_ (_04221_, _02220_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55568_ (_04222_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04212_);
  nor _55569_ (_04223_, _04222_, _04221_);
  and _55570_ (_04224_, _04223_, _04220_);
  nor _55571_ (_04225_, _04223_, _04220_);
  nor _55572_ (_04226_, _04225_, _04224_);
  not _55573_ (_04227_, _04226_);
  nor _55574_ (_04228_, _02239_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55575_ (_04229_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04212_);
  nor _55576_ (_04230_, _04229_, _04228_);
  and _55577_ (_04231_, _04230_, _04224_);
  nor _55578_ (_04232_, _04230_, _04224_);
  nor _55579_ (_04233_, _04232_, _04231_);
  and _55580_ (_04234_, _04233_, _04227_);
  and _55581_ (_04235_, _04234_, _04219_);
  and _55582_ (_04236_, _04235_, _04210_);
  not _55583_ (_04237_, _00312_);
  nor _55584_ (_04238_, _04217_, _04214_);
  and _55585_ (_04239_, _04238_, _04234_);
  and _55586_ (_04240_, _04239_, _04237_);
  or _55587_ (_04241_, _04240_, _04236_);
  not _55588_ (_04242_, _00353_);
  and _55589_ (_04243_, _04218_, _04214_);
  and _55590_ (_04244_, _04243_, _04234_);
  and _55591_ (_04245_, _04244_, _04242_);
  not _55592_ (_04246_, _00035_);
  nor _55593_ (_04247_, _04233_, _04226_);
  and _55594_ (_04248_, _04247_, _04219_);
  and _55595_ (_04249_, _04248_, _04246_);
  or _55596_ (_04251_, _04249_, _04245_);
  or _55597_ (_04252_, _04251_, _04241_);
  not _55598_ (_04253_, _43980_);
  and _55599_ (_04254_, _04247_, _04238_);
  and _55600_ (_04255_, _04254_, _04253_);
  not _55601_ (_04256_, _44021_);
  and _55602_ (_04257_, _04247_, _04243_);
  and _55603_ (_04258_, _04257_, _04256_);
  or _55604_ (_04259_, _04258_, _04255_);
  not _55605_ (_04260_, _00476_);
  and _55606_ (_04261_, _04230_, _04226_);
  and _55607_ (_04262_, _04261_, _04238_);
  and _55608_ (_04263_, _04262_, _04260_);
  not _55609_ (_04264_, _00230_);
  not _55610_ (_04265_, _04230_);
  and _55611_ (_04266_, _04265_, _04226_);
  and _55612_ (_04267_, _04266_, _04219_);
  and _55613_ (_04268_, _04267_, _04264_);
  or _55614_ (_04269_, _04268_, _04263_);
  not _55615_ (_04270_, _00517_);
  and _55616_ (_04271_, _04261_, _04243_);
  and _55617_ (_04272_, _04271_, _04270_);
  not _55618_ (_04273_, _00117_);
  and _55619_ (_04274_, _04266_, _04238_);
  and _55620_ (_04275_, _04274_, _04273_);
  or _55621_ (_04276_, _04275_, _04272_);
  or _55622_ (_04277_, _04276_, _04269_);
  not _55623_ (_04278_, _00076_);
  and _55624_ (_04279_, _04232_, _04220_);
  and _55625_ (_04280_, _04279_, _04278_);
  not _55626_ (_04281_, _00271_);
  and _55627_ (_04282_, _04265_, _04224_);
  and _55628_ (_04283_, _04282_, _04281_);
  and _55629_ (_04284_, _04223_, _04219_);
  and _55630_ (_04285_, _04284_, _04230_);
  and _55631_ (_04286_, _04285_, _00567_);
  not _55632_ (_04287_, _43939_);
  and _55633_ (_04288_, _04231_, _04287_);
  or _55634_ (_04289_, _04288_, _04286_);
  or _55635_ (_04290_, _04289_, _04283_);
  or _55636_ (_04291_, _04290_, _04280_);
  not _55637_ (_04292_, _00435_);
  and _55638_ (_04293_, _04261_, _04220_);
  and _55639_ (_04294_, _04293_, _04292_);
  not _55640_ (_04295_, _00189_);
  and _55641_ (_04296_, _04266_, _04243_);
  and _55642_ (_04297_, _04296_, _04295_);
  or _55643_ (_04298_, _04297_, _04294_);
  or _55644_ (_04299_, _04298_, _04291_);
  or _55645_ (_04300_, _04299_, _04277_);
  or _55646_ (_04301_, _04300_, _04259_);
  or _55647_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04301_, _04252_);
  and _55648_ (_04302_, _04235_, _04292_);
  and _55649_ (_04303_, _04239_, _04242_);
  or _55650_ (_04304_, _04303_, _04302_);
  and _55651_ (_04305_, _04244_, _04210_);
  and _55652_ (_04306_, _04248_, _04278_);
  or _55653_ (_04307_, _04306_, _04305_);
  or _55654_ (_04308_, _04307_, _04304_);
  and _55655_ (_04309_, _04296_, _04264_);
  and _55656_ (_04310_, _04274_, _04295_);
  or _55657_ (_04311_, _04310_, _04309_);
  and _55658_ (_04312_, _04262_, _04270_);
  and _55659_ (_04313_, _04267_, _04281_);
  or _55660_ (_04314_, _04313_, _04312_);
  or _55661_ (_04315_, _04314_, _04311_);
  and _55662_ (_04316_, _04279_, _04273_);
  and _55663_ (_04317_, _04231_, _04253_);
  and _55664_ (_04318_, _04282_, _04237_);
  and _55665_ (_04319_, _04285_, _04287_);
  or _55666_ (_04320_, _04319_, _04318_);
  or _55667_ (_04321_, _04320_, _04317_);
  or _55668_ (_04322_, _04321_, _04316_);
  and _55669_ (_04323_, _04271_, _00567_);
  and _55670_ (_04324_, _04293_, _04260_);
  or _55671_ (_04325_, _04324_, _04323_);
  or _55672_ (_04326_, _04325_, _04322_);
  or _55673_ (_04327_, _04326_, _04315_);
  and _55674_ (_04328_, _04257_, _04246_);
  and _55675_ (_04329_, _04254_, _04256_);
  or _55676_ (_04330_, _04329_, _04328_);
  or _55677_ (_04331_, _04330_, _04327_);
  or _55678_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04331_, _04308_);
  and _55679_ (_04332_, _04239_, _04210_);
  and _55680_ (_04333_, _04248_, _04273_);
  or _55681_ (_04334_, _04333_, _04332_);
  and _55682_ (_04335_, _04244_, _04292_);
  and _55683_ (_04336_, _04235_, _04260_);
  or _55684_ (_04337_, _04336_, _04335_);
  or _55685_ (_04338_, _04337_, _04334_);
  and _55686_ (_04339_, _04254_, _04246_);
  and _55687_ (_04340_, _04257_, _04278_);
  or _55688_ (_04341_, _04340_, _04339_);
  and _55689_ (_04342_, _04262_, _00567_);
  and _55690_ (_04343_, _04267_, _04237_);
  or _55691_ (_04344_, _04343_, _04342_);
  and _55692_ (_04345_, _04293_, _04270_);
  and _55693_ (_04346_, _04274_, _04264_);
  or _55694_ (_04347_, _04346_, _04345_);
  or _55695_ (_04348_, _04347_, _04344_);
  and _55696_ (_04350_, _04279_, _04295_);
  and _55697_ (_04351_, _04285_, _04253_);
  and _55698_ (_04352_, _04282_, _04242_);
  and _55699_ (_04353_, _04231_, _04256_);
  or _55700_ (_04354_, _04353_, _04352_);
  or _55701_ (_04355_, _04354_, _04351_);
  or _55702_ (_04356_, _04355_, _04350_);
  and _55703_ (_04357_, _04296_, _04281_);
  and _55704_ (_04358_, _04271_, _04287_);
  or _55705_ (_04359_, _04358_, _04357_);
  or _55706_ (_04360_, _04359_, _04356_);
  or _55707_ (_04361_, _04360_, _04348_);
  or _55708_ (_04362_, _04361_, _04341_);
  or _55709_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04362_, _04338_);
  and _55710_ (_04363_, _04231_, _00567_);
  and _55711_ (_04364_, _04248_, _04256_);
  and _55712_ (_04365_, _04254_, _04287_);
  or _55713_ (_04366_, _04365_, _04364_);
  and _55714_ (_04367_, _04257_, _04253_);
  and _55715_ (_04368_, _04267_, _04295_);
  and _55716_ (_04369_, _04296_, _04273_);
  or _55717_ (_04370_, _04369_, _04368_);
  and _55718_ (_04371_, _04274_, _04278_);
  and _55719_ (_04372_, _04279_, _04246_);
  or _55720_ (_04373_, _04372_, _04371_);
  or _55721_ (_04374_, _04373_, _04370_);
  or _55722_ (_04375_, _04374_, _04367_);
  or _55723_ (_04376_, _04375_, _04366_);
  and _55724_ (_04377_, _04271_, _04260_);
  and _55725_ (_04378_, _04285_, _04270_);
  or _55726_ (_04379_, _04378_, _04377_);
  and _55727_ (_04380_, _04293_, _04210_);
  and _55728_ (_04381_, _04262_, _04292_);
  or _55729_ (_04382_, _04381_, _04380_);
  or _55730_ (_04383_, _04382_, _04379_);
  and _55731_ (_04384_, _04235_, _04242_);
  and _55732_ (_04385_, _04244_, _04237_);
  or _55733_ (_04386_, _04385_, _04384_);
  and _55734_ (_04387_, _04239_, _04281_);
  and _55735_ (_04388_, _04282_, _04264_);
  or _55736_ (_04389_, _04388_, _04387_);
  or _55737_ (_04390_, _04389_, _04386_);
  or _55738_ (_04391_, _04390_, _04383_);
  or _55739_ (_04392_, _04391_, _04376_);
  or _55740_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04392_, _04363_);
  not _55741_ (_04393_, _00399_);
  and _55742_ (_04394_, _04239_, _04393_);
  not _55743_ (_04395_, _00440_);
  and _55744_ (_04396_, _04244_, _04395_);
  or _55745_ (_04397_, _04396_, _04394_);
  not _55746_ (_04398_, _00481_);
  and _55747_ (_04399_, _04235_, _04398_);
  not _55748_ (_04400_, _00122_);
  and _55749_ (_04401_, _04248_, _04400_);
  or _55750_ (_04402_, _04401_, _04399_);
  or _55751_ (_04403_, _04402_, _04397_);
  not _55752_ (_04404_, _00081_);
  and _55753_ (_04405_, _04257_, _04404_);
  not _55754_ (_04406_, _00040_);
  and _55755_ (_04407_, _04254_, _04406_);
  or _55756_ (_04408_, _04407_, _04405_);
  not _55757_ (_04409_, _00317_);
  and _55758_ (_04410_, _04267_, _04409_);
  not _55759_ (_04411_, _00276_);
  and _55760_ (_04412_, _04296_, _04411_);
  or _55761_ (_04413_, _04412_, _04410_);
  not _55762_ (_04414_, _00235_);
  and _55763_ (_04415_, _04274_, _04414_);
  not _55764_ (_04416_, _43944_);
  and _55765_ (_04417_, _04271_, _04416_);
  or _55766_ (_04418_, _04417_, _04415_);
  or _55767_ (_04419_, _04418_, _04413_);
  not _55768_ (_04420_, _00194_);
  and _55769_ (_04421_, _04279_, _04420_);
  not _55770_ (_04422_, _44026_);
  and _55771_ (_04423_, _04231_, _04422_);
  not _55772_ (_04424_, _00358_);
  and _55773_ (_04425_, _04282_, _04424_);
  not _55774_ (_04426_, _43985_);
  and _55775_ (_04427_, _04285_, _04426_);
  or _55776_ (_04428_, _04427_, _04425_);
  or _55777_ (_04429_, _04428_, _04423_);
  or _55778_ (_04430_, _04429_, _04421_);
  and _55779_ (_04431_, _04262_, _00575_);
  not _55780_ (_04432_, _00522_);
  and _55781_ (_04433_, _04293_, _04432_);
  or _55782_ (_04434_, _04433_, _04431_);
  or _55783_ (_04435_, _04434_, _04430_);
  or _55784_ (_04436_, _04435_, _04419_);
  or _55785_ (_04437_, _04436_, _04408_);
  or _55786_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04437_, _04403_);
  not _55787_ (_04438_, _00404_);
  and _55788_ (_04439_, _04239_, _04438_);
  not _55789_ (_04440_, _00445_);
  and _55790_ (_04441_, _04244_, _04440_);
  or _55791_ (_04442_, _04441_, _04439_);
  not _55792_ (_04443_, _00486_);
  and _55793_ (_04444_, _04235_, _04443_);
  not _55794_ (_04445_, _00127_);
  and _55795_ (_04446_, _04248_, _04445_);
  or _55796_ (_04448_, _04446_, _04444_);
  or _55797_ (_04449_, _04448_, _04442_);
  not _55798_ (_04450_, _00086_);
  and _55799_ (_04451_, _04257_, _04450_);
  not _55800_ (_04452_, _00045_);
  and _55801_ (_04453_, _04254_, _04452_);
  or _55802_ (_04454_, _04453_, _04451_);
  not _55803_ (_04455_, _00322_);
  and _55804_ (_04456_, _04267_, _04455_);
  not _55805_ (_04457_, _00281_);
  and _55806_ (_04458_, _04296_, _04457_);
  or _55807_ (_04459_, _04458_, _04456_);
  not _55808_ (_04460_, _00240_);
  and _55809_ (_04461_, _04274_, _04460_);
  not _55810_ (_04462_, _43949_);
  and _55811_ (_04463_, _04271_, _04462_);
  or _55812_ (_04464_, _04463_, _04461_);
  or _55813_ (_04465_, _04464_, _04459_);
  not _55814_ (_04466_, _00199_);
  and _55815_ (_04467_, _04279_, _04466_);
  not _55816_ (_04468_, _00004_);
  and _55817_ (_04469_, _04231_, _04468_);
  not _55818_ (_04470_, _00363_);
  and _55819_ (_04471_, _04282_, _04470_);
  not _55820_ (_04472_, _43990_);
  and _55821_ (_04473_, _04285_, _04472_);
  or _55822_ (_04474_, _04473_, _04471_);
  or _55823_ (_04475_, _04474_, _04469_);
  or _55824_ (_04476_, _04475_, _04467_);
  and _55825_ (_04477_, _04262_, _00583_);
  not _55826_ (_04478_, _00527_);
  and _55827_ (_04479_, _04293_, _04478_);
  or _55828_ (_04480_, _04479_, _04477_);
  or _55829_ (_04481_, _04480_, _04476_);
  or _55830_ (_04482_, _04481_, _04465_);
  or _55831_ (_04483_, _04482_, _04454_);
  or _55832_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04483_, _04449_);
  not _55833_ (_04484_, _00409_);
  and _55834_ (_04485_, _04239_, _04484_);
  not _55835_ (_04486_, _00450_);
  and _55836_ (_04487_, _04244_, _04486_);
  or _55837_ (_04488_, _04487_, _04485_);
  not _55838_ (_04489_, _00491_);
  and _55839_ (_04490_, _04235_, _04489_);
  not _55840_ (_04491_, _00134_);
  and _55841_ (_04492_, _04248_, _04491_);
  or _55842_ (_04493_, _04492_, _04490_);
  or _55843_ (_04494_, _04493_, _04488_);
  not _55844_ (_04495_, _00091_);
  and _55845_ (_04496_, _04257_, _04495_);
  not _55846_ (_04497_, _00050_);
  and _55847_ (_04498_, _04254_, _04497_);
  or _55848_ (_04499_, _04498_, _04496_);
  not _55849_ (_04500_, _00327_);
  and _55850_ (_04501_, _04267_, _04500_);
  not _55851_ (_04502_, _00286_);
  and _55852_ (_04503_, _04296_, _04502_);
  or _55853_ (_04504_, _04503_, _04501_);
  not _55854_ (_04505_, _00245_);
  and _55855_ (_04506_, _04274_, _04505_);
  not _55856_ (_04507_, _43954_);
  and _55857_ (_04508_, _04271_, _04507_);
  or _55858_ (_04509_, _04508_, _04506_);
  or _55859_ (_04510_, _04509_, _04504_);
  not _55860_ (_04511_, _00204_);
  and _55861_ (_04512_, _04279_, _04511_);
  not _55862_ (_04513_, _00009_);
  and _55863_ (_04514_, _04231_, _04513_);
  not _55864_ (_04515_, _00368_);
  and _55865_ (_04516_, _04282_, _04515_);
  not _55866_ (_04517_, _43995_);
  and _55867_ (_04518_, _04285_, _04517_);
  or _55868_ (_04519_, _04518_, _04516_);
  or _55869_ (_04520_, _04519_, _04514_);
  or _55870_ (_04521_, _04520_, _04512_);
  and _55871_ (_04522_, _04262_, _00591_);
  not _55872_ (_04523_, _00532_);
  and _55873_ (_04524_, _04293_, _04523_);
  or _55874_ (_04525_, _04524_, _04522_);
  or _55875_ (_04526_, _04525_, _04521_);
  or _55876_ (_04527_, _04526_, _04510_);
  or _55877_ (_04528_, _04527_, _04499_);
  or _55878_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04528_, _04494_);
  not _55879_ (_04529_, _00455_);
  and _55880_ (_04530_, _04244_, _04529_);
  not _55881_ (_04531_, _00145_);
  and _55882_ (_04532_, _04248_, _04531_);
  or _55883_ (_04533_, _04532_, _04530_);
  not _55884_ (_04534_, _00414_);
  and _55885_ (_04535_, _04239_, _04534_);
  not _55886_ (_04536_, _00496_);
  and _55887_ (_04537_, _04235_, _04536_);
  or _55888_ (_04538_, _04537_, _04535_);
  or _55889_ (_04539_, _04538_, _04533_);
  not _55890_ (_04540_, _00096_);
  and _55891_ (_04541_, _04257_, _04540_);
  not _55892_ (_04542_, _00055_);
  and _55893_ (_04543_, _04254_, _04542_);
  or _55894_ (_04544_, _04543_, _04541_);
  not _55895_ (_04545_, _00332_);
  and _55896_ (_04547_, _04267_, _04545_);
  not _55897_ (_04548_, _00291_);
  and _55898_ (_04549_, _04296_, _04548_);
  or _55899_ (_04550_, _04549_, _04547_);
  not _55900_ (_04551_, _00537_);
  and _55901_ (_04552_, _04293_, _04551_);
  not _55902_ (_04553_, _43959_);
  and _55903_ (_04554_, _04271_, _04553_);
  or _55904_ (_04555_, _04554_, _04552_);
  or _55905_ (_04556_, _04555_, _04550_);
  not _55906_ (_04557_, _00209_);
  and _55907_ (_04558_, _04279_, _04557_);
  not _55908_ (_04559_, _00014_);
  and _55909_ (_04560_, _04231_, _04559_);
  not _55910_ (_04561_, _00373_);
  and _55911_ (_04562_, _04282_, _04561_);
  not _55912_ (_04563_, _44000_);
  and _55913_ (_04564_, _04285_, _04563_);
  or _55914_ (_04565_, _04564_, _04562_);
  or _55915_ (_04566_, _04565_, _04560_);
  or _55916_ (_04567_, _04566_, _04558_);
  and _55917_ (_04568_, _04262_, _00597_);
  not _55918_ (_04569_, _00250_);
  and _55919_ (_04570_, _04274_, _04569_);
  or _55920_ (_04571_, _04570_, _04568_);
  or _55921_ (_04572_, _04571_, _04567_);
  or _55922_ (_04573_, _04572_, _04556_);
  or _55923_ (_04574_, _04573_, _04544_);
  or _55924_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04574_, _04539_);
  not _55925_ (_04575_, _00460_);
  and _55926_ (_04576_, _04244_, _04575_);
  not _55927_ (_04577_, _00156_);
  and _55928_ (_04578_, _04248_, _04577_);
  or _55929_ (_04579_, _04578_, _04576_);
  not _55930_ (_04580_, _00419_);
  and _55931_ (_04581_, _04239_, _04580_);
  not _55932_ (_04582_, _00501_);
  and _55933_ (_04583_, _04235_, _04582_);
  or _55934_ (_04584_, _04583_, _04581_);
  or _55935_ (_04585_, _04584_, _04579_);
  not _55936_ (_04586_, _00101_);
  and _55937_ (_04587_, _04257_, _04586_);
  not _55938_ (_04588_, _00060_);
  and _55939_ (_04589_, _04254_, _04588_);
  or _55940_ (_04590_, _04589_, _04587_);
  not _55941_ (_04591_, _00337_);
  and _55942_ (_04592_, _04267_, _04591_);
  not _55943_ (_04593_, _00296_);
  and _55944_ (_04594_, _04296_, _04593_);
  or _55945_ (_04595_, _04594_, _04592_);
  not _55946_ (_04596_, _00542_);
  and _55947_ (_04597_, _04293_, _04596_);
  not _55948_ (_04598_, _43964_);
  and _55949_ (_04599_, _04271_, _04598_);
  or _55950_ (_04600_, _04599_, _04597_);
  or _55951_ (_04601_, _04600_, _04595_);
  not _55952_ (_04602_, _00214_);
  and _55953_ (_04603_, _04279_, _04602_);
  not _55954_ (_04604_, _00378_);
  and _55955_ (_04605_, _04282_, _04604_);
  not _55956_ (_04606_, _44005_);
  and _55957_ (_04607_, _04285_, _04606_);
  not _55958_ (_04608_, _00019_);
  and _55959_ (_04609_, _04231_, _04608_);
  or _55960_ (_04610_, _04609_, _04607_);
  or _55961_ (_04611_, _04610_, _04605_);
  or _55962_ (_04612_, _04611_, _04603_);
  and _55963_ (_04613_, _04262_, _00602_);
  not _55964_ (_04614_, _00255_);
  and _55965_ (_04615_, _04274_, _04614_);
  or _55966_ (_04616_, _04615_, _04613_);
  or _55967_ (_04617_, _04616_, _04612_);
  or _55968_ (_04618_, _04617_, _04601_);
  or _55969_ (_04619_, _04618_, _04590_);
  or _55970_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _04619_, _04585_);
  not _55971_ (_04620_, _00424_);
  and _55972_ (_04621_, _04239_, _04620_);
  not _55973_ (_04622_, _00465_);
  and _55974_ (_04623_, _04244_, _04622_);
  or _55975_ (_04624_, _04623_, _04621_);
  not _55976_ (_04625_, _00506_);
  and _55977_ (_04626_, _04235_, _04625_);
  not _55978_ (_04627_, _00167_);
  and _55979_ (_04628_, _04248_, _04627_);
  or _55980_ (_04629_, _04628_, _04626_);
  or _55981_ (_04630_, _04629_, _04624_);
  not _55982_ (_04631_, _00106_);
  and _55983_ (_04632_, _04257_, _04631_);
  not _55984_ (_04633_, _00065_);
  and _55985_ (_04634_, _04254_, _04633_);
  or _55986_ (_04635_, _04634_, _04632_);
  not _55987_ (_04636_, _00342_);
  and _55988_ (_04637_, _04267_, _04636_);
  not _55989_ (_04638_, _00301_);
  and _55990_ (_04639_, _04296_, _04638_);
  or _55991_ (_04640_, _04639_, _04637_);
  not _55992_ (_04641_, _00260_);
  and _55993_ (_04642_, _04274_, _04641_);
  not _55994_ (_04643_, _43969_);
  and _55995_ (_04644_, _04271_, _04643_);
  or _55996_ (_04646_, _04644_, _04642_);
  or _55997_ (_04647_, _04646_, _04640_);
  not _55998_ (_04648_, _00219_);
  and _55999_ (_04649_, _04279_, _04648_);
  not _56000_ (_04650_, _00024_);
  and _56001_ (_04651_, _04231_, _04650_);
  not _56002_ (_04652_, _00383_);
  and _56003_ (_04653_, _04282_, _04652_);
  not _56004_ (_04654_, _44010_);
  and _56005_ (_04655_, _04285_, _04654_);
  or _56006_ (_04656_, _04655_, _04653_);
  or _56007_ (_04657_, _04656_, _04651_);
  or _56008_ (_04658_, _04657_, _04649_);
  and _56009_ (_04659_, _04262_, _00607_);
  not _56010_ (_04660_, _00550_);
  and _56011_ (_04661_, _04293_, _04660_);
  or _56012_ (_04662_, _04661_, _04659_);
  or _56013_ (_04663_, _04662_, _04658_);
  or _56014_ (_04664_, _04663_, _04647_);
  or _56015_ (_04665_, _04664_, _04635_);
  or _56016_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _04665_, _04630_);
  not _56017_ (_04666_, _00429_);
  and _56018_ (_04667_, _04239_, _04666_);
  not _56019_ (_04668_, _00470_);
  and _56020_ (_04669_, _04244_, _04668_);
  or _56021_ (_04670_, _04669_, _04667_);
  not _56022_ (_04671_, _00511_);
  and _56023_ (_04672_, _04235_, _04671_);
  not _56024_ (_04673_, _00178_);
  and _56025_ (_04674_, _04248_, _04673_);
  or _56026_ (_04675_, _04674_, _04672_);
  or _56027_ (_04676_, _04675_, _04670_);
  not _56028_ (_04677_, _00111_);
  and _56029_ (_04678_, _04257_, _04677_);
  not _56030_ (_04679_, _00070_);
  and _56031_ (_04680_, _04254_, _04679_);
  or _56032_ (_04681_, _04680_, _04678_);
  not _56033_ (_04682_, _00347_);
  and _56034_ (_04683_, _04267_, _04682_);
  not _56035_ (_04684_, _00306_);
  and _56036_ (_04685_, _04296_, _04684_);
  or _56037_ (_04686_, _04685_, _04683_);
  not _56038_ (_04687_, _00265_);
  and _56039_ (_04688_, _04274_, _04687_);
  not _56040_ (_04689_, _43974_);
  and _56041_ (_04690_, _04271_, _04689_);
  or _56042_ (_04691_, _04690_, _04688_);
  or _56043_ (_04692_, _04691_, _04686_);
  not _56044_ (_04693_, _00224_);
  and _56045_ (_04694_, _04279_, _04693_);
  not _56046_ (_04695_, _00029_);
  and _56047_ (_04696_, _04231_, _04695_);
  not _56048_ (_04697_, _00388_);
  and _56049_ (_04698_, _04282_, _04697_);
  not _56050_ (_04699_, _44015_);
  and _56051_ (_04700_, _04285_, _04699_);
  or _56052_ (_04701_, _04700_, _04698_);
  or _56053_ (_04702_, _04701_, _04696_);
  or _56054_ (_04703_, _04702_, _04694_);
  and _56055_ (_04704_, _04262_, _00612_);
  not _56056_ (_04705_, _00558_);
  and _56057_ (_04706_, _04293_, _04705_);
  or _56058_ (_04707_, _04706_, _04704_);
  or _56059_ (_04708_, _04707_, _04703_);
  or _56060_ (_04709_, _04708_, _04692_);
  or _56061_ (_04710_, _04709_, _04681_);
  or _56062_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _04710_, _04676_);
  and _56063_ (_04711_, _04235_, _04395_);
  and _56064_ (_04712_, _04244_, _04393_);
  or _56065_ (_04713_, _04712_, _04711_);
  and _56066_ (_04714_, _04239_, _04424_);
  and _56067_ (_04715_, _04248_, _04404_);
  or _56068_ (_04716_, _04715_, _04714_);
  or _56069_ (_04717_, _04716_, _04713_);
  and _56070_ (_04718_, _04296_, _04414_);
  and _56071_ (_04719_, _04274_, _04420_);
  or _56072_ (_04720_, _04719_, _04718_);
  and _56073_ (_04721_, _04262_, _04432_);
  and _56074_ (_04722_, _04267_, _04411_);
  or _56075_ (_04723_, _04722_, _04721_);
  or _56076_ (_04724_, _04723_, _04720_);
  and _56077_ (_04725_, _04279_, _04400_);
  and _56078_ (_04726_, _04231_, _04426_);
  and _56079_ (_04727_, _04282_, _04409_);
  and _56080_ (_04728_, _04285_, _04416_);
  or _56081_ (_04729_, _04728_, _04727_);
  or _56082_ (_04730_, _04729_, _04726_);
  or _56083_ (_04731_, _04730_, _04725_);
  and _56084_ (_04732_, _04271_, _00575_);
  and _56085_ (_04733_, _04293_, _04398_);
  or _56086_ (_04734_, _04733_, _04732_);
  or _56087_ (_04735_, _04734_, _04731_);
  or _56088_ (_04736_, _04735_, _04724_);
  and _56089_ (_04737_, _04257_, _04406_);
  and _56090_ (_04738_, _04254_, _04422_);
  or _56091_ (_04739_, _04738_, _04737_);
  or _56092_ (_04740_, _04739_, _04736_);
  or _56093_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _04740_, _04717_);
  and _56094_ (_04741_, _04244_, _04438_);
  and _56095_ (_04742_, _04239_, _04470_);
  or _56096_ (_04743_, _04742_, _04741_);
  and _56097_ (_04744_, _04235_, _04440_);
  and _56098_ (_04745_, _04248_, _04450_);
  or _56099_ (_04746_, _04745_, _04744_);
  or _56100_ (_04747_, _04746_, _04743_);
  and _56101_ (_04748_, _04296_, _04460_);
  and _56102_ (_04749_, _04274_, _04466_);
  or _56103_ (_04750_, _04749_, _04748_);
  and _56104_ (_04751_, _04271_, _00583_);
  and _56105_ (_04752_, _04262_, _04478_);
  or _56106_ (_04753_, _04752_, _04751_);
  or _56107_ (_04754_, _04753_, _04750_);
  and _56108_ (_04755_, _04279_, _04445_);
  and _56109_ (_04756_, _04231_, _04472_);
  and _56110_ (_04757_, _04282_, _04455_);
  and _56111_ (_04758_, _04285_, _04462_);
  or _56112_ (_04759_, _04758_, _04757_);
  or _56113_ (_04760_, _04759_, _04756_);
  or _56114_ (_04761_, _04760_, _04755_);
  and _56115_ (_04762_, _04293_, _04443_);
  and _56116_ (_04763_, _04267_, _04457_);
  or _56117_ (_04764_, _04763_, _04762_);
  or _56118_ (_04765_, _04764_, _04761_);
  or _56119_ (_04766_, _04765_, _04754_);
  and _56120_ (_04767_, _04257_, _04452_);
  and _56121_ (_04768_, _04254_, _04468_);
  or _56122_ (_04769_, _04768_, _04767_);
  or _56123_ (_04770_, _04769_, _04766_);
  or _56124_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _04770_, _04747_);
  and _56125_ (_04771_, _04235_, _04486_);
  and _56126_ (_04772_, _04244_, _04484_);
  or _56127_ (_04773_, _04772_, _04771_);
  and _56128_ (_04774_, _04239_, _04515_);
  and _56129_ (_04775_, _04248_, _04495_);
  or _56130_ (_04776_, _04775_, _04774_);
  or _56131_ (_04777_, _04776_, _04773_);
  and _56132_ (_04778_, _04296_, _04505_);
  and _56133_ (_04779_, _04274_, _04511_);
  or _56134_ (_04780_, _04779_, _04778_);
  and _56135_ (_04781_, _04262_, _04523_);
  and _56136_ (_04782_, _04267_, _04502_);
  or _56137_ (_04783_, _04782_, _04781_);
  or _56138_ (_04784_, _04783_, _04780_);
  and _56139_ (_04785_, _04279_, _04491_);
  and _56140_ (_04786_, _04231_, _04517_);
  and _56141_ (_04787_, _04282_, _04500_);
  and _56142_ (_04788_, _04285_, _04507_);
  or _56143_ (_04789_, _04788_, _04787_);
  or _56144_ (_04790_, _04789_, _04786_);
  or _56145_ (_04791_, _04790_, _04785_);
  and _56146_ (_04792_, _04271_, _00591_);
  and _56147_ (_04793_, _04293_, _04489_);
  or _56148_ (_04794_, _04793_, _04792_);
  or _56149_ (_04795_, _04794_, _04791_);
  or _56150_ (_04796_, _04795_, _04784_);
  and _56151_ (_04797_, _04257_, _04497_);
  and _56152_ (_04798_, _04254_, _04513_);
  or _56153_ (_04799_, _04798_, _04797_);
  or _56154_ (_04800_, _04799_, _04796_);
  or _56155_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _04800_, _04777_);
  and _56156_ (_04801_, _04244_, _04534_);
  and _56157_ (_04802_, _04235_, _04529_);
  or _56158_ (_04803_, _04802_, _04801_);
  and _56159_ (_04804_, _04239_, _04561_);
  and _56160_ (_04805_, _04248_, _04540_);
  or _56161_ (_04806_, _04805_, _04804_);
  or _56162_ (_04807_, _04806_, _04803_);
  and _56163_ (_04808_, _04271_, _00597_);
  and _56164_ (_04809_, _04267_, _04548_);
  or _56165_ (_04810_, _04809_, _04808_);
  and _56166_ (_04811_, _04293_, _04536_);
  and _56167_ (_04812_, _04274_, _04557_);
  or _56168_ (_04813_, _04812_, _04811_);
  or _56169_ (_04814_, _04813_, _04810_);
  and _56170_ (_04815_, _04279_, _04531_);
  and _56171_ (_04816_, _04282_, _04545_);
  and _56172_ (_04817_, _04285_, _04553_);
  and _56173_ (_04818_, _04231_, _04563_);
  or _56174_ (_04819_, _04818_, _04817_);
  or _56175_ (_04820_, _04819_, _04816_);
  or _56176_ (_04821_, _04820_, _04815_);
  and _56177_ (_04822_, _04262_, _04551_);
  and _56178_ (_04823_, _04296_, _04569_);
  or _56179_ (_04824_, _04823_, _04822_);
  or _56180_ (_04825_, _04824_, _04821_);
  or _56181_ (_04826_, _04825_, _04814_);
  and _56182_ (_04827_, _04257_, _04542_);
  and _56183_ (_04828_, _04254_, _04559_);
  or _56184_ (_04829_, _04828_, _04827_);
  or _56185_ (_04830_, _04829_, _04826_);
  or _56186_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _04830_, _04807_);
  and _56187_ (_04831_, _04235_, _04575_);
  and _56188_ (_04832_, _04239_, _04604_);
  or _56189_ (_04833_, _04832_, _04831_);
  and _56190_ (_04834_, _04244_, _04580_);
  and _56191_ (_04835_, _04248_, _04586_);
  or _56192_ (_04836_, _04835_, _04834_);
  or _56193_ (_04837_, _04836_, _04833_);
  and _56194_ (_04838_, _04296_, _04614_);
  and _56195_ (_04839_, _04274_, _04602_);
  or _56196_ (_04840_, _04839_, _04838_);
  and _56197_ (_04841_, _04262_, _04596_);
  and _56198_ (_04842_, _04267_, _04593_);
  or _56199_ (_04843_, _04842_, _04841_);
  or _56200_ (_04844_, _04843_, _04840_);
  and _56201_ (_04845_, _04279_, _04577_);
  and _56202_ (_04846_, _04231_, _04606_);
  and _56203_ (_04847_, _04282_, _04591_);
  and _56204_ (_04848_, _04285_, _04598_);
  or _56205_ (_04849_, _04848_, _04847_);
  or _56206_ (_04850_, _04849_, _04846_);
  or _56207_ (_04851_, _04850_, _04845_);
  and _56208_ (_04852_, _04271_, _00602_);
  and _56209_ (_04853_, _04293_, _04582_);
  or _56210_ (_04854_, _04853_, _04852_);
  or _56211_ (_04855_, _04854_, _04851_);
  or _56212_ (_04856_, _04855_, _04844_);
  and _56213_ (_04857_, _04257_, _04588_);
  and _56214_ (_04858_, _04254_, _04608_);
  or _56215_ (_04859_, _04858_, _04857_);
  or _56216_ (_04860_, _04859_, _04856_);
  or _56217_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _04860_, _04837_);
  and _56218_ (_04861_, _04244_, _04620_);
  and _56219_ (_04862_, _04235_, _04622_);
  or _56220_ (_04863_, _04862_, _04861_);
  and _56221_ (_04864_, _04239_, _04652_);
  and _56222_ (_04865_, _04248_, _04631_);
  or _56223_ (_04866_, _04865_, _04864_);
  or _56224_ (_04867_, _04866_, _04863_);
  and _56225_ (_04868_, _04296_, _04641_);
  and _56226_ (_04869_, _04274_, _04648_);
  or _56227_ (_04870_, _04869_, _04868_);
  and _56228_ (_04871_, _04271_, _00607_);
  and _56229_ (_04872_, _04293_, _04625_);
  or _56230_ (_04873_, _04872_, _04871_);
  or _56231_ (_04874_, _04873_, _04870_);
  and _56232_ (_04875_, _04279_, _04627_);
  and _56233_ (_04876_, _04285_, _04643_);
  and _56234_ (_04877_, _04282_, _04636_);
  and _56235_ (_04878_, _04231_, _04654_);
  or _56236_ (_04879_, _04878_, _04877_);
  or _56237_ (_04880_, _04879_, _04876_);
  or _56238_ (_04881_, _04880_, _04875_);
  and _56239_ (_04882_, _04262_, _04660_);
  and _56240_ (_04883_, _04267_, _04638_);
  or _56241_ (_04884_, _04883_, _04882_);
  or _56242_ (_04885_, _04884_, _04881_);
  or _56243_ (_04886_, _04885_, _04874_);
  and _56244_ (_04887_, _04257_, _04633_);
  and _56245_ (_04888_, _04254_, _04650_);
  or _56246_ (_04889_, _04888_, _04887_);
  or _56247_ (_04890_, _04889_, _04886_);
  or _56248_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _04890_, _04867_);
  and _56249_ (_04891_, _04235_, _04668_);
  and _56250_ (_04892_, _04239_, _04697_);
  or _56251_ (_04893_, _04892_, _04891_);
  and _56252_ (_04894_, _04244_, _04666_);
  and _56253_ (_04895_, _04248_, _04677_);
  or _56254_ (_04896_, _04895_, _04894_);
  or _56255_ (_04897_, _04896_, _04893_);
  and _56256_ (_04898_, _04296_, _04687_);
  and _56257_ (_04899_, _04274_, _04693_);
  or _56258_ (_04900_, _04899_, _04898_);
  and _56259_ (_04901_, _04262_, _04705_);
  and _56260_ (_04902_, _04267_, _04684_);
  or _56261_ (_04903_, _04902_, _04901_);
  or _56262_ (_04904_, _04903_, _04900_);
  and _56263_ (_04905_, _04279_, _04673_);
  and _56264_ (_04906_, _04231_, _04699_);
  and _56265_ (_04907_, _04282_, _04682_);
  and _56266_ (_04908_, _04285_, _04689_);
  or _56267_ (_04909_, _04908_, _04907_);
  or _56268_ (_04910_, _04909_, _04906_);
  or _56269_ (_04911_, _04910_, _04905_);
  and _56270_ (_04912_, _04271_, _00612_);
  and _56271_ (_04913_, _04293_, _04671_);
  or _56272_ (_04914_, _04913_, _04912_);
  or _56273_ (_04915_, _04914_, _04911_);
  or _56274_ (_04916_, _04915_, _04904_);
  and _56275_ (_04917_, _04257_, _04679_);
  and _56276_ (_04918_, _04254_, _04695_);
  or _56277_ (_04919_, _04918_, _04917_);
  or _56278_ (_04920_, _04919_, _04916_);
  or _56279_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _04920_, _04897_);
  and _56280_ (_04921_, _04235_, _04393_);
  and _56281_ (_04922_, _04239_, _04409_);
  or _56282_ (_04923_, _04922_, _04921_);
  and _56283_ (_04924_, _04244_, _04424_);
  and _56284_ (_04925_, _04248_, _04406_);
  or _56285_ (_04926_, _04925_, _04924_);
  or _56286_ (_04927_, _04926_, _04923_);
  and _56287_ (_04928_, _04254_, _04426_);
  and _56288_ (_04929_, _04257_, _04422_);
  or _56289_ (_04930_, _04929_, _04928_);
  and _56290_ (_04931_, _04274_, _04400_);
  and _56291_ (_04932_, _04296_, _04420_);
  or _56292_ (_04933_, _04932_, _04931_);
  and _56293_ (_04934_, _04262_, _04398_);
  and _56294_ (_04935_, _04267_, _04414_);
  or _56295_ (_04936_, _04935_, _04934_);
  or _56296_ (_04937_, _04936_, _04933_);
  and _56297_ (_04938_, _04279_, _04404_);
  and _56298_ (_04939_, _04231_, _04416_);
  and _56299_ (_04940_, _04285_, _00575_);
  and _56300_ (_04941_, _04282_, _04411_);
  or _56301_ (_04942_, _04941_, _04940_);
  or _56302_ (_04943_, _04942_, _04939_);
  or _56303_ (_04944_, _04943_, _04938_);
  and _56304_ (_04945_, _04271_, _04432_);
  and _56305_ (_04946_, _04293_, _04395_);
  or _56306_ (_04947_, _04946_, _04945_);
  or _56307_ (_04948_, _04947_, _04944_);
  or _56308_ (_04949_, _04948_, _04937_);
  or _56309_ (_04950_, _04949_, _04930_);
  or _56310_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _04950_, _04927_);
  and _56311_ (_04951_, _04239_, _04455_);
  and _56312_ (_04952_, _04244_, _04470_);
  or _56313_ (_04953_, _04952_, _04951_);
  and _56314_ (_04954_, _04235_, _04438_);
  and _56315_ (_04955_, _04248_, _04452_);
  or _56316_ (_04956_, _04955_, _04954_);
  or _56317_ (_04957_, _04956_, _04953_);
  and _56318_ (_04958_, _04254_, _04472_);
  and _56319_ (_04959_, _04257_, _04468_);
  or _56320_ (_04960_, _04959_, _04958_);
  and _56321_ (_04961_, _04262_, _04443_);
  and _56322_ (_04962_, _04271_, _04478_);
  or _56323_ (_04963_, _04962_, _04961_);
  and _56324_ (_04964_, _04274_, _04445_);
  and _56325_ (_04965_, _04296_, _04466_);
  or _56326_ (_04966_, _04965_, _04964_);
  or _56327_ (_04967_, _04966_, _04963_);
  and _56328_ (_04968_, _04279_, _04450_);
  and _56329_ (_04969_, _04285_, _00583_);
  and _56330_ (_04970_, _04282_, _04457_);
  and _56331_ (_04971_, _04231_, _04462_);
  or _56332_ (_04972_, _04971_, _04970_);
  or _56333_ (_04973_, _04972_, _04969_);
  or _56334_ (_04974_, _04973_, _04968_);
  and _56335_ (_04975_, _04293_, _04440_);
  and _56336_ (_04976_, _04267_, _04460_);
  or _56337_ (_04977_, _04976_, _04975_);
  or _56338_ (_04978_, _04977_, _04974_);
  or _56339_ (_04979_, _04978_, _04967_);
  or _56340_ (_04980_, _04979_, _04960_);
  or _56341_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _04980_, _04957_);
  and _56342_ (_04981_, _04244_, _04515_);
  and _56343_ (_04982_, _04239_, _04500_);
  or _56344_ (_04983_, _04982_, _04981_);
  and _56345_ (_04984_, _04235_, _04484_);
  and _56346_ (_04985_, _04248_, _04497_);
  or _56347_ (_04986_, _04985_, _04984_);
  or _56348_ (_04987_, _04986_, _04983_);
  and _56349_ (_04988_, _04254_, _04517_);
  and _56350_ (_04989_, _04257_, _04513_);
  or _56351_ (_04990_, _04989_, _04988_);
  and _56352_ (_04991_, _04267_, _04505_);
  and _56353_ (_04992_, _04274_, _04491_);
  or _56354_ (_04993_, _04992_, _04991_);
  and _56355_ (_04994_, _04293_, _04486_);
  and _56356_ (_04995_, _04296_, _04511_);
  or _56357_ (_04996_, _04995_, _04994_);
  or _56358_ (_04997_, _04996_, _04993_);
  and _56359_ (_04998_, _04271_, _04523_);
  and _56360_ (_04999_, _04262_, _04489_);
  or _56361_ (_05000_, _04999_, _04998_);
  and _56362_ (_05001_, _04279_, _04495_);
  and _56363_ (_05002_, _04231_, _04507_);
  and _56364_ (_05003_, _04285_, _00591_);
  and _56365_ (_05004_, _04282_, _04502_);
  or _56366_ (_05005_, _05004_, _05003_);
  or _56367_ (_05006_, _05005_, _05002_);
  or _56368_ (_05007_, _05006_, _05001_);
  or _56369_ (_05008_, _05007_, _05000_);
  or _56370_ (_05009_, _05008_, _04997_);
  or _56371_ (_05010_, _05009_, _04990_);
  or _56372_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05010_, _04987_);
  and _56373_ (_05011_, _04239_, _04545_);
  and _56374_ (_05012_, _04244_, _04561_);
  or _56375_ (_05013_, _05012_, _05011_);
  and _56376_ (_05014_, _04235_, _04534_);
  and _56377_ (_05015_, _04248_, _04542_);
  or _56378_ (_05016_, _05015_, _05014_);
  or _56379_ (_05017_, _05016_, _05013_);
  and _56380_ (_05018_, _04254_, _04563_);
  and _56381_ (_05019_, _04257_, _04559_);
  or _56382_ (_05020_, _05019_, _05018_);
  and _56383_ (_05021_, _04262_, _04536_);
  and _56384_ (_05022_, _04271_, _04551_);
  or _56385_ (_05023_, _05022_, _05021_);
  and _56386_ (_05024_, _04274_, _04531_);
  and _56387_ (_05025_, _04296_, _04557_);
  or _56388_ (_05026_, _05025_, _05024_);
  or _56389_ (_05027_, _05026_, _05023_);
  and _56390_ (_05028_, _04279_, _04540_);
  and _56391_ (_05029_, _04285_, _00597_);
  and _56392_ (_05030_, _04282_, _04548_);
  and _56393_ (_05031_, _04231_, _04553_);
  or _56394_ (_05032_, _05031_, _05030_);
  or _56395_ (_05033_, _05032_, _05029_);
  or _56396_ (_05034_, _05033_, _05028_);
  and _56397_ (_05035_, _04293_, _04529_);
  and _56398_ (_05036_, _04267_, _04569_);
  or _56399_ (_05037_, _05036_, _05035_);
  or _56400_ (_05038_, _05037_, _05034_);
  or _56401_ (_05039_, _05038_, _05027_);
  or _56402_ (_05040_, _05039_, _05020_);
  or _56403_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05040_, _05017_);
  and _56404_ (_05041_, _04235_, _04580_);
  and _56405_ (_05042_, _04239_, _04591_);
  or _56406_ (_05043_, _05042_, _05041_);
  and _56407_ (_05044_, _04244_, _04604_);
  and _56408_ (_05045_, _04248_, _04588_);
  or _56409_ (_05046_, _05045_, _05044_);
  or _56410_ (_05047_, _05046_, _05043_);
  and _56411_ (_05048_, _04254_, _04606_);
  and _56412_ (_05049_, _04257_, _04608_);
  or _56413_ (_05050_, _05049_, _05048_);
  and _56414_ (_05051_, _04274_, _04577_);
  and _56415_ (_05052_, _04296_, _04602_);
  or _56416_ (_05053_, _05052_, _05051_);
  and _56417_ (_05054_, _04262_, _04582_);
  and _56418_ (_05055_, _04267_, _04614_);
  or _56419_ (_05056_, _05055_, _05054_);
  or _56420_ (_05057_, _05056_, _05053_);
  and _56421_ (_05058_, _04279_, _04586_);
  and _56422_ (_05059_, _04231_, _04598_);
  and _56423_ (_05060_, _04285_, _00602_);
  and _56424_ (_05061_, _04282_, _04593_);
  or _56425_ (_05062_, _05061_, _05060_);
  or _56426_ (_05063_, _05062_, _05059_);
  or _56427_ (_05064_, _05063_, _05058_);
  and _56428_ (_05065_, _04271_, _04596_);
  and _56429_ (_05066_, _04293_, _04575_);
  or _56430_ (_05067_, _05066_, _05065_);
  or _56431_ (_05068_, _05067_, _05064_);
  or _56432_ (_05069_, _05068_, _05057_);
  or _56433_ (_05070_, _05069_, _05050_);
  or _56434_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05070_, _05047_);
  and _56435_ (_05071_, _04235_, _04620_);
  and _56436_ (_05072_, _04244_, _04652_);
  or _56437_ (_05073_, _05072_, _05071_);
  and _56438_ (_05074_, _04239_, _04636_);
  and _56439_ (_05075_, _04248_, _04633_);
  or _56440_ (_05076_, _05075_, _05074_);
  or _56441_ (_05077_, _05076_, _05073_);
  and _56442_ (_05078_, _04254_, _04654_);
  and _56443_ (_05079_, _04257_, _04650_);
  or _56444_ (_05080_, _05079_, _05078_);
  and _56445_ (_05081_, _04274_, _04627_);
  and _56446_ (_05082_, _04296_, _04648_);
  or _56447_ (_05083_, _05082_, _05081_);
  and _56448_ (_05084_, _04262_, _04625_);
  and _56449_ (_05086_, _04267_, _04641_);
  or _56450_ (_05088_, _05086_, _05084_);
  or _56451_ (_05090_, _05088_, _05083_);
  and _56452_ (_05092_, _04279_, _04631_);
  and _56453_ (_05094_, _04231_, _04643_);
  and _56454_ (_05096_, _04285_, _00607_);
  and _56455_ (_05098_, _04282_, _04638_);
  or _56456_ (_05099_, _05098_, _05096_);
  or _56457_ (_05100_, _05099_, _05094_);
  or _56458_ (_05101_, _05100_, _05092_);
  and _56459_ (_05102_, _04271_, _04660_);
  and _56460_ (_05103_, _04293_, _04622_);
  or _56461_ (_05104_, _05103_, _05102_);
  or _56462_ (_05106_, _05104_, _05101_);
  or _56463_ (_05107_, _05106_, _05090_);
  or _56464_ (_05109_, _05107_, _05080_);
  or _56465_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05109_, _05077_);
  and _56466_ (_05110_, _04235_, _04666_);
  and _56467_ (_05112_, _04244_, _04697_);
  or _56468_ (_05113_, _05112_, _05110_);
  and _56469_ (_05114_, _04239_, _04682_);
  and _56470_ (_05116_, _04248_, _04679_);
  or _56471_ (_05117_, _05116_, _05114_);
  or _56472_ (_05118_, _05117_, _05113_);
  and _56473_ (_05120_, _04254_, _04699_);
  and _56474_ (_05121_, _04257_, _04695_);
  or _56475_ (_05122_, _05121_, _05120_);
  and _56476_ (_05124_, _04274_, _04673_);
  and _56477_ (_05125_, _04296_, _04693_);
  or _56478_ (_05126_, _05125_, _05124_);
  and _56479_ (_05128_, _04262_, _04671_);
  and _56480_ (_05129_, _04267_, _04687_);
  or _56481_ (_05130_, _05129_, _05128_);
  or _56482_ (_05132_, _05130_, _05126_);
  and _56483_ (_05133_, _04279_, _04677_);
  and _56484_ (_05134_, _04231_, _04689_);
  and _56485_ (_05136_, _04285_, _00612_);
  and _56486_ (_05137_, _04282_, _04684_);
  or _56487_ (_05138_, _05137_, _05136_);
  or _56488_ (_05139_, _05138_, _05134_);
  or _56489_ (_05140_, _05139_, _05133_);
  and _56490_ (_05141_, _04271_, _04705_);
  and _56491_ (_05142_, _04293_, _04668_);
  or _56492_ (_05143_, _05142_, _05141_);
  or _56493_ (_05144_, _05143_, _05140_);
  or _56494_ (_05145_, _05144_, _05132_);
  or _56495_ (_05146_, _05145_, _05122_);
  or _56496_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05146_, _05118_);
  and _56497_ (_05147_, _04244_, _04409_);
  and _56498_ (_05148_, _04235_, _04424_);
  or _56499_ (_05149_, _05148_, _05147_);
  and _56500_ (_05150_, _04239_, _04411_);
  and _56501_ (_05151_, _04248_, _04422_);
  or _56502_ (_05152_, _05151_, _05150_);
  or _56503_ (_05153_, _05152_, _05149_);
  and _56504_ (_05154_, _04271_, _04398_);
  and _56505_ (_05155_, _04274_, _04404_);
  or _56506_ (_05157_, _05155_, _05154_);
  and _56507_ (_05158_, _04293_, _04393_);
  and _56508_ (_05160_, _04267_, _04420_);
  or _56509_ (_05161_, _05160_, _05158_);
  or _56510_ (_05162_, _05161_, _05157_);
  and _56511_ (_05164_, _04279_, _04406_);
  and _56512_ (_05165_, _04231_, _00575_);
  and _56513_ (_05166_, _04285_, _04432_);
  and _56514_ (_05168_, _04282_, _04414_);
  or _56515_ (_05169_, _05168_, _05166_);
  or _56516_ (_05170_, _05169_, _05165_);
  or _56517_ (_05172_, _05170_, _05164_);
  and _56518_ (_05173_, _04262_, _04395_);
  and _56519_ (_05174_, _04296_, _04400_);
  or _56520_ (_05176_, _05174_, _05173_);
  or _56521_ (_05177_, _05176_, _05172_);
  or _56522_ (_05178_, _05177_, _05162_);
  and _56523_ (_05180_, _04254_, _04416_);
  and _56524_ (_05181_, _04257_, _04426_);
  or _56525_ (_05182_, _05181_, _05180_);
  or _56526_ (_05184_, _05182_, _05178_);
  or _56527_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _05184_, _05153_);
  and _56528_ (_05185_, _04231_, _00583_);
  and _56529_ (_05187_, _04248_, _04468_);
  and _56530_ (_05188_, _04254_, _04462_);
  or _56531_ (_05189_, _05188_, _05187_);
  and _56532_ (_05190_, _04257_, _04472_);
  and _56533_ (_05191_, _04267_, _04466_);
  and _56534_ (_05192_, _04296_, _04445_);
  or _56535_ (_05193_, _05192_, _05191_);
  and _56536_ (_05194_, _04274_, _04450_);
  and _56537_ (_05195_, _04279_, _04452_);
  or _56538_ (_05196_, _05195_, _05194_);
  or _56539_ (_05197_, _05196_, _05193_);
  or _56540_ (_05198_, _05197_, _05190_);
  or _56541_ (_05199_, _05198_, _05189_);
  and _56542_ (_05200_, _04271_, _04443_);
  and _56543_ (_05201_, _04285_, _04478_);
  or _56544_ (_05202_, _05201_, _05200_);
  and _56545_ (_05203_, _04293_, _04438_);
  and _56546_ (_05204_, _04262_, _04440_);
  or _56547_ (_05205_, _05204_, _05203_);
  or _56548_ (_05206_, _05205_, _05202_);
  and _56549_ (_05207_, _04235_, _04470_);
  and _56550_ (_05209_, _04244_, _04455_);
  or _56551_ (_05210_, _05209_, _05207_);
  and _56552_ (_05212_, _04239_, _04457_);
  and _56553_ (_05213_, _04282_, _04460_);
  or _56554_ (_05214_, _05213_, _05212_);
  or _56555_ (_05216_, _05214_, _05210_);
  or _56556_ (_05217_, _05216_, _05206_);
  or _56557_ (_05218_, _05217_, _05199_);
  or _56558_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _05218_, _05185_);
  and _56559_ (_05220_, _04244_, _04500_);
  and _56560_ (_05221_, _04235_, _04515_);
  or _56561_ (_05223_, _05221_, _05220_);
  and _56562_ (_05224_, _04239_, _04502_);
  and _56563_ (_05225_, _04248_, _04513_);
  or _56564_ (_05227_, _05225_, _05224_);
  or _56565_ (_05228_, _05227_, _05223_);
  and _56566_ (_05229_, _04267_, _04511_);
  and _56567_ (_05231_, _04274_, _04495_);
  or _56568_ (_05232_, _05231_, _05229_);
  and _56569_ (_05233_, _04293_, _04484_);
  and _56570_ (_05235_, _04296_, _04491_);
  or _56571_ (_05236_, _05235_, _05233_);
  or _56572_ (_05237_, _05236_, _05232_);
  and _56573_ (_05239_, _04279_, _04497_);
  and _56574_ (_05240_, _04231_, _00591_);
  and _56575_ (_05241_, _04285_, _04523_);
  and _56576_ (_05242_, _04282_, _04505_);
  or _56577_ (_05243_, _05242_, _05241_);
  or _56578_ (_05244_, _05243_, _05240_);
  or _56579_ (_05245_, _05244_, _05239_);
  and _56580_ (_05246_, _04271_, _04489_);
  and _56581_ (_05247_, _04262_, _04486_);
  or _56582_ (_05248_, _05247_, _05246_);
  or _56583_ (_05249_, _05248_, _05245_);
  or _56584_ (_05250_, _05249_, _05237_);
  and _56585_ (_05251_, _04254_, _04507_);
  and _56586_ (_05252_, _04257_, _04517_);
  or _56587_ (_05253_, _05252_, _05251_);
  or _56588_ (_05254_, _05253_, _05250_);
  or _56589_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _05254_, _05228_);
  and _56590_ (_05255_, _04244_, _04545_);
  and _56591_ (_05256_, _04235_, _04561_);
  or _56592_ (_05257_, _05256_, _05255_);
  and _56593_ (_05258_, _04239_, _04548_);
  and _56594_ (_05260_, _04248_, _04559_);
  or _56595_ (_05261_, _05260_, _05258_);
  or _56596_ (_05263_, _05261_, _05257_);
  and _56597_ (_05264_, _04271_, _04536_);
  and _56598_ (_05265_, _04274_, _04540_);
  or _56599_ (_05267_, _05265_, _05264_);
  and _56600_ (_05268_, _04293_, _04534_);
  and _56601_ (_05269_, _04267_, _04557_);
  or _56602_ (_05271_, _05269_, _05268_);
  or _56603_ (_05272_, _05271_, _05267_);
  and _56604_ (_05273_, _04279_, _04542_);
  and _56605_ (_05275_, _04231_, _00597_);
  and _56606_ (_05276_, _04285_, _04551_);
  and _56607_ (_05277_, _04282_, _04569_);
  or _56608_ (_05279_, _05277_, _05276_);
  or _56609_ (_05280_, _05279_, _05275_);
  or _56610_ (_05281_, _05280_, _05273_);
  and _56611_ (_05283_, _04262_, _04529_);
  and _56612_ (_05284_, _04296_, _04531_);
  or _56613_ (_05285_, _05284_, _05283_);
  or _56614_ (_05287_, _05285_, _05281_);
  or _56615_ (_05288_, _05287_, _05272_);
  and _56616_ (_05289_, _04254_, _04553_);
  and _56617_ (_05291_, _04257_, _04563_);
  or _56618_ (_05292_, _05291_, _05289_);
  or _56619_ (_05293_, _05292_, _05288_);
  or _56620_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _05293_, _05263_);
  and _56621_ (_05294_, _04231_, _00602_);
  and _56622_ (_05295_, _04248_, _04608_);
  and _56623_ (_05296_, _04254_, _04598_);
  or _56624_ (_05297_, _05296_, _05295_);
  and _56625_ (_05298_, _04257_, _04606_);
  and _56626_ (_05299_, _04267_, _04602_);
  and _56627_ (_05300_, _04296_, _04577_);
  or _56628_ (_05301_, _05300_, _05299_);
  and _56629_ (_05302_, _04279_, _04588_);
  and _56630_ (_05303_, _04274_, _04586_);
  or _56631_ (_05304_, _05303_, _05302_);
  or _56632_ (_05305_, _05304_, _05301_);
  or _56633_ (_05306_, _05305_, _05298_);
  or _56634_ (_05307_, _05306_, _05297_);
  and _56635_ (_05308_, _04262_, _04575_);
  and _56636_ (_05309_, _04293_, _04580_);
  or _56637_ (_05310_, _05309_, _05308_);
  and _56638_ (_05312_, _04271_, _04582_);
  and _56639_ (_05313_, _04285_, _04596_);
  or _56640_ (_05315_, _05313_, _05312_);
  or _56641_ (_05316_, _05315_, _05310_);
  and _56642_ (_05317_, _04235_, _04604_);
  and _56643_ (_05319_, _04244_, _04591_);
  or _56644_ (_05320_, _05319_, _05317_);
  and _56645_ (_05321_, _04239_, _04593_);
  and _56646_ (_05323_, _04282_, _04614_);
  or _56647_ (_05324_, _05323_, _05321_);
  or _56648_ (_05325_, _05324_, _05320_);
  or _56649_ (_05327_, _05325_, _05316_);
  or _56650_ (_05328_, _05327_, _05307_);
  or _56651_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _05328_, _05294_);
  and _56652_ (_05330_, _04235_, _04652_);
  and _56653_ (_05331_, _04244_, _04636_);
  or _56654_ (_05332_, _05331_, _05330_);
  and _56655_ (_05334_, _04239_, _04638_);
  and _56656_ (_05335_, _04248_, _04650_);
  or _56657_ (_05336_, _05335_, _05334_);
  or _56658_ (_05338_, _05336_, _05332_);
  and _56659_ (_05339_, _04254_, _04643_);
  and _56660_ (_05340_, _04257_, _04654_);
  or _56661_ (_05342_, _05340_, _05339_);
  and _56662_ (_05343_, _04271_, _04625_);
  and _56663_ (_05344_, _04296_, _04627_);
  or _56664_ (_05345_, _05344_, _05343_);
  and _56665_ (_05346_, _04267_, _04648_);
  and _56666_ (_05347_, _04274_, _04631_);
  or _56667_ (_05348_, _05347_, _05346_);
  or _56668_ (_05349_, _05348_, _05345_);
  and _56669_ (_05350_, _04262_, _04622_);
  and _56670_ (_05351_, _04293_, _04620_);
  or _56671_ (_05352_, _05351_, _05350_);
  and _56672_ (_05353_, _04279_, _04633_);
  and _56673_ (_05354_, _04282_, _04641_);
  and _56674_ (_05355_, _04231_, _00607_);
  and _56675_ (_05356_, _04285_, _04660_);
  or _56676_ (_05357_, _05356_, _05355_);
  or _56677_ (_05358_, _05357_, _05354_);
  or _56678_ (_05359_, _05358_, _05353_);
  or _56679_ (_05360_, _05359_, _05352_);
  or _56680_ (_05361_, _05360_, _05349_);
  or _56681_ (_05362_, _05361_, _05342_);
  or _56682_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _05362_, _05338_);
  and _56683_ (_05364_, _04244_, _04682_);
  and _56684_ (_05366_, _04235_, _04697_);
  or _56685_ (_05367_, _05366_, _05364_);
  and _56686_ (_05368_, _04239_, _04684_);
  and _56687_ (_05370_, _04248_, _04695_);
  or _56688_ (_05371_, _05370_, _05368_);
  or _56689_ (_05372_, _05371_, _05367_);
  and _56690_ (_05374_, _04271_, _04671_);
  and _56691_ (_05375_, _04274_, _04677_);
  or _56692_ (_05376_, _05375_, _05374_);
  and _56693_ (_05378_, _04293_, _04666_);
  and _56694_ (_05379_, _04267_, _04693_);
  or _56695_ (_05380_, _05379_, _05378_);
  or _56696_ (_05382_, _05380_, _05376_);
  and _56697_ (_05383_, _04279_, _04679_);
  and _56698_ (_05384_, _04231_, _00612_);
  and _56699_ (_05386_, _04285_, _04705_);
  and _56700_ (_05387_, _04282_, _04687_);
  or _56701_ (_05388_, _05387_, _05386_);
  or _56702_ (_05390_, _05388_, _05384_);
  or _56703_ (_05391_, _05390_, _05383_);
  and _56704_ (_05392_, _04262_, _04668_);
  and _56705_ (_05394_, _04296_, _04673_);
  or _56706_ (_05395_, _05394_, _05392_);
  or _56707_ (_05396_, _05395_, _05391_);
  or _56708_ (_05397_, _05396_, _05382_);
  and _56709_ (_05398_, _04254_, _04689_);
  and _56710_ (_05399_, _04257_, _04699_);
  or _56711_ (_05400_, _05399_, _05398_);
  or _56712_ (_05401_, _05400_, _05397_);
  or _56713_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _05401_, _05372_);
  nand _56714_ (_05402_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not _56715_ (_05403_, \oc8051_golden_model_1.PC [3]);
  or _56716_ (_05404_, \oc8051_golden_model_1.PC [2], _05403_);
  or _56717_ (_05405_, _05404_, _05402_);
  or _56718_ (_05406_, _05405_, _00429_);
  not _56719_ (_05407_, \oc8051_golden_model_1.PC [1]);
  or _56720_ (_05408_, _05407_, \oc8051_golden_model_1.PC [0]);
  or _56721_ (_05409_, _05408_, _05404_);
  or _56722_ (_05410_, _05409_, _00388_);
  and _56723_ (_05411_, _05410_, _05406_);
  not _56724_ (_05412_, \oc8051_golden_model_1.PC [2]);
  or _56725_ (_05413_, _05412_, \oc8051_golden_model_1.PC [3]);
  or _56726_ (_05415_, _05413_, _05402_);
  or _56727_ (_05416_, _05415_, _00265_);
  or _56728_ (_05418_, _05413_, _05408_);
  or _56729_ (_05419_, _05418_, _00224_);
  and _56730_ (_05420_, _05419_, _05416_);
  and _56731_ (_05422_, _05420_, _05411_);
  and _56732_ (_05423_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  and _56733_ (_05424_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and _56734_ (_05426_, _05424_, _05423_);
  nand _56735_ (_05427_, _05426_, _00612_);
  nand _56736_ (_05428_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _56737_ (_05430_, _05428_, _05408_);
  or _56738_ (_05431_, _05430_, _00558_);
  and _56739_ (_05432_, _05431_, _05427_);
  or _56740_ (_05434_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _56741_ (_05435_, _05434_, _05402_);
  or _56742_ (_05436_, _05435_, _00070_);
  or _56743_ (_05438_, _05434_, _05408_);
  or _56744_ (_05439_, _05438_, _00029_);
  and _56745_ (_05440_, _05439_, _05436_);
  and _56746_ (_05442_, _05440_, _05432_);
  and _56747_ (_05443_, _05442_, _05422_);
  not _56748_ (_05444_, \oc8051_golden_model_1.PC [0]);
  or _56749_ (_05446_, \oc8051_golden_model_1.PC [1], _05444_);
  or _56750_ (_05447_, _05446_, _05428_);
  or _56751_ (_05448_, _05447_, _00511_);
  or _56752_ (_05449_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or _56753_ (_05450_, _05449_, _05428_);
  or _56754_ (_05451_, _05450_, _00470_);
  and _56755_ (_05452_, _05451_, _05448_);
  or _56756_ (_05453_, _05434_, _05449_);
  or _56757_ (_05454_, _05453_, _43974_);
  or _56758_ (_05455_, _05434_, _05446_);
  or _56759_ (_05456_, _05455_, _44015_);
  and _56760_ (_05457_, _05456_, _05454_);
  and _56761_ (_05458_, _05457_, _05452_);
  or _56762_ (_05459_, _05446_, _05404_);
  or _56763_ (_05460_, _05459_, _00347_);
  or _56764_ (_05461_, _05449_, _05404_);
  or _56765_ (_05462_, _05461_, _00306_);
  and _56766_ (_05463_, _05462_, _05460_);
  or _56767_ (_05464_, _05446_, _05413_);
  or _56768_ (_05465_, _05464_, _00178_);
  or _56769_ (_05466_, _05449_, _05413_);
  or _56770_ (_05468_, _05466_, _00111_);
  and _56771_ (_05469_, _05468_, _05465_);
  and _56772_ (_05471_, _05469_, _05463_);
  and _56773_ (_05472_, _05471_, _05458_);
  and _56774_ (_05473_, _05472_, _05443_);
  or _56775_ (_05475_, _05405_, _00394_);
  or _56776_ (_05476_, _05409_, _00353_);
  and _56777_ (_05477_, _05476_, _05475_);
  or _56778_ (_05479_, _05415_, _00230_);
  or _56779_ (_05480_, _05418_, _00189_);
  and _56780_ (_05481_, _05480_, _05479_);
  and _56781_ (_05483_, _05481_, _05477_);
  nand _56782_ (_05484_, _05426_, _00567_);
  or _56783_ (_05485_, _05430_, _00517_);
  and _56784_ (_05487_, _05485_, _05484_);
  or _56785_ (_05488_, _05435_, _00035_);
  or _56786_ (_05489_, _05438_, _44021_);
  and _56787_ (_05491_, _05489_, _05488_);
  and _56788_ (_05492_, _05491_, _05487_);
  and _56789_ (_05493_, _05492_, _05483_);
  or _56790_ (_05495_, _05447_, _00476_);
  or _56791_ (_05496_, _05450_, _00435_);
  and _56792_ (_05497_, _05496_, _05495_);
  or _56793_ (_05499_, _05453_, _43939_);
  or _56794_ (_05500_, _05455_, _43980_);
  and _56795_ (_05501_, _05500_, _05499_);
  and _56796_ (_05502_, _05501_, _05497_);
  or _56797_ (_05503_, _05459_, _00312_);
  or _56798_ (_05504_, _05461_, _00271_);
  and _56799_ (_05505_, _05504_, _05503_);
  or _56800_ (_05506_, _05464_, _00117_);
  or _56801_ (_05507_, _05466_, _00076_);
  and _56802_ (_05508_, _05507_, _05506_);
  and _56803_ (_05509_, _05508_, _05505_);
  and _56804_ (_05510_, _05509_, _05502_);
  and _56805_ (_05511_, _05510_, _05493_);
  and _56806_ (_05512_, _05511_, _05473_);
  or _56807_ (_05513_, _05405_, _00419_);
  or _56808_ (_05514_, _05409_, _00378_);
  and _56809_ (_05515_, _05514_, _05513_);
  or _56810_ (_05516_, _05415_, _00255_);
  or _56811_ (_05517_, _05418_, _00214_);
  and _56812_ (_05518_, _05517_, _05516_);
  and _56813_ (_05519_, _05518_, _05515_);
  nand _56814_ (_05521_, _05426_, _00602_);
  or _56815_ (_05522_, _05430_, _00542_);
  and _56816_ (_05524_, _05522_, _05521_);
  or _56817_ (_05525_, _05435_, _00060_);
  or _56818_ (_05526_, _05438_, _00019_);
  and _56819_ (_05528_, _05526_, _05525_);
  and _56820_ (_05529_, _05528_, _05524_);
  and _56821_ (_05530_, _05529_, _05519_);
  or _56822_ (_05532_, _05447_, _00501_);
  or _56823_ (_05533_, _05450_, _00460_);
  and _56824_ (_05534_, _05533_, _05532_);
  or _56825_ (_05536_, _05453_, _43964_);
  or _56826_ (_05537_, _05455_, _44005_);
  and _56827_ (_05538_, _05537_, _05536_);
  and _56828_ (_05540_, _05538_, _05534_);
  or _56829_ (_05541_, _05459_, _00337_);
  or _56830_ (_05542_, _05461_, _00296_);
  and _56831_ (_05544_, _05542_, _05541_);
  or _56832_ (_05545_, _05464_, _00156_);
  or _56833_ (_05546_, _05466_, _00101_);
  and _56834_ (_05548_, _05546_, _05545_);
  and _56835_ (_05549_, _05548_, _05544_);
  and _56836_ (_05550_, _05549_, _05540_);
  and _56837_ (_05552_, _05550_, _05530_);
  or _56838_ (_05553_, _05405_, _00424_);
  or _56839_ (_05554_, _05409_, _00383_);
  and _56840_ (_05555_, _05554_, _05553_);
  or _56841_ (_05556_, _05415_, _00260_);
  or _56842_ (_05557_, _05418_, _00219_);
  and _56843_ (_05558_, _05557_, _05556_);
  and _56844_ (_05559_, _05558_, _05555_);
  nand _56845_ (_05560_, _05426_, _00607_);
  or _56846_ (_05561_, _05430_, _00550_);
  and _56847_ (_05562_, _05561_, _05560_);
  or _56848_ (_05563_, _05435_, _00065_);
  or _56849_ (_05564_, _05438_, _00024_);
  and _56850_ (_05565_, _05564_, _05563_);
  and _56851_ (_05566_, _05565_, _05562_);
  and _56852_ (_05567_, _05566_, _05559_);
  or _56853_ (_05568_, _05447_, _00506_);
  or _56854_ (_05569_, _05450_, _00465_);
  and _56855_ (_05570_, _05569_, _05568_);
  or _56856_ (_05571_, _05453_, _43969_);
  or _56857_ (_05572_, _05455_, _44010_);
  and _56858_ (_05574_, _05572_, _05571_);
  and _56859_ (_05575_, _05574_, _05570_);
  or _56860_ (_05577_, _05459_, _00342_);
  or _56861_ (_05578_, _05461_, _00301_);
  and _56862_ (_05579_, _05578_, _05577_);
  or _56863_ (_05581_, _05464_, _00167_);
  or _56864_ (_05582_, _05466_, _00106_);
  and _56865_ (_05583_, _05582_, _05581_);
  and _56866_ (_05585_, _05583_, _05579_);
  and _56867_ (_05586_, _05585_, _05575_);
  nand _56868_ (_05587_, _05586_, _05567_);
  or _56869_ (_05589_, _05587_, _05552_);
  not _56870_ (_05590_, _05589_);
  and _56871_ (_05591_, _05590_, _05512_);
  or _56872_ (_05593_, _05405_, _00409_);
  or _56873_ (_05594_, _05409_, _00368_);
  and _56874_ (_05595_, _05594_, _05593_);
  or _56875_ (_05597_, _05415_, _00245_);
  or _56876_ (_05598_, _05418_, _00204_);
  and _56877_ (_05599_, _05598_, _05597_);
  and _56878_ (_05601_, _05599_, _05595_);
  nand _56879_ (_05602_, _05426_, _00591_);
  or _56880_ (_05603_, _05430_, _00532_);
  and _56881_ (_05605_, _05603_, _05602_);
  or _56882_ (_05606_, _05435_, _00050_);
  or _56883_ (_05607_, _05438_, _00009_);
  and _56884_ (_05608_, _05607_, _05606_);
  and _56885_ (_05609_, _05608_, _05605_);
  and _56886_ (_05610_, _05609_, _05601_);
  or _56887_ (_05611_, _05447_, _00491_);
  or _56888_ (_05612_, _05450_, _00450_);
  and _56889_ (_05613_, _05612_, _05611_);
  or _56890_ (_05614_, _05453_, _43954_);
  or _56891_ (_05615_, _05455_, _43995_);
  and _56892_ (_05616_, _05615_, _05614_);
  and _56893_ (_05617_, _05616_, _05613_);
  or _56894_ (_05618_, _05459_, _00327_);
  or _56895_ (_05619_, _05461_, _00286_);
  and _56896_ (_05620_, _05619_, _05618_);
  or _56897_ (_05621_, _05464_, _00134_);
  or _56898_ (_05622_, _05466_, _00091_);
  and _56899_ (_05623_, _05622_, _05621_);
  and _56900_ (_05624_, _05623_, _05620_);
  and _56901_ (_05625_, _05624_, _05617_);
  nand _56902_ (_05627_, _05625_, _05610_);
  or _56903_ (_05628_, _05405_, _00414_);
  or _56904_ (_05630_, _05409_, _00373_);
  and _56905_ (_05631_, _05630_, _05628_);
  or _56906_ (_05632_, _05415_, _00250_);
  or _56907_ (_05634_, _05418_, _00209_);
  and _56908_ (_05635_, _05634_, _05632_);
  and _56909_ (_05636_, _05635_, _05631_);
  nand _56910_ (_05638_, _05426_, _00597_);
  or _56911_ (_05639_, _05430_, _00537_);
  and _56912_ (_05640_, _05639_, _05638_);
  or _56913_ (_05642_, _05435_, _00055_);
  or _56914_ (_05643_, _05438_, _00014_);
  and _56915_ (_05644_, _05643_, _05642_);
  and _56916_ (_05646_, _05644_, _05640_);
  and _56917_ (_05647_, _05646_, _05636_);
  or _56918_ (_05648_, _05447_, _00496_);
  or _56919_ (_05650_, _05450_, _00455_);
  and _56920_ (_05651_, _05650_, _05648_);
  or _56921_ (_05652_, _05453_, _43959_);
  or _56922_ (_05654_, _05455_, _44000_);
  and _56923_ (_05655_, _05654_, _05652_);
  and _56924_ (_05656_, _05655_, _05651_);
  or _56925_ (_05658_, _05459_, _00332_);
  or _56926_ (_05659_, _05461_, _00291_);
  and _56927_ (_05660_, _05659_, _05658_);
  or _56928_ (_05661_, _05464_, _00145_);
  or _56929_ (_05662_, _05466_, _00096_);
  and _56930_ (_05663_, _05662_, _05661_);
  and _56931_ (_05664_, _05663_, _05660_);
  and _56932_ (_05665_, _05664_, _05656_);
  nand _56933_ (_05666_, _05665_, _05647_);
  or _56934_ (_05667_, _05666_, _05627_);
  not _56935_ (_05668_, _05667_);
  or _56936_ (_05669_, _05405_, _00399_);
  or _56937_ (_05670_, _05409_, _00358_);
  and _56938_ (_05671_, _05670_, _05669_);
  or _56939_ (_05672_, _05415_, _00235_);
  or _56940_ (_05673_, _05418_, _00194_);
  and _56941_ (_05674_, _05673_, _05672_);
  and _56942_ (_05675_, _05674_, _05671_);
  nand _56943_ (_05676_, _05426_, _00575_);
  or _56944_ (_05677_, _05430_, _00522_);
  and _56945_ (_05678_, _05677_, _05676_);
  or _56946_ (_05680_, _05435_, _00040_);
  or _56947_ (_05681_, _05438_, _44026_);
  and _56948_ (_05683_, _05681_, _05680_);
  and _56949_ (_05684_, _05683_, _05678_);
  and _56950_ (_05685_, _05684_, _05675_);
  or _56951_ (_05687_, _05447_, _00481_);
  or _56952_ (_05688_, _05450_, _00440_);
  and _56953_ (_05689_, _05688_, _05687_);
  or _56954_ (_05691_, _05453_, _43944_);
  or _56955_ (_05692_, _05455_, _43985_);
  and _56956_ (_05693_, _05692_, _05691_);
  and _56957_ (_05695_, _05693_, _05689_);
  or _56958_ (_05696_, _05459_, _00317_);
  or _56959_ (_05697_, _05461_, _00276_);
  and _56960_ (_05699_, _05697_, _05696_);
  or _56961_ (_05700_, _05464_, _00122_);
  or _56962_ (_05701_, _05466_, _00081_);
  and _56963_ (_05703_, _05701_, _05700_);
  and _56964_ (_05704_, _05703_, _05699_);
  and _56965_ (_05705_, _05704_, _05695_);
  and _56966_ (_05707_, _05705_, _05685_);
  or _56967_ (_05708_, _05405_, _00404_);
  or _56968_ (_05709_, _05409_, _00363_);
  and _56969_ (_05711_, _05709_, _05708_);
  or _56970_ (_05712_, _05415_, _00240_);
  or _56971_ (_05713_, _05418_, _00199_);
  and _56972_ (_05714_, _05713_, _05712_);
  and _56973_ (_05715_, _05714_, _05711_);
  nand _56974_ (_05716_, _05426_, _00583_);
  or _56975_ (_05717_, _05430_, _00527_);
  and _56976_ (_05718_, _05717_, _05716_);
  or _56977_ (_05719_, _05435_, _00045_);
  or _56978_ (_05720_, _05438_, _00004_);
  and _56979_ (_05721_, _05720_, _05719_);
  and _56980_ (_05722_, _05721_, _05718_);
  and _56981_ (_05723_, _05722_, _05715_);
  or _56982_ (_05724_, _05447_, _00486_);
  or _56983_ (_05725_, _05450_, _00445_);
  and _56984_ (_05726_, _05725_, _05724_);
  or _56985_ (_05727_, _05453_, _43949_);
  or _56986_ (_05728_, _05455_, _43990_);
  and _56987_ (_05729_, _05728_, _05727_);
  and _56988_ (_05730_, _05729_, _05726_);
  or _56989_ (_05731_, _05459_, _00322_);
  or _56990_ (_05733_, _05461_, _00281_);
  and _56991_ (_05734_, _05733_, _05731_);
  or _56992_ (_05736_, _05464_, _00127_);
  or _56993_ (_05737_, _05466_, _00086_);
  and _56994_ (_05738_, _05737_, _05736_);
  and _56995_ (_05740_, _05738_, _05734_);
  and _56996_ (_05741_, _05740_, _05730_);
  nand _56997_ (_05742_, _05741_, _05723_);
  not _56998_ (_05744_, _05742_);
  and _56999_ (_05745_, _05744_, _05707_);
  and _57000_ (_05746_, _05745_, _05668_);
  and _57001_ (_05748_, _05746_, _05591_);
  not _57002_ (_05749_, _05748_);
  or _57003_ (_05750_, _05742_, _05707_);
  or _57004_ (_05752_, _05750_, _05667_);
  and _57005_ (_05753_, _05586_, _05567_);
  or _57006_ (_05754_, _05753_, _05552_);
  nand _57007_ (_05756_, _05472_, _05443_);
  or _57008_ (_05757_, _05511_, _05756_);
  or _57009_ (_05758_, _05757_, _05754_);
  or _57010_ (_05760_, _05758_, _05752_);
  or _57011_ (_05761_, _05511_, _05473_);
  or _57012_ (_05762_, _05761_, _05589_);
  or _57013_ (_05764_, _05762_, _05752_);
  and _57014_ (_05765_, _05764_, _05760_);
  nand _57015_ (_05766_, _05550_, _05530_);
  or _57016_ (_05767_, _05587_, _05766_);
  or _57017_ (_05768_, _05767_, _05761_);
  or _57018_ (_05769_, _05768_, _05752_);
  or _57019_ (_05770_, _05753_, _05766_);
  or _57020_ (_05771_, _05770_, _05761_);
  or _57021_ (_05772_, _05771_, _05752_);
  and _57022_ (_05773_, _05772_, _05769_);
  or _57023_ (_05774_, _05770_, _05757_);
  or _57024_ (_05775_, _05774_, _05752_);
  or _57025_ (_05776_, _05761_, _05754_);
  or _57026_ (_05777_, _05776_, _05752_);
  and _57027_ (_05778_, _05777_, _05775_);
  and _57028_ (_05779_, _05778_, _05773_);
  and _57029_ (_05780_, _05779_, _05765_);
  nor _57030_ (_05781_, _05767_, _05757_);
  not _57031_ (_05782_, _05750_);
  not _57032_ (_05783_, _05666_);
  and _57033_ (_05784_, _05783_, _05627_);
  and _57034_ (_05786_, _05784_, _05782_);
  and _57035_ (_05787_, _05786_, _05781_);
  not _57036_ (_05789_, _05752_);
  nor _57037_ (_05790_, _05757_, _05589_);
  and _57038_ (_05791_, _05790_, _05789_);
  nor _57039_ (_05793_, _05791_, _05787_);
  and _57040_ (_05794_, _05793_, _05780_);
  or _57041_ (_05795_, _05794_, \oc8051_golden_model_1.PC [0]);
  not _57042_ (_05797_, _05781_);
  or _57043_ (_05798_, _05744_, _05707_);
  or _57044_ (_05799_, _05798_, _05667_);
  nor _57045_ (_05801_, _05799_, _05797_);
  not _57046_ (_05802_, _05801_);
  not _57047_ (_05803_, _05790_);
  or _57048_ (_05805_, _05799_, _05803_);
  and _57049_ (_05806_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _57050_ (_05807_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _57051_ (_05809_, _05807_, _05806_);
  or _57052_ (_05810_, _05809_, _05805_);
  and _57053_ (_05811_, _05805_, \oc8051_golden_model_1.PC [0]);
  nand _57054_ (_05813_, _05811_, _05780_);
  nand _57055_ (_05814_, _05813_, _05810_);
  nand _57056_ (_05815_, _05814_, _05793_);
  and _57057_ (_05817_, _05815_, _05802_);
  nand _57058_ (_05818_, _05817_, _05795_);
  not _57059_ (_05819_, _05767_);
  and _57060_ (_05820_, _05819_, _05512_);
  and _57061_ (_05821_, _05820_, _05789_);
  not _57062_ (_05822_, _05821_);
  and _57063_ (_05823_, _05789_, _05591_);
  not _57064_ (_05824_, _05512_);
  nor _57065_ (_05825_, _05770_, _05824_);
  and _57066_ (_05826_, _05825_, _05789_);
  nor _57067_ (_05827_, _05826_, _05823_);
  and _57068_ (_05828_, _05827_, _05822_);
  and _57069_ (_05829_, _05781_, _05789_);
  not _57070_ (_05830_, _05829_);
  and _57071_ (_05831_, _05511_, _05756_);
  not _57072_ (_05832_, _05831_);
  or _57073_ (_05833_, _05832_, _05770_);
  or _57074_ (_05834_, _05833_, _05752_);
  or _57075_ (_05835_, _05832_, _05754_);
  or _57076_ (_05836_, _05835_, _05752_);
  and _57077_ (_05837_, _05836_, _05834_);
  and _57078_ (_05839_, _05837_, _05830_);
  and _57079_ (_05840_, _05831_, _05819_);
  and _57080_ (_05842_, _05840_, _05789_);
  not _57081_ (_05843_, _05842_);
  or _57082_ (_05844_, _05754_, _05824_);
  or _57083_ (_05846_, _05844_, _05752_);
  or _57084_ (_05847_, _05832_, _05589_);
  or _57085_ (_05848_, _05847_, _05752_);
  and _57086_ (_05850_, _05848_, _05846_);
  and _57087_ (_05851_, _05850_, _05843_);
  and _57088_ (_05852_, _05851_, _05839_);
  and _57089_ (_05854_, _05852_, _05828_);
  not _57090_ (_05855_, \oc8051_golden_model_1.ACC [0]);
  and _57091_ (_05856_, _05855_, \oc8051_golden_model_1.PC [0]);
  and _57092_ (_05858_, \oc8051_golden_model_1.ACC [0], _05444_);
  or _57093_ (_05859_, _05858_, _05802_);
  or _57094_ (_05860_, _05859_, _05856_);
  and _57095_ (_05862_, _05860_, _05854_);
  nand _57096_ (_05863_, _05862_, _05818_);
  nor _57097_ (_05864_, _05854_, \oc8051_golden_model_1.PC [0]);
  not _57098_ (_05866_, _05864_);
  and _57099_ (_05867_, _05866_, _05863_);
  or _57100_ (_05868_, _05794_, \oc8051_golden_model_1.PC [1]);
  not _57101_ (_05870_, _05805_);
  and _57102_ (_05871_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _57103_ (_05872_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _57104_ (_05873_, _05872_, _05871_);
  and _57105_ (_05874_, _05873_, _05806_);
  nor _57106_ (_05875_, _05873_, _05806_);
  nor _57107_ (_05876_, _05875_, _05874_);
  and _57108_ (_05877_, _05876_, _05870_);
  and _57109_ (_05878_, _05446_, _05408_);
  not _57110_ (_05879_, _05878_);
  and _57111_ (_05880_, _05879_, _05805_);
  and _57112_ (_05881_, _05880_, _05780_);
  or _57113_ (_05882_, _05881_, _05877_);
  and _57114_ (_05883_, _05854_, _05793_);
  nand _57115_ (_05884_, _05883_, _05882_);
  nand _57116_ (_05885_, _05884_, _05868_);
  nand _57117_ (_05886_, _05885_, _05802_);
  not _57118_ (_05887_, \oc8051_golden_model_1.ACC [1]);
  nor _57119_ (_05888_, _05878_, _05887_);
  and _57120_ (_05889_, _05878_, _05887_);
  nor _57121_ (_05890_, _05889_, _05888_);
  and _57122_ (_05892_, _05890_, _05858_);
  nor _57123_ (_05893_, _05890_, _05858_);
  nor _57124_ (_05895_, _05893_, _05892_);
  and _57125_ (_05896_, _05895_, _05801_);
  nor _57126_ (_05897_, _05854_, \oc8051_golden_model_1.PC [1]);
  nor _57127_ (_05899_, _05897_, _05896_);
  and _57128_ (_05900_, _05899_, _05886_);
  or _57129_ (_05901_, _05900_, _05867_);
  nor _57130_ (_05903_, _05892_, _05888_);
  and _57131_ (_05904_, _05423_, \oc8051_golden_model_1.PC [2]);
  and _57132_ (_05905_, _05402_, _05412_);
  nor _57133_ (_05907_, _05905_, _05904_);
  and _57134_ (_05908_, _05907_, \oc8051_golden_model_1.ACC [2]);
  nor _57135_ (_05909_, _05907_, \oc8051_golden_model_1.ACC [2]);
  nor _57136_ (_05911_, _05909_, _05908_);
  not _57137_ (_05912_, _05911_);
  and _57138_ (_05913_, _05912_, _05903_);
  nor _57139_ (_05915_, _05912_, _05903_);
  nor _57140_ (_05916_, _05915_, _05913_);
  and _57141_ (_05917_, _05916_, _05801_);
  and _57142_ (_05919_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _57143_ (_05920_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _57144_ (_05921_, _05920_, _05919_);
  not _57145_ (_05923_, _05921_);
  or _57146_ (_05924_, _05923_, _05780_);
  nand _57147_ (_05925_, _05907_, _05780_);
  nand _57148_ (_05926_, _05925_, _05924_);
  nand _57149_ (_05927_, _05926_, _05805_);
  nor _57150_ (_05928_, _05874_, _05871_);
  and _57151_ (_05929_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _57152_ (_05930_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _57153_ (_05931_, _05930_, _05929_);
  not _57154_ (_05932_, _05931_);
  nor _57155_ (_05933_, _05932_, _05928_);
  and _57156_ (_05934_, _05932_, _05928_);
  nor _57157_ (_05935_, _05934_, _05933_);
  not _57158_ (_05936_, _05935_);
  or _57159_ (_05937_, _05936_, _05805_);
  and _57160_ (_05938_, _05937_, _05793_);
  nand _57161_ (_05939_, _05938_, _05927_);
  or _57162_ (_05940_, _05921_, _05793_);
  and _57163_ (_05941_, _05940_, _05802_);
  and _57164_ (_05942_, _05941_, _05939_);
  or _57165_ (_05943_, _05942_, _05917_);
  nand _57166_ (_05944_, _05943_, _05854_);
  nor _57167_ (_05945_, _05923_, _05854_);
  not _57168_ (_05946_, _05945_);
  and _57169_ (_05947_, _05946_, _05944_);
  nor _57170_ (_05948_, _05915_, _05908_);
  not _57171_ (_05949_, _05415_);
  nor _57172_ (_05950_, _05904_, _05403_);
  nor _57173_ (_05951_, _05950_, _05949_);
  nor _57174_ (_05952_, _05951_, \oc8051_golden_model_1.ACC [3]);
  and _57175_ (_05953_, _05951_, \oc8051_golden_model_1.ACC [3]);
  nor _57176_ (_05954_, _05953_, _05952_);
  and _57177_ (_05955_, _05954_, _05948_);
  nor _57178_ (_05956_, _05954_, _05948_);
  nor _57179_ (_05957_, _05956_, _05955_);
  and _57180_ (_05958_, _05957_, _05801_);
  and _57181_ (_05959_, _05805_, _05951_);
  nand _57182_ (_05960_, _05959_, _05780_);
  nor _57183_ (_05961_, _05933_, _05929_);
  and _57184_ (_05962_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _57185_ (_05963_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _57186_ (_05964_, _05963_, _05962_);
  not _57187_ (_05965_, _05964_);
  nor _57188_ (_05966_, _05965_, _05961_);
  and _57189_ (_05967_, _05965_, _05961_);
  nor _57190_ (_05968_, _05967_, _05966_);
  or _57191_ (_05969_, _05968_, _05805_);
  nand _57192_ (_05970_, _05969_, _05960_);
  nand _57193_ (_05971_, _05970_, _05793_);
  and _57194_ (_05972_, _05424_, \oc8051_golden_model_1.PC [1]);
  nor _57195_ (_05973_, _05919_, \oc8051_golden_model_1.PC [3]);
  nor _57196_ (_05974_, _05973_, _05972_);
  or _57197_ (_05975_, _05974_, _05794_);
  and _57198_ (_05976_, _05975_, _05971_);
  nand _57199_ (_05977_, _05976_, _05802_);
  nand _57200_ (_05978_, _05977_, _05854_);
  nor _57201_ (_05979_, _05978_, _05958_);
  nor _57202_ (_05980_, _05974_, _05854_);
  or _57203_ (_05981_, _05980_, _05979_);
  or _57204_ (_05982_, _05981_, _05947_);
  or _57205_ (_05983_, _05982_, _05901_);
  or _57206_ (_05984_, _05983_, _00517_);
  nand _57207_ (_05985_, _05866_, _05863_);
  nand _57208_ (_05986_, _05899_, _05886_);
  or _57209_ (_05987_, _05986_, _05985_);
  or _57210_ (_05988_, _05987_, _05982_);
  or _57211_ (_05989_, _05988_, _00476_);
  and _57212_ (_05990_, _05989_, _05984_);
  or _57213_ (_05991_, _05900_, _05985_);
  nor _57214_ (_05992_, _05980_, _05979_);
  or _57215_ (_05993_, _05992_, _05947_);
  or _57216_ (_05994_, _05993_, _05991_);
  or _57217_ (_05995_, _05994_, _00230_);
  nand _57218_ (_05996_, _05946_, _05944_);
  or _57219_ (_05997_, _05992_, _05996_);
  or _57220_ (_05998_, _05997_, _05991_);
  or _57221_ (_05999_, _05998_, _00035_);
  and _57222_ (_06000_, _05999_, _05995_);
  and _57223_ (_06001_, _06000_, _05990_);
  or _57224_ (_06002_, _05997_, _05901_);
  or _57225_ (_06003_, _06002_, _44021_);
  or _57226_ (_06004_, _05997_, _05987_);
  or _57227_ (_06005_, _06004_, _43980_);
  and _57228_ (_06006_, _06005_, _06003_);
  or _57229_ (_06007_, _05993_, _05901_);
  or _57230_ (_06008_, _06007_, _00189_);
  or _57231_ (_06009_, _05986_, _05867_);
  or _57232_ (_06010_, _06009_, _05993_);
  or _57233_ (_06011_, _06010_, _00076_);
  and _57234_ (_06012_, _06011_, _06008_);
  and _57235_ (_06013_, _06012_, _06006_);
  and _57236_ (_06014_, _06013_, _06001_);
  or _57237_ (_06015_, _05981_, _05996_);
  or _57238_ (_06016_, _06015_, _05901_);
  or _57239_ (_06017_, _06016_, _00353_);
  or _57240_ (_06018_, _06015_, _06009_);
  or _57241_ (_06019_, _06018_, _00271_);
  and _57242_ (_06020_, _06019_, _06017_);
  nor _57243_ (_06021_, _05991_, _05982_);
  nand _57244_ (_06022_, _06021_, _00567_);
  or _57245_ (_06023_, _06009_, _05982_);
  or _57246_ (_06024_, _06023_, _00435_);
  and _57247_ (_06025_, _06024_, _06022_);
  and _57248_ (_06026_, _06025_, _06020_);
  or _57249_ (_06027_, _05993_, _05987_);
  or _57250_ (_06028_, _06027_, _00117_);
  or _57251_ (_06029_, _06009_, _05997_);
  or _57252_ (_06030_, _06029_, _43939_);
  and _57253_ (_06031_, _06030_, _06028_);
  or _57254_ (_06032_, _06015_, _05991_);
  or _57255_ (_06033_, _06032_, _00394_);
  or _57256_ (_06034_, _06015_, _05987_);
  or _57257_ (_06035_, _06034_, _00312_);
  and _57258_ (_06036_, _06035_, _06033_);
  and _57259_ (_06037_, _06036_, _06031_);
  and _57260_ (_06038_, _06037_, _06026_);
  nand _57261_ (_06039_, _06038_, _06014_);
  nand _57262_ (_06040_, _06021_, _00597_);
  or _57263_ (_06041_, _05998_, _00055_);
  and _57264_ (_06042_, _06041_, _06040_);
  or _57265_ (_06043_, _05983_, _00537_);
  or _57266_ (_06044_, _06034_, _00332_);
  and _57267_ (_06045_, _06044_, _06043_);
  and _57268_ (_06046_, _06045_, _06042_);
  or _57269_ (_06047_, _06032_, _00414_);
  or _57270_ (_06048_, _05994_, _00250_);
  and _57271_ (_06049_, _06048_, _06047_);
  or _57272_ (_06050_, _06007_, _00209_);
  or _57273_ (_06051_, _06004_, _44000_);
  and _57274_ (_06052_, _06051_, _06050_);
  and _57275_ (_06053_, _06052_, _06049_);
  and _57276_ (_06054_, _06053_, _06046_);
  or _57277_ (_06055_, _05988_, _00496_);
  or _57278_ (_06056_, _06023_, _00455_);
  and _57279_ (_06057_, _06056_, _06055_);
  or _57280_ (_06058_, _06018_, _00291_);
  or _57281_ (_06059_, _06027_, _00145_);
  and _57282_ (_06060_, _06059_, _06058_);
  and _57283_ (_06061_, _06060_, _06057_);
  or _57284_ (_06062_, _06016_, _00373_);
  or _57285_ (_06063_, _06002_, _00014_);
  and _57286_ (_06064_, _06063_, _06062_);
  or _57287_ (_06065_, _06010_, _00096_);
  or _57288_ (_06066_, _06029_, _43959_);
  and _57289_ (_06067_, _06066_, _06065_);
  and _57290_ (_06068_, _06067_, _06064_);
  and _57291_ (_06069_, _06068_, _06061_);
  and _57292_ (_06070_, _06069_, _06054_);
  or _57293_ (_06071_, _06070_, _06039_);
  nor _57294_ (_06072_, _06071_, _05749_);
  nor _57295_ (_06073_, _06039_, _05749_);
  not _57296_ (_06074_, _06073_);
  nor _57297_ (_06075_, _05846_, \oc8051_golden_model_1.SP [0]);
  not _57298_ (_06076_, _05836_);
  or _57299_ (_06077_, _06007_, _00194_);
  or _57300_ (_06078_, _06027_, _00122_);
  and _57301_ (_06079_, _06078_, _06077_);
  or _57302_ (_06080_, _05998_, _00040_);
  or _57303_ (_06081_, _06002_, _44026_);
  and _57304_ (_06082_, _06081_, _06080_);
  and _57305_ (_06083_, _06082_, _06079_);
  or _57306_ (_06084_, _06034_, _00317_);
  or _57307_ (_06085_, _06018_, _00276_);
  and _57308_ (_06086_, _06085_, _06084_);
  or _57309_ (_06087_, _05988_, _00481_);
  or _57310_ (_06088_, _06023_, _00440_);
  and _57311_ (_06089_, _06088_, _06087_);
  and _57312_ (_06090_, _06089_, _06086_);
  and _57313_ (_06091_, _06090_, _06083_);
  or _57314_ (_06092_, _06029_, _43944_);
  or _57315_ (_06093_, _06004_, _43985_);
  and _57316_ (_06094_, _06093_, _06092_);
  or _57317_ (_06095_, _05994_, _00235_);
  or _57318_ (_06096_, _06010_, _00081_);
  and _57319_ (_06097_, _06096_, _06095_);
  and _57320_ (_06098_, _06097_, _06094_);
  nand _57321_ (_06099_, _06021_, _00575_);
  or _57322_ (_06100_, _05983_, _00522_);
  and _57323_ (_06101_, _06100_, _06099_);
  or _57324_ (_06102_, _06032_, _00399_);
  or _57325_ (_06103_, _06016_, _00358_);
  and _57326_ (_06104_, _06103_, _06102_);
  and _57327_ (_06105_, _06104_, _06101_);
  and _57328_ (_06106_, _06105_, _06098_);
  and _57329_ (_06107_, _06106_, _06091_);
  not _57330_ (_06108_, _06107_);
  not _57331_ (_06109_, _05835_);
  and _57332_ (_06110_, _06109_, _05786_);
  not _57333_ (_06111_, _06110_);
  nor _57334_ (_06112_, _06111_, _06039_);
  and _57335_ (_06113_, _06112_, _06108_);
  not _57336_ (_06114_, _05787_);
  and _57337_ (_06115_, _05784_, _05742_);
  and _57338_ (_06116_, _06115_, _05781_);
  not _57339_ (_06117_, _06116_);
  nor _57340_ (_06118_, _05783_, _05627_);
  and _57341_ (_06119_, _06118_, _05744_);
  and _57342_ (_06120_, _06119_, _05781_);
  not _57343_ (_06121_, _06120_);
  and _57344_ (_06122_, _05666_, _05627_);
  and _57345_ (_06123_, _06122_, _05782_);
  and _57346_ (_06124_, _06122_, _05742_);
  or _57347_ (_06125_, _06124_, _06123_);
  and _57348_ (_06126_, _06125_, _05781_);
  and _57349_ (_06127_, _06122_, _05745_);
  and _57350_ (_06128_, _06118_, _05742_);
  nor _57351_ (_06129_, _06128_, _06127_);
  nor _57352_ (_06130_, _06129_, _05797_);
  nor _57353_ (_06131_, _06130_, _06126_);
  and _57354_ (_06132_, _06131_, _06121_);
  and _57355_ (_06133_, _06132_, _06117_);
  and _57356_ (_06134_, _06133_, _06114_);
  nor _57357_ (_06135_, _06134_, _06039_);
  and _57358_ (_06136_, _06135_, _06107_);
  and _57359_ (_06137_, _05742_, _05707_);
  and _57360_ (_06138_, _06137_, _05668_);
  and _57361_ (_06139_, _06138_, _05790_);
  not _57362_ (_06140_, _06139_);
  nor _57363_ (_06141_, _06140_, _06071_);
  not _57364_ (_06142_, \oc8051_golden_model_1.SP [0]);
  nor _57365_ (_06143_, _05760_, _06142_);
  not _57366_ (_06144_, _05758_);
  and _57367_ (_06145_, _06138_, _06144_);
  not _57368_ (_06146_, _06145_);
  nor _57369_ (_06147_, _06146_, _06071_);
  nor _57370_ (_06148_, _06146_, _06039_);
  not _57371_ (_06149_, _06148_);
  not _57372_ (_06150_, _05768_);
  and _57373_ (_06151_, _06150_, _05746_);
  and _57374_ (_06152_, _06138_, _06150_);
  not _57375_ (_06153_, _06152_);
  nor _57376_ (_06154_, _06153_, _06071_);
  not _57377_ (_06155_, _05762_);
  and _57378_ (_06156_, _06138_, _06155_);
  not _57379_ (_06157_, _06156_);
  or _57380_ (_06158_, _06157_, _06071_);
  nor _57381_ (_06159_, _06157_, _06039_);
  and _57382_ (_06160_, _05786_, _06155_);
  not _57383_ (_06161_, _06160_);
  nor _57384_ (_06162_, _06161_, _06039_);
  and _57385_ (_06163_, _06162_, _06108_);
  not _57386_ (_06164_, _05777_);
  and _57387_ (_06165_, _05825_, _05746_);
  not _57388_ (_06166_, _06165_);
  and _57389_ (_06167_, _06138_, _05825_);
  not _57390_ (_06168_, _06167_);
  and _57391_ (_06169_, _05825_, _05786_);
  and _57392_ (_06170_, _06169_, _06070_);
  not _57393_ (_06171_, _06169_);
  not _57394_ (_06172_, _06039_);
  and _57395_ (_06173_, _06021_, _00612_);
  nor _57396_ (_06174_, _06027_, _00178_);
  nor _57397_ (_06175_, _06174_, _06173_);
  nor _57398_ (_06176_, _05983_, _00558_);
  nor _57399_ (_06177_, _06018_, _00306_);
  nor _57400_ (_06178_, _06177_, _06176_);
  and _57401_ (_06179_, _06178_, _06175_);
  nor _57402_ (_06180_, _06004_, _44015_);
  nor _57403_ (_06181_, _06002_, _00029_);
  nor _57404_ (_06182_, _06181_, _06180_);
  nor _57405_ (_06183_, _06032_, _00429_);
  nor _57406_ (_06184_, _05998_, _00070_);
  nor _57407_ (_06185_, _06184_, _06183_);
  and _57408_ (_06186_, _06185_, _06182_);
  and _57409_ (_06187_, _06186_, _06179_);
  nor _57410_ (_06188_, _05988_, _00511_);
  nor _57411_ (_06189_, _06023_, _00470_);
  nor _57412_ (_06190_, _06189_, _06188_);
  nor _57413_ (_06191_, _06034_, _00347_);
  nor _57414_ (_06192_, _05994_, _00265_);
  nor _57415_ (_06193_, _06192_, _06191_);
  and _57416_ (_06194_, _06193_, _06190_);
  nor _57417_ (_06195_, _06016_, _00388_);
  nor _57418_ (_06196_, _06007_, _00224_);
  nor _57419_ (_06197_, _06196_, _06195_);
  nor _57420_ (_06198_, _06010_, _00111_);
  nor _57421_ (_06199_, _06029_, _43974_);
  nor _57422_ (_06200_, _06199_, _06198_);
  and _57423_ (_06201_, _06200_, _06197_);
  and _57424_ (_06202_, _06201_, _06194_);
  and _57425_ (_06203_, _06202_, _06187_);
  and _57426_ (_06204_, _06203_, _06172_);
  and _57427_ (_06205_, _06070_, _06039_);
  or _57428_ (_06206_, _06205_, _06204_);
  not _57429_ (_06207_, _06206_);
  and _57430_ (_06208_, _06138_, _06109_);
  and _57431_ (_06209_, _06138_, _05781_);
  nor _57432_ (_06210_, _06209_, _06208_);
  nor _57433_ (_06211_, _06210_, _06207_);
  and _57434_ (_06212_, _06144_, _05746_);
  nor _57435_ (_06213_, _06145_, _06212_);
  or _57436_ (_06214_, _06213_, _06206_);
  and _57437_ (_06215_, _06206_, _06156_);
  not _57438_ (_06216_, \oc8051_golden_model_1.SP [3]);
  and _57439_ (_06217_, _06155_, _05746_);
  and _57440_ (_06218_, _06217_, _06216_);
  or _57441_ (_06219_, _06218_, _06215_);
  and _57442_ (_06220_, _05786_, _06150_);
  nor _57443_ (_06221_, _06217_, _06156_);
  not _57444_ (_06222_, _05771_);
  and _57445_ (_06223_, _05786_, _06222_);
  nor _57446_ (_06224_, _06223_, _06160_);
  nand _57447_ (_06225_, _06224_, \oc8051_golden_model_1.PSW [3]);
  and _57448_ (_06226_, _06225_, _06221_);
  or _57449_ (_06227_, _06226_, _06220_);
  not _57450_ (_06228_, _06070_);
  not _57451_ (_06229_, _06220_);
  nand _57452_ (_06230_, _06224_, _06229_);
  nand _57453_ (_06231_, _06230_, _06228_);
  and _57454_ (_06232_, _06231_, _06227_);
  or _57455_ (_06233_, _06232_, _06152_);
  or _57456_ (_06234_, _06233_, _06219_);
  or _57457_ (_06235_, _06206_, _06153_);
  and _57458_ (_06236_, _05786_, _06144_);
  nor _57459_ (_06237_, _06236_, _06151_);
  and _57460_ (_06238_, _06237_, _06235_);
  and _57461_ (_06239_, _06238_, _06234_);
  not _57462_ (_06240_, _06213_);
  nor _57463_ (_06241_, _06237_, _06228_);
  or _57464_ (_06242_, _06241_, _06240_);
  or _57465_ (_06243_, _06242_, _06239_);
  and _57466_ (_06244_, _06243_, _06214_);
  not _57467_ (_06245_, _05774_);
  and _57468_ (_06246_, _06125_, _06245_);
  not _57469_ (_06247_, _06246_);
  and _57470_ (_06248_, _06127_, _06245_);
  and _57471_ (_06249_, _06118_, _06245_);
  nor _57472_ (_06250_, _06249_, _06248_);
  and _57473_ (_06251_, _06250_, _06247_);
  not _57474_ (_06252_, _06251_);
  or _57475_ (_06253_, _06252_, _06244_);
  and _57476_ (_06254_, _06245_, _05746_);
  and _57477_ (_06255_, _06138_, _06245_);
  nor _57478_ (_06256_, _06255_, _06254_);
  or _57479_ (_06257_, _06251_, _06070_);
  and _57480_ (_06258_, _06257_, _06256_);
  and _57481_ (_06259_, _06258_, _06253_);
  and _57482_ (_06260_, _05790_, _05786_);
  not _57483_ (_06261_, _06256_);
  and _57484_ (_06262_, _06261_, _06206_);
  or _57485_ (_06263_, _06262_, _06260_);
  or _57486_ (_06264_, _06263_, _06259_);
  not _57487_ (_06265_, _06260_);
  or _57488_ (_06266_, _06265_, _06070_);
  and _57489_ (_06267_, _06266_, _06140_);
  and _57490_ (_06268_, _06267_, _06264_);
  and _57491_ (_06269_, _06206_, _06139_);
  or _57492_ (_06270_, _06269_, _05787_);
  or _57493_ (_06271_, _06270_, _06268_);
  and _57494_ (_06272_, _06123_, _06144_);
  and _57495_ (_06273_, _06118_, _05745_);
  and _57496_ (_06274_, _06273_, _06144_);
  nor _57497_ (_06275_, _06274_, _06272_);
  not _57498_ (_06276_, _05707_);
  and _57499_ (_06277_, _06124_, _06276_);
  and _57500_ (_06278_, _06277_, _06144_);
  nor _57501_ (_06279_, _06278_, _06160_);
  and _57502_ (_06280_, _06279_, _06275_);
  and _57503_ (_06281_, _06137_, _05784_);
  and _57504_ (_06282_, _06281_, _06144_);
  not _57505_ (_06283_, _05798_);
  and _57506_ (_06284_, _06283_, _05784_);
  and _57507_ (_06285_, _06284_, _06144_);
  nor _57508_ (_06286_, _06285_, _06282_);
  and _57509_ (_06287_, _06286_, _06280_);
  and _57510_ (_06288_, _06118_, _05782_);
  and _57511_ (_06289_, _06288_, _06144_);
  nor _57512_ (_06290_, _06129_, _05758_);
  nor _57513_ (_06291_, _06290_, _06289_);
  and _57514_ (_06292_, _06291_, _06287_);
  and _57515_ (_06293_, _05790_, _05746_);
  and _57516_ (_06294_, _05784_, _05745_);
  and _57517_ (_06295_, _06294_, _06144_);
  nor _57518_ (_06296_, _06295_, _06293_);
  nor _57519_ (_06297_, _05833_, _05799_);
  nor _57520_ (_06298_, _06297_, _06110_);
  and _57521_ (_06299_, _06298_, _06296_);
  not _57522_ (_06300_, _05844_);
  and _57523_ (_06301_, _06300_, _05746_);
  not _57524_ (_06302_, _05799_);
  and _57525_ (_06303_, _05840_, _06302_);
  nor _57526_ (_06304_, _06303_, _06301_);
  and _57527_ (_06305_, _06138_, _05820_);
  nor _57528_ (_06306_, _05847_, _05799_);
  nor _57529_ (_06307_, _06306_, _06305_);
  and _57530_ (_06308_, _06307_, _06304_);
  and _57531_ (_06309_, _06308_, _06299_);
  and _57532_ (_06310_, _06138_, _05591_);
  nor _57533_ (_06311_, _06310_, _05748_);
  and _57534_ (_06312_, _06311_, _06166_);
  and _57535_ (_06313_, _06122_, _06137_);
  and _57536_ (_06314_, _06313_, _06144_);
  nor _57537_ (_06315_, _06314_, _06236_);
  and _57538_ (_06316_, _06315_, _06312_);
  and _57539_ (_06317_, _06316_, _06309_);
  and _57540_ (_06318_, _06317_, _06292_);
  nor _57541_ (_06319_, _06318_, _05923_);
  and _57542_ (_06320_, _06318_, _05907_);
  nor _57543_ (_06321_, _06320_, _06319_);
  not _57544_ (_06322_, _05974_);
  nor _57545_ (_06323_, _06318_, _06322_);
  not _57546_ (_06324_, _05951_);
  and _57547_ (_06325_, _06318_, _06324_);
  nor _57548_ (_06326_, _06325_, _06323_);
  nor _57549_ (_06327_, _06326_, _06321_);
  nor _57550_ (_06328_, _06318_, _05444_);
  and _57551_ (_06329_, _06318_, _05444_);
  nor _57552_ (_06330_, _06329_, _06328_);
  not _57553_ (_06331_, _06330_);
  nor _57554_ (_06332_, _06329_, _05407_);
  and _57555_ (_06333_, _06329_, _05407_);
  nor _57556_ (_06334_, _06333_, _06332_);
  and _57557_ (_06335_, _06334_, _06331_);
  and _57558_ (_06336_, _06335_, _06327_);
  and _57559_ (_06337_, _06336_, _00597_);
  nor _57560_ (_06338_, _06334_, _06330_);
  and _57561_ (_06339_, _06326_, _06321_);
  and _57562_ (_06340_, _06339_, _06338_);
  and _57563_ (_06341_, _06340_, _04563_);
  nor _57564_ (_06342_, _06341_, _06337_);
  not _57565_ (_06343_, _06321_);
  nor _57566_ (_06344_, _06326_, _06343_);
  and _57567_ (_06345_, _06344_, _06335_);
  and _57568_ (_06346_, _06345_, _04534_);
  nor _57569_ (_06347_, _06334_, _06331_);
  and _57570_ (_06348_, _06339_, _06347_);
  and _57571_ (_06349_, _06348_, _04553_);
  nor _57572_ (_06350_, _06349_, _06346_);
  and _57573_ (_06351_, _06350_, _06342_);
  and _57574_ (_06352_, _06344_, _06338_);
  and _57575_ (_06353_, _06352_, _04545_);
  and _57576_ (_06354_, _06334_, _06330_);
  and _57577_ (_06355_, _06339_, _06354_);
  and _57578_ (_06356_, _06355_, _04559_);
  nor _57579_ (_06357_, _06356_, _06353_);
  and _57580_ (_06358_, _06326_, _06343_);
  and _57581_ (_06359_, _06358_, _06335_);
  and _57582_ (_06360_, _06359_, _04569_);
  and _57583_ (_06361_, _06358_, _06347_);
  and _57584_ (_06362_, _06361_, _04540_);
  nor _57585_ (_06363_, _06362_, _06360_);
  and _57586_ (_06364_, _06363_, _06357_);
  and _57587_ (_06365_, _06364_, _06351_);
  and _57588_ (_06366_, _06358_, _06338_);
  and _57589_ (_06367_, _06366_, _04531_);
  and _57590_ (_06368_, _06339_, _06335_);
  and _57591_ (_06369_, _06368_, _04542_);
  nor _57592_ (_06370_, _06369_, _06367_);
  and _57593_ (_06371_, _06338_, _06327_);
  and _57594_ (_06372_, _06371_, _04536_);
  and _57595_ (_06373_, _06344_, _06354_);
  and _57596_ (_06374_, _06373_, _04561_);
  nor _57597_ (_06375_, _06374_, _06372_);
  and _57598_ (_06376_, _06375_, _06370_);
  and _57599_ (_06377_, _06354_, _06327_);
  and _57600_ (_06378_, _06377_, _04551_);
  and _57601_ (_06379_, _06347_, _06344_);
  and _57602_ (_06380_, _06379_, _04548_);
  nor _57603_ (_06381_, _06380_, _06378_);
  and _57604_ (_06382_, _06347_, _06327_);
  and _57605_ (_06383_, _06382_, _04529_);
  and _57606_ (_06384_, _06358_, _06354_);
  and _57607_ (_06385_, _06384_, _04557_);
  nor _57608_ (_06386_, _06385_, _06383_);
  and _57609_ (_06387_, _06386_, _06381_);
  and _57610_ (_06388_, _06387_, _06376_);
  and _57611_ (_06389_, _06388_, _06365_);
  or _57612_ (_06390_, _06389_, _06114_);
  and _57613_ (_06391_, _06390_, _06210_);
  and _57614_ (_06392_, _06391_, _06271_);
  or _57615_ (_06393_, _06392_, _06211_);
  and _57616_ (_06394_, _05840_, _05786_);
  not _57617_ (_06395_, _06394_);
  and _57618_ (_06396_, _06138_, _05840_);
  nor _57619_ (_06397_, _06396_, _06303_);
  and _57620_ (_06398_, _06397_, _06395_);
  not _57621_ (_06399_, _05833_);
  and _57622_ (_06400_, _06399_, _05786_);
  not _57623_ (_06401_, _06400_);
  and _57624_ (_06402_, _06138_, _06399_);
  nor _57625_ (_06403_, _06402_, _06297_);
  and _57626_ (_06404_, _06403_, _06401_);
  and _57627_ (_06405_, _06404_, _06398_);
  and _57628_ (_06406_, _06300_, _05786_);
  not _57629_ (_06407_, _06406_);
  not _57630_ (_06408_, _05847_);
  and _57631_ (_06409_, _06408_, _05786_);
  not _57632_ (_06410_, _06409_);
  and _57633_ (_06411_, _06138_, _06408_);
  nor _57634_ (_06412_, _06411_, _06306_);
  and _57635_ (_06413_, _06412_, _06410_);
  and _57636_ (_06414_, _06413_, _06407_);
  and _57637_ (_06415_, _06414_, _06405_);
  and _57638_ (_06416_, _06415_, _06393_);
  and _57639_ (_06417_, _06138_, _06300_);
  nor _57640_ (_06418_, _06415_, _06228_);
  or _57641_ (_06419_, _06418_, _06417_);
  or _57642_ (_06420_, _06419_, _06416_);
  not _57643_ (_06421_, _06301_);
  nand _57644_ (_06422_, _06417_, \oc8051_golden_model_1.SP [3]);
  and _57645_ (_06423_, _06422_, _06421_);
  and _57646_ (_06424_, _06423_, _06420_);
  and _57647_ (_06425_, _06301_, _06206_);
  or _57648_ (_06426_, _06425_, _06424_);
  and _57649_ (_06427_, _06426_, _06171_);
  nor _57650_ (_06428_, _06427_, _06170_);
  and _57651_ (_06429_, _06428_, _06168_);
  and _57652_ (_06430_, _06167_, \oc8051_golden_model_1.SP [3]);
  or _57653_ (_06431_, _06430_, _06429_);
  and _57654_ (_06432_, _06431_, _06166_);
  and _57655_ (_06433_, _05786_, _05591_);
  nor _57656_ (_06434_, _06206_, _06166_);
  or _57657_ (_06435_, _06434_, _06433_);
  or _57658_ (_06436_, _06435_, _06432_);
  nand _57659_ (_06437_, _06433_, _06070_);
  and _57660_ (_06438_, _06437_, _06436_);
  nor _57661_ (_06439_, _06438_, _05748_);
  and _57662_ (_06440_, _05820_, _05786_);
  and _57663_ (_06441_, _06206_, _05748_);
  or _57664_ (_06442_, _06441_, _06440_);
  nor _57665_ (_06443_, _06442_, _06439_);
  not _57666_ (_06444_, _06440_);
  nor _57667_ (_06445_, _06444_, _06070_);
  nor _57668_ (_06446_, _06445_, _06443_);
  and _57669_ (_06447_, _06021_, _00607_);
  nor _57670_ (_06448_, _06004_, _44010_);
  nor _57671_ (_06449_, _06448_, _06447_);
  nor _57672_ (_06450_, _06016_, _00383_);
  nor _57673_ (_06451_, _06029_, _43969_);
  nor _57674_ (_06452_, _06451_, _06450_);
  and _57675_ (_06453_, _06452_, _06449_);
  nor _57676_ (_06454_, _06018_, _00301_);
  nor _57677_ (_06455_, _06002_, _00024_);
  nor _57678_ (_06456_, _06455_, _06454_);
  nor _57679_ (_06457_, _05994_, _00260_);
  nor _57680_ (_06458_, _06010_, _00106_);
  nor _57681_ (_06459_, _06458_, _06457_);
  and _57682_ (_06460_, _06459_, _06456_);
  and _57683_ (_06461_, _06460_, _06453_);
  nor _57684_ (_06462_, _06027_, _00167_);
  nor _57685_ (_06463_, _05998_, _00065_);
  nor _57686_ (_06464_, _06463_, _06462_);
  nor _57687_ (_06465_, _05983_, _00550_);
  nor _57688_ (_06466_, _06032_, _00424_);
  nor _57689_ (_06467_, _06466_, _06465_);
  and _57690_ (_06468_, _06467_, _06464_);
  nor _57691_ (_06469_, _06023_, _00465_);
  nor _57692_ (_06470_, _06034_, _00342_);
  nor _57693_ (_06471_, _06470_, _06469_);
  nor _57694_ (_06472_, _05988_, _00506_);
  nor _57695_ (_06473_, _06007_, _00219_);
  nor _57696_ (_06474_, _06473_, _06472_);
  and _57697_ (_06475_, _06474_, _06471_);
  and _57698_ (_06476_, _06475_, _06468_);
  and _57699_ (_06477_, _06476_, _06461_);
  nor _57700_ (_06478_, _06477_, _06039_);
  not _57701_ (_06479_, _06478_);
  nor _57702_ (_06480_, _06165_, _06152_);
  and _57703_ (_06481_, _06480_, _06421_);
  and _57704_ (_06482_, _06256_, _06213_);
  nor _57705_ (_06483_, _06139_, _05748_);
  and _57706_ (_06484_, _06483_, _06210_);
  and _57707_ (_06485_, _06484_, _06482_);
  and _57708_ (_06486_, _06485_, _06481_);
  nor _57709_ (_06487_, _06486_, _06479_);
  not _57710_ (_06488_, _06487_);
  and _57711_ (_06489_, _06478_, _06156_);
  not _57712_ (_06490_, _06489_);
  and _57713_ (_06491_, _06359_, _04505_);
  and _57714_ (_06492_, _06368_, _04497_);
  nor _57715_ (_06493_, _06492_, _06491_);
  and _57716_ (_06494_, _06382_, _04486_);
  and _57717_ (_06495_, _06352_, _04500_);
  nor _57718_ (_06496_, _06495_, _06494_);
  and _57719_ (_06497_, _06496_, _06493_);
  and _57720_ (_06498_, _06384_, _04511_);
  and _57721_ (_06499_, _06361_, _04495_);
  nor _57722_ (_06500_, _06499_, _06498_);
  and _57723_ (_06501_, _06366_, _04491_);
  and _57724_ (_06502_, _06348_, _04507_);
  nor _57725_ (_06503_, _06502_, _06501_);
  and _57726_ (_06504_, _06503_, _06500_);
  and _57727_ (_06505_, _06504_, _06497_);
  and _57728_ (_06506_, _06336_, _00591_);
  and _57729_ (_06507_, _06377_, _04523_);
  nor _57730_ (_06508_, _06507_, _06506_);
  and _57731_ (_06509_, _06371_, _04489_);
  and _57732_ (_06510_, _06345_, _04484_);
  nor _57733_ (_06511_, _06510_, _06509_);
  and _57734_ (_06512_, _06511_, _06508_);
  and _57735_ (_06513_, _06355_, _04513_);
  and _57736_ (_06514_, _06340_, _04517_);
  nor _57737_ (_06515_, _06514_, _06513_);
  and _57738_ (_06516_, _06373_, _04515_);
  and _57739_ (_06517_, _06379_, _04502_);
  nor _57740_ (_06518_, _06517_, _06516_);
  and _57741_ (_06519_, _06518_, _06515_);
  and _57742_ (_06520_, _06519_, _06512_);
  and _57743_ (_06521_, _06520_, _06505_);
  nor _57744_ (_06522_, _06521_, _06114_);
  and _57745_ (_06523_, _06124_, _06300_);
  and _57746_ (_06524_, _06124_, _05840_);
  nor _57747_ (_06525_, _06524_, _06523_);
  and _57748_ (_06526_, _06124_, _05781_);
  not _57749_ (_06527_, _06526_);
  and _57750_ (_06528_, _06527_, _06525_);
  and _57751_ (_06529_, _06124_, _06150_);
  and _57752_ (_06530_, _06124_, _05591_);
  nor _57753_ (_06531_, _06530_, _06529_);
  and _57754_ (_06532_, _06167_, \oc8051_golden_model_1.SP [2]);
  and _57755_ (_06533_, _06122_, _05744_);
  and _57756_ (_06534_, _06533_, _05825_);
  nor _57757_ (_06535_, _06534_, _06532_);
  and _57758_ (_06536_, _06127_, _05790_);
  not _57759_ (_06537_, _06536_);
  and _57760_ (_06538_, _06533_, _06150_);
  and _57761_ (_06539_, _06122_, _05820_);
  nor _57762_ (_06540_, _06539_, _06538_);
  and _57763_ (_06541_, _06540_, _06537_);
  and _57764_ (_06542_, _06541_, _06535_);
  and _57765_ (_06543_, _06542_, _06531_);
  and _57766_ (_06544_, _06543_, _06528_);
  and _57767_ (_06545_, _06124_, _06222_);
  and _57768_ (_06546_, _06124_, _06155_);
  nor _57769_ (_06547_, _06546_, _06545_);
  and _57770_ (_06548_, _06124_, _05790_);
  and _57771_ (_06549_, _06124_, _06144_);
  nor _57772_ (_06550_, _06549_, _06548_);
  and _57773_ (_06551_, _06550_, _06547_);
  and _57774_ (_06552_, _06124_, _05825_);
  not _57775_ (_06553_, _06552_);
  and _57776_ (_06554_, _06533_, _06408_);
  and _57777_ (_06555_, _06533_, _05840_);
  nor _57778_ (_06556_, _06555_, _06554_);
  and _57779_ (_06557_, _06124_, _06408_);
  and _57780_ (_06558_, _06125_, _06399_);
  nor _57781_ (_06559_, _06558_, _06557_);
  and _57782_ (_06560_, _06559_, _06556_);
  and _57783_ (_06561_, _06560_, _06553_);
  and _57784_ (_06562_, _06127_, _05591_);
  and _57785_ (_06563_, _06123_, _05591_);
  nor _57786_ (_06564_, _06563_, _06562_);
  not _57787_ (_06565_, _06564_);
  not _57788_ (_06566_, \oc8051_golden_model_1.SP [2]);
  nor _57789_ (_06567_, _06217_, _06417_);
  nor _57790_ (_06568_, _06567_, _06566_);
  nor _57791_ (_06569_, _06568_, _06565_);
  and _57792_ (_06570_, _06569_, _06561_);
  and _57793_ (_06571_, _06127_, _05781_);
  and _57794_ (_06572_, _06127_, _06222_);
  nor _57795_ (_06573_, _06572_, _06571_);
  and _57796_ (_06574_, _06127_, _06399_);
  or _57797_ (_06575_, _05790_, _05781_);
  and _57798_ (_06576_, _06575_, _06123_);
  nor _57799_ (_06577_, _06576_, _06574_);
  and _57800_ (_06578_, _06577_, _06573_);
  and _57801_ (_06579_, _06127_, _06144_);
  nor _57802_ (_06580_, _06272_, _06579_);
  and _57803_ (_06581_, _06123_, _06222_);
  not _57804_ (_06582_, _06581_);
  and _57805_ (_06583_, _06533_, _06300_);
  and _57806_ (_06584_, _06533_, _06155_);
  nor _57807_ (_06585_, _06584_, _06583_);
  and _57808_ (_06586_, _06585_, _06582_);
  and _57809_ (_06587_, _06586_, _06580_);
  and _57810_ (_06588_, _06587_, _06578_);
  and _57811_ (_06589_, _06588_, _06570_);
  and _57812_ (_06590_, _06589_, _06551_);
  and _57813_ (_06591_, _06590_, _06544_);
  not _57814_ (_06592_, _06591_);
  nor _57815_ (_06593_, _06592_, _06522_);
  not _57816_ (_06594_, _06593_);
  nor _57817_ (_06595_, _06023_, _00450_);
  nor _57818_ (_06596_, _05994_, _00245_);
  nor _57819_ (_06597_, _06596_, _06595_);
  nor _57820_ (_06598_, _06007_, _00204_);
  nor _57821_ (_06599_, _06029_, _43954_);
  nor _57822_ (_06600_, _06599_, _06598_);
  and _57823_ (_06601_, _06600_, _06597_);
  nor _57824_ (_06602_, _06032_, _00409_);
  nor _57825_ (_06603_, _05998_, _00050_);
  nor _57826_ (_06604_, _06603_, _06602_);
  nor _57827_ (_06605_, _06016_, _00368_);
  nor _57828_ (_06606_, _06018_, _00286_);
  nor _57829_ (_06607_, _06606_, _06605_);
  and _57830_ (_06608_, _06607_, _06604_);
  and _57831_ (_06609_, _06608_, _06601_);
  nor _57832_ (_06610_, _06027_, _00134_);
  nor _57833_ (_06611_, _06010_, _00091_);
  nor _57834_ (_06612_, _06611_, _06610_);
  and _57835_ (_06613_, _06021_, _00591_);
  nor _57836_ (_06614_, _06004_, _43995_);
  nor _57837_ (_06615_, _06614_, _06613_);
  and _57838_ (_06616_, _06615_, _06612_);
  nor _57839_ (_06617_, _05983_, _00532_);
  nor _57840_ (_06618_, _06002_, _00009_);
  nor _57841_ (_06619_, _06618_, _06617_);
  nor _57842_ (_06620_, _05988_, _00491_);
  nor _57843_ (_06621_, _06034_, _00327_);
  nor _57844_ (_06622_, _06621_, _06620_);
  and _57845_ (_06623_, _06622_, _06619_);
  and _57846_ (_06624_, _06623_, _06616_);
  and _57847_ (_06625_, _06624_, _06609_);
  not _57848_ (_06626_, _06625_);
  nand _57849_ (_06627_, _06265_, _06237_);
  nor _57850_ (_06628_, _06627_, _06230_);
  nand _57851_ (_06629_, _06628_, _06251_);
  nor _57852_ (_06630_, _06440_, _06433_);
  and _57853_ (_06631_, _06630_, _06171_);
  nand _57854_ (_06632_, _06631_, _06415_);
  or _57855_ (_06633_, _06632_, _06629_);
  and _57856_ (_06634_, _06633_, _06626_);
  nor _57857_ (_06635_, _06634_, _06594_);
  and _57858_ (_06636_, _06635_, _06490_);
  and _57859_ (_06637_, _06636_, _06488_);
  not _57860_ (_06638_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor _57861_ (_06639_, _06444_, _06107_);
  not _57862_ (_06640_, _06639_);
  nor _57863_ (_06641_, _06265_, _06107_);
  nor _57864_ (_06642_, _06256_, _06071_);
  not _57865_ (_06643_, _06236_);
  nor _57866_ (_06644_, _06643_, _06107_);
  or _57867_ (_06645_, _06229_, _06107_);
  nor _57868_ (_06646_, _06224_, _06107_);
  and _57869_ (_06647_, _06281_, _06155_);
  nand _57870_ (_06648_, _05707_, _05666_);
  nor _57871_ (_06649_, _06648_, _05762_);
  nor _57872_ (_06650_, _06649_, _06647_);
  not _57873_ (_06651_, _05776_);
  and _57874_ (_06652_, _06281_, _06651_);
  and _57875_ (_06653_, _06313_, _06222_);
  nor _57876_ (_06654_, _06653_, _06652_);
  nor _57877_ (_06655_, _06572_, _06160_);
  and _57878_ (_06656_, _06655_, _06654_);
  nor _57879_ (_06657_, _06281_, _05786_);
  or _57880_ (_06658_, _06657_, _05771_);
  nand _57881_ (_06659_, _06118_, _05707_);
  nor _57882_ (_06660_, _06659_, _05771_);
  not _57883_ (_06661_, _06660_);
  and _57884_ (_06662_, _06661_, _06658_);
  and _57885_ (_06663_, _06662_, _06656_);
  and _57886_ (_06665_, _06663_, _06650_);
  or _57887_ (_06666_, _06665_, _06646_);
  nand _57888_ (_06667_, _06666_, _06157_);
  nand _57889_ (_06668_, _06158_, _06667_);
  and _57890_ (_06669_, _06217_, _06142_);
  nor _57891_ (_06670_, _06669_, _06220_);
  not _57892_ (_06671_, _06670_);
  and _57893_ (_06672_, _06122_, _05707_);
  not _57894_ (_06673_, _06672_);
  not _57895_ (_06674_, _06281_);
  and _57896_ (_06675_, _06659_, _06674_);
  and _57897_ (_06676_, _06675_, _06673_);
  nor _57898_ (_06677_, _06676_, _05768_);
  nor _57899_ (_06678_, _06677_, _06671_);
  nand _57900_ (_06679_, _06678_, _06668_);
  nand _57901_ (_06680_, _06679_, _06645_);
  and _57902_ (_06681_, _06680_, _06153_);
  or _57903_ (_06682_, _06154_, _06681_);
  and _57904_ (_06683_, _06151_, _06107_);
  and _57905_ (_06684_, _06118_, _06137_);
  and _57906_ (_06685_, _06684_, _06144_);
  nor _57907_ (_06686_, _06274_, _06685_);
  and _57908_ (_06687_, _06115_, _06144_);
  and _57909_ (_06688_, _06687_, _05707_);
  nor _57910_ (_06689_, _06688_, _06579_);
  and _57911_ (_06690_, _06689_, _06686_);
  and _57912_ (_06691_, _06690_, _06315_);
  not _57913_ (_06692_, _06691_);
  nor _57914_ (_06693_, _06692_, _06683_);
  and _57915_ (_06694_, _06693_, _06682_);
  or _57916_ (_06695_, _06694_, _06644_);
  nand _57917_ (_06696_, _06695_, _06213_);
  nor _57918_ (_06697_, _06213_, _06071_);
  nor _57919_ (_06698_, _06697_, _06252_);
  nand _57920_ (_06699_, _06698_, _06696_);
  and _57921_ (_06700_, _06252_, _06107_);
  and _57922_ (_06701_, _06115_, _06245_);
  and _57923_ (_06702_, _06701_, _05707_);
  nor _57924_ (_06703_, _06702_, _06261_);
  not _57925_ (_06704_, _06703_);
  nor _57926_ (_06705_, _06704_, _06700_);
  and _57927_ (_06706_, _06705_, _06699_);
  or _57928_ (_06707_, _06706_, _06642_);
  nor _57929_ (_06708_, _06536_, _06260_);
  and _57930_ (_06709_, _06281_, _05790_);
  not _57931_ (_06710_, _06709_);
  and _57932_ (_06711_, _06137_, _05666_);
  nor _57933_ (_06712_, _06273_, _06711_);
  or _57934_ (_06713_, _06712_, _05803_);
  and _57935_ (_06714_, _06713_, _06710_);
  and _57936_ (_06715_, _06714_, _06708_);
  and _57937_ (_06716_, _06715_, _06707_);
  or _57938_ (_06717_, _06716_, _06641_);
  and _57939_ (_06718_, _06717_, _06140_);
  or _57940_ (_06719_, _06718_, _06141_);
  nor _57941_ (_06720_, _06684_, _06127_);
  or _57942_ (_06721_, _06720_, _05797_);
  not _57943_ (_06722_, _06313_);
  nor _57944_ (_06723_, _06281_, _06273_);
  and _57945_ (_06724_, _06723_, _06722_);
  or _57946_ (_06725_, _06724_, _05797_);
  and _57947_ (_06726_, _06725_, _06721_);
  and _57948_ (_06727_, _06726_, _06719_);
  and _57949_ (_06728_, _06336_, _00575_);
  and _57950_ (_06729_, _06345_, _04393_);
  nor _57951_ (_06730_, _06729_, _06728_);
  and _57952_ (_06731_, _06384_, _04420_);
  and _57953_ (_06732_, _06348_, _04416_);
  nor _57954_ (_06733_, _06732_, _06731_);
  and _57955_ (_06734_, _06733_, _06730_);
  and _57956_ (_06735_, _06373_, _04424_);
  and _57957_ (_06736_, _06352_, _04409_);
  nor _57958_ (_06737_, _06736_, _06735_);
  and _57959_ (_06738_, _06371_, _04398_);
  and _57960_ (_06739_, _06382_, _04395_);
  nor _57961_ (_06740_, _06739_, _06738_);
  and _57962_ (_06741_, _06740_, _06737_);
  and _57963_ (_06742_, _06741_, _06734_);
  and _57964_ (_06743_, _06361_, _04404_);
  and _57965_ (_06744_, _06368_, _04406_);
  nor _57966_ (_06745_, _06744_, _06743_);
  and _57967_ (_06746_, _06359_, _04414_);
  and _57968_ (_06747_, _06366_, _04400_);
  nor _57969_ (_06748_, _06747_, _06746_);
  and _57970_ (_06749_, _06748_, _06745_);
  and _57971_ (_06750_, _06355_, _04422_);
  and _57972_ (_06751_, _06340_, _04426_);
  nor _57973_ (_06752_, _06751_, _06750_);
  and _57974_ (_06753_, _06377_, _04432_);
  and _57975_ (_06754_, _06379_, _04411_);
  nor _57976_ (_06755_, _06754_, _06753_);
  and _57977_ (_06756_, _06755_, _06752_);
  and _57978_ (_06757_, _06756_, _06749_);
  and _57979_ (_06758_, _06757_, _06742_);
  and _57980_ (_06759_, _06758_, _05787_);
  nor _57981_ (_06760_, _06759_, _06209_);
  and _57982_ (_06761_, _06760_, _06727_);
  not _57983_ (_06762_, _06209_);
  nor _57984_ (_06763_, _06762_, _06071_);
  or _57985_ (_06764_, _06763_, _06761_);
  and _57986_ (_06765_, _06281_, _06109_);
  nor _57987_ (_06766_, _06765_, _06208_);
  and _57988_ (_06767_, _06766_, _06764_);
  not _57989_ (_06768_, _06208_);
  nor _57990_ (_06769_, _06768_, _06071_);
  or _57991_ (_06770_, _06769_, _06767_);
  and _57992_ (_06771_, _06273_, _06399_);
  nor _57993_ (_06772_, _06771_, _06574_);
  and _57994_ (_06773_, _06281_, _06399_);
  and _57995_ (_06774_, _06711_, _06399_);
  nor _57996_ (_06775_, _06774_, _06773_);
  and _57997_ (_06776_, _06775_, _06772_);
  and _57998_ (_06777_, _06776_, _06770_);
  nor _57999_ (_06778_, _06404_, _06108_);
  nor _58000_ (_06779_, _06676_, _05847_);
  nor _58001_ (_06780_, _06779_, _06778_);
  and _58002_ (_06781_, _06780_, _06777_);
  nor _58003_ (_06782_, _06413_, _06108_);
  not _58004_ (_06783_, _05840_);
  nor _58005_ (_06784_, _06676_, _06783_);
  nor _58006_ (_06785_, _06784_, _06782_);
  and _58007_ (_06786_, _06785_, _06781_);
  nor _58008_ (_06787_, _06398_, _06108_);
  nor _58009_ (_06788_, _06722_, _05844_);
  nor _58010_ (_06789_, _06788_, _06406_);
  and _58011_ (_06790_, _06273_, _06300_);
  not _58012_ (_06791_, _06790_);
  and _58013_ (_06792_, _06281_, _06300_);
  not _58014_ (_06793_, _06792_);
  and _58015_ (_06794_, _06127_, _06300_);
  and _58016_ (_06795_, _06684_, _06300_);
  nor _58017_ (_06796_, _06795_, _06794_);
  and _58018_ (_06797_, _06796_, _06793_);
  and _58019_ (_06798_, _06797_, _06791_);
  and _58020_ (_06799_, _06798_, _06789_);
  not _58021_ (_06800_, _06799_);
  nor _58022_ (_06801_, _06800_, _06787_);
  and _58023_ (_06802_, _06801_, _06786_);
  nor _58024_ (_06803_, _06407_, _06107_);
  or _58025_ (_06804_, _06803_, _06802_);
  and _58026_ (_06805_, _06417_, _06142_);
  nor _58027_ (_06806_, _06805_, _06301_);
  and _58028_ (_06807_, _06806_, _06804_);
  nor _58029_ (_06808_, _06421_, _06071_);
  or _58030_ (_06809_, _06808_, _06807_);
  and _58031_ (_06810_, _06127_, _05825_);
  not _58032_ (_06811_, _05825_);
  and _58033_ (_06812_, _06712_, _06657_);
  nor _58034_ (_06813_, _06812_, _06811_);
  nor _58035_ (_06814_, _06813_, _06810_);
  and _58036_ (_06815_, _06814_, _06809_);
  nor _58037_ (_06816_, _06171_, _06107_);
  or _58038_ (_06817_, _06816_, _06815_);
  and _58039_ (_06818_, _06167_, _06142_);
  nor _58040_ (_06819_, _06818_, _06165_);
  and _58041_ (_06820_, _06819_, _06817_);
  nor _58042_ (_06821_, _06166_, _06071_);
  nor _58043_ (_06822_, _06821_, _06820_);
  not _58044_ (_06823_, _05591_);
  nor _58045_ (_06824_, _06127_, _05786_);
  and _58046_ (_06825_, _06824_, _06722_);
  and _58047_ (_06826_, _06825_, _06675_);
  nor _58048_ (_06827_, _06826_, _06823_);
  nor _58049_ (_06828_, _06827_, _06822_);
  not _58050_ (_06829_, _06433_);
  nor _58051_ (_06830_, _06829_, _06107_);
  or _58052_ (_06831_, _06830_, _06828_);
  and _58053_ (_06832_, _06831_, _05749_);
  or _58054_ (_06833_, _06832_, _06072_);
  and _58055_ (_06834_, _06281_, _05820_);
  not _58056_ (_06835_, _06834_);
  and _58057_ (_06836_, _06273_, _05820_);
  nor _58058_ (_06837_, _06836_, _06440_);
  and _58059_ (_06838_, _06837_, _06835_);
  and _58060_ (_06839_, _06684_, _05820_);
  and _58061_ (_06840_, _06672_, _05820_);
  nor _58062_ (_06841_, _06840_, _06839_);
  and _58063_ (_06842_, _06841_, _06838_);
  nand _58064_ (_06843_, _06842_, _06833_);
  nand _58065_ (_06844_, _06843_, _06640_);
  or _58066_ (_06845_, _06844_, _06638_);
  nor _58067_ (_06846_, _06004_, _44005_);
  nor _58068_ (_06847_, _06002_, _00019_);
  nor _58069_ (_06848_, _06847_, _06846_);
  nor _58070_ (_06849_, _05983_, _00542_);
  nor _58071_ (_06850_, _06007_, _00214_);
  nor _58072_ (_06851_, _06850_, _06849_);
  and _58073_ (_06852_, _06851_, _06848_);
  nor _58074_ (_06853_, _05998_, _00060_);
  nor _58075_ (_06854_, _06010_, _00101_);
  nor _58076_ (_06855_, _06854_, _06853_);
  nor _58077_ (_06856_, _06032_, _00419_);
  nor _58078_ (_06857_, _06018_, _00296_);
  nor _58079_ (_06858_, _06857_, _06856_);
  and _58080_ (_06859_, _06858_, _06855_);
  and _58081_ (_06860_, _06859_, _06852_);
  nor _58082_ (_06861_, _06023_, _00460_);
  nor _58083_ (_06862_, _06034_, _00337_);
  nor _58084_ (_06863_, _06862_, _06861_);
  and _58085_ (_06864_, _06021_, _00602_);
  nor _58086_ (_06865_, _05988_, _00501_);
  nor _58087_ (_06866_, _06865_, _06864_);
  and _58088_ (_06867_, _06866_, _06863_);
  nor _58089_ (_06868_, _06016_, _00378_);
  nor _58090_ (_06869_, _06029_, _43964_);
  nor _58091_ (_06870_, _06869_, _06868_);
  nor _58092_ (_06871_, _05994_, _00255_);
  nor _58093_ (_06872_, _06027_, _00156_);
  nor _58094_ (_06873_, _06872_, _06871_);
  and _58095_ (_06874_, _06873_, _06870_);
  and _58096_ (_06875_, _06874_, _06867_);
  and _58097_ (_06876_, _06875_, _06860_);
  nor _58098_ (_06877_, _06876_, _06039_);
  and _58099_ (_06878_, _06486_, _06157_);
  not _58100_ (_06879_, _06878_);
  and _58101_ (_06880_, _06879_, _06877_);
  not _58102_ (_06881_, _06880_);
  and _58103_ (_06882_, _06021_, _00583_);
  nor _58104_ (_06883_, _05998_, _00045_);
  nor _58105_ (_06884_, _06883_, _06882_);
  nor _58106_ (_06885_, _05983_, _00527_);
  nor _58107_ (_06886_, _06034_, _00322_);
  nor _58108_ (_06887_, _06886_, _06885_);
  and _58109_ (_06888_, _06887_, _06884_);
  nor _58110_ (_06889_, _06027_, _00127_);
  nor _58111_ (_06890_, _06007_, _00199_);
  nor _58112_ (_06891_, _06890_, _06889_);
  nor _58113_ (_06892_, _06032_, _00404_);
  nor _58114_ (_06893_, _05994_, _00240_);
  nor _58115_ (_06894_, _06893_, _06892_);
  and _58116_ (_06895_, _06894_, _06891_);
  and _58117_ (_06896_, _06895_, _06888_);
  nor _58118_ (_06897_, _05988_, _00486_);
  nor _58119_ (_06898_, _06023_, _00445_);
  nor _58120_ (_06899_, _06898_, _06897_);
  nor _58121_ (_06900_, _06018_, _00281_);
  nor _58122_ (_06901_, _06002_, _00004_);
  nor _58123_ (_06902_, _06901_, _06900_);
  and _58124_ (_06903_, _06902_, _06899_);
  nor _58125_ (_06904_, _06016_, _00363_);
  nor _58126_ (_06905_, _06010_, _00086_);
  nor _58127_ (_06906_, _06905_, _06904_);
  nor _58128_ (_06907_, _06029_, _43949_);
  nor _58129_ (_06908_, _06004_, _43990_);
  nor _58130_ (_06909_, _06908_, _06907_);
  and _58131_ (_06910_, _06909_, _06906_);
  and _58132_ (_06911_, _06910_, _06903_);
  and _58133_ (_06912_, _06911_, _06896_);
  not _58134_ (_06913_, _06912_);
  and _58135_ (_06914_, _06913_, _06633_);
  and _58136_ (_06915_, _06359_, _04460_);
  and _58137_ (_06916_, _06368_, _04452_);
  nor _58138_ (_06917_, _06916_, _06915_);
  and _58139_ (_06918_, _06373_, _04470_);
  and _58140_ (_06919_, _06379_, _04457_);
  nor _58141_ (_06920_, _06919_, _06918_);
  and _58142_ (_06921_, _06920_, _06917_);
  and _58143_ (_06922_, _06384_, _04466_);
  and _58144_ (_06923_, _06366_, _04445_);
  nor _58145_ (_06924_, _06923_, _06922_);
  and _58146_ (_06925_, _06355_, _04468_);
  and _58147_ (_06926_, _06340_, _04472_);
  nor _58148_ (_06927_, _06926_, _06925_);
  and _58149_ (_06928_, _06927_, _06924_);
  and _58150_ (_06929_, _06928_, _06921_);
  and _58151_ (_06930_, _06382_, _04440_);
  and _58152_ (_06931_, _06345_, _04438_);
  nor _58153_ (_06932_, _06931_, _06930_);
  and _58154_ (_06933_, _06377_, _04478_);
  and _58155_ (_06934_, _06352_, _04455_);
  nor _58156_ (_06935_, _06934_, _06933_);
  and _58157_ (_06936_, _06935_, _06932_);
  and _58158_ (_06937_, _06361_, _04450_);
  and _58159_ (_06938_, _06348_, _04462_);
  nor _58160_ (_06939_, _06938_, _06937_);
  and _58161_ (_06940_, _06336_, _00583_);
  and _58162_ (_06941_, _06371_, _04443_);
  nor _58163_ (_06942_, _06941_, _06940_);
  and _58164_ (_06943_, _06942_, _06939_);
  and _58165_ (_06944_, _06943_, _06936_);
  and _58166_ (_06945_, _06944_, _06929_);
  nor _58167_ (_06946_, _06945_, _06114_);
  and _58168_ (_06947_, _06217_, \oc8051_golden_model_1.SP [1]);
  not _58169_ (_06948_, _06128_);
  nor _58170_ (_06949_, _05820_, _06150_);
  nor _58171_ (_06950_, _06949_, _06948_);
  nor _58172_ (_06951_, _06950_, _06947_);
  and _58173_ (_06952_, _06684_, _05825_);
  and _58174_ (_06953_, _06539_, _05742_);
  nor _58175_ (_06954_, _06953_, _06952_);
  and _58176_ (_06955_, _06954_, _06951_);
  and _58177_ (_06956_, _06124_, _06399_);
  and _58178_ (_06957_, _06118_, _06283_);
  and _58179_ (_06958_, _06957_, _05825_);
  or _58180_ (_06959_, _06958_, _06557_);
  nor _58181_ (_06960_, _06959_, _06956_);
  and _58182_ (_06961_, _06960_, _06553_);
  and _58183_ (_06962_, _06961_, _06955_);
  and _58184_ (_06963_, _06531_, _06528_);
  and _58185_ (_06964_, _06963_, _06962_);
  and _58186_ (_06965_, _06128_, _06408_);
  and _58187_ (_06966_, _05771_, _05758_);
  and _58188_ (_06967_, _05833_, _05797_);
  and _58189_ (_06968_, _06967_, _06966_);
  nor _58190_ (_06969_, _06968_, _06948_);
  nor _58191_ (_06970_, _06969_, _06965_);
  and _58192_ (_06971_, _06128_, _05790_);
  and _58193_ (_06972_, _06128_, _05591_);
  nor _58194_ (_06973_, _06972_, _06971_);
  and _58195_ (_06974_, _06973_, _06970_);
  and _58196_ (_06975_, _06128_, _05840_);
  and _58197_ (_06976_, _06128_, _06300_);
  nor _58198_ (_06977_, _06976_, _06975_);
  and _58199_ (_06978_, _06128_, _06155_);
  not _58200_ (_06979_, \oc8051_golden_model_1.SP [1]);
  nor _58201_ (_06980_, _06417_, _06167_);
  nor _58202_ (_06981_, _06980_, _06979_);
  nor _58203_ (_06982_, _06981_, _06978_);
  and _58204_ (_06983_, _06982_, _06977_);
  and _58205_ (_06984_, _06983_, _06974_);
  and _58206_ (_06985_, _06984_, _06551_);
  and _58207_ (_06986_, _06985_, _06964_);
  not _58208_ (_06987_, _06986_);
  nor _58209_ (_06988_, _06987_, _06946_);
  not _58210_ (_06989_, _06988_);
  nor _58211_ (_06990_, _06989_, _06914_);
  and _58212_ (_06991_, _06990_, _06881_);
  not _58213_ (_06992_, \oc8051_golden_model_1.IRAM[1] [0]);
  and _58214_ (_06993_, _06843_, _06640_);
  or _58215_ (_06994_, _06993_, _06992_);
  and _58216_ (_06995_, _06994_, _06991_);
  nand _58217_ (_06996_, _06995_, _06845_);
  not _58218_ (_06997_, \oc8051_golden_model_1.IRAM[3] [0]);
  or _58219_ (_06998_, _06993_, _06997_);
  not _58220_ (_06999_, _06991_);
  not _58221_ (_07000_, \oc8051_golden_model_1.IRAM[2] [0]);
  or _58222_ (_07001_, _06844_, _07000_);
  and _58223_ (_07002_, _07001_, _06999_);
  nand _58224_ (_07003_, _07002_, _06998_);
  nand _58225_ (_07004_, _07003_, _06996_);
  nand _58226_ (_07005_, _07004_, _06637_);
  not _58227_ (_07006_, _06637_);
  not _58228_ (_07007_, \oc8051_golden_model_1.IRAM[7] [0]);
  or _58229_ (_07008_, _06993_, _07007_);
  not _58230_ (_07009_, \oc8051_golden_model_1.IRAM[6] [0]);
  or _58231_ (_07010_, _06844_, _07009_);
  and _58232_ (_07011_, _07010_, _06999_);
  nand _58233_ (_07012_, _07011_, _07008_);
  not _58234_ (_07013_, \oc8051_golden_model_1.IRAM[4] [0]);
  or _58235_ (_07014_, _06844_, _07013_);
  not _58236_ (_07015_, \oc8051_golden_model_1.IRAM[5] [0]);
  or _58237_ (_07016_, _06993_, _07015_);
  and _58238_ (_07017_, _07016_, _06991_);
  nand _58239_ (_07018_, _07017_, _07014_);
  nand _58240_ (_07019_, _07018_, _07012_);
  nand _58241_ (_07020_, _07019_, _07006_);
  nand _58242_ (_07021_, _07020_, _07005_);
  nand _58243_ (_07022_, _07021_, _06446_);
  not _58244_ (_07023_, _06446_);
  nand _58245_ (_07024_, _06844_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _58246_ (_07025_, _06993_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _58247_ (_07026_, _07025_, _06999_);
  nand _58248_ (_07027_, _07026_, _07024_);
  nand _58249_ (_07028_, _06993_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand _58250_ (_07029_, _06844_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _58251_ (_07030_, _07029_, _06991_);
  nand _58252_ (_07031_, _07030_, _07028_);
  nand _58253_ (_07032_, _07031_, _07027_);
  nand _58254_ (_07033_, _07032_, _06637_);
  not _58255_ (_07034_, \oc8051_golden_model_1.IRAM[15] [0]);
  or _58256_ (_07035_, _06993_, _07034_);
  nand _58257_ (_07036_, _06993_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _58258_ (_07037_, _07036_, _06999_);
  nand _58259_ (_07038_, _07037_, _07035_);
  not _58260_ (_07039_, \oc8051_golden_model_1.IRAM[12] [0]);
  or _58261_ (_07040_, _06844_, _07039_);
  not _58262_ (_07041_, \oc8051_golden_model_1.IRAM[13] [0]);
  or _58263_ (_07042_, _06993_, _07041_);
  and _58264_ (_07043_, _07042_, _06991_);
  nand _58265_ (_07044_, _07043_, _07040_);
  nand _58266_ (_07045_, _07044_, _07038_);
  nand _58267_ (_07046_, _07045_, _07006_);
  nand _58268_ (_07047_, _07046_, _07033_);
  nand _58269_ (_07048_, _07047_, _07023_);
  and _58270_ (_07049_, _07048_, _07022_);
  and _58271_ (_07050_, _07049_, _06164_);
  nor _58272_ (_07051_, _06294_, _05789_);
  and _58273_ (_07052_, _07051_, _06723_);
  nor _58274_ (_07053_, _07052_, _05776_);
  not _58275_ (_07054_, _07053_);
  nor _58276_ (_07055_, _07054_, _07050_);
  and _58277_ (_07056_, _06277_, _06222_);
  not _58278_ (_07057_, _07056_);
  nor _58279_ (_07058_, _07057_, _06039_);
  and _58280_ (_07059_, _07058_, _06107_);
  nor _58281_ (_07060_, _07059_, _07055_);
  and _58282_ (_07061_, _06581_, \oc8051_golden_model_1.SP [0]);
  nor _58283_ (_07062_, _07061_, _06649_);
  and _58284_ (_07063_, _07062_, _07060_);
  and _58285_ (_07064_, _06115_, _06155_);
  not _58286_ (_07065_, _07064_);
  nor _58287_ (_07066_, _07065_, _07049_);
  nor _58288_ (_07067_, _07066_, _06162_);
  and _58289_ (_07068_, _07067_, _07063_);
  nor _58290_ (_07069_, _07068_, _06163_);
  nor _58291_ (_07070_, _07069_, _06159_);
  not _58292_ (_07071_, _07070_);
  and _58293_ (_07072_, _07071_, _06158_);
  nor _58294_ (_07073_, _05764_, _06142_);
  nor _58295_ (_07074_, _07073_, _07072_);
  not _58296_ (_07075_, _06217_);
  nor _58297_ (_07076_, _07075_, _06039_);
  and _58298_ (_07077_, _07076_, _06107_);
  nor _58299_ (_07078_, _06648_, _05768_);
  nor _58300_ (_07079_, _07078_, _07077_);
  and _58301_ (_07080_, _07079_, _07074_);
  and _58302_ (_07081_, _06115_, _06150_);
  not _58303_ (_07082_, _07081_);
  nor _58304_ (_07083_, _07082_, _07049_);
  not _58305_ (_07084_, _07083_);
  and _58306_ (_07085_, _07084_, _07080_);
  nor _58307_ (_07086_, _06153_, _06039_);
  nor _58308_ (_07087_, _06229_, _06039_);
  and _58309_ (_07088_, _07087_, _06107_);
  nor _58310_ (_07089_, _07088_, _07086_);
  and _58311_ (_07090_, _07089_, _07085_);
  nor _58312_ (_07091_, _07090_, _06154_);
  or _58313_ (_07092_, _07091_, _06151_);
  nand _58314_ (_07093_, _06151_, _06142_);
  nand _58315_ (_07094_, _07093_, _07092_);
  and _58316_ (_07095_, _07094_, _06149_);
  nor _58317_ (_07096_, _07095_, _06147_);
  and _58318_ (_07097_, _06313_, _06245_);
  or _58319_ (_07098_, _06248_, _07097_);
  nor _58320_ (_07099_, _06659_, _05774_);
  or _58321_ (_07100_, _07099_, _07098_);
  or _58322_ (_07101_, _07100_, _07096_);
  nor _58323_ (_07102_, _07101_, _06143_);
  nor _58324_ (_07103_, _06140_, _06039_);
  not _58325_ (_07104_, _06701_);
  nor _58326_ (_07105_, _07049_, _07104_);
  nor _58327_ (_07106_, _07105_, _07103_);
  and _58328_ (_07107_, _07106_, _07102_);
  nor _58329_ (_07108_, _07107_, _06141_);
  nor _58330_ (_07109_, _07108_, _05791_);
  and _58331_ (_07110_, _05791_, _06142_);
  nor _58332_ (_07111_, _07110_, _07109_);
  nor _58333_ (_07112_, _06648_, _05835_);
  or _58334_ (_07113_, _07112_, _07111_);
  nor _58335_ (_07114_, _07113_, _06136_);
  and _58336_ (_07115_, _06115_, _06109_);
  not _58337_ (_07116_, _07115_);
  nor _58338_ (_07117_, _07116_, _07049_);
  nor _58339_ (_07118_, _07117_, _06112_);
  and _58340_ (_07119_, _07118_, _07114_);
  nor _58341_ (_07120_, _07119_, _06113_);
  nor _58342_ (_07121_, _07120_, _06076_);
  nor _58343_ (_07122_, _05836_, \oc8051_golden_model_1.SP [0]);
  nor _58344_ (_07123_, _07122_, _07121_);
  not _58345_ (_07124_, _05848_);
  not _58346_ (_07125_, _06402_);
  nor _58347_ (_07126_, _07125_, _06039_);
  not _58348_ (_07127_, _06297_);
  nor _58349_ (_07128_, _07127_, _06039_);
  nor _58350_ (_07129_, _07128_, _07126_);
  not _58351_ (_07130_, _06411_);
  nor _58352_ (_07131_, _07130_, _06039_);
  not _58353_ (_07132_, _06306_);
  nor _58354_ (_07133_, _07132_, _06039_);
  nor _58355_ (_07134_, _07133_, _07131_);
  and _58356_ (_07135_, _07134_, _07129_);
  nor _58357_ (_07136_, _07135_, _06108_);
  nor _58358_ (_07137_, _07136_, _07124_);
  not _58359_ (_07138_, _07137_);
  nor _58360_ (_07139_, _07138_, _07123_);
  nor _58361_ (_07140_, _05848_, \oc8051_golden_model_1.SP [0]);
  nor _58362_ (_07141_, _07140_, _07139_);
  not _58363_ (_07142_, _05846_);
  nor _58364_ (_07143_, _06397_, _06039_);
  and _58365_ (_07144_, _07143_, _06107_);
  nor _58366_ (_07145_, _07144_, _07142_);
  not _58367_ (_07146_, _07145_);
  nor _58368_ (_07147_, _07146_, _07141_);
  nor _58369_ (_07148_, _07147_, _06075_);
  not _58370_ (_07149_, _06648_);
  and _58371_ (_07150_, _07149_, _05591_);
  nor _58372_ (_07151_, _07150_, _07148_);
  nor _58373_ (_07152_, _06829_, _06039_);
  and _58374_ (_07153_, _06115_, _05591_);
  not _58375_ (_07154_, _07153_);
  nor _58376_ (_07155_, _07154_, _07049_);
  nor _58377_ (_07156_, _07155_, _07152_);
  and _58378_ (_07157_, _07156_, _07151_);
  and _58379_ (_07158_, _07152_, _06108_);
  nor _58380_ (_07159_, _07158_, _07157_);
  nor _58381_ (_07160_, _06310_, _05823_);
  nor _58382_ (_07161_, _07160_, _06142_);
  nor _58383_ (_07162_, _07161_, _07159_);
  and _58384_ (_07163_, _07162_, _06074_);
  nor _58385_ (_07164_, _07163_, _06072_);
  and _58386_ (_07165_, _07149_, _05820_);
  nor _58387_ (_07166_, _07165_, _07164_);
  nor _58388_ (_07167_, _06444_, _06039_);
  and _58389_ (_07168_, _06115_, _05820_);
  not _58390_ (_07169_, _07168_);
  nor _58391_ (_07170_, _07169_, _07049_);
  nor _58392_ (_07171_, _07170_, _07167_);
  and _58393_ (_07172_, _07171_, _07166_);
  and _58394_ (_07173_, _07167_, _06108_);
  nor _58395_ (_07174_, _07173_, _07172_);
  and _58396_ (_07175_, _07167_, _06913_);
  and _58397_ (_07176_, _06877_, _05748_);
  and _58398_ (_07177_, _06979_, \oc8051_golden_model_1.SP [0]);
  and _58399_ (_07178_, \oc8051_golden_model_1.SP [1], _06142_);
  nor _58400_ (_07179_, _07178_, _07177_);
  nor _58401_ (_07180_, _07179_, _05846_);
  and _58402_ (_07181_, _06913_, _06112_);
  and _58403_ (_07182_, _06135_, _06912_);
  and _58404_ (_07183_, _06273_, _06109_);
  and _58405_ (_07184_, _06127_, _06109_);
  nor _58406_ (_07185_, _07184_, _07183_);
  not _58407_ (_07186_, _07185_);
  nor _58408_ (_07187_, _07186_, _07182_);
  and _58409_ (_07188_, _06877_, _06139_);
  not _58410_ (_07189_, _07179_);
  and _58411_ (_07190_, _07189_, _06151_);
  not _58412_ (_07191_, _06151_);
  and _58413_ (_07192_, _06115_, _06651_);
  not _58414_ (_07193_, \oc8051_golden_model_1.IRAM[0] [1]);
  or _58415_ (_07194_, _06844_, _07193_);
  not _58416_ (_07195_, \oc8051_golden_model_1.IRAM[1] [1]);
  or _58417_ (_07196_, _06993_, _07195_);
  and _58418_ (_07197_, _07196_, _06991_);
  nand _58419_ (_07198_, _07197_, _07194_);
  not _58420_ (_07199_, \oc8051_golden_model_1.IRAM[3] [1]);
  or _58421_ (_07200_, _06993_, _07199_);
  not _58422_ (_07201_, \oc8051_golden_model_1.IRAM[2] [1]);
  or _58423_ (_07202_, _06844_, _07201_);
  and _58424_ (_07203_, _07202_, _06999_);
  nand _58425_ (_07204_, _07203_, _07200_);
  nand _58426_ (_07205_, _07204_, _07198_);
  nand _58427_ (_07206_, _07205_, _06637_);
  not _58428_ (_07207_, \oc8051_golden_model_1.IRAM[7] [1]);
  or _58429_ (_07208_, _06993_, _07207_);
  not _58430_ (_07209_, \oc8051_golden_model_1.IRAM[6] [1]);
  or _58431_ (_07210_, _06844_, _07209_);
  and _58432_ (_07211_, _07210_, _06999_);
  nand _58433_ (_07212_, _07211_, _07208_);
  not _58434_ (_07213_, \oc8051_golden_model_1.IRAM[4] [1]);
  or _58435_ (_07214_, _06844_, _07213_);
  not _58436_ (_07215_, \oc8051_golden_model_1.IRAM[5] [1]);
  or _58437_ (_07216_, _06993_, _07215_);
  and _58438_ (_07217_, _07216_, _06991_);
  nand _58439_ (_07218_, _07217_, _07214_);
  nand _58440_ (_07219_, _07218_, _07212_);
  nand _58441_ (_07220_, _07219_, _07006_);
  nand _58442_ (_07221_, _07220_, _07206_);
  nand _58443_ (_07222_, _07221_, _06446_);
  not _58444_ (_07223_, \oc8051_golden_model_1.IRAM[11] [1]);
  or _58445_ (_07224_, _06993_, _07223_);
  not _58446_ (_07225_, \oc8051_golden_model_1.IRAM[10] [1]);
  or _58447_ (_07226_, _06844_, _07225_);
  and _58448_ (_07227_, _07226_, _06999_);
  nand _58449_ (_07228_, _07227_, _07224_);
  not _58450_ (_07229_, \oc8051_golden_model_1.IRAM[8] [1]);
  or _58451_ (_07230_, _06844_, _07229_);
  not _58452_ (_07231_, \oc8051_golden_model_1.IRAM[9] [1]);
  or _58453_ (_07232_, _06993_, _07231_);
  and _58454_ (_07233_, _07232_, _06991_);
  nand _58455_ (_07234_, _07233_, _07230_);
  nand _58456_ (_07235_, _07234_, _07228_);
  nand _58457_ (_07236_, _07235_, _06637_);
  not _58458_ (_07237_, \oc8051_golden_model_1.IRAM[15] [1]);
  or _58459_ (_07238_, _06993_, _07237_);
  nand _58460_ (_07239_, _06993_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _58461_ (_07240_, _07239_, _06999_);
  nand _58462_ (_07241_, _07240_, _07238_);
  not _58463_ (_07242_, \oc8051_golden_model_1.IRAM[12] [1]);
  or _58464_ (_07243_, _06844_, _07242_);
  not _58465_ (_07244_, \oc8051_golden_model_1.IRAM[13] [1]);
  or _58466_ (_07245_, _06993_, _07244_);
  and _58467_ (_07246_, _07245_, _06991_);
  nand _58468_ (_07247_, _07246_, _07243_);
  nand _58469_ (_07248_, _07247_, _07241_);
  nand _58470_ (_07249_, _07248_, _07006_);
  nand _58471_ (_07250_, _07249_, _07236_);
  nand _58472_ (_07251_, _07250_, _07023_);
  nand _58473_ (_07252_, _07251_, _07222_);
  and _58474_ (_07253_, _07252_, _06164_);
  or _58475_ (_07254_, _07253_, _07192_);
  and _58476_ (_07255_, _07058_, _06912_);
  nor _58477_ (_07256_, _07255_, _07254_);
  and _58478_ (_07257_, _07179_, _06581_);
  not _58479_ (_07258_, _07257_);
  and _58480_ (_07259_, _06119_, _06155_);
  nor _58481_ (_07260_, _07259_, _06584_);
  and _58482_ (_07261_, _07260_, _07258_);
  and _58483_ (_07262_, _07261_, _07256_);
  and _58484_ (_07263_, _07252_, _07064_);
  nor _58485_ (_07264_, _07263_, _06162_);
  and _58486_ (_07265_, _07264_, _07262_);
  and _58487_ (_07266_, _06913_, _06162_);
  nor _58488_ (_07267_, _07266_, _07265_);
  and _58489_ (_07268_, _06876_, _06159_);
  nor _58490_ (_07269_, _07268_, _07267_);
  or _58491_ (_07270_, _07189_, _05764_);
  nand _58492_ (_07271_, _07270_, _07269_);
  and _58493_ (_07272_, _07076_, _06912_);
  and _58494_ (_07273_, _06119_, _06150_);
  nor _58495_ (_07274_, _07273_, _06538_);
  not _58496_ (_07275_, _07274_);
  nor _58497_ (_07276_, _07275_, _07272_);
  not _58498_ (_07277_, _07276_);
  nor _58499_ (_07278_, _07277_, _07271_);
  and _58500_ (_07279_, _07252_, _07081_);
  nor _58501_ (_07280_, _07279_, _07087_);
  and _58502_ (_07281_, _07280_, _07278_);
  and _58503_ (_07282_, _07087_, _06913_);
  nor _58504_ (_07283_, _07282_, _07281_);
  and _58505_ (_07284_, _06876_, _07086_);
  nor _58506_ (_07285_, _07284_, _07283_);
  and _58507_ (_07286_, _07285_, _07191_);
  nor _58508_ (_07287_, _07286_, _07190_);
  and _58509_ (_07288_, _06148_, _06876_);
  or _58510_ (_07289_, _07288_, _07287_);
  nor _58511_ (_07290_, _07189_, _05760_);
  and _58512_ (_07291_, _05744_, _05666_);
  and _58513_ (_07292_, _07291_, _06245_);
  or _58514_ (_07293_, _07292_, _07290_);
  nor _58515_ (_07294_, _07293_, _07289_);
  and _58516_ (_07295_, _07252_, _06701_);
  nor _58517_ (_07296_, _07295_, _07103_);
  and _58518_ (_07297_, _07296_, _07294_);
  nor _58519_ (_07298_, _07297_, _07188_);
  nor _58520_ (_07299_, _07298_, _05791_);
  and _58521_ (_07300_, _07189_, _05791_);
  nor _58522_ (_07301_, _07300_, _07299_);
  or _58523_ (_07302_, _06288_, _06123_);
  and _58524_ (_07303_, _07302_, _06109_);
  nor _58525_ (_07304_, _07303_, _07301_);
  and _58526_ (_07305_, _07304_, _07187_);
  and _58527_ (_07306_, _07251_, _07222_);
  nor _58528_ (_07307_, _07306_, _07116_);
  nor _58529_ (_07308_, _07307_, _06112_);
  and _58530_ (_07309_, _07308_, _07305_);
  nor _58531_ (_07310_, _07309_, _07181_);
  nor _58532_ (_07311_, _07310_, _06076_);
  nor _58533_ (_07312_, _07179_, _05836_);
  nor _58534_ (_07313_, _07312_, _07311_);
  nor _58535_ (_07314_, _07135_, _06913_);
  nor _58536_ (_07315_, _07314_, _07124_);
  not _58537_ (_07316_, _07315_);
  nor _58538_ (_07317_, _07316_, _07313_);
  nor _58539_ (_07318_, _07179_, _05848_);
  nor _58540_ (_07319_, _07318_, _07317_);
  and _58541_ (_07320_, _07143_, _06912_);
  nor _58542_ (_07321_, _07320_, _07142_);
  not _58543_ (_07322_, _07321_);
  nor _58544_ (_07323_, _07322_, _07319_);
  nor _58545_ (_07324_, _07323_, _07180_);
  and _58546_ (_07325_, _06119_, _05591_);
  not _58547_ (_07326_, _07325_);
  and _58548_ (_07327_, _07326_, _06564_);
  not _58549_ (_07328_, _07327_);
  nor _58550_ (_07329_, _07328_, _07324_);
  and _58551_ (_07330_, _07252_, _07153_);
  nor _58552_ (_07331_, _07330_, _07152_);
  and _58553_ (_07332_, _07331_, _07329_);
  and _58554_ (_07333_, _07152_, _06913_);
  nor _58555_ (_07334_, _07333_, _07332_);
  nor _58556_ (_07335_, _07189_, _07160_);
  nor _58557_ (_07336_, _07335_, _06073_);
  not _58558_ (_07337_, _07336_);
  nor _58559_ (_07338_, _07337_, _07334_);
  nor _58560_ (_07339_, _07338_, _07176_);
  and _58561_ (_07340_, _07291_, _05820_);
  nor _58562_ (_07341_, _07340_, _07339_);
  and _58563_ (_07342_, _07252_, _07168_);
  nor _58564_ (_07343_, _07342_, _07167_);
  and _58565_ (_07344_, _07343_, _07341_);
  nor _58566_ (_07345_, _07344_, _07175_);
  not _58567_ (_07346_, _00000_);
  nor _58568_ (_07347_, _07076_, _06159_);
  nor _58569_ (_07348_, _07058_, _06162_);
  and _58570_ (_07349_, _07348_, _07347_);
  not _58571_ (_07350_, _06112_);
  and _58572_ (_07351_, _06125_, _06109_);
  not _58573_ (_07352_, _07351_);
  nor _58574_ (_07353_, _06972_, _06562_);
  and _58575_ (_07354_, _07353_, _06531_);
  and _58576_ (_07355_, _07354_, _07352_);
  nor _58577_ (_07356_, _06563_, _06248_);
  not _58578_ (_07357_, _06950_);
  and _58579_ (_07358_, _07357_, _06540_);
  and _58580_ (_07359_, _07358_, _07356_);
  and _58581_ (_07360_, _05836_, _05764_);
  and _58582_ (_07361_, _07360_, _06582_);
  and _58583_ (_07362_, _07160_, _05850_);
  and _58584_ (_07363_, _07362_, _07361_);
  and _58585_ (_07364_, _07363_, _07359_);
  nor _58586_ (_07365_, _06119_, _06115_);
  nor _58587_ (_07366_, _07365_, _05768_);
  and _58588_ (_07367_, _06249_, _05742_);
  nor _58589_ (_07368_, _07367_, _07366_);
  not _58590_ (_07369_, _05745_);
  and _58591_ (_07370_, _06118_, _06109_);
  and _58592_ (_07371_, _07370_, _07369_);
  nor _58593_ (_07372_, _07365_, _05776_);
  nor _58594_ (_07373_, _07372_, _07371_);
  and _58595_ (_07374_, _07373_, _07368_);
  and _58596_ (_07375_, _07374_, _06247_);
  and _58597_ (_07376_, _07375_, _07364_);
  and _58598_ (_07377_, _06122_, _06155_);
  not _58599_ (_07378_, _07377_);
  and _58600_ (_07379_, _06294_, _06651_);
  and _58601_ (_07380_, _05786_, _06651_);
  nor _58602_ (_07381_, _07380_, _07379_);
  nand _58603_ (_07382_, _07381_, _05777_);
  nor _58604_ (_07383_, _07382_, _07186_);
  and _58605_ (_07384_, _07383_, _07378_);
  nor _58606_ (_07385_, _06701_, _06151_);
  nor _58607_ (_07386_, _07115_, _07064_);
  and _58608_ (_07387_, _07386_, _07385_);
  not _58609_ (_07388_, _05760_);
  nor _58610_ (_07389_, _05791_, _07388_);
  nor _58611_ (_07390_, _07168_, _07153_);
  and _58612_ (_07391_, _07390_, _07389_);
  and _58613_ (_07392_, _07391_, _07387_);
  not _58614_ (_07393_, _06978_);
  and _58615_ (_07394_, _06119_, _05820_);
  nor _58616_ (_07395_, _07394_, _07259_);
  and _58617_ (_07396_, _06119_, _06245_);
  nor _58618_ (_07397_, _07396_, _07325_);
  and _58619_ (_07398_, _07397_, _07395_);
  and _58620_ (_07399_, _07398_, _07393_);
  and _58621_ (_07400_, _07399_, _07392_);
  and _58622_ (_07401_, _07400_, _07384_);
  and _58623_ (_07402_, _07401_, _07376_);
  and _58624_ (_07403_, _07402_, _07355_);
  and _58625_ (_07404_, _07403_, _07350_);
  nor _58626_ (_07405_, _07087_, _07086_);
  and _58627_ (_07406_, _07405_, _07404_);
  and _58628_ (_07407_, _07406_, _07349_);
  not _58629_ (_07408_, _06135_);
  nor _58630_ (_07409_, _07167_, _06073_);
  and _58631_ (_07410_, _07409_, _07408_);
  nor _58632_ (_07411_, _06148_, _07103_);
  nor _58633_ (_07412_, _07152_, _07143_);
  and _58634_ (_07413_, _07412_, _07411_);
  and _58635_ (_07414_, _07413_, _07410_);
  and _58636_ (_07415_, _07414_, _07135_);
  and _58637_ (_07416_, _07415_, _07407_);
  nor _58638_ (_07417_, _07416_, _07346_);
  not _58639_ (_07418_, _07417_);
  nor _58640_ (_07419_, _07418_, _07345_);
  not _58641_ (_07420_, _07419_);
  nor _58642_ (_07421_, _07420_, _07174_);
  not _58643_ (_07422_, \oc8051_golden_model_1.IRAM[0] [3]);
  or _58644_ (_07423_, _06844_, _07422_);
  not _58645_ (_07424_, \oc8051_golden_model_1.IRAM[1] [3]);
  or _58646_ (_07425_, _06993_, _07424_);
  and _58647_ (_07426_, _07425_, _06991_);
  nand _58648_ (_07427_, _07426_, _07423_);
  not _58649_ (_07428_, \oc8051_golden_model_1.IRAM[3] [3]);
  or _58650_ (_07429_, _06993_, _07428_);
  not _58651_ (_07430_, \oc8051_golden_model_1.IRAM[2] [3]);
  or _58652_ (_07431_, _06844_, _07430_);
  and _58653_ (_07432_, _07431_, _06999_);
  nand _58654_ (_07433_, _07432_, _07429_);
  nand _58655_ (_07434_, _07433_, _07427_);
  nand _58656_ (_07435_, _07434_, _06637_);
  not _58657_ (_07436_, \oc8051_golden_model_1.IRAM[7] [3]);
  or _58658_ (_07437_, _06993_, _07436_);
  not _58659_ (_07438_, \oc8051_golden_model_1.IRAM[6] [3]);
  or _58660_ (_07439_, _06844_, _07438_);
  and _58661_ (_07440_, _07439_, _06999_);
  nand _58662_ (_07441_, _07440_, _07437_);
  not _58663_ (_07442_, \oc8051_golden_model_1.IRAM[4] [3]);
  or _58664_ (_07443_, _06844_, _07442_);
  not _58665_ (_07444_, \oc8051_golden_model_1.IRAM[5] [3]);
  or _58666_ (_07445_, _06993_, _07444_);
  and _58667_ (_07446_, _07445_, _06991_);
  nand _58668_ (_07447_, _07446_, _07443_);
  nand _58669_ (_07448_, _07447_, _07441_);
  nand _58670_ (_07449_, _07448_, _07006_);
  nand _58671_ (_07450_, _07449_, _07435_);
  nand _58672_ (_07451_, _07450_, _06446_);
  nand _58673_ (_07452_, _06844_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _58674_ (_07453_, _06993_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _58675_ (_07454_, _07453_, _06999_);
  nand _58676_ (_07455_, _07454_, _07452_);
  nand _58677_ (_07456_, _06993_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand _58678_ (_07457_, _06844_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _58679_ (_07458_, _07457_, _06991_);
  nand _58680_ (_07459_, _07458_, _07456_);
  nand _58681_ (_07460_, _07459_, _07455_);
  nand _58682_ (_07461_, _07460_, _06637_);
  nand _58683_ (_07462_, _06844_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _58684_ (_07463_, _06993_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _58685_ (_07464_, _07463_, _06999_);
  nand _58686_ (_07465_, _07464_, _07462_);
  nand _58687_ (_07466_, _06993_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand _58688_ (_07467_, _06844_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _58689_ (_07468_, _07467_, _06991_);
  nand _58690_ (_07469_, _07468_, _07466_);
  nand _58691_ (_07470_, _07469_, _07465_);
  nand _58692_ (_07471_, _07470_, _07006_);
  nand _58693_ (_07472_, _07471_, _07461_);
  nand _58694_ (_07473_, _07472_, _07023_);
  nand _58695_ (_07474_, _07473_, _07451_);
  and _58696_ (_07475_, _07474_, _07168_);
  and _58697_ (_07476_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _58698_ (_07477_, _07476_, \oc8051_golden_model_1.SP [2]);
  nor _58699_ (_07478_, _07477_, \oc8051_golden_model_1.SP [3]);
  and _58700_ (_07479_, _07477_, \oc8051_golden_model_1.SP [3]);
  nor _58701_ (_07480_, _07479_, _07478_);
  and _58702_ (_07481_, _07480_, _05791_);
  not _58703_ (_07482_, _06203_);
  and _58704_ (_07483_, _07103_, _07482_);
  and _58705_ (_07484_, _07480_, _07388_);
  not _58706_ (_07485_, _05764_);
  and _58707_ (_07486_, _06203_, _06159_);
  and _58708_ (_07487_, _07480_, _06581_);
  and _58709_ (_07488_, _07474_, _06164_);
  nor _58710_ (_07489_, _06164_, \oc8051_golden_model_1.PSW [3]);
  nor _58711_ (_07490_, _07489_, _07058_);
  not _58712_ (_07491_, _07490_);
  nor _58713_ (_07492_, _07491_, _07488_);
  and _58714_ (_07493_, _07058_, _06228_);
  nor _58715_ (_07494_, _07493_, _07492_);
  nor _58716_ (_07495_, _07494_, _06581_);
  or _58717_ (_07496_, _07495_, _07064_);
  nor _58718_ (_07497_, _07496_, _07487_);
  and _58719_ (_07498_, _07474_, _07064_);
  nor _58720_ (_07499_, _07498_, _06162_);
  not _58721_ (_07500_, _07499_);
  nor _58722_ (_07501_, _07500_, _07497_);
  nor _58723_ (_07502_, _06161_, _06071_);
  or _58724_ (_07503_, _07502_, _06159_);
  nor _58725_ (_07504_, _07503_, _07501_);
  nor _58726_ (_07505_, _07504_, _07486_);
  nor _58727_ (_07506_, _07505_, _07485_);
  nor _58728_ (_07507_, _07480_, _05764_);
  nor _58729_ (_07508_, _07507_, _07076_);
  not _58730_ (_07509_, _07508_);
  nor _58731_ (_07510_, _07509_, _07506_);
  and _58732_ (_07511_, _07076_, _06228_);
  nor _58733_ (_07512_, _07511_, _07081_);
  not _58734_ (_07513_, _07512_);
  nor _58735_ (_07514_, _07513_, _07510_);
  and _58736_ (_07515_, _07474_, _07081_);
  nor _58737_ (_07516_, _07515_, _07087_);
  not _58738_ (_07517_, _07516_);
  nor _58739_ (_07518_, _07517_, _07514_);
  and _58740_ (_07519_, _07087_, _06228_);
  or _58741_ (_07520_, _07519_, _07086_);
  nor _58742_ (_07521_, _07520_, _07518_);
  and _58743_ (_07522_, _06203_, _07086_);
  nor _58744_ (_07523_, _07522_, _07521_);
  and _58745_ (_07524_, _07523_, _07191_);
  and _58746_ (_07525_, _07480_, _06151_);
  nor _58747_ (_07526_, _07525_, _07524_);
  nor _58748_ (_07527_, _07526_, _06148_);
  nor _58749_ (_07528_, _06149_, _06206_);
  or _58750_ (_07529_, _07528_, _07527_);
  and _58751_ (_07530_, _07529_, _05760_);
  or _58752_ (_07531_, _07530_, _06701_);
  nor _58753_ (_07532_, _07531_, _07484_);
  and _58754_ (_07533_, _07474_, _06701_);
  nor _58755_ (_07534_, _07533_, _07103_);
  not _58756_ (_07535_, _07534_);
  nor _58757_ (_07536_, _07535_, _07532_);
  nor _58758_ (_07537_, _07536_, _07483_);
  nor _58759_ (_07538_, _07537_, _05791_);
  or _58760_ (_07539_, _07538_, _06135_);
  nor _58761_ (_07540_, _07539_, _07481_);
  and _58762_ (_07541_, _06135_, _06070_);
  or _58763_ (_07542_, _07541_, _07540_);
  and _58764_ (_07543_, _07542_, _07116_);
  and _58765_ (_07544_, _07473_, _07451_);
  nor _58766_ (_07545_, _07544_, _07116_);
  nor _58767_ (_07546_, _07545_, _06112_);
  not _58768_ (_07547_, _07546_);
  nor _58769_ (_07548_, _07547_, _07543_);
  nor _58770_ (_07549_, _06111_, _06071_);
  nor _58771_ (_07550_, _07549_, _07548_);
  nor _58772_ (_07551_, _07550_, _06076_);
  and _58773_ (_07552_, _07480_, _06076_);
  not _58774_ (_07553_, _07552_);
  and _58775_ (_07554_, _07553_, _07135_);
  not _58776_ (_07555_, _07554_);
  nor _58777_ (_07556_, _07555_, _07551_);
  nor _58778_ (_07557_, _07135_, _06228_);
  nor _58779_ (_07558_, _07557_, _07124_);
  not _58780_ (_07559_, _07558_);
  nor _58781_ (_07560_, _07559_, _07556_);
  and _58782_ (_07561_, _07480_, _07124_);
  nor _58783_ (_07562_, _07561_, _07143_);
  not _58784_ (_07563_, _07562_);
  nor _58785_ (_07564_, _07563_, _07560_);
  and _58786_ (_07565_, _07143_, _06070_);
  nor _58787_ (_07566_, _07565_, _07142_);
  not _58788_ (_07567_, _07566_);
  nor _58789_ (_07568_, _07567_, _07564_);
  and _58790_ (_07569_, _07480_, _07142_);
  nor _58791_ (_07570_, _07569_, _07153_);
  not _58792_ (_07571_, _07570_);
  nor _58793_ (_07572_, _07571_, _07568_);
  and _58794_ (_07573_, _07474_, _07153_);
  nor _58795_ (_07574_, _07573_, _07152_);
  not _58796_ (_07575_, _07574_);
  nor _58797_ (_07576_, _07575_, _07572_);
  not _58798_ (_07577_, _07160_);
  and _58799_ (_07578_, _07152_, _06228_);
  nor _58800_ (_07579_, _07578_, _07577_);
  not _58801_ (_07580_, _07579_);
  nor _58802_ (_07581_, _07580_, _07576_);
  nor _58803_ (_07582_, _07480_, _07160_);
  nor _58804_ (_07583_, _07582_, _06073_);
  not _58805_ (_07584_, _07583_);
  nor _58806_ (_07585_, _07584_, _07581_);
  and _58807_ (_07586_, _06073_, _07482_);
  nor _58808_ (_07587_, _07586_, _07168_);
  not _58809_ (_07588_, _07587_);
  nor _58810_ (_07589_, _07588_, _07585_);
  or _58811_ (_07590_, _07589_, _07167_);
  nor _58812_ (_07591_, _07590_, _07475_);
  and _58813_ (_07592_, _07167_, _06228_);
  nor _58814_ (_07593_, _07592_, _07591_);
  and _58815_ (_07594_, _06478_, _05748_);
  nor _58816_ (_07595_, _07476_, \oc8051_golden_model_1.SP [2]);
  nor _58817_ (_07596_, _07595_, _07477_);
  not _58818_ (_07597_, _07596_);
  nor _58819_ (_07598_, _07597_, _05846_);
  and _58820_ (_07599_, _06626_, _06112_);
  and _58821_ (_07600_, _06478_, _06139_);
  and _58822_ (_07601_, _07596_, _06151_);
  and _58823_ (_07602_, _06626_, _06162_);
  not _58824_ (_07603_, \oc8051_golden_model_1.IRAM[0] [2]);
  or _58825_ (_07604_, _06844_, _07603_);
  not _58826_ (_07605_, \oc8051_golden_model_1.IRAM[1] [2]);
  or _58827_ (_07606_, _06993_, _07605_);
  and _58828_ (_07607_, _07606_, _06991_);
  nand _58829_ (_07608_, _07607_, _07604_);
  not _58830_ (_07609_, \oc8051_golden_model_1.IRAM[3] [2]);
  or _58831_ (_07610_, _06993_, _07609_);
  not _58832_ (_07611_, \oc8051_golden_model_1.IRAM[2] [2]);
  or _58833_ (_07612_, _06844_, _07611_);
  and _58834_ (_07613_, _07612_, _06999_);
  nand _58835_ (_07614_, _07613_, _07610_);
  nand _58836_ (_07615_, _07614_, _07608_);
  nand _58837_ (_07616_, _07615_, _06637_);
  not _58838_ (_07617_, \oc8051_golden_model_1.IRAM[7] [2]);
  or _58839_ (_07618_, _06993_, _07617_);
  not _58840_ (_07619_, \oc8051_golden_model_1.IRAM[6] [2]);
  or _58841_ (_07620_, _06844_, _07619_);
  and _58842_ (_07621_, _07620_, _06999_);
  nand _58843_ (_07622_, _07621_, _07618_);
  not _58844_ (_07623_, \oc8051_golden_model_1.IRAM[4] [2]);
  or _58845_ (_07624_, _06844_, _07623_);
  not _58846_ (_07625_, \oc8051_golden_model_1.IRAM[5] [2]);
  or _58847_ (_07626_, _06993_, _07625_);
  and _58848_ (_07627_, _07626_, _06991_);
  nand _58849_ (_07628_, _07627_, _07624_);
  nand _58850_ (_07629_, _07628_, _07622_);
  nand _58851_ (_07630_, _07629_, _07006_);
  nand _58852_ (_07631_, _07630_, _07616_);
  nand _58853_ (_07632_, _07631_, _06446_);
  not _58854_ (_07633_, \oc8051_golden_model_1.IRAM[11] [2]);
  or _58855_ (_07634_, _06993_, _07633_);
  not _58856_ (_07635_, \oc8051_golden_model_1.IRAM[10] [2]);
  or _58857_ (_07636_, _06844_, _07635_);
  and _58858_ (_07637_, _07636_, _06999_);
  nand _58859_ (_07638_, _07637_, _07634_);
  nand _58860_ (_07639_, _06993_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand _58861_ (_07640_, _06844_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _58862_ (_07641_, _07640_, _06991_);
  nand _58863_ (_07642_, _07641_, _07639_);
  nand _58864_ (_07643_, _07642_, _07638_);
  nand _58865_ (_07644_, _07643_, _06637_);
  nand _58866_ (_07645_, _06844_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _58867_ (_07646_, _06993_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _58868_ (_07647_, _07646_, _06999_);
  nand _58869_ (_07648_, _07647_, _07645_);
  nand _58870_ (_07649_, _06993_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand _58871_ (_07650_, _06844_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _58872_ (_07651_, _07650_, _06991_);
  nand _58873_ (_07652_, _07651_, _07649_);
  nand _58874_ (_07653_, _07652_, _07648_);
  nand _58875_ (_07654_, _07653_, _07006_);
  nand _58876_ (_07655_, _07654_, _07644_);
  nand _58877_ (_07656_, _07655_, _07023_);
  nand _58878_ (_07657_, _07656_, _07632_);
  or _58879_ (_07658_, _07657_, _05752_);
  and _58880_ (_07659_, _07658_, _07382_);
  and _58881_ (_07660_, _07058_, _06625_);
  nor _58882_ (_07661_, _07660_, _07659_);
  and _58883_ (_07662_, _07597_, _06581_);
  not _58884_ (_07663_, _07662_);
  and _58885_ (_07664_, _06273_, _06155_);
  and _58886_ (_07665_, _06288_, _06155_);
  or _58887_ (_07666_, _07665_, _06978_);
  nor _58888_ (_07667_, _07666_, _07664_);
  and _58889_ (_07668_, _07667_, _07663_);
  and _58890_ (_07669_, _07668_, _07661_);
  and _58891_ (_07670_, _07657_, _07064_);
  nor _58892_ (_07671_, _07670_, _06162_);
  and _58893_ (_07672_, _07671_, _07669_);
  nor _58894_ (_07673_, _07672_, _07602_);
  nor _58895_ (_07674_, _07673_, _06159_);
  nor _58896_ (_07675_, _07674_, _06489_);
  nor _58897_ (_07676_, _07596_, _05764_);
  nor _58898_ (_07677_, _07676_, _07675_);
  and _58899_ (_07678_, _06118_, _06150_);
  and _58900_ (_07679_, _07076_, _06625_);
  nor _58901_ (_07680_, _07679_, _07678_);
  and _58902_ (_07681_, _07680_, _07677_);
  and _58903_ (_07682_, _07657_, _07081_);
  nor _58904_ (_07683_, _07682_, _07087_);
  and _58905_ (_07684_, _07683_, _07681_);
  and _58906_ (_07685_, _07087_, _06626_);
  nor _58907_ (_07686_, _07685_, _07684_);
  and _58908_ (_07687_, _06477_, _07086_);
  nor _58909_ (_07688_, _07687_, _07686_);
  and _58910_ (_07689_, _07688_, _07191_);
  nor _58911_ (_07690_, _07689_, _07601_);
  and _58912_ (_07691_, _06148_, _06477_);
  or _58913_ (_07692_, _07691_, _07690_);
  nor _58914_ (_07693_, _07596_, _05760_);
  nor _58915_ (_07694_, _07693_, _06249_);
  not _58916_ (_07695_, _07694_);
  nor _58917_ (_07696_, _07695_, _07692_);
  and _58918_ (_07697_, _07657_, _06701_);
  nor _58919_ (_07698_, _07697_, _07103_);
  and _58920_ (_07699_, _07698_, _07696_);
  nor _58921_ (_07700_, _07699_, _07600_);
  nor _58922_ (_07701_, _07700_, _05791_);
  and _58923_ (_07702_, _07596_, _05791_);
  nor _58924_ (_07703_, _07702_, _07701_);
  and _58925_ (_07704_, _06135_, _06625_);
  nor _58926_ (_07705_, _07704_, _07370_);
  not _58927_ (_07706_, _07705_);
  nor _58928_ (_07707_, _07706_, _07703_);
  and _58929_ (_07708_, _07656_, _07632_);
  nor _58930_ (_07709_, _07708_, _07116_);
  nor _58931_ (_07710_, _07709_, _06112_);
  and _58932_ (_07711_, _07710_, _07707_);
  nor _58933_ (_07712_, _07711_, _07599_);
  nor _58934_ (_07713_, _07712_, _06076_);
  nor _58935_ (_07714_, _07597_, _05836_);
  nor _58936_ (_07715_, _07714_, _07713_);
  nor _58937_ (_07716_, _07135_, _06626_);
  nor _58938_ (_07717_, _07716_, _07124_);
  not _58939_ (_07718_, _07717_);
  nor _58940_ (_07719_, _07718_, _07715_);
  nor _58941_ (_07720_, _07597_, _05848_);
  nor _58942_ (_07721_, _07720_, _07719_);
  and _58943_ (_07722_, _07143_, _06625_);
  nor _58944_ (_07723_, _07722_, _07142_);
  not _58945_ (_07724_, _07723_);
  nor _58946_ (_07725_, _07724_, _07721_);
  nor _58947_ (_07726_, _07725_, _07598_);
  nor _58948_ (_07727_, _07325_, _06972_);
  not _58949_ (_07728_, _07727_);
  nor _58950_ (_07729_, _07728_, _07726_);
  and _58951_ (_07730_, _07657_, _07153_);
  nor _58952_ (_07731_, _07730_, _07152_);
  and _58953_ (_07732_, _07731_, _07729_);
  and _58954_ (_07733_, _07152_, _06626_);
  nor _58955_ (_07734_, _07733_, _07732_);
  nor _58956_ (_07735_, _07596_, _07160_);
  nor _58957_ (_07736_, _07735_, _06073_);
  not _58958_ (_07737_, _07736_);
  nor _58959_ (_07738_, _07737_, _07734_);
  nor _58960_ (_07739_, _07738_, _07594_);
  and _58961_ (_07740_, _06118_, _05820_);
  nor _58962_ (_07741_, _07740_, _07739_);
  and _58963_ (_07742_, _07657_, _07168_);
  nor _58964_ (_07743_, _07742_, _07167_);
  and _58965_ (_07744_, _07743_, _07741_);
  and _58966_ (_07745_, _07167_, _06626_);
  nor _58967_ (_07746_, _07745_, _07744_);
  nor _58968_ (_07747_, _07746_, _07418_);
  not _58969_ (_07748_, _07747_);
  nor _58970_ (_07749_, _07748_, _07593_);
  and _58971_ (_07750_, _07749_, _07421_);
  or _58972_ (_07751_, _07750_, \oc8051_golden_model_1.IRAM[15] [7]);
  and _58973_ (_07752_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _58974_ (_07753_, _07752_, _06142_);
  nor _58975_ (_07754_, _07596_, _07178_);
  nor _58976_ (_07755_, _07754_, _07753_);
  and _58977_ (_07756_, _07752_, \oc8051_golden_model_1.SP [3]);
  and _58978_ (_07757_, _07756_, _06142_);
  nor _58979_ (_07758_, _07753_, _07480_);
  nor _58980_ (_07759_, _07758_, _07757_);
  and _58981_ (_07760_, _07389_, _07360_);
  and _58982_ (_07761_, _07160_, _06582_);
  and _58983_ (_07762_, _07761_, _05850_);
  and _58984_ (_07763_, _07762_, _07760_);
  nor _58985_ (_07764_, _07763_, _07346_);
  and _58986_ (_07765_, _07764_, _07759_);
  and _58987_ (_07766_, _07765_, _07755_);
  and _58988_ (_07767_, _07766_, _07177_);
  not _58989_ (_07768_, _07767_);
  and _58990_ (_07769_, _07768_, _07751_);
  not _58991_ (_07770_, _07750_);
  and _58992_ (_07771_, _06912_, _06107_);
  and _58993_ (_07772_, _07771_, _06625_);
  and _58994_ (_07773_, _07772_, _06228_);
  and _58995_ (_07774_, _06203_, _06039_);
  not _58996_ (_07775_, _06876_);
  and _58997_ (_07776_, _07775_, _06477_);
  and _58998_ (_07777_, _07776_, _07774_);
  and _58999_ (_07778_, _07777_, _07773_);
  and _59000_ (_07779_, _07778_, \oc8051_golden_model_1.SCON [7]);
  and _59001_ (_07780_, _06912_, _06108_);
  and _59002_ (_07781_, _07780_, _06625_);
  and _59003_ (_07782_, _07781_, _06228_);
  and _59004_ (_07783_, _07782_, _07777_);
  and _59005_ (_07784_, _07783_, \oc8051_golden_model_1.SBUF [7]);
  or _59006_ (_07785_, _07784_, _07779_);
  and _59007_ (_07786_, _07774_, _06477_);
  and _59008_ (_07787_, _07786_, _06876_);
  and _59009_ (_07788_, _07787_, _07773_);
  and _59010_ (_07789_, _07788_, \oc8051_golden_model_1.TCON [7]);
  nand _59011_ (_07790_, _07772_, _06070_);
  nor _59012_ (_07791_, _06203_, _06172_);
  and _59013_ (_07792_, _07791_, _07776_);
  not _59014_ (_07793_, _07792_);
  nor _59015_ (_07794_, _07793_, _07790_);
  and _59016_ (_07795_, _07794_, \oc8051_golden_model_1.PSW [7]);
  or _59017_ (_07796_, _07795_, _07789_);
  or _59018_ (_07797_, _07796_, _07785_);
  not _59019_ (_07798_, _07787_);
  nand _59020_ (_07799_, _06625_, _06228_);
  nor _59021_ (_07800_, _06912_, _06108_);
  not _59022_ (_07801_, _07800_);
  or _59023_ (_07802_, _07801_, _07799_);
  nor _59024_ (_07803_, _07802_, _07798_);
  and _59025_ (_07804_, _07803_, \oc8051_golden_model_1.TL0 [7]);
  not _59026_ (_07805_, _06477_);
  and _59027_ (_07806_, _06876_, _07805_);
  and _59028_ (_07807_, _07806_, _07791_);
  not _59029_ (_07808_, _07807_);
  nor _59030_ (_07809_, _07808_, _07790_);
  and _59031_ (_07810_, _07809_, \oc8051_golden_model_1.ACC [7]);
  or _59032_ (_07811_, _07810_, _07804_);
  and _59033_ (_07812_, _07787_, _07782_);
  and _59034_ (_07813_, _07812_, \oc8051_golden_model_1.TMOD [7]);
  not _59035_ (_07814_, _07780_);
  or _59036_ (_07815_, _06625_, _06070_);
  or _59037_ (_07816_, _07815_, _07814_);
  nor _59038_ (_07817_, _07816_, _07798_);
  and _59039_ (_07818_, _07817_, \oc8051_golden_model_1.TH1 [7]);
  or _59040_ (_07819_, _07818_, _07813_);
  or _59041_ (_07820_, _07819_, _07811_);
  not _59042_ (_07821_, _07771_);
  or _59043_ (_07822_, _07815_, _07821_);
  nor _59044_ (_07823_, _07822_, _07798_);
  and _59045_ (_07824_, _07823_, \oc8051_golden_model_1.TH0 [7]);
  and _59046_ (_07825_, _07806_, _07774_);
  and _59047_ (_07826_, _07825_, _07773_);
  and _59048_ (_07827_, _07826_, \oc8051_golden_model_1.IE [7]);
  nor _59049_ (_07828_, _06876_, _06477_);
  and _59050_ (_07829_, _07828_, _07774_);
  and _59051_ (_07830_, _07829_, _07773_);
  and _59052_ (_07831_, _07830_, \oc8051_golden_model_1.IP [7]);
  or _59053_ (_07832_, _07831_, _07827_);
  or _59054_ (_07833_, _07832_, _07824_);
  nor _59055_ (_07834_, _06912_, _06107_);
  not _59056_ (_07835_, _07834_);
  or _59057_ (_07836_, _07835_, _07799_);
  nor _59058_ (_07837_, _07836_, _07798_);
  and _59059_ (_07838_, _07837_, \oc8051_golden_model_1.TL1 [7]);
  and _59060_ (_07839_, _07828_, _07791_);
  not _59061_ (_07840_, _07839_);
  nor _59062_ (_07841_, _07840_, _07790_);
  and _59063_ (_07842_, _07841_, \oc8051_golden_model_1.B [7]);
  or _59064_ (_07843_, _07842_, _07838_);
  or _59065_ (_07844_, _07843_, _07833_);
  or _59066_ (_07845_, _07844_, _07820_);
  or _59067_ (_07846_, _07845_, _07797_);
  and _59068_ (_07847_, _07787_, _06070_);
  and _59069_ (_07848_, _07800_, _06625_);
  and _59070_ (_07849_, _07848_, _07847_);
  and _59071_ (_07850_, _07849_, \oc8051_golden_model_1.DPL [7]);
  and _59072_ (_07851_, _07834_, _06625_);
  and _59073_ (_07852_, _07851_, _07847_);
  and _59074_ (_07853_, _07852_, \oc8051_golden_model_1.DPH [7]);
  or _59075_ (_07854_, _07853_, _07850_);
  and _59076_ (_07855_, _07834_, _06626_);
  and _59077_ (_07856_, _07855_, _07847_);
  and _59078_ (_07857_, _07856_, \oc8051_golden_model_1.PCON [7]);
  and _59079_ (_07858_, _07847_, _07781_);
  and _59080_ (_07859_, _07858_, \oc8051_golden_model_1.SP [7]);
  or _59081_ (_07860_, _07859_, _07857_);
  or _59082_ (_07861_, _07860_, _07854_);
  or _59083_ (_07862_, _07861_, _07846_);
  not _59084_ (_07863_, \oc8051_golden_model_1.IRAM[0] [7]);
  or _59085_ (_07864_, _06844_, _07863_);
  not _59086_ (_07865_, \oc8051_golden_model_1.IRAM[1] [7]);
  or _59087_ (_07866_, _06993_, _07865_);
  and _59088_ (_07867_, _07866_, _06991_);
  nand _59089_ (_07868_, _07867_, _07864_);
  not _59090_ (_07869_, \oc8051_golden_model_1.IRAM[3] [7]);
  or _59091_ (_07870_, _06993_, _07869_);
  not _59092_ (_07871_, \oc8051_golden_model_1.IRAM[2] [7]);
  or _59093_ (_07872_, _06844_, _07871_);
  and _59094_ (_07873_, _07872_, _06999_);
  nand _59095_ (_07874_, _07873_, _07870_);
  nand _59096_ (_07875_, _07874_, _07868_);
  nand _59097_ (_07876_, _07875_, _06637_);
  not _59098_ (_07877_, \oc8051_golden_model_1.IRAM[7] [7]);
  or _59099_ (_07878_, _06993_, _07877_);
  not _59100_ (_07879_, \oc8051_golden_model_1.IRAM[6] [7]);
  or _59101_ (_07880_, _06844_, _07879_);
  and _59102_ (_07881_, _07880_, _06999_);
  nand _59103_ (_07882_, _07881_, _07878_);
  not _59104_ (_07883_, \oc8051_golden_model_1.IRAM[4] [7]);
  or _59105_ (_07884_, _06844_, _07883_);
  not _59106_ (_07885_, \oc8051_golden_model_1.IRAM[5] [7]);
  or _59107_ (_07886_, _06993_, _07885_);
  and _59108_ (_07887_, _07886_, _06991_);
  nand _59109_ (_07888_, _07887_, _07884_);
  nand _59110_ (_07889_, _07888_, _07882_);
  nand _59111_ (_07890_, _07889_, _07006_);
  nand _59112_ (_07891_, _07890_, _07876_);
  nand _59113_ (_07892_, _07891_, _06446_);
  not _59114_ (_07893_, \oc8051_golden_model_1.IRAM[11] [7]);
  or _59115_ (_07894_, _06993_, _07893_);
  not _59116_ (_07895_, \oc8051_golden_model_1.IRAM[10] [7]);
  or _59117_ (_07896_, _06844_, _07895_);
  and _59118_ (_07897_, _07896_, _06999_);
  nand _59119_ (_07898_, _07897_, _07894_);
  not _59120_ (_07899_, \oc8051_golden_model_1.IRAM[8] [7]);
  or _59121_ (_07900_, _06844_, _07899_);
  not _59122_ (_07901_, \oc8051_golden_model_1.IRAM[9] [7]);
  or _59123_ (_07902_, _06993_, _07901_);
  and _59124_ (_07903_, _07902_, _06991_);
  nand _59125_ (_07904_, _07903_, _07900_);
  nand _59126_ (_07905_, _07904_, _07898_);
  nand _59127_ (_07906_, _07905_, _06637_);
  not _59128_ (_07907_, \oc8051_golden_model_1.IRAM[15] [7]);
  or _59129_ (_07908_, _06993_, _07907_);
  not _59130_ (_07909_, \oc8051_golden_model_1.IRAM[14] [7]);
  or _59131_ (_07910_, _06844_, _07909_);
  and _59132_ (_07911_, _07910_, _06999_);
  nand _59133_ (_07912_, _07911_, _07908_);
  not _59134_ (_07913_, \oc8051_golden_model_1.IRAM[12] [7]);
  or _59135_ (_07914_, _06844_, _07913_);
  not _59136_ (_07915_, \oc8051_golden_model_1.IRAM[13] [7]);
  or _59137_ (_07916_, _06993_, _07915_);
  and _59138_ (_07917_, _07916_, _06991_);
  nand _59139_ (_07918_, _07917_, _07914_);
  nand _59140_ (_07919_, _07918_, _07912_);
  nand _59141_ (_07920_, _07919_, _07006_);
  nand _59142_ (_07921_, _07920_, _07906_);
  nand _59143_ (_07922_, _07921_, _07023_);
  and _59144_ (_07923_, _07922_, _07892_);
  and _59145_ (_07924_, _07923_, _06172_);
  nor _59146_ (_07925_, _07924_, _07862_);
  not _59147_ (_07926_, _07925_);
  and _59148_ (_07927_, _07837_, \oc8051_golden_model_1.TL1 [6]);
  and _59149_ (_07928_, _07817_, \oc8051_golden_model_1.TH1 [6]);
  or _59150_ (_07929_, _07928_, _07927_);
  and _59151_ (_07930_, _07788_, \oc8051_golden_model_1.TCON [6]);
  and _59152_ (_07931_, _07812_, \oc8051_golden_model_1.TMOD [6]);
  or _59153_ (_07932_, _07931_, _07930_);
  or _59154_ (_07933_, _07932_, _07929_);
  and _59155_ (_07934_, _07803_, \oc8051_golden_model_1.TL0 [6]);
  and _59156_ (_07935_, _07778_, \oc8051_golden_model_1.SCON [6]);
  or _59157_ (_07936_, _07935_, _07934_);
  and _59158_ (_07937_, _07823_, \oc8051_golden_model_1.TH0 [6]);
  and _59159_ (_07938_, _07794_, \oc8051_golden_model_1.PSW [6]);
  or _59160_ (_07939_, _07938_, _07937_);
  or _59161_ (_07940_, _07939_, _07936_);
  and _59162_ (_07941_, _07841_, \oc8051_golden_model_1.B [6]);
  and _59163_ (_07942_, _07826_, \oc8051_golden_model_1.IE [6]);
  and _59164_ (_07943_, _07830_, \oc8051_golden_model_1.IP [6]);
  or _59165_ (_07944_, _07943_, _07942_);
  or _59166_ (_07945_, _07944_, _07941_);
  and _59167_ (_07946_, _07783_, \oc8051_golden_model_1.SBUF [6]);
  and _59168_ (_07947_, _07809_, \oc8051_golden_model_1.ACC [6]);
  or _59169_ (_07948_, _07947_, _07946_);
  or _59170_ (_07949_, _07948_, _07945_);
  or _59171_ (_07950_, _07949_, _07940_);
  or _59172_ (_07951_, _07950_, _07933_);
  and _59173_ (_07952_, _07856_, \oc8051_golden_model_1.PCON [6]);
  and _59174_ (_07953_, _07852_, \oc8051_golden_model_1.DPH [6]);
  or _59175_ (_07954_, _07953_, _07952_);
  and _59176_ (_07955_, _07849_, \oc8051_golden_model_1.DPL [6]);
  and _59177_ (_07956_, _07858_, \oc8051_golden_model_1.SP [6]);
  or _59178_ (_07957_, _07956_, _07955_);
  or _59179_ (_07958_, _07957_, _07954_);
  or _59180_ (_07959_, _07958_, _07951_);
  not _59181_ (_07960_, \oc8051_golden_model_1.IRAM[0] [6]);
  or _59182_ (_07961_, _06844_, _07960_);
  not _59183_ (_07962_, \oc8051_golden_model_1.IRAM[1] [6]);
  or _59184_ (_07963_, _06993_, _07962_);
  and _59185_ (_07964_, _07963_, _06991_);
  nand _59186_ (_07965_, _07964_, _07961_);
  not _59187_ (_07966_, \oc8051_golden_model_1.IRAM[3] [6]);
  or _59188_ (_07967_, _06993_, _07966_);
  not _59189_ (_07968_, \oc8051_golden_model_1.IRAM[2] [6]);
  or _59190_ (_07969_, _06844_, _07968_);
  and _59191_ (_07970_, _07969_, _06999_);
  nand _59192_ (_07971_, _07970_, _07967_);
  nand _59193_ (_07972_, _07971_, _07965_);
  nand _59194_ (_07973_, _07972_, _06637_);
  not _59195_ (_07974_, \oc8051_golden_model_1.IRAM[7] [6]);
  or _59196_ (_07975_, _06993_, _07974_);
  not _59197_ (_07976_, \oc8051_golden_model_1.IRAM[6] [6]);
  or _59198_ (_07977_, _06844_, _07976_);
  and _59199_ (_07978_, _07977_, _06999_);
  nand _59200_ (_07979_, _07978_, _07975_);
  not _59201_ (_07980_, \oc8051_golden_model_1.IRAM[4] [6]);
  or _59202_ (_07981_, _06844_, _07980_);
  not _59203_ (_07982_, \oc8051_golden_model_1.IRAM[5] [6]);
  or _59204_ (_07983_, _06993_, _07982_);
  and _59205_ (_07984_, _07983_, _06991_);
  nand _59206_ (_07985_, _07984_, _07981_);
  nand _59207_ (_07986_, _07985_, _07979_);
  nand _59208_ (_07987_, _07986_, _07006_);
  nand _59209_ (_07988_, _07987_, _07973_);
  nand _59210_ (_07989_, _07988_, _06446_);
  nand _59211_ (_07990_, _06844_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _59212_ (_07991_, _06993_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _59213_ (_07992_, _07991_, _06999_);
  nand _59214_ (_07993_, _07992_, _07990_);
  nand _59215_ (_07994_, _06993_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand _59216_ (_07995_, _06844_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _59217_ (_07996_, _07995_, _06991_);
  nand _59218_ (_07997_, _07996_, _07994_);
  nand _59219_ (_07998_, _07997_, _07993_);
  nand _59220_ (_07999_, _07998_, _06637_);
  nand _59221_ (_08000_, _06844_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _59222_ (_08001_, _06993_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _59223_ (_08002_, _08001_, _06999_);
  nand _59224_ (_08003_, _08002_, _08000_);
  nand _59225_ (_08004_, _06993_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand _59226_ (_08005_, _06844_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _59227_ (_08006_, _08005_, _06991_);
  nand _59228_ (_08007_, _08006_, _08004_);
  nand _59229_ (_08008_, _08007_, _08003_);
  nand _59230_ (_08009_, _08008_, _07006_);
  nand _59231_ (_08010_, _08009_, _07999_);
  nand _59232_ (_08011_, _08010_, _07023_);
  and _59233_ (_08012_, _08011_, _07989_);
  and _59234_ (_08013_, _08012_, _06172_);
  nor _59235_ (_08014_, _08013_, _07959_);
  not _59236_ (_08015_, _08014_);
  and _59237_ (_08016_, _07788_, \oc8051_golden_model_1.TCON [5]);
  and _59238_ (_08017_, _07812_, \oc8051_golden_model_1.TMOD [5]);
  or _59239_ (_08018_, _08017_, _08016_);
  and _59240_ (_08019_, _07778_, \oc8051_golden_model_1.SCON [5]);
  and _59241_ (_08020_, _07794_, \oc8051_golden_model_1.PSW [5]);
  or _59242_ (_08021_, _08020_, _08019_);
  or _59243_ (_08022_, _08021_, _08018_);
  and _59244_ (_08023_, _07817_, \oc8051_golden_model_1.TH1 [5]);
  and _59245_ (_08024_, _07783_, \oc8051_golden_model_1.SBUF [5]);
  or _59246_ (_08025_, _08024_, _08023_);
  and _59247_ (_08026_, _07803_, \oc8051_golden_model_1.TL0 [5]);
  and _59248_ (_08027_, _07837_, \oc8051_golden_model_1.TL1 [5]);
  or _59249_ (_08028_, _08027_, _08026_);
  or _59250_ (_08029_, _08028_, _08025_);
  and _59251_ (_08030_, _07841_, \oc8051_golden_model_1.B [5]);
  and _59252_ (_08031_, _07826_, \oc8051_golden_model_1.IE [5]);
  and _59253_ (_08032_, _07830_, \oc8051_golden_model_1.IP [5]);
  or _59254_ (_08033_, _08032_, _08031_);
  or _59255_ (_08034_, _08033_, _08030_);
  and _59256_ (_08035_, _07823_, \oc8051_golden_model_1.TH0 [5]);
  and _59257_ (_08036_, _07809_, \oc8051_golden_model_1.ACC [5]);
  or _59258_ (_08037_, _08036_, _08035_);
  or _59259_ (_08038_, _08037_, _08034_);
  or _59260_ (_08039_, _08038_, _08029_);
  or _59261_ (_08040_, _08039_, _08022_);
  and _59262_ (_08041_, _07849_, \oc8051_golden_model_1.DPL [5]);
  and _59263_ (_08042_, _07852_, \oc8051_golden_model_1.DPH [5]);
  or _59264_ (_08043_, _08042_, _08041_);
  and _59265_ (_08044_, _07856_, \oc8051_golden_model_1.PCON [5]);
  and _59266_ (_08045_, _07858_, \oc8051_golden_model_1.SP [5]);
  or _59267_ (_08046_, _08045_, _08044_);
  or _59268_ (_08047_, _08046_, _08043_);
  or _59269_ (_08048_, _08047_, _08040_);
  not _59270_ (_08049_, \oc8051_golden_model_1.IRAM[0] [5]);
  or _59271_ (_08050_, _06844_, _08049_);
  not _59272_ (_08051_, \oc8051_golden_model_1.IRAM[1] [5]);
  or _59273_ (_08052_, _06993_, _08051_);
  and _59274_ (_08053_, _08052_, _06991_);
  nand _59275_ (_08054_, _08053_, _08050_);
  not _59276_ (_08055_, \oc8051_golden_model_1.IRAM[3] [5]);
  or _59277_ (_08056_, _06993_, _08055_);
  not _59278_ (_08057_, \oc8051_golden_model_1.IRAM[2] [5]);
  or _59279_ (_08058_, _06844_, _08057_);
  and _59280_ (_08059_, _08058_, _06999_);
  nand _59281_ (_08060_, _08059_, _08056_);
  nand _59282_ (_08061_, _08060_, _08054_);
  nand _59283_ (_08062_, _08061_, _06637_);
  not _59284_ (_08063_, \oc8051_golden_model_1.IRAM[7] [5]);
  or _59285_ (_08064_, _06993_, _08063_);
  not _59286_ (_08065_, \oc8051_golden_model_1.IRAM[6] [5]);
  or _59287_ (_08066_, _06844_, _08065_);
  and _59288_ (_08067_, _08066_, _06999_);
  nand _59289_ (_08068_, _08067_, _08064_);
  not _59290_ (_08069_, \oc8051_golden_model_1.IRAM[4] [5]);
  or _59291_ (_08070_, _06844_, _08069_);
  not _59292_ (_08071_, \oc8051_golden_model_1.IRAM[5] [5]);
  or _59293_ (_08072_, _06993_, _08071_);
  and _59294_ (_08073_, _08072_, _06991_);
  nand _59295_ (_08074_, _08073_, _08070_);
  nand _59296_ (_08075_, _08074_, _08068_);
  nand _59297_ (_08076_, _08075_, _07006_);
  nand _59298_ (_08077_, _08076_, _08062_);
  nand _59299_ (_08078_, _08077_, _06446_);
  nand _59300_ (_08079_, _06844_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _59301_ (_08080_, _06993_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _59302_ (_08081_, _08080_, _06999_);
  nand _59303_ (_08082_, _08081_, _08079_);
  nand _59304_ (_08083_, _06993_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand _59305_ (_08084_, _06844_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _59306_ (_08085_, _08084_, _06991_);
  nand _59307_ (_08086_, _08085_, _08083_);
  nand _59308_ (_08087_, _08086_, _08082_);
  nand _59309_ (_08088_, _08087_, _06637_);
  nand _59310_ (_08089_, _06844_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _59311_ (_08090_, _06993_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _59312_ (_08091_, _08090_, _06999_);
  nand _59313_ (_08092_, _08091_, _08089_);
  nand _59314_ (_08093_, _06993_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand _59315_ (_08094_, _06844_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _59316_ (_08095_, _08094_, _06991_);
  nand _59317_ (_08096_, _08095_, _08093_);
  nand _59318_ (_08097_, _08096_, _08092_);
  nand _59319_ (_08098_, _08097_, _07006_);
  nand _59320_ (_08099_, _08098_, _08088_);
  nand _59321_ (_08100_, _08099_, _07023_);
  and _59322_ (_08101_, _08100_, _08078_);
  and _59323_ (_08102_, _08101_, _06172_);
  nor _59324_ (_08103_, _08102_, _08048_);
  not _59325_ (_08104_, _08103_);
  and _59326_ (_08105_, _07788_, \oc8051_golden_model_1.TCON [3]);
  and _59327_ (_08106_, _07812_, \oc8051_golden_model_1.TMOD [3]);
  or _59328_ (_08107_, _08106_, _08105_);
  and _59329_ (_08108_, _07778_, \oc8051_golden_model_1.SCON [3]);
  and _59330_ (_08109_, _07794_, \oc8051_golden_model_1.PSW [3]);
  or _59331_ (_08110_, _08109_, _08108_);
  or _59332_ (_08111_, _08110_, _08107_);
  and _59333_ (_08112_, _07823_, \oc8051_golden_model_1.TH0 [3]);
  and _59334_ (_08113_, _07837_, \oc8051_golden_model_1.TL1 [3]);
  or _59335_ (_08114_, _08113_, _08112_);
  and _59336_ (_08115_, _07803_, \oc8051_golden_model_1.TL0 [3]);
  and _59337_ (_08116_, _07817_, \oc8051_golden_model_1.TH1 [3]);
  or _59338_ (_08117_, _08116_, _08115_);
  or _59339_ (_08118_, _08117_, _08114_);
  and _59340_ (_08119_, _07841_, \oc8051_golden_model_1.B [3]);
  and _59341_ (_08120_, _07826_, \oc8051_golden_model_1.IE [3]);
  and _59342_ (_08121_, _07830_, \oc8051_golden_model_1.IP [3]);
  or _59343_ (_08122_, _08121_, _08120_);
  or _59344_ (_08123_, _08122_, _08119_);
  and _59345_ (_08124_, _07783_, \oc8051_golden_model_1.SBUF [3]);
  and _59346_ (_08125_, _07809_, \oc8051_golden_model_1.ACC [3]);
  or _59347_ (_08126_, _08125_, _08124_);
  or _59348_ (_08127_, _08126_, _08123_);
  or _59349_ (_08128_, _08127_, _08118_);
  or _59350_ (_08129_, _08128_, _08111_);
  and _59351_ (_08130_, _07856_, \oc8051_golden_model_1.PCON [3]);
  and _59352_ (_08131_, _07858_, \oc8051_golden_model_1.SP [3]);
  or _59353_ (_08132_, _08131_, _08130_);
  and _59354_ (_08133_, _07849_, \oc8051_golden_model_1.DPL [3]);
  and _59355_ (_08134_, _07852_, \oc8051_golden_model_1.DPH [3]);
  or _59356_ (_08135_, _08134_, _08133_);
  or _59357_ (_08136_, _08135_, _08132_);
  or _59358_ (_08137_, _08136_, _08129_);
  and _59359_ (_08138_, _07544_, _06172_);
  nor _59360_ (_08139_, _08138_, _08137_);
  not _59361_ (_08140_, _08139_);
  and _59362_ (_08141_, _07778_, \oc8051_golden_model_1.SCON [1]);
  and _59363_ (_08142_, _07783_, \oc8051_golden_model_1.SBUF [1]);
  or _59364_ (_08143_, _08142_, _08141_);
  and _59365_ (_08144_, _07788_, \oc8051_golden_model_1.TCON [1]);
  and _59366_ (_08145_, _07794_, \oc8051_golden_model_1.PSW [1]);
  or _59367_ (_08146_, _08145_, _08144_);
  or _59368_ (_08147_, _08146_, _08143_);
  and _59369_ (_08148_, _07841_, \oc8051_golden_model_1.B [1]);
  and _59370_ (_08149_, _07809_, \oc8051_golden_model_1.ACC [1]);
  or _59371_ (_08150_, _08149_, _08148_);
  and _59372_ (_08151_, _07823_, \oc8051_golden_model_1.TH0 [1]);
  and _59373_ (_08152_, _07837_, \oc8051_golden_model_1.TL1 [1]);
  or _59374_ (_08153_, _08152_, _08151_);
  or _59375_ (_08154_, _08153_, _08150_);
  and _59376_ (_08155_, _07817_, \oc8051_golden_model_1.TH1 [1]);
  and _59377_ (_08156_, _07826_, \oc8051_golden_model_1.IE [1]);
  and _59378_ (_08157_, _07830_, \oc8051_golden_model_1.IP [1]);
  or _59379_ (_08158_, _08157_, _08156_);
  or _59380_ (_08159_, _08158_, _08155_);
  and _59381_ (_08160_, _07812_, \oc8051_golden_model_1.TMOD [1]);
  and _59382_ (_08161_, _07803_, \oc8051_golden_model_1.TL0 [1]);
  or _59383_ (_08162_, _08161_, _08160_);
  or _59384_ (_08163_, _08162_, _08159_);
  or _59385_ (_08164_, _08163_, _08154_);
  or _59386_ (_08165_, _08164_, _08147_);
  and _59387_ (_08166_, _07858_, \oc8051_golden_model_1.SP [1]);
  and _59388_ (_08167_, _07852_, \oc8051_golden_model_1.DPH [1]);
  or _59389_ (_08168_, _08167_, _08166_);
  and _59390_ (_08169_, _07849_, \oc8051_golden_model_1.DPL [1]);
  and _59391_ (_08170_, _07856_, \oc8051_golden_model_1.PCON [1]);
  or _59392_ (_08171_, _08170_, _08169_);
  or _59393_ (_08172_, _08171_, _08168_);
  or _59394_ (_08173_, _08172_, _08165_);
  and _59395_ (_08174_, _07306_, _06172_);
  nor _59396_ (_08175_, _08174_, _08173_);
  not _59397_ (_08176_, _08175_);
  and _59398_ (_08177_, _07788_, \oc8051_golden_model_1.TCON [0]);
  and _59399_ (_08178_, _07778_, \oc8051_golden_model_1.SCON [0]);
  or _59400_ (_08179_, _08178_, _08177_);
  and _59401_ (_08180_, _07783_, \oc8051_golden_model_1.SBUF [0]);
  and _59402_ (_08181_, _07809_, \oc8051_golden_model_1.ACC [0]);
  or _59403_ (_08182_, _08181_, _08180_);
  or _59404_ (_08183_, _08182_, _08179_);
  and _59405_ (_08184_, _07812_, \oc8051_golden_model_1.TMOD [0]);
  and _59406_ (_08185_, _07803_, \oc8051_golden_model_1.TL0 [0]);
  or _59407_ (_08186_, _08185_, _08184_);
  and _59408_ (_08187_, _07823_, \oc8051_golden_model_1.TH0 [0]);
  and _59409_ (_08188_, _07837_, \oc8051_golden_model_1.TL1 [0]);
  or _59410_ (_08189_, _08188_, _08187_);
  or _59411_ (_08190_, _08189_, _08186_);
  and _59412_ (_08191_, _07794_, \oc8051_golden_model_1.PSW [0]);
  and _59413_ (_08192_, _07826_, \oc8051_golden_model_1.IE [0]);
  and _59414_ (_08193_, _07830_, \oc8051_golden_model_1.IP [0]);
  or _59415_ (_08194_, _08193_, _08192_);
  or _59416_ (_08195_, _08194_, _08191_);
  and _59417_ (_08196_, _07817_, \oc8051_golden_model_1.TH1 [0]);
  and _59418_ (_08197_, _07841_, \oc8051_golden_model_1.B [0]);
  or _59419_ (_08198_, _08197_, _08196_);
  or _59420_ (_08199_, _08198_, _08195_);
  or _59421_ (_08200_, _08199_, _08190_);
  or _59422_ (_08201_, _08200_, _08183_);
  and _59423_ (_08202_, _07849_, \oc8051_golden_model_1.DPL [0]);
  and _59424_ (_08203_, _07852_, \oc8051_golden_model_1.DPH [0]);
  or _59425_ (_08204_, _08203_, _08202_);
  and _59426_ (_08205_, _07856_, \oc8051_golden_model_1.PCON [0]);
  and _59427_ (_08206_, _07858_, \oc8051_golden_model_1.SP [0]);
  or _59428_ (_08207_, _08206_, _08205_);
  or _59429_ (_08208_, _08207_, _08204_);
  or _59430_ (_08209_, _08208_, _08201_);
  and _59431_ (_08210_, _07049_, _06172_);
  or _59432_ (_08211_, _08210_, _08209_);
  and _59433_ (_08212_, _08211_, _08176_);
  and _59434_ (_08213_, _07837_, \oc8051_golden_model_1.TL1 [2]);
  and _59435_ (_08214_, _07817_, \oc8051_golden_model_1.TH1 [2]);
  or _59436_ (_08215_, _08214_, _08213_);
  and _59437_ (_08216_, _07788_, \oc8051_golden_model_1.TCON [2]);
  and _59438_ (_08217_, _07812_, \oc8051_golden_model_1.TMOD [2]);
  or _59439_ (_08218_, _08217_, _08216_);
  or _59440_ (_08219_, _08218_, _08215_);
  and _59441_ (_08220_, _07803_, \oc8051_golden_model_1.TL0 [2]);
  and _59442_ (_08221_, _07809_, \oc8051_golden_model_1.ACC [2]);
  or _59443_ (_08222_, _08221_, _08220_);
  and _59444_ (_08223_, _07823_, \oc8051_golden_model_1.TH0 [2]);
  and _59445_ (_08224_, _07841_, \oc8051_golden_model_1.B [2]);
  or _59446_ (_08225_, _08224_, _08223_);
  or _59447_ (_08226_, _08225_, _08222_);
  and _59448_ (_08227_, _07783_, \oc8051_golden_model_1.SBUF [2]);
  and _59449_ (_08228_, _07826_, \oc8051_golden_model_1.IE [2]);
  and _59450_ (_08229_, _07830_, \oc8051_golden_model_1.IP [2]);
  or _59451_ (_08230_, _08229_, _08228_);
  or _59452_ (_08231_, _08230_, _08227_);
  and _59453_ (_08232_, _07778_, \oc8051_golden_model_1.SCON [2]);
  and _59454_ (_08233_, _07794_, \oc8051_golden_model_1.PSW [2]);
  or _59455_ (_08234_, _08233_, _08232_);
  or _59456_ (_08235_, _08234_, _08231_);
  or _59457_ (_08236_, _08235_, _08226_);
  or _59458_ (_08237_, _08236_, _08219_);
  and _59459_ (_08238_, _07849_, \oc8051_golden_model_1.DPL [2]);
  and _59460_ (_08239_, _07852_, \oc8051_golden_model_1.DPH [2]);
  or _59461_ (_08240_, _08239_, _08238_);
  and _59462_ (_08241_, _07856_, \oc8051_golden_model_1.PCON [2]);
  and _59463_ (_08242_, _07858_, \oc8051_golden_model_1.SP [2]);
  or _59464_ (_08243_, _08242_, _08241_);
  or _59465_ (_08244_, _08243_, _08240_);
  or _59466_ (_08245_, _08244_, _08237_);
  and _59467_ (_08246_, _07708_, _06172_);
  nor _59468_ (_08247_, _08246_, _08245_);
  not _59469_ (_08248_, _08247_);
  and _59470_ (_08249_, _08248_, _08212_);
  and _59471_ (_08250_, _08249_, _08140_);
  and _59472_ (_08251_, _07788_, \oc8051_golden_model_1.TCON [4]);
  and _59473_ (_08252_, _07778_, \oc8051_golden_model_1.SCON [4]);
  or _59474_ (_08253_, _08252_, _08251_);
  and _59475_ (_08254_, _07794_, \oc8051_golden_model_1.PSW [4]);
  and _59476_ (_08255_, _07809_, \oc8051_golden_model_1.ACC [4]);
  or _59477_ (_08256_, _08255_, _08254_);
  or _59478_ (_08257_, _08256_, _08253_);
  and _59479_ (_08258_, _07812_, \oc8051_golden_model_1.TMOD [4]);
  and _59480_ (_08259_, _07803_, \oc8051_golden_model_1.TL0 [4]);
  or _59481_ (_08260_, _08259_, _08258_);
  and _59482_ (_08261_, _07823_, \oc8051_golden_model_1.TH0 [4]);
  and _59483_ (_08262_, _07837_, \oc8051_golden_model_1.TL1 [4]);
  or _59484_ (_08263_, _08262_, _08261_);
  or _59485_ (_08264_, _08263_, _08260_);
  and _59486_ (_08265_, _07783_, \oc8051_golden_model_1.SBUF [4]);
  and _59487_ (_08266_, _07826_, \oc8051_golden_model_1.IE [4]);
  and _59488_ (_08267_, _07830_, \oc8051_golden_model_1.IP [4]);
  or _59489_ (_08268_, _08267_, _08266_);
  or _59490_ (_08269_, _08268_, _08265_);
  and _59491_ (_08270_, _07817_, \oc8051_golden_model_1.TH1 [4]);
  and _59492_ (_08271_, _07841_, \oc8051_golden_model_1.B [4]);
  or _59493_ (_08272_, _08271_, _08270_);
  or _59494_ (_08273_, _08272_, _08269_);
  or _59495_ (_08274_, _08273_, _08264_);
  or _59496_ (_08275_, _08274_, _08257_);
  and _59497_ (_08276_, _07849_, \oc8051_golden_model_1.DPL [4]);
  and _59498_ (_08277_, _07852_, \oc8051_golden_model_1.DPH [4]);
  or _59499_ (_08278_, _08277_, _08276_);
  and _59500_ (_08279_, _07856_, \oc8051_golden_model_1.PCON [4]);
  and _59501_ (_08280_, _07858_, \oc8051_golden_model_1.SP [4]);
  or _59502_ (_08281_, _08280_, _08279_);
  or _59503_ (_08282_, _08281_, _08278_);
  or _59504_ (_08283_, _08282_, _08275_);
  not _59505_ (_08284_, \oc8051_golden_model_1.IRAM[0] [4]);
  or _59506_ (_08285_, _06844_, _08284_);
  not _59507_ (_08286_, \oc8051_golden_model_1.IRAM[1] [4]);
  or _59508_ (_08287_, _06993_, _08286_);
  and _59509_ (_08288_, _08287_, _06991_);
  nand _59510_ (_08289_, _08288_, _08285_);
  not _59511_ (_08290_, \oc8051_golden_model_1.IRAM[3] [4]);
  or _59512_ (_08291_, _06993_, _08290_);
  not _59513_ (_08292_, \oc8051_golden_model_1.IRAM[2] [4]);
  or _59514_ (_08293_, _06844_, _08292_);
  and _59515_ (_08294_, _08293_, _06999_);
  nand _59516_ (_08295_, _08294_, _08291_);
  nand _59517_ (_08296_, _08295_, _08289_);
  nand _59518_ (_08297_, _08296_, _06637_);
  not _59519_ (_08298_, \oc8051_golden_model_1.IRAM[7] [4]);
  or _59520_ (_08299_, _06993_, _08298_);
  not _59521_ (_08300_, \oc8051_golden_model_1.IRAM[6] [4]);
  or _59522_ (_08301_, _06844_, _08300_);
  and _59523_ (_08302_, _08301_, _06999_);
  nand _59524_ (_08303_, _08302_, _08299_);
  not _59525_ (_08304_, \oc8051_golden_model_1.IRAM[4] [4]);
  or _59526_ (_08305_, _06844_, _08304_);
  not _59527_ (_08306_, \oc8051_golden_model_1.IRAM[5] [4]);
  or _59528_ (_08307_, _06993_, _08306_);
  and _59529_ (_08308_, _08307_, _06991_);
  nand _59530_ (_08309_, _08308_, _08305_);
  nand _59531_ (_08310_, _08309_, _08303_);
  nand _59532_ (_08311_, _08310_, _07006_);
  nand _59533_ (_08312_, _08311_, _08297_);
  nand _59534_ (_08313_, _08312_, _06446_);
  nand _59535_ (_08314_, _06844_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _59536_ (_08315_, _06993_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _59537_ (_08316_, _08315_, _06999_);
  nand _59538_ (_08317_, _08316_, _08314_);
  nand _59539_ (_08318_, _06993_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand _59540_ (_08319_, _06844_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _59541_ (_08320_, _08319_, _06991_);
  nand _59542_ (_08321_, _08320_, _08318_);
  nand _59543_ (_08322_, _08321_, _08317_);
  nand _59544_ (_08323_, _08322_, _06637_);
  nand _59545_ (_08324_, _06844_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _59546_ (_08325_, _06993_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _59547_ (_08326_, _08325_, _06999_);
  nand _59548_ (_08327_, _08326_, _08324_);
  nand _59549_ (_08328_, _06993_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand _59550_ (_08329_, _06844_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _59551_ (_08330_, _08329_, _06991_);
  nand _59552_ (_08331_, _08330_, _08328_);
  nand _59553_ (_08332_, _08331_, _08327_);
  nand _59554_ (_08333_, _08332_, _07006_);
  nand _59555_ (_08334_, _08333_, _08323_);
  nand _59556_ (_08335_, _08334_, _07023_);
  and _59557_ (_08336_, _08335_, _08313_);
  and _59558_ (_08337_, _08336_, _06172_);
  nor _59559_ (_08338_, _08337_, _08283_);
  not _59560_ (_08339_, _08338_);
  and _59561_ (_08340_, _08339_, _08250_);
  and _59562_ (_08341_, _08340_, _08104_);
  and _59563_ (_08342_, _08341_, _08015_);
  nor _59564_ (_08343_, _08342_, _07926_);
  and _59565_ (_08344_, _08342_, _07926_);
  nor _59566_ (_08345_, _08344_, _08343_);
  and _59567_ (_08346_, _08345_, _07167_);
  nand _59568_ (_08347_, _08011_, _07989_);
  nand _59569_ (_08348_, _08100_, _08078_);
  nand _59570_ (_08349_, _08335_, _08313_);
  and _59571_ (_08350_, _08349_, _08348_);
  and _59572_ (_08351_, _07657_, _07474_);
  nor _59573_ (_08352_, _07306_, _07049_);
  and _59574_ (_08353_, _08352_, _08351_);
  and _59575_ (_08354_, _08353_, _08350_);
  and _59576_ (_08355_, _08354_, _08347_);
  or _59577_ (_08356_, _08355_, _07923_);
  nand _59578_ (_08357_, _08355_, _07923_);
  and _59579_ (_08358_, _08357_, _08356_);
  and _59580_ (_08359_, _06125_, _05591_);
  not _59581_ (_08360_, _08359_);
  and _59582_ (_08361_, _08360_, _07353_);
  and _59583_ (_08362_, _08361_, _07326_);
  or _59584_ (_08363_, _08362_, _08358_);
  not _59585_ (_08364_, _07131_);
  and _59586_ (_08365_, _06366_, _04273_);
  and _59587_ (_08366_, _06368_, _04246_);
  nor _59588_ (_08367_, _08366_, _08365_);
  and _59589_ (_08368_, _06377_, _04270_);
  and _59590_ (_08369_, _06382_, _04292_);
  nor _59591_ (_08370_, _08369_, _08368_);
  and _59592_ (_08371_, _08370_, _08367_);
  and _59593_ (_08372_, _06355_, _04256_);
  and _59594_ (_08373_, _06340_, _04253_);
  nor _59595_ (_08374_, _08373_, _08372_);
  and _59596_ (_08375_, _06384_, _04295_);
  and _59597_ (_08376_, _06361_, _04278_);
  nor _59598_ (_08377_, _08376_, _08375_);
  and _59599_ (_08378_, _08377_, _08374_);
  and _59600_ (_08379_, _08378_, _08371_);
  and _59601_ (_08380_, _06373_, _04242_);
  and _59602_ (_08381_, _06379_, _04281_);
  nor _59603_ (_08382_, _08381_, _08380_);
  and _59604_ (_08383_, _06336_, _00567_);
  and _59605_ (_08384_, _06371_, _04260_);
  nor _59606_ (_08385_, _08384_, _08383_);
  and _59607_ (_08386_, _08385_, _08382_);
  and _59608_ (_08387_, _06359_, _04264_);
  and _59609_ (_08388_, _06348_, _04287_);
  nor _59610_ (_08389_, _08388_, _08387_);
  and _59611_ (_08390_, _06345_, _04210_);
  and _59612_ (_08391_, _06352_, _04237_);
  nor _59613_ (_08392_, _08391_, _08390_);
  and _59614_ (_08393_, _08392_, _08389_);
  and _59615_ (_08394_, _08393_, _08386_);
  and _59616_ (_08395_, _08394_, _08379_);
  nor _59617_ (_08396_, _08395_, _07925_);
  and _59618_ (_08397_, _08396_, _07133_);
  not _59619_ (_08398_, _07086_);
  not _59620_ (_08399_, _07855_);
  not _59621_ (_08400_, _06071_);
  nor _59622_ (_08401_, _06877_, _08400_);
  and _59623_ (_08402_, _08401_, _06479_);
  and _59624_ (_08403_, _08402_, _06206_);
  and _59625_ (_08404_, _08403_, _07792_);
  nand _59626_ (_08405_, _08404_, \oc8051_golden_model_1.PSW [7]);
  and _59627_ (_08406_, _08402_, _06207_);
  and _59628_ (_08407_, _08406_, _07787_);
  nand _59629_ (_08408_, _08407_, \oc8051_golden_model_1.TCON [7]);
  and _59630_ (_08409_, _08403_, _07807_);
  nand _59631_ (_08410_, _08409_, \oc8051_golden_model_1.ACC [7]);
  and _59632_ (_08411_, _08410_, _08408_);
  nand _59633_ (_08412_, _08411_, _08405_);
  and _59634_ (_08413_, _08406_, _07777_);
  nand _59635_ (_08414_, _08413_, \oc8051_golden_model_1.SCON [7]);
  and _59636_ (_08415_, _08406_, _07829_);
  nand _59637_ (_08416_, _08415_, \oc8051_golden_model_1.IP [7]);
  nand _59638_ (_08417_, _08416_, _08414_);
  and _59639_ (_08418_, _08406_, _07825_);
  nand _59640_ (_08419_, _08418_, \oc8051_golden_model_1.IE [7]);
  and _59641_ (_08420_, _08403_, _07839_);
  nand _59642_ (_08421_, _08420_, \oc8051_golden_model_1.B [7]);
  nand _59643_ (_08422_, _08421_, _08419_);
  or _59644_ (_08423_, _08422_, _08417_);
  or _59645_ (_08424_, _08423_, _08412_);
  or _59646_ (_08425_, _08424_, _07924_);
  and _59647_ (_08426_, _08425_, _08399_);
  or _59648_ (_08427_, _08426_, _08398_);
  not _59649_ (_08428_, _06159_);
  not _59650_ (_08429_, _06162_);
  not _59651_ (_08430_, \oc8051_golden_model_1.ACC [7]);
  nor _59652_ (_08431_, _06581_, _08430_);
  and _59653_ (_08432_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and _59654_ (_08433_, _08432_, \oc8051_golden_model_1.PC [6]);
  and _59655_ (_08434_, _08433_, _05972_);
  and _59656_ (_08435_, _08434_, \oc8051_golden_model_1.PC [7]);
  nor _59657_ (_08436_, _08434_, \oc8051_golden_model_1.PC [7]);
  nor _59658_ (_08437_, _08436_, _08435_);
  and _59659_ (_08438_, _08437_, _06581_);
  or _59660_ (_08439_, _08438_, _08431_);
  not _59661_ (_08440_, _06129_);
  nor _59662_ (_08441_, _08440_, _06125_);
  nor _59663_ (_08442_, _08441_, _05762_);
  nor _59664_ (_08443_, _08442_, _07259_);
  and _59665_ (_08444_, _08443_, _08439_);
  not _59666_ (_08445_, _08443_);
  and _59667_ (_08446_, _08445_, _08358_);
  or _59668_ (_08447_, _08446_, _08444_);
  and _59669_ (_08448_, _08447_, _07065_);
  nor _59670_ (_08449_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _59671_ (_08450_, _08449_, _06566_);
  nor _59672_ (_08451_, _08450_, _06216_);
  nor _59673_ (_08452_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _59674_ (_08453_, _08452_, _06216_);
  and _59675_ (_08454_, _08453_, _06142_);
  nor _59676_ (_08455_, _08454_, _08451_);
  nor _59677_ (_08456_, _08455_, _06980_);
  not _59678_ (_08457_, _08456_);
  or _59679_ (_08458_, _07544_, _06701_);
  not _59680_ (_08459_, _06980_);
  and _59681_ (_08460_, _06701_, _06070_);
  nor _59682_ (_08461_, _08460_, _08459_);
  nand _59683_ (_08462_, _08461_, _08458_);
  and _59684_ (_08463_, _08462_, _08457_);
  nor _59685_ (_08464_, _08449_, _06566_);
  nor _59686_ (_08465_, _08464_, _08450_);
  nor _59687_ (_08466_, _08465_, _06980_);
  not _59688_ (_08467_, _08466_);
  or _59689_ (_08468_, _07708_, _06701_);
  and _59690_ (_08469_, _06701_, _06625_);
  nor _59691_ (_08470_, _08469_, _08459_);
  nand _59692_ (_08471_, _08470_, _08468_);
  and _59693_ (_08472_, _08471_, _08467_);
  or _59694_ (_08473_, _07049_, _06701_);
  and _59695_ (_08474_, _06701_, _06107_);
  nor _59696_ (_08475_, _08474_, _08459_);
  nand _59697_ (_08476_, _08475_, _08473_);
  nor _59698_ (_08477_, _06980_, \oc8051_golden_model_1.SP [0]);
  not _59699_ (_08478_, _08477_);
  nand _59700_ (_08479_, _08478_, _08476_);
  or _59701_ (_08480_, _08479_, _07863_);
  nor _59702_ (_08481_, _07179_, _06980_);
  not _59703_ (_08482_, _08481_);
  and _59704_ (_08483_, _07306_, _07104_);
  nor _59705_ (_08484_, _06912_, _07104_);
  or _59706_ (_08485_, _08484_, _08459_);
  or _59707_ (_08486_, _08485_, _08483_);
  nand _59708_ (_08487_, _08486_, _08482_);
  and _59709_ (_08488_, _08478_, _08476_);
  or _59710_ (_08489_, _08488_, _07865_);
  and _59711_ (_08490_, _08489_, _08487_);
  nand _59712_ (_08491_, _08490_, _08480_);
  or _59713_ (_08492_, _08479_, _07871_);
  and _59714_ (_08493_, _08486_, _08482_);
  or _59715_ (_08494_, _08488_, _07869_);
  and _59716_ (_08495_, _08494_, _08493_);
  nand _59717_ (_08496_, _08495_, _08492_);
  nand _59718_ (_08497_, _08496_, _08491_);
  nand _59719_ (_08498_, _08497_, _08472_);
  not _59720_ (_08499_, _08472_);
  or _59721_ (_08500_, _08479_, _07883_);
  or _59722_ (_08501_, _08488_, _07885_);
  and _59723_ (_08502_, _08501_, _08487_);
  nand _59724_ (_08503_, _08502_, _08500_);
  or _59725_ (_08504_, _08479_, _07879_);
  or _59726_ (_08505_, _08488_, _07877_);
  and _59727_ (_08506_, _08505_, _08493_);
  nand _59728_ (_08507_, _08506_, _08504_);
  nand _59729_ (_08508_, _08507_, _08503_);
  nand _59730_ (_08509_, _08508_, _08499_);
  nand _59731_ (_08510_, _08509_, _08498_);
  nand _59732_ (_08511_, _08510_, _08463_);
  not _59733_ (_08512_, _08463_);
  or _59734_ (_08513_, _08479_, _07895_);
  or _59735_ (_08514_, _08488_, _07893_);
  and _59736_ (_08515_, _08514_, _08493_);
  nand _59737_ (_08516_, _08515_, _08513_);
  or _59738_ (_08517_, _08479_, _07899_);
  or _59739_ (_08518_, _08488_, _07901_);
  and _59740_ (_08519_, _08518_, _08487_);
  nand _59741_ (_08520_, _08519_, _08517_);
  nand _59742_ (_08521_, _08520_, _08516_);
  nand _59743_ (_08522_, _08521_, _08472_);
  or _59744_ (_08523_, _08479_, _07913_);
  or _59745_ (_08524_, _08488_, _07915_);
  and _59746_ (_08525_, _08524_, _08487_);
  nand _59747_ (_08526_, _08525_, _08523_);
  or _59748_ (_08527_, _08479_, _07909_);
  or _59749_ (_08528_, _08488_, _07907_);
  and _59750_ (_08529_, _08528_, _08493_);
  nand _59751_ (_08530_, _08529_, _08527_);
  nand _59752_ (_08531_, _08530_, _08526_);
  nand _59753_ (_08532_, _08531_, _08499_);
  nand _59754_ (_08533_, _08532_, _08522_);
  nand _59755_ (_08534_, _08533_, _08512_);
  and _59756_ (_08535_, _08534_, _08511_);
  and _59757_ (_08536_, _08535_, _07064_);
  or _59758_ (_08537_, _08536_, _08448_);
  and _59759_ (_08538_, _08537_, _08429_);
  and _59760_ (_08539_, _08338_, _08103_);
  not _59761_ (_08540_, _08211_);
  and _59762_ (_08541_, _08540_, _08175_);
  and _59763_ (_08542_, _08247_, _08139_);
  and _59764_ (_08543_, _08542_, _08541_);
  and _59765_ (_08544_, _08543_, _08539_);
  and _59766_ (_08545_, _08544_, _08014_);
  or _59767_ (_08546_, _08545_, _07926_);
  nand _59768_ (_08547_, _08545_, _07926_);
  and _59769_ (_08548_, _08547_, _08546_);
  and _59770_ (_08549_, _08548_, _06162_);
  or _59771_ (_08550_, _08549_, _08538_);
  and _59772_ (_08551_, _08550_, _08428_);
  or _59773_ (_08552_, _08425_, _07855_);
  and _59774_ (_08553_, _08552_, _06159_);
  or _59775_ (_08554_, _08553_, _07485_);
  or _59776_ (_08555_, _08554_, _08551_);
  nor _59777_ (_08556_, _08437_, _05764_);
  nor _59778_ (_08557_, _08556_, _07076_);
  and _59779_ (_08558_, _08557_, _08555_);
  and _59780_ (_08559_, _07923_, _07076_);
  or _59781_ (_08560_, _08559_, _07086_);
  or _59782_ (_08561_, _08560_, _08558_);
  and _59783_ (_08562_, _08561_, _08427_);
  or _59784_ (_08563_, _08562_, _06151_);
  nand _59785_ (_08564_, _07925_, _06151_);
  and _59786_ (_08565_, _08564_, _06149_);
  and _59787_ (_08566_, _08565_, _08563_);
  and _59788_ (_08567_, _08425_, _07855_);
  not _59789_ (_08568_, _08567_);
  and _59790_ (_08569_, _08568_, _08552_);
  and _59791_ (_08570_, _08569_, _06148_);
  or _59792_ (_08571_, _08570_, _08566_);
  and _59793_ (_08572_, _08571_, _05760_);
  not _59794_ (_08573_, _08437_);
  or _59795_ (_08574_, _08573_, _05760_);
  nand _59796_ (_08575_, _08574_, _06251_);
  or _59797_ (_08576_, _08575_, _08572_);
  nand _59798_ (_08577_, _07925_, _06252_);
  and _59799_ (_08578_, _08577_, _08576_);
  or _59800_ (_08579_, _08578_, _06701_);
  not _59801_ (_08580_, _07103_);
  and _59802_ (_08581_, _08535_, _06172_);
  or _59803_ (_08582_, _07862_, _07104_);
  or _59804_ (_08583_, _08582_, _08581_);
  and _59805_ (_08584_, _08583_, _08580_);
  and _59806_ (_08585_, _08584_, _08579_);
  and _59807_ (_08586_, _07855_, \oc8051_golden_model_1.PSW [7]);
  or _59808_ (_08587_, _08586_, _08426_);
  and _59809_ (_08588_, _08587_, _07103_);
  or _59810_ (_08589_, _08588_, _05791_);
  or _59811_ (_08590_, _08589_, _08585_);
  nor _59812_ (_08591_, _06132_, _06039_);
  and _59813_ (_08592_, _08573_, _05791_);
  nor _59814_ (_08593_, _08592_, _08591_);
  and _59815_ (_08594_, _08593_, _08590_);
  nor _59816_ (_08595_, _06117_, _06039_);
  and _59817_ (_08596_, _07923_, _08591_);
  or _59818_ (_08597_, _08596_, _08595_);
  or _59819_ (_08598_, _08597_, _08594_);
  nor _59820_ (_08599_, _06039_, _06114_);
  not _59821_ (_08600_, _08599_);
  not _59822_ (_08601_, _08595_);
  or _59823_ (_08602_, _08535_, _08601_);
  and _59824_ (_08603_, _08602_, _08600_);
  and _59825_ (_08604_, _08603_, _08598_);
  and _59826_ (_08605_, _08395_, _07923_);
  and _59827_ (_08606_, _06945_, _06758_);
  not _59828_ (_08607_, _08395_);
  and _59829_ (_08608_, _06359_, _04687_);
  and _59830_ (_08609_, _06368_, _04679_);
  nor _59831_ (_08610_, _08609_, _08608_);
  and _59832_ (_08611_, _06371_, _04671_);
  and _59833_ (_08612_, _06382_, _04668_);
  nor _59834_ (_08613_, _08612_, _08611_);
  and _59835_ (_08614_, _08613_, _08610_);
  and _59836_ (_08615_, _06384_, _04693_);
  and _59837_ (_08616_, _06366_, _04673_);
  nor _59838_ (_08617_, _08616_, _08615_);
  and _59839_ (_08618_, _06355_, _04695_);
  and _59840_ (_08619_, _06340_, _04699_);
  nor _59841_ (_08620_, _08619_, _08618_);
  and _59842_ (_08621_, _08620_, _08617_);
  and _59843_ (_08622_, _08621_, _08614_);
  and _59844_ (_08623_, _06345_, _04666_);
  and _59845_ (_08624_, _06373_, _04697_);
  nor _59846_ (_08625_, _08624_, _08623_);
  and _59847_ (_08626_, _06336_, _00612_);
  and _59848_ (_08627_, _06352_, _04682_);
  nor _59849_ (_08628_, _08627_, _08626_);
  and _59850_ (_08629_, _08628_, _08625_);
  and _59851_ (_08630_, _06361_, _04677_);
  and _59852_ (_08631_, _06348_, _04689_);
  nor _59853_ (_08632_, _08631_, _08630_);
  and _59854_ (_08633_, _06377_, _04705_);
  and _59855_ (_08634_, _06379_, _04684_);
  nor _59856_ (_08635_, _08634_, _08633_);
  and _59857_ (_08636_, _08635_, _08632_);
  and _59858_ (_08637_, _08636_, _08629_);
  and _59859_ (_08638_, _08637_, _08622_);
  and _59860_ (_08639_, _08638_, _08607_);
  and _59861_ (_08640_, _06359_, _04614_);
  and _59862_ (_08641_, _06368_, _04588_);
  nor _59863_ (_08642_, _08641_, _08640_);
  and _59864_ (_08643_, _06377_, _04596_);
  and _59865_ (_08644_, _06352_, _04591_);
  nor _59866_ (_08645_, _08644_, _08643_);
  and _59867_ (_08646_, _08645_, _08642_);
  and _59868_ (_08647_, _06355_, _04608_);
  and _59869_ (_08648_, _06340_, _04606_);
  nor _59870_ (_08649_, _08648_, _08647_);
  and _59871_ (_08650_, _06384_, _04602_);
  and _59872_ (_08651_, _06361_, _04586_);
  nor _59873_ (_08652_, _08651_, _08650_);
  and _59874_ (_08653_, _08652_, _08649_);
  and _59875_ (_08654_, _08653_, _08646_);
  and _59876_ (_08655_, _06382_, _04575_);
  and _59877_ (_08656_, _06345_, _04580_);
  nor _59878_ (_08657_, _08656_, _08655_);
  and _59879_ (_08658_, _06336_, _00602_);
  and _59880_ (_08659_, _06371_, _04582_);
  nor _59881_ (_08660_, _08659_, _08658_);
  and _59882_ (_08661_, _08660_, _08657_);
  and _59883_ (_08662_, _06366_, _04577_);
  and _59884_ (_08663_, _06348_, _04598_);
  nor _59885_ (_08664_, _08663_, _08662_);
  and _59886_ (_08665_, _06373_, _04604_);
  and _59887_ (_08666_, _06379_, _04593_);
  nor _59888_ (_08667_, _08666_, _08665_);
  and _59889_ (_08668_, _08667_, _08664_);
  and _59890_ (_08669_, _08668_, _08661_);
  and _59891_ (_08670_, _08669_, _08654_);
  and _59892_ (_08671_, _06359_, _04641_);
  and _59893_ (_08672_, _06340_, _04654_);
  nor _59894_ (_08673_, _08672_, _08671_);
  and _59895_ (_08674_, _06379_, _04638_);
  and _59896_ (_08675_, _06355_, _04650_);
  nor _59897_ (_08676_, _08675_, _08674_);
  and _59898_ (_08677_, _08676_, _08673_);
  and _59899_ (_08678_, _06345_, _04620_);
  and _59900_ (_08679_, _06348_, _04643_);
  nor _59901_ (_08680_, _08679_, _08678_);
  and _59902_ (_08681_, _06371_, _04625_);
  and _59903_ (_08682_, _06382_, _04622_);
  nor _59904_ (_08683_, _08682_, _08681_);
  and _59905_ (_08684_, _08683_, _08680_);
  and _59906_ (_08685_, _08684_, _08677_);
  and _59907_ (_08686_, _06377_, _04660_);
  and _59908_ (_08687_, _06368_, _04633_);
  nor _59909_ (_08688_, _08687_, _08686_);
  and _59910_ (_08689_, _06352_, _04636_);
  and _59911_ (_08690_, _06384_, _04648_);
  nor _59912_ (_08691_, _08690_, _08689_);
  and _59913_ (_08692_, _08691_, _08688_);
  and _59914_ (_08693_, _06373_, _04652_);
  and _59915_ (_08694_, _06361_, _04631_);
  nor _59916_ (_08695_, _08694_, _08693_);
  and _59917_ (_08696_, _06336_, _00607_);
  and _59918_ (_08697_, _06366_, _04627_);
  nor _59919_ (_08698_, _08697_, _08696_);
  and _59920_ (_08699_, _08698_, _08695_);
  and _59921_ (_08700_, _08699_, _08692_);
  and _59922_ (_08701_, _08700_, _08685_);
  and _59923_ (_08702_, _08701_, _08670_);
  and _59924_ (_08703_, _08702_, _08639_);
  nor _59925_ (_08704_, _06521_, _06389_);
  and _59926_ (_08705_, _08704_, _08703_);
  and _59927_ (_08706_, _08705_, _08606_);
  and _59928_ (_08707_, _08706_, \oc8051_golden_model_1.TH0 [7]);
  not _59929_ (_08708_, _06758_);
  and _59930_ (_08709_, _06945_, _08708_);
  and _59931_ (_08710_, _08709_, _08705_);
  and _59932_ (_08711_, _08710_, \oc8051_golden_model_1.TH1 [7]);
  not _59933_ (_08712_, _06389_);
  and _59934_ (_08713_, _06521_, _08712_);
  and _59935_ (_08714_, _08713_, _08606_);
  not _59936_ (_08715_, _08670_);
  and _59937_ (_08716_, _08701_, _08715_);
  and _59938_ (_08717_, _08716_, _08639_);
  and _59939_ (_08718_, _08717_, _08714_);
  and _59940_ (_08719_, _08718_, \oc8051_golden_model_1.SCON [7]);
  or _59941_ (_08720_, _08719_, _08711_);
  or _59942_ (_08721_, _08720_, _08707_);
  nor _59943_ (_08722_, _06945_, _06758_);
  and _59944_ (_08723_, _08722_, _08703_);
  and _59945_ (_08724_, _08723_, _08713_);
  and _59946_ (_08725_, _08724_, \oc8051_golden_model_1.TL1 [7]);
  and _59947_ (_08726_, _08714_, _08703_);
  and _59948_ (_08727_, _08726_, \oc8051_golden_model_1.TCON [7]);
  or _59949_ (_08728_, _08727_, _08725_);
  or _59950_ (_08729_, _08728_, _08721_);
  and _59951_ (_08730_, _06521_, _06389_);
  and _59952_ (_08731_, _08730_, _08606_);
  nor _59953_ (_08732_, _08638_, _08395_);
  and _59954_ (_08733_, _08732_, _08731_);
  and _59955_ (_08734_, _08716_, _08733_);
  and _59956_ (_08735_, _08734_, \oc8051_golden_model_1.PSW [7]);
  not _59957_ (_08736_, _08701_);
  and _59958_ (_08737_, _08736_, _08670_);
  and _59959_ (_08738_, _08733_, _08737_);
  and _59960_ (_08739_, _08738_, \oc8051_golden_model_1.ACC [7]);
  nor _59961_ (_08740_, _08701_, _08670_);
  and _59962_ (_08741_, _08733_, _08740_);
  and _59963_ (_08742_, _08741_, \oc8051_golden_model_1.B [7]);
  or _59964_ (_08743_, _08742_, _08739_);
  or _59965_ (_08744_, _08743_, _08735_);
  and _59966_ (_08745_, _08740_, _08639_);
  and _59967_ (_08746_, _08745_, _08714_);
  and _59968_ (_08747_, _08746_, \oc8051_golden_model_1.IP [7]);
  and _59969_ (_08748_, _08737_, _08639_);
  and _59970_ (_08749_, _08748_, _08714_);
  and _59971_ (_08750_, _08749_, \oc8051_golden_model_1.IE [7]);
  and _59972_ (_08751_, _08713_, _08709_);
  and _59973_ (_08752_, _08751_, _08717_);
  and _59974_ (_08753_, _08752_, \oc8051_golden_model_1.SBUF [7]);
  or _59975_ (_08754_, _08753_, _08750_);
  or _59976_ (_08755_, _08754_, _08747_);
  or _59977_ (_08756_, _08755_, _08744_);
  and _59978_ (_08757_, _08730_, _08703_);
  and _59979_ (_08758_, _08757_, _08709_);
  and _59980_ (_08759_, _08758_, \oc8051_golden_model_1.SP [7]);
  and _59981_ (_08760_, _08730_, _08723_);
  and _59982_ (_08761_, _08760_, \oc8051_golden_model_1.DPH [7]);
  or _59983_ (_08762_, _08761_, _08759_);
  not _59984_ (_08763_, _06945_);
  and _59985_ (_08764_, _08763_, _06758_);
  and _59986_ (_08765_, _08757_, _08764_);
  and _59987_ (_08766_, _08765_, \oc8051_golden_model_1.DPL [7]);
  or _59988_ (_08767_, _08766_, _08762_);
  not _59989_ (_08768_, _06521_);
  and _59990_ (_08769_, _08768_, _06389_);
  and _59991_ (_08770_, _08769_, _08723_);
  and _59992_ (_08771_, _08770_, \oc8051_golden_model_1.PCON [7]);
  and _59993_ (_08772_, _08713_, _08703_);
  and _59994_ (_08773_, _08772_, _08764_);
  and _59995_ (_08774_, _08773_, \oc8051_golden_model_1.TL0 [7]);
  and _59996_ (_08775_, _08751_, _08703_);
  and _59997_ (_08776_, _08775_, \oc8051_golden_model_1.TMOD [7]);
  or _59998_ (_08777_, _08776_, _08774_);
  or _59999_ (_08778_, _08777_, _08771_);
  or _60000_ (_08779_, _08778_, _08767_);
  or _60001_ (_08780_, _08779_, _08756_);
  or _60002_ (_08781_, _08780_, _08729_);
  or _60003_ (_08782_, _08781_, _08605_);
  and _60004_ (_08783_, _08782_, _08599_);
  not _60005_ (_08784_, _07184_);
  nor _60006_ (_08785_, _07115_, _07370_);
  and _60007_ (_08786_, _08785_, _08784_);
  and _60008_ (_08787_, _08786_, _07352_);
  not _60009_ (_08788_, _08787_);
  or _60010_ (_08789_, _08788_, _08783_);
  or _60011_ (_08790_, _08789_, _08604_);
  nor _60012_ (_08791_, _08787_, _06039_);
  nor _60013_ (_08792_, _08791_, _06112_);
  and _60014_ (_08793_, _08792_, _08790_);
  and _60015_ (_08794_, _08607_, _06112_);
  or _60016_ (_08795_, _08794_, _06076_);
  or _60017_ (_08796_, _08795_, _08793_);
  nor _60018_ (_08797_, _08437_, _05836_);
  nor _60019_ (_08798_, _08797_, _07128_);
  and _60020_ (_08799_, _08798_, _08796_);
  not _60021_ (_08800_, _08396_);
  nand _60022_ (_08801_, _08395_, _07925_);
  and _60023_ (_08802_, _08801_, _08800_);
  nor _60024_ (_08803_, _08802_, _07126_);
  nor _60025_ (_08804_, _08803_, _07129_);
  or _60026_ (_08805_, _08804_, _08799_);
  not _60027_ (_08806_, _07133_);
  not _60028_ (_08807_, _07126_);
  nor _60029_ (_08808_, _07925_, _08430_);
  and _60030_ (_08809_, _07925_, _08430_);
  nor _60031_ (_08810_, _08809_, _08808_);
  or _60032_ (_08811_, _08810_, _08807_);
  and _60033_ (_08812_, _08811_, _08806_);
  and _60034_ (_08813_, _08812_, _08805_);
  or _60035_ (_08814_, _08813_, _08397_);
  and _60036_ (_08815_, _08814_, _08364_);
  and _60037_ (_08816_, _08808_, _07131_);
  or _60038_ (_08817_, _08816_, _07124_);
  or _60039_ (_08818_, _08817_, _08815_);
  not _60040_ (_08819_, _06303_);
  nor _60041_ (_08820_, _08819_, _06039_);
  nor _60042_ (_08821_, _08437_, _05848_);
  nor _60043_ (_08822_, _08821_, _08820_);
  and _60044_ (_08823_, _08822_, _08818_);
  not _60045_ (_08824_, _06396_);
  nor _60046_ (_08825_, _08824_, _06039_);
  and _60047_ (_08826_, _08801_, _08820_);
  or _60048_ (_08827_, _08826_, _08825_);
  or _60049_ (_08828_, _08827_, _08823_);
  nand _60050_ (_08829_, _08809_, _08825_);
  and _60051_ (_08830_, _08829_, _05846_);
  and _60052_ (_08831_, _08830_, _08828_);
  or _60053_ (_08832_, _08573_, _05846_);
  nand _60054_ (_08833_, _08832_, _08362_);
  or _60055_ (_08834_, _08833_, _08831_);
  and _60056_ (_08835_, _08834_, _08363_);
  or _60057_ (_08836_, _08835_, _07153_);
  not _60058_ (_08837_, _07152_);
  nand _60059_ (_08838_, _08534_, _08511_);
  or _60060_ (_08839_, _08479_, _07960_);
  or _60061_ (_08840_, _08488_, _07962_);
  and _60062_ (_08841_, _08840_, _08487_);
  nand _60063_ (_08842_, _08841_, _08839_);
  or _60064_ (_08843_, _08479_, _07968_);
  or _60065_ (_08844_, _08488_, _07966_);
  and _60066_ (_08845_, _08844_, _08493_);
  nand _60067_ (_08846_, _08845_, _08843_);
  nand _60068_ (_08847_, _08846_, _08842_);
  nand _60069_ (_08848_, _08847_, _08472_);
  or _60070_ (_08849_, _08479_, _07980_);
  or _60071_ (_08850_, _08488_, _07982_);
  and _60072_ (_08851_, _08850_, _08487_);
  nand _60073_ (_08852_, _08851_, _08849_);
  or _60074_ (_08853_, _08479_, _07976_);
  or _60075_ (_08854_, _08488_, _07974_);
  and _60076_ (_08855_, _08854_, _08493_);
  nand _60077_ (_08856_, _08855_, _08853_);
  nand _60078_ (_08857_, _08856_, _08852_);
  nand _60079_ (_08858_, _08857_, _08499_);
  and _60080_ (_08859_, _08858_, _08463_);
  and _60081_ (_08860_, _08859_, _08848_);
  or _60082_ (_08861_, _08479_, \oc8051_golden_model_1.IRAM[10] [6]);
  or _60083_ (_08862_, _08488_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _60084_ (_08863_, _08862_, _08861_);
  nand _60085_ (_08864_, _08863_, _08493_);
  or _60086_ (_08865_, _08479_, \oc8051_golden_model_1.IRAM[8] [6]);
  or _60087_ (_08866_, _08488_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand _60088_ (_08867_, _08866_, _08865_);
  nand _60089_ (_08868_, _08867_, _08487_);
  nand _60090_ (_08869_, _08868_, _08864_);
  nand _60091_ (_08870_, _08869_, _08472_);
  or _60092_ (_08871_, _08479_, \oc8051_golden_model_1.IRAM[14] [6]);
  or _60093_ (_08872_, _08488_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _60094_ (_08873_, _08872_, _08871_);
  nand _60095_ (_08874_, _08873_, _08493_);
  or _60096_ (_08875_, _08479_, \oc8051_golden_model_1.IRAM[12] [6]);
  or _60097_ (_08876_, _08488_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand _60098_ (_08877_, _08876_, _08875_);
  nand _60099_ (_08878_, _08877_, _08487_);
  nand _60100_ (_08879_, _08878_, _08874_);
  nand _60101_ (_08880_, _08879_, _08499_);
  and _60102_ (_08881_, _08880_, _08512_);
  and _60103_ (_08882_, _08881_, _08870_);
  nor _60104_ (_08883_, _08882_, _08860_);
  or _60105_ (_08884_, _08479_, _08049_);
  or _60106_ (_08885_, _08488_, _08051_);
  and _60107_ (_08886_, _08885_, _08487_);
  nand _60108_ (_08887_, _08886_, _08884_);
  or _60109_ (_08888_, _08479_, _08057_);
  or _60110_ (_08889_, _08488_, _08055_);
  and _60111_ (_08890_, _08889_, _08493_);
  nand _60112_ (_08891_, _08890_, _08888_);
  nand _60113_ (_08892_, _08891_, _08887_);
  nand _60114_ (_08893_, _08892_, _08472_);
  or _60115_ (_08894_, _08479_, _08069_);
  or _60116_ (_08895_, _08488_, _08071_);
  and _60117_ (_08896_, _08895_, _08487_);
  nand _60118_ (_08897_, _08896_, _08894_);
  or _60119_ (_08898_, _08479_, _08065_);
  or _60120_ (_08899_, _08488_, _08063_);
  and _60121_ (_08900_, _08899_, _08493_);
  nand _60122_ (_08901_, _08900_, _08898_);
  nand _60123_ (_08902_, _08901_, _08897_);
  nand _60124_ (_08903_, _08902_, _08499_);
  and _60125_ (_08904_, _08903_, _08463_);
  and _60126_ (_08906_, _08904_, _08893_);
  or _60127_ (_08907_, _08479_, \oc8051_golden_model_1.IRAM[10] [5]);
  or _60128_ (_08908_, _08488_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _60129_ (_08909_, _08908_, _08907_);
  nand _60130_ (_08910_, _08909_, _08493_);
  or _60131_ (_08911_, _08479_, \oc8051_golden_model_1.IRAM[8] [5]);
  or _60132_ (_08912_, _08488_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand _60133_ (_08913_, _08912_, _08911_);
  nand _60134_ (_08914_, _08913_, _08487_);
  nand _60135_ (_08915_, _08914_, _08910_);
  nand _60136_ (_08917_, _08915_, _08472_);
  or _60137_ (_08918_, _08479_, \oc8051_golden_model_1.IRAM[14] [5]);
  or _60138_ (_08919_, _08488_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _60139_ (_08920_, _08919_, _08918_);
  nand _60140_ (_08921_, _08920_, _08493_);
  or _60141_ (_08922_, _08479_, \oc8051_golden_model_1.IRAM[12] [5]);
  or _60142_ (_08923_, _08488_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand _60143_ (_08924_, _08923_, _08922_);
  nand _60144_ (_08925_, _08924_, _08487_);
  nand _60145_ (_08926_, _08925_, _08921_);
  nand _60146_ (_08928_, _08926_, _08499_);
  and _60147_ (_08929_, _08928_, _08512_);
  and _60148_ (_08930_, _08929_, _08917_);
  nor _60149_ (_08931_, _08930_, _08906_);
  or _60150_ (_08932_, _08479_, _08284_);
  or _60151_ (_08933_, _08488_, _08286_);
  and _60152_ (_08934_, _08933_, _08487_);
  nand _60153_ (_08935_, _08934_, _08932_);
  or _60154_ (_08936_, _08479_, _08292_);
  or _60155_ (_08937_, _08488_, _08290_);
  and _60156_ (_08939_, _08937_, _08493_);
  nand _60157_ (_08940_, _08939_, _08936_);
  nand _60158_ (_08941_, _08940_, _08935_);
  nand _60159_ (_08942_, _08941_, _08472_);
  or _60160_ (_08943_, _08479_, _08304_);
  or _60161_ (_08944_, _08488_, _08306_);
  and _60162_ (_08945_, _08944_, _08487_);
  nand _60163_ (_08946_, _08945_, _08943_);
  or _60164_ (_08947_, _08479_, _08300_);
  or _60165_ (_08948_, _08488_, _08298_);
  and _60166_ (_08950_, _08948_, _08493_);
  nand _60167_ (_08951_, _08950_, _08947_);
  nand _60168_ (_08952_, _08951_, _08946_);
  nand _60169_ (_08953_, _08952_, _08499_);
  and _60170_ (_08954_, _08953_, _08463_);
  and _60171_ (_08955_, _08954_, _08942_);
  or _60172_ (_08956_, _08479_, \oc8051_golden_model_1.IRAM[10] [4]);
  or _60173_ (_08957_, _08488_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _60174_ (_08958_, _08957_, _08956_);
  nand _60175_ (_08959_, _08958_, _08493_);
  or _60176_ (_08961_, _08479_, \oc8051_golden_model_1.IRAM[8] [4]);
  or _60177_ (_08962_, _08488_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand _60178_ (_08963_, _08962_, _08961_);
  nand _60179_ (_08964_, _08963_, _08487_);
  nand _60180_ (_08965_, _08964_, _08959_);
  nand _60181_ (_08966_, _08965_, _08472_);
  or _60182_ (_08967_, _08479_, \oc8051_golden_model_1.IRAM[14] [4]);
  or _60183_ (_08968_, _08488_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _60184_ (_08969_, _08968_, _08967_);
  nand _60185_ (_08970_, _08969_, _08493_);
  or _60186_ (_08972_, _08479_, \oc8051_golden_model_1.IRAM[12] [4]);
  or _60187_ (_08973_, _08488_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand _60188_ (_08974_, _08973_, _08972_);
  nand _60189_ (_08975_, _08974_, _08487_);
  nand _60190_ (_08976_, _08975_, _08970_);
  nand _60191_ (_08977_, _08976_, _08499_);
  and _60192_ (_08978_, _08977_, _08512_);
  and _60193_ (_08979_, _08978_, _08966_);
  nor _60194_ (_08980_, _08979_, _08955_);
  or _60195_ (_08981_, _08479_, _07422_);
  or _60196_ (_08982_, _08488_, _07424_);
  and _60197_ (_08983_, _08982_, _08487_);
  nand _60198_ (_08984_, _08983_, _08981_);
  or _60199_ (_08985_, _08479_, _07430_);
  or _60200_ (_08986_, _08488_, _07428_);
  and _60201_ (_08987_, _08986_, _08493_);
  nand _60202_ (_08988_, _08987_, _08985_);
  nand _60203_ (_08989_, _08988_, _08984_);
  nand _60204_ (_08990_, _08989_, _08472_);
  or _60205_ (_08991_, _08479_, _07442_);
  or _60206_ (_08992_, _08488_, _07444_);
  and _60207_ (_08993_, _08992_, _08487_);
  nand _60208_ (_08994_, _08993_, _08991_);
  or _60209_ (_08995_, _08479_, _07438_);
  or _60210_ (_08996_, _08488_, _07436_);
  and _60211_ (_08997_, _08996_, _08493_);
  nand _60212_ (_08998_, _08997_, _08995_);
  nand _60213_ (_08999_, _08998_, _08994_);
  nand _60214_ (_09000_, _08999_, _08499_);
  and _60215_ (_09001_, _09000_, _08463_);
  and _60216_ (_09002_, _09001_, _08990_);
  or _60217_ (_09003_, _08479_, \oc8051_golden_model_1.IRAM[10] [3]);
  or _60218_ (_09004_, _08488_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _60219_ (_09005_, _09004_, _09003_);
  nand _60220_ (_09006_, _09005_, _08493_);
  or _60221_ (_09007_, _08479_, \oc8051_golden_model_1.IRAM[8] [3]);
  or _60222_ (_09008_, _08488_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand _60223_ (_09009_, _09008_, _09007_);
  nand _60224_ (_09010_, _09009_, _08487_);
  nand _60225_ (_09011_, _09010_, _09006_);
  nand _60226_ (_09012_, _09011_, _08472_);
  or _60227_ (_09013_, _08479_, \oc8051_golden_model_1.IRAM[14] [3]);
  or _60228_ (_09014_, _08488_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _60229_ (_09015_, _09014_, _09013_);
  nand _60230_ (_09016_, _09015_, _08493_);
  or _60231_ (_09017_, _08479_, \oc8051_golden_model_1.IRAM[12] [3]);
  or _60232_ (_09018_, _08488_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand _60233_ (_09019_, _09018_, _09017_);
  nand _60234_ (_09020_, _09019_, _08487_);
  nand _60235_ (_09021_, _09020_, _09016_);
  nand _60236_ (_09022_, _09021_, _08499_);
  and _60237_ (_09023_, _09022_, _08512_);
  and _60238_ (_09024_, _09023_, _09012_);
  nor _60239_ (_09025_, _09024_, _09002_);
  or _60240_ (_09026_, _08479_, _07603_);
  or _60241_ (_09027_, _08488_, _07605_);
  and _60242_ (_09028_, _09027_, _08487_);
  nand _60243_ (_09029_, _09028_, _09026_);
  or _60244_ (_09030_, _08479_, _07611_);
  or _60245_ (_09031_, _08488_, _07609_);
  and _60246_ (_09032_, _09031_, _08493_);
  nand _60247_ (_09033_, _09032_, _09030_);
  nand _60248_ (_09034_, _09033_, _09029_);
  nand _60249_ (_09035_, _09034_, _08472_);
  or _60250_ (_09036_, _08479_, _07623_);
  or _60251_ (_09037_, _08488_, _07625_);
  and _60252_ (_09038_, _09037_, _08487_);
  nand _60253_ (_09039_, _09038_, _09036_);
  or _60254_ (_09040_, _08479_, _07619_);
  or _60255_ (_09041_, _08488_, _07617_);
  and _60256_ (_09042_, _09041_, _08493_);
  nand _60257_ (_09043_, _09042_, _09040_);
  nand _60258_ (_09044_, _09043_, _09039_);
  nand _60259_ (_09045_, _09044_, _08499_);
  and _60260_ (_09046_, _09045_, _08463_);
  and _60261_ (_09047_, _09046_, _09035_);
  or _60262_ (_09048_, _08479_, \oc8051_golden_model_1.IRAM[10] [2]);
  or _60263_ (_09049_, _08488_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _60264_ (_09050_, _09049_, _09048_);
  nand _60265_ (_09051_, _09050_, _08493_);
  or _60266_ (_09052_, _08479_, \oc8051_golden_model_1.IRAM[8] [2]);
  or _60267_ (_09053_, _08488_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand _60268_ (_09054_, _09053_, _09052_);
  nand _60269_ (_09055_, _09054_, _08487_);
  nand _60270_ (_09056_, _09055_, _09051_);
  nand _60271_ (_09057_, _09056_, _08472_);
  or _60272_ (_09058_, _08479_, \oc8051_golden_model_1.IRAM[14] [2]);
  or _60273_ (_09059_, _08488_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _60274_ (_09060_, _09059_, _09058_);
  nand _60275_ (_09061_, _09060_, _08493_);
  or _60276_ (_09062_, _08479_, \oc8051_golden_model_1.IRAM[12] [2]);
  or _60277_ (_09063_, _08488_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand _60278_ (_09064_, _09063_, _09062_);
  nand _60279_ (_09065_, _09064_, _08487_);
  nand _60280_ (_09066_, _09065_, _09061_);
  nand _60281_ (_09067_, _09066_, _08499_);
  and _60282_ (_09068_, _09067_, _08512_);
  and _60283_ (_09069_, _09068_, _09057_);
  nor _60284_ (_09070_, _09069_, _09047_);
  or _60285_ (_09071_, _08479_, _07193_);
  or _60286_ (_09072_, _08488_, _07195_);
  and _60287_ (_09073_, _09072_, _08487_);
  nand _60288_ (_09074_, _09073_, _09071_);
  or _60289_ (_09075_, _08479_, _07201_);
  or _60290_ (_09076_, _08488_, _07199_);
  and _60291_ (_09077_, _09076_, _08493_);
  nand _60292_ (_09078_, _09077_, _09075_);
  nand _60293_ (_09079_, _09078_, _09074_);
  nand _60294_ (_09080_, _09079_, _08472_);
  or _60295_ (_09081_, _08479_, _07213_);
  or _60296_ (_09082_, _08488_, _07215_);
  and _60297_ (_09083_, _09082_, _08487_);
  nand _60298_ (_09084_, _09083_, _09081_);
  or _60299_ (_09085_, _08479_, _07209_);
  or _60300_ (_09086_, _08488_, _07207_);
  and _60301_ (_09087_, _09086_, _08493_);
  nand _60302_ (_09088_, _09087_, _09085_);
  nand _60303_ (_09089_, _09088_, _09084_);
  nand _60304_ (_09090_, _09089_, _08499_);
  and _60305_ (_09091_, _09090_, _08463_);
  and _60306_ (_09092_, _09091_, _09080_);
  or _60307_ (_09093_, _08479_, \oc8051_golden_model_1.IRAM[10] [1]);
  or _60308_ (_09094_, _08488_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _60309_ (_09095_, _09094_, _09093_);
  nand _60310_ (_09096_, _09095_, _08493_);
  or _60311_ (_09097_, _08479_, \oc8051_golden_model_1.IRAM[8] [1]);
  or _60312_ (_09098_, _08488_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand _60313_ (_09099_, _09098_, _09097_);
  nand _60314_ (_09100_, _09099_, _08487_);
  nand _60315_ (_09101_, _09100_, _09096_);
  nand _60316_ (_09102_, _09101_, _08472_);
  or _60317_ (_09103_, _08479_, \oc8051_golden_model_1.IRAM[14] [1]);
  or _60318_ (_09104_, _08488_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _60319_ (_09105_, _09104_, _09103_);
  nand _60320_ (_09106_, _09105_, _08493_);
  or _60321_ (_09107_, _08479_, \oc8051_golden_model_1.IRAM[12] [1]);
  or _60322_ (_09108_, _08488_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand _60323_ (_09109_, _09108_, _09107_);
  nand _60324_ (_09110_, _09109_, _08487_);
  nand _60325_ (_09111_, _09110_, _09106_);
  nand _60326_ (_09112_, _09111_, _08499_);
  and _60327_ (_09113_, _09112_, _08512_);
  and _60328_ (_09114_, _09113_, _09102_);
  or _60329_ (_09115_, _09114_, _09092_);
  or _60330_ (_09116_, _08479_, _06638_);
  or _60331_ (_09117_, _08488_, _06992_);
  and _60332_ (_09118_, _09117_, _08487_);
  nand _60333_ (_09119_, _09118_, _09116_);
  or _60334_ (_09120_, _08479_, _07000_);
  or _60335_ (_09121_, _08488_, _06997_);
  and _60336_ (_09122_, _09121_, _08493_);
  nand _60337_ (_09123_, _09122_, _09120_);
  nand _60338_ (_09124_, _09123_, _09119_);
  nand _60339_ (_09125_, _09124_, _08472_);
  or _60340_ (_09126_, _08479_, _07013_);
  or _60341_ (_09127_, _08488_, _07015_);
  and _60342_ (_09128_, _09127_, _08487_);
  nand _60343_ (_09129_, _09128_, _09126_);
  or _60344_ (_09130_, _08479_, _07009_);
  or _60345_ (_09131_, _08488_, _07007_);
  and _60346_ (_09132_, _09131_, _08493_);
  nand _60347_ (_09133_, _09132_, _09130_);
  nand _60348_ (_09134_, _09133_, _09129_);
  nand _60349_ (_09135_, _09134_, _08499_);
  and _60350_ (_09136_, _09135_, _08463_);
  and _60351_ (_09137_, _09136_, _09125_);
  or _60352_ (_09138_, _08479_, \oc8051_golden_model_1.IRAM[10] [0]);
  or _60353_ (_09139_, _08488_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _60354_ (_09140_, _09139_, _09138_);
  nand _60355_ (_09141_, _09140_, _08493_);
  or _60356_ (_09142_, _08479_, \oc8051_golden_model_1.IRAM[8] [0]);
  or _60357_ (_09143_, _08488_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand _60358_ (_09144_, _09143_, _09142_);
  nand _60359_ (_09145_, _09144_, _08487_);
  nand _60360_ (_09146_, _09145_, _09141_);
  nand _60361_ (_09147_, _09146_, _08472_);
  or _60362_ (_09148_, _08479_, \oc8051_golden_model_1.IRAM[14] [0]);
  or _60363_ (_09149_, _08488_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand _60364_ (_09150_, _09149_, _09148_);
  nand _60365_ (_09151_, _09150_, _08493_);
  or _60366_ (_09152_, _08479_, \oc8051_golden_model_1.IRAM[12] [0]);
  or _60367_ (_09153_, _08488_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand _60368_ (_09154_, _09153_, _09152_);
  nand _60369_ (_09155_, _09154_, _08487_);
  nand _60370_ (_09156_, _09155_, _09151_);
  nand _60371_ (_09157_, _09156_, _08499_);
  and _60372_ (_09158_, _09157_, _08512_);
  and _60373_ (_09159_, _09158_, _09147_);
  or _60374_ (_09160_, _09159_, _09137_);
  nor _60375_ (_09161_, _09160_, _09115_);
  and _60376_ (_09162_, _09161_, _09070_);
  and _60377_ (_09163_, _09162_, _09025_);
  and _60378_ (_09164_, _09163_, _08980_);
  and _60379_ (_09165_, _09164_, _08931_);
  and _60380_ (_09166_, _09165_, _08883_);
  nor _60381_ (_09167_, _09166_, _08838_);
  and _60382_ (_09168_, _09166_, _08838_);
  or _60383_ (_09169_, _09168_, _09167_);
  or _60384_ (_09170_, _09169_, _07154_);
  and _60385_ (_09171_, _09170_, _08837_);
  and _60386_ (_09172_, _09171_, _08836_);
  and _60387_ (_09173_, _08548_, _07152_);
  or _60388_ (_09174_, _09173_, _06310_);
  or _60389_ (_09175_, _09174_, _09172_);
  and _60390_ (_09176_, _05449_, _05424_);
  and _60391_ (_09177_, _09176_, _08433_);
  and _60392_ (_09178_, _09177_, \oc8051_golden_model_1.PC [7]);
  nor _60393_ (_09179_, _09177_, \oc8051_golden_model_1.PC [7]);
  nor _60394_ (_09180_, _09179_, _09178_);
  not _60395_ (_09181_, _09180_);
  nand _60396_ (_09182_, _09181_, _06310_);
  and _60397_ (_09183_, _09182_, _09175_);
  or _60398_ (_09184_, _09183_, _05823_);
  and _60399_ (_09185_, _08573_, _05823_);
  nor _60400_ (_09186_, _09185_, _06073_);
  and _60401_ (_09187_, _09186_, _09184_);
  and _60402_ (_09188_, _08426_, _06073_);
  and _60403_ (_09189_, _05820_, _05666_);
  nor _60404_ (_09190_, _09189_, _09188_);
  not _60405_ (_09191_, _09190_);
  nor _60406_ (_09192_, _09191_, _09187_);
  not _60407_ (_09193_, _09189_);
  nand _60408_ (_09194_, _07922_, _07892_);
  and _60409_ (_09195_, _07306_, _07049_);
  and _60410_ (_09196_, _09195_, _07708_);
  and _60411_ (_09197_, _09196_, _07544_);
  and _60412_ (_09198_, _09197_, _08336_);
  and _60413_ (_09199_, _09198_, _08101_);
  and _60414_ (_09200_, _09199_, _08012_);
  nor _60415_ (_09201_, _09200_, _09194_);
  and _60416_ (_09202_, _09200_, _09194_);
  or _60417_ (_09203_, _09202_, _09201_);
  nor _60418_ (_09204_, _09203_, _09193_);
  nor _60419_ (_09205_, _09204_, _09192_);
  nor _60420_ (_09206_, _09205_, _07168_);
  or _60421_ (_09207_, _08882_, _08860_);
  or _60422_ (_09208_, _08930_, _08906_);
  or _60423_ (_09209_, _08979_, _08955_);
  or _60424_ (_09210_, _09024_, _09002_);
  or _60425_ (_09211_, _09069_, _09047_);
  and _60426_ (_09212_, _09160_, _09115_);
  and _60427_ (_09213_, _09212_, _09211_);
  and _60428_ (_09214_, _09213_, _09210_);
  and _60429_ (_09215_, _09214_, _09209_);
  and _60430_ (_09216_, _09215_, _09208_);
  and _60431_ (_09217_, _09216_, _09207_);
  nor _60432_ (_09218_, _09217_, _08838_);
  and _60433_ (_09219_, _09217_, _08838_);
  or _60434_ (_09220_, _09219_, _09218_);
  nor _60435_ (_09221_, _09220_, _07169_);
  nor _60436_ (_09222_, _09221_, _07167_);
  not _60437_ (_09223_, _09222_);
  nor _60438_ (_09224_, _09223_, _09206_);
  nor _60439_ (_09225_, _09224_, _08346_);
  nor _60440_ (_09226_, _09225_, _07418_);
  or _60441_ (_09227_, _09226_, _07770_);
  and _60442_ (_09228_, _09227_, _07769_);
  not _60443_ (_09229_, \oc8051_golden_model_1.PC [15]);
  and _60444_ (_09230_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and _60445_ (_09231_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and _60446_ (_09232_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and _60447_ (_09233_, _09232_, _09231_);
  and _60448_ (_09234_, _09233_, _09178_);
  and _60449_ (_09235_, _09234_, _09230_);
  and _60450_ (_09236_, _09235_, \oc8051_golden_model_1.PC [14]);
  and _60451_ (_09237_, _09236_, _09229_);
  nor _60452_ (_09238_, _09236_, _09229_);
  or _60453_ (_09239_, _09238_, _09237_);
  not _60454_ (_09240_, _09239_);
  nand _60455_ (_09241_, _09240_, _06310_);
  and _60456_ (_09242_, _09231_, \oc8051_golden_model_1.PC [10]);
  and _60457_ (_09243_, _09242_, _08435_);
  and _60458_ (_09244_, _09243_, \oc8051_golden_model_1.PC [11]);
  and _60459_ (_09245_, _09244_, \oc8051_golden_model_1.PC [12]);
  and _60460_ (_09246_, _09245_, \oc8051_golden_model_1.PC [13]);
  and _60461_ (_09247_, _09246_, \oc8051_golden_model_1.PC [14]);
  nor _60462_ (_09248_, _09247_, \oc8051_golden_model_1.PC [15]);
  and _60463_ (_09249_, _09231_, _08435_);
  and _60464_ (_09250_, _09249_, \oc8051_golden_model_1.PC [10]);
  and _60465_ (_09251_, _09250_, \oc8051_golden_model_1.PC [11]);
  and _60466_ (_09252_, _09251_, \oc8051_golden_model_1.PC [12]);
  and _60467_ (_09253_, _09252_, \oc8051_golden_model_1.PC [13]);
  and _60468_ (_09254_, _09253_, \oc8051_golden_model_1.PC [14]);
  and _60469_ (_09255_, _09254_, \oc8051_golden_model_1.PC [15]);
  nor _60470_ (_09256_, _09255_, _09248_);
  or _60471_ (_09257_, _09256_, _06310_);
  and _60472_ (_09258_, _09257_, _09241_);
  and _60473_ (_09259_, _09258_, _07764_);
  and _60474_ (_09260_, _09259_, _07767_);
  or _60475_ (_40979_, _09260_, _09228_);
  not _60476_ (_09261_, \oc8051_golden_model_1.B [7]);
  nor _60477_ (_09262_, _01317_, _09261_);
  nor _60478_ (_09263_, _07841_, _09261_);
  and _60479_ (_09264_, _07923_, _07841_);
  or _60480_ (_09265_, _09264_, _09263_);
  or _60481_ (_09266_, _09265_, _06132_);
  nor _60482_ (_09267_, _08420_, _09261_);
  and _60483_ (_09268_, _08426_, _08420_);
  or _60484_ (_09269_, _09268_, _09267_);
  and _60485_ (_09270_, _09269_, _06152_);
  and _60486_ (_09271_, _08548_, _07841_);
  or _60487_ (_09272_, _09271_, _09263_);
  or _60488_ (_09273_, _09272_, _06161_);
  and _60489_ (_09274_, _07841_, \oc8051_golden_model_1.ACC [7]);
  or _60490_ (_09275_, _09274_, _09263_);
  and _60491_ (_09276_, _09275_, _07056_);
  nor _60492_ (_09277_, _07056_, _09261_);
  or _60493_ (_09278_, _09277_, _06160_);
  or _60494_ (_09279_, _09278_, _09276_);
  and _60495_ (_09280_, _09279_, _06157_);
  and _60496_ (_09281_, _09280_, _09273_);
  and _60497_ (_09282_, _08552_, _08420_);
  or _60498_ (_09283_, _09282_, _09267_);
  and _60499_ (_09284_, _09283_, _06156_);
  or _60500_ (_09285_, _09284_, _06217_);
  or _60501_ (_09286_, _09285_, _09281_);
  or _60502_ (_09287_, _09265_, _07075_);
  and _60503_ (_09288_, _09287_, _09286_);
  or _60504_ (_09289_, _09288_, _06220_);
  or _60505_ (_09290_, _09275_, _06229_);
  and _60506_ (_09291_, _09290_, _06153_);
  and _60507_ (_09292_, _09291_, _09289_);
  or _60508_ (_09293_, _09292_, _09270_);
  and _60509_ (_09294_, _09293_, _06146_);
  and _60510_ (_09295_, _06294_, _06245_);
  or _60511_ (_09296_, _09267_, _08568_);
  and _60512_ (_09297_, _09283_, _06145_);
  and _60513_ (_09298_, _09297_, _09296_);
  or _60514_ (_09299_, _09298_, _09295_);
  or _60515_ (_09300_, _09299_, _09294_);
  not _60516_ (_09301_, _09295_);
  and _60517_ (_09302_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and _60518_ (_09303_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and _60519_ (_09304_, _09303_, _09302_);
  and _60520_ (_09305_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and _60521_ (_09306_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and _60522_ (_09307_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor _60523_ (_09308_, _09307_, _09306_);
  nor _60524_ (_09309_, _09308_, _09304_);
  and _60525_ (_09310_, _09309_, _09305_);
  nor _60526_ (_09311_, _09310_, _09304_);
  and _60527_ (_09312_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and _60528_ (_09313_, _09312_, _09306_);
  and _60529_ (_09314_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor _60530_ (_09315_, _09314_, _09302_);
  nor _60531_ (_09316_, _09315_, _09313_);
  not _60532_ (_09317_, _09316_);
  nor _60533_ (_09318_, _09317_, _09311_);
  and _60534_ (_09319_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and _60535_ (_09320_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and _60536_ (_09321_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and _60537_ (_09322_, _09321_, _09320_);
  nor _60538_ (_09323_, _09321_, _09320_);
  nor _60539_ (_09324_, _09323_, _09322_);
  and _60540_ (_09325_, _09324_, _09319_);
  nor _60541_ (_09326_, _09324_, _09319_);
  nor _60542_ (_09327_, _09326_, _09325_);
  and _60543_ (_09328_, _09317_, _09311_);
  nor _60544_ (_09329_, _09328_, _09318_);
  and _60545_ (_09330_, _09329_, _09327_);
  nor _60546_ (_09331_, _09330_, _09318_);
  not _60547_ (_09332_, _09306_);
  and _60548_ (_09333_, _09312_, _09332_);
  and _60549_ (_09334_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and _60550_ (_09335_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and _60551_ (_09336_, _09335_, _09320_);
  and _60552_ (_09337_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  and _60553_ (_09338_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor _60554_ (_09339_, _09338_, _09337_);
  nor _60555_ (_09340_, _09339_, _09336_);
  and _60556_ (_09341_, _09340_, _09334_);
  nor _60557_ (_09342_, _09340_, _09334_);
  nor _60558_ (_09343_, _09342_, _09341_);
  and _60559_ (_09344_, _09343_, _09333_);
  nor _60560_ (_09345_, _09343_, _09333_);
  nor _60561_ (_09346_, _09345_, _09344_);
  not _60562_ (_09347_, _09346_);
  nor _60563_ (_09348_, _09347_, _09331_);
  and _60564_ (_09349_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and _60565_ (_09350_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and _60566_ (_09351_, _09350_, _09349_);
  nor _60567_ (_09352_, _09325_, _09322_);
  and _60568_ (_09353_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and _60569_ (_09354_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and _60570_ (_09355_, _09354_, _09353_);
  nor _60571_ (_09356_, _09354_, _09353_);
  nor _60572_ (_09357_, _09356_, _09355_);
  not _60573_ (_09358_, _09357_);
  nor _60574_ (_09359_, _09358_, _09352_);
  and _60575_ (_09360_, _09358_, _09352_);
  nor _60576_ (_09361_, _09360_, _09359_);
  and _60577_ (_09362_, _09361_, _09351_);
  nor _60578_ (_09363_, _09361_, _09351_);
  nor _60579_ (_09364_, _09363_, _09362_);
  and _60580_ (_09365_, _09347_, _09331_);
  nor _60581_ (_09366_, _09365_, _09348_);
  and _60582_ (_09367_, _09366_, _09364_);
  nor _60583_ (_09368_, _09367_, _09348_);
  nor _60584_ (_09369_, _09341_, _09336_);
  and _60585_ (_09370_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and _60586_ (_09371_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and _60587_ (_09372_, _09371_, _09370_);
  nor _60588_ (_09373_, _09371_, _09370_);
  nor _60589_ (_09374_, _09373_, _09372_);
  not _60590_ (_09375_, _09374_);
  nor _60591_ (_09376_, _09375_, _09369_);
  and _60592_ (_09377_, _09375_, _09369_);
  nor _60593_ (_09378_, _09377_, _09376_);
  and _60594_ (_09379_, _09378_, _09355_);
  nor _60595_ (_09380_, _09378_, _09355_);
  nor _60596_ (_09381_, _09380_, _09379_);
  nor _60597_ (_09382_, _09344_, _09313_);
  and _60598_ (_09383_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  and _60599_ (_09384_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and _60600_ (_09385_, _09384_, _09335_);
  nor _60601_ (_09386_, _09384_, _09335_);
  nor _60602_ (_09387_, _09386_, _09385_);
  and _60603_ (_09388_, _09387_, _09383_);
  nor _60604_ (_09389_, _09387_, _09383_);
  nor _60605_ (_09390_, _09389_, _09388_);
  not _60606_ (_09391_, _09390_);
  nor _60607_ (_09392_, _09391_, _09382_);
  and _60608_ (_09393_, _09391_, _09382_);
  nor _60609_ (_09394_, _09393_, _09392_);
  and _60610_ (_09395_, _09394_, _09381_);
  nor _60611_ (_09396_, _09394_, _09381_);
  nor _60612_ (_09397_, _09396_, _09395_);
  not _60613_ (_09398_, _09397_);
  nor _60614_ (_09399_, _09398_, _09368_);
  nor _60615_ (_09400_, _09362_, _09359_);
  not _60616_ (_09401_, _09400_);
  and _60617_ (_09402_, _09398_, _09368_);
  nor _60618_ (_09403_, _09402_, _09399_);
  and _60619_ (_09404_, _09403_, _09401_);
  nor _60620_ (_09405_, _09404_, _09399_);
  nor _60621_ (_09406_, _09379_, _09376_);
  not _60622_ (_09407_, _09406_);
  nor _60623_ (_09408_, _09395_, _09392_);
  not _60624_ (_09409_, _09408_);
  and _60625_ (_09410_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and _60626_ (_09411_, _09410_, _09335_);
  and _60627_ (_09412_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and _60628_ (_09413_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor _60629_ (_09414_, _09413_, _09412_);
  nor _60630_ (_09415_, _09414_, _09411_);
  nor _60631_ (_09416_, _09388_, _09385_);
  and _60632_ (_09417_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and _60633_ (_09418_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and _60634_ (_09419_, _09418_, _09417_);
  nor _60635_ (_09420_, _09418_, _09417_);
  nor _60636_ (_09421_, _09420_, _09419_);
  not _60637_ (_09422_, _09421_);
  nor _60638_ (_09423_, _09422_, _09416_);
  and _60639_ (_09424_, _09422_, _09416_);
  nor _60640_ (_09425_, _09424_, _09423_);
  and _60641_ (_09426_, _09425_, _09372_);
  nor _60642_ (_09427_, _09425_, _09372_);
  nor _60643_ (_09428_, _09427_, _09426_);
  and _60644_ (_09429_, _09428_, _09415_);
  nor _60645_ (_09430_, _09428_, _09415_);
  nor _60646_ (_09431_, _09430_, _09429_);
  and _60647_ (_09432_, _09431_, _09409_);
  nor _60648_ (_09433_, _09431_, _09409_);
  nor _60649_ (_09434_, _09433_, _09432_);
  and _60650_ (_09435_, _09434_, _09407_);
  nor _60651_ (_09436_, _09434_, _09407_);
  nor _60652_ (_09437_, _09436_, _09435_);
  not _60653_ (_09438_, _09437_);
  nor _60654_ (_09439_, _09438_, _09405_);
  nor _60655_ (_09440_, _09435_, _09432_);
  nor _60656_ (_09441_, _09426_, _09423_);
  not _60657_ (_09442_, _09441_);
  and _60658_ (_09443_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and _60659_ (_09444_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and _60660_ (_09445_, _09444_, _09443_);
  nor _60661_ (_09446_, _09444_, _09443_);
  nor _60662_ (_09447_, _09446_, _09445_);
  and _60663_ (_09448_, _09447_, _09411_);
  nor _60664_ (_09449_, _09447_, _09411_);
  nor _60665_ (_09450_, _09449_, _09448_);
  and _60666_ (_09451_, _09450_, _09419_);
  nor _60667_ (_09452_, _09450_, _09419_);
  nor _60668_ (_09453_, _09452_, _09451_);
  and _60669_ (_09454_, _09453_, _09410_);
  nor _60670_ (_09455_, _09453_, _09410_);
  nor _60671_ (_09456_, _09455_, _09454_);
  and _60672_ (_09457_, _09456_, _09429_);
  nor _60673_ (_09458_, _09456_, _09429_);
  nor _60674_ (_09459_, _09458_, _09457_);
  and _60675_ (_09460_, _09459_, _09442_);
  nor _60676_ (_09461_, _09459_, _09442_);
  nor _60677_ (_09462_, _09461_, _09460_);
  not _60678_ (_09463_, _09462_);
  nor _60679_ (_09464_, _09463_, _09440_);
  and _60680_ (_09465_, _09463_, _09440_);
  nor _60681_ (_09466_, _09465_, _09464_);
  and _60682_ (_09467_, _09466_, _09439_);
  nor _60683_ (_09468_, _09460_, _09457_);
  nor _60684_ (_09469_, _09451_, _09448_);
  not _60685_ (_09470_, _09469_);
  and _60686_ (_09471_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and _60687_ (_09472_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and _60688_ (_09473_, _09472_, _09471_);
  nor _60689_ (_09474_, _09472_, _09471_);
  nor _60690_ (_09475_, _09474_, _09473_);
  and _60691_ (_09476_, _09475_, _09445_);
  nor _60692_ (_09477_, _09475_, _09445_);
  nor _60693_ (_09478_, _09477_, _09476_);
  and _60694_ (_09479_, _09478_, _09454_);
  nor _60695_ (_09480_, _09478_, _09454_);
  nor _60696_ (_09481_, _09480_, _09479_);
  and _60697_ (_09482_, _09481_, _09470_);
  nor _60698_ (_09483_, _09481_, _09470_);
  nor _60699_ (_09484_, _09483_, _09482_);
  not _60700_ (_09485_, _09484_);
  nor _60701_ (_09486_, _09485_, _09468_);
  and _60702_ (_09487_, _09485_, _09468_);
  nor _60703_ (_09488_, _09487_, _09486_);
  and _60704_ (_09489_, _09488_, _09464_);
  nor _60705_ (_09490_, _09488_, _09464_);
  nor _60706_ (_09491_, _09490_, _09489_);
  and _60707_ (_09492_, _09491_, _09467_);
  nor _60708_ (_09493_, _09491_, _09467_);
  and _60709_ (_09494_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and _60710_ (_09495_, _09494_, _09306_);
  and _60711_ (_09496_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and _60712_ (_09497_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor _60713_ (_09498_, _09497_, _09303_);
  nor _60714_ (_09499_, _09498_, _09495_);
  and _60715_ (_09500_, _09499_, _09496_);
  nor _60716_ (_09501_, _09500_, _09495_);
  not _60717_ (_09502_, _09501_);
  nor _60718_ (_09503_, _09309_, _09305_);
  nor _60719_ (_09504_, _09503_, _09310_);
  and _60720_ (_09505_, _09504_, _09502_);
  and _60721_ (_09506_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and _60722_ (_09507_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and _60723_ (_09508_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and _60724_ (_09509_, _09508_, _09507_);
  nor _60725_ (_09510_, _09508_, _09507_);
  nor _60726_ (_09511_, _09510_, _09509_);
  and _60727_ (_09512_, _09511_, _09506_);
  nor _60728_ (_09513_, _09511_, _09506_);
  nor _60729_ (_09514_, _09513_, _09512_);
  nor _60730_ (_09515_, _09504_, _09502_);
  nor _60731_ (_09516_, _09515_, _09505_);
  and _60732_ (_09517_, _09516_, _09514_);
  nor _60733_ (_09518_, _09517_, _09505_);
  nor _60734_ (_09519_, _09329_, _09327_);
  nor _60735_ (_09520_, _09519_, _09330_);
  not _60736_ (_09522_, _09520_);
  nor _60737_ (_09523_, _09522_, _09518_);
  and _60738_ (_09524_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and _60739_ (_09525_, _09524_, _09350_);
  nor _60740_ (_09526_, _09512_, _09509_);
  nor _60741_ (_09527_, _09350_, _09349_);
  nor _60742_ (_09528_, _09527_, _09351_);
  not _60743_ (_09529_, _09528_);
  nor _60744_ (_09530_, _09529_, _09526_);
  and _60745_ (_09531_, _09529_, _09526_);
  nor _60746_ (_09532_, _09531_, _09530_);
  and _60747_ (_09533_, _09532_, _09525_);
  nor _60748_ (_09534_, _09532_, _09525_);
  nor _60749_ (_09535_, _09534_, _09533_);
  and _60750_ (_09536_, _09522_, _09518_);
  nor _60751_ (_09537_, _09536_, _09523_);
  and _60752_ (_09538_, _09537_, _09535_);
  nor _60753_ (_09539_, _09538_, _09523_);
  nor _60754_ (_09540_, _09366_, _09364_);
  nor _60755_ (_09541_, _09540_, _09367_);
  not _60756_ (_09543_, _09541_);
  nor _60757_ (_09544_, _09543_, _09539_);
  nor _60758_ (_09545_, _09533_, _09530_);
  not _60759_ (_09546_, _09545_);
  and _60760_ (_09547_, _09543_, _09539_);
  nor _60761_ (_09548_, _09547_, _09544_);
  and _60762_ (_09549_, _09548_, _09546_);
  nor _60763_ (_09550_, _09549_, _09544_);
  nor _60764_ (_09551_, _09403_, _09401_);
  nor _60765_ (_09552_, _09551_, _09404_);
  not _60766_ (_09553_, _09552_);
  nor _60767_ (_09554_, _09553_, _09550_);
  and _60768_ (_09555_, _09438_, _09405_);
  nor _60769_ (_09556_, _09555_, _09439_);
  and _60770_ (_09557_, _09556_, _09554_);
  nor _60771_ (_09558_, _09466_, _09439_);
  nor _60772_ (_09559_, _09558_, _09467_);
  nand _60773_ (_09560_, _09559_, _09557_);
  and _60774_ (_09561_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and _60775_ (_09562_, _09561_, _09494_);
  and _60776_ (_09563_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor _60777_ (_09564_, _09561_, _09494_);
  nor _60778_ (_09565_, _09564_, _09562_);
  and _60779_ (_09566_, _09565_, _09563_);
  nor _60780_ (_09567_, _09566_, _09562_);
  not _60781_ (_09568_, _09567_);
  nor _60782_ (_09569_, _09499_, _09496_);
  nor _60783_ (_09570_, _09569_, _09500_);
  and _60784_ (_09571_, _09570_, _09568_);
  and _60785_ (_09572_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and _60786_ (_09573_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and _60787_ (_09574_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and _60788_ (_09575_, _09574_, _09573_);
  nor _60789_ (_09576_, _09574_, _09573_);
  nor _60790_ (_09577_, _09576_, _09575_);
  and _60791_ (_09578_, _09577_, _09572_);
  nor _60792_ (_09579_, _09577_, _09572_);
  nor _60793_ (_09580_, _09579_, _09578_);
  nor _60794_ (_09581_, _09570_, _09568_);
  nor _60795_ (_09582_, _09581_, _09571_);
  and _60796_ (_09583_, _09582_, _09580_);
  nor _60797_ (_09584_, _09583_, _09571_);
  not _60798_ (_09585_, _09584_);
  nor _60799_ (_09586_, _09516_, _09514_);
  nor _60800_ (_09587_, _09586_, _09517_);
  and _60801_ (_09588_, _09587_, _09585_);
  nor _60802_ (_09589_, _09578_, _09575_);
  and _60803_ (_09590_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and _60804_ (_09591_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor _60805_ (_09592_, _09591_, _09590_);
  nor _60806_ (_09593_, _09592_, _09525_);
  not _60807_ (_09594_, _09593_);
  nor _60808_ (_09595_, _09594_, _09589_);
  and _60809_ (_09596_, _09594_, _09589_);
  nor _60810_ (_09597_, _09596_, _09595_);
  nor _60811_ (_09598_, _09587_, _09585_);
  nor _60812_ (_09599_, _09598_, _09588_);
  and _60813_ (_09600_, _09599_, _09597_);
  nor _60814_ (_09601_, _09600_, _09588_);
  nor _60815_ (_09602_, _09537_, _09535_);
  nor _60816_ (_09603_, _09602_, _09538_);
  not _60817_ (_09604_, _09603_);
  nor _60818_ (_09605_, _09604_, _09601_);
  and _60819_ (_09606_, _09604_, _09601_);
  nor _60820_ (_09607_, _09606_, _09605_);
  and _60821_ (_09608_, _09607_, _09595_);
  nor _60822_ (_09609_, _09608_, _09605_);
  nor _60823_ (_09610_, _09548_, _09546_);
  nor _60824_ (_09611_, _09610_, _09549_);
  not _60825_ (_09612_, _09611_);
  nor _60826_ (_09613_, _09612_, _09609_);
  and _60827_ (_09614_, _09553_, _09550_);
  nor _60828_ (_09615_, _09614_, _09554_);
  and _60829_ (_09616_, _09615_, _09613_);
  nor _60830_ (_09617_, _09556_, _09554_);
  nor _60831_ (_09618_, _09617_, _09557_);
  and _60832_ (_09619_, _09618_, _09616_);
  nor _60833_ (_09620_, _09618_, _09616_);
  nor _60834_ (_09621_, _09620_, _09619_);
  and _60835_ (_09622_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and _60836_ (_09623_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and _60837_ (_09624_, _09623_, _09622_);
  and _60838_ (_09625_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor _60839_ (_09626_, _09623_, _09622_);
  nor _60840_ (_09627_, _09626_, _09624_);
  and _60841_ (_09628_, _09627_, _09625_);
  nor _60842_ (_09629_, _09628_, _09624_);
  not _60843_ (_09630_, _09629_);
  nor _60844_ (_09631_, _09565_, _09563_);
  nor _60845_ (_09632_, _09631_, _09566_);
  and _60846_ (_09633_, _09632_, _09630_);
  and _60847_ (_09634_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and _60848_ (_09635_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and _60849_ (_09636_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and _60850_ (_09637_, _09636_, _09635_);
  nor _60851_ (_09638_, _09636_, _09635_);
  nor _60852_ (_09639_, _09638_, _09637_);
  and _60853_ (_09640_, _09639_, _09634_);
  nor _60854_ (_09641_, _09639_, _09634_);
  nor _60855_ (_09642_, _09641_, _09640_);
  nor _60856_ (_09643_, _09632_, _09630_);
  nor _60857_ (_09644_, _09643_, _09633_);
  and _60858_ (_09645_, _09644_, _09642_);
  nor _60859_ (_09646_, _09645_, _09633_);
  not _60860_ (_09647_, _09646_);
  nor _60861_ (_09648_, _09582_, _09580_);
  nor _60862_ (_09649_, _09648_, _09583_);
  and _60863_ (_09650_, _09649_, _09647_);
  not _60864_ (_09651_, _09524_);
  nor _60865_ (_09652_, _09640_, _09637_);
  nor _60866_ (_09653_, _09652_, _09651_);
  and _60867_ (_09654_, _09652_, _09651_);
  nor _60868_ (_09655_, _09654_, _09653_);
  nor _60869_ (_09656_, _09649_, _09647_);
  nor _60870_ (_09657_, _09656_, _09650_);
  and _60871_ (_09658_, _09657_, _09655_);
  nor _60872_ (_09659_, _09658_, _09650_);
  not _60873_ (_09660_, _09659_);
  nor _60874_ (_09661_, _09599_, _09597_);
  nor _60875_ (_09662_, _09661_, _09600_);
  and _60876_ (_09663_, _09662_, _09660_);
  nor _60877_ (_09664_, _09662_, _09660_);
  nor _60878_ (_09665_, _09664_, _09663_);
  and _60879_ (_09666_, _09665_, _09653_);
  nor _60880_ (_09667_, _09666_, _09663_);
  nor _60881_ (_09668_, _09607_, _09595_);
  nor _60882_ (_09669_, _09668_, _09608_);
  not _60883_ (_09670_, _09669_);
  nor _60884_ (_09671_, _09670_, _09667_);
  and _60885_ (_09672_, _09612_, _09609_);
  nor _60886_ (_09673_, _09672_, _09613_);
  and _60887_ (_09674_, _09673_, _09671_);
  nor _60888_ (_09675_, _09615_, _09613_);
  nor _60889_ (_09676_, _09675_, _09616_);
  nand _60890_ (_09677_, _09676_, _09674_);
  or _60891_ (_09678_, _09676_, _09674_);
  and _60892_ (_09679_, _09678_, _09677_);
  and _60893_ (_09680_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and _60894_ (_09681_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and _60895_ (_09682_, _09681_, _09680_);
  and _60896_ (_09683_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor _60897_ (_09684_, _09681_, _09680_);
  nor _60898_ (_09685_, _09684_, _09682_);
  and _60899_ (_09686_, _09685_, _09683_);
  nor _60900_ (_09687_, _09686_, _09682_);
  not _60901_ (_09688_, _09687_);
  nor _60902_ (_09689_, _09627_, _09625_);
  nor _60903_ (_09690_, _09689_, _09628_);
  and _60904_ (_09691_, _09690_, _09688_);
  and _60905_ (_09692_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and _60906_ (_09693_, _09692_, _09636_);
  and _60907_ (_09694_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and _60908_ (_09695_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor _60909_ (_09696_, _09695_, _09694_);
  nor _60910_ (_09698_, _09696_, _09693_);
  nor _60911_ (_09699_, _09690_, _09688_);
  nor _60912_ (_09701_, _09699_, _09691_);
  and _60913_ (_09702_, _09701_, _09698_);
  nor _60914_ (_09704_, _09702_, _09691_);
  not _60915_ (_09705_, _09704_);
  nor _60916_ (_09707_, _09644_, _09642_);
  nor _60917_ (_09708_, _09707_, _09645_);
  and _60918_ (_09710_, _09708_, _09705_);
  nor _60919_ (_09711_, _09708_, _09705_);
  nor _60920_ (_09713_, _09711_, _09710_);
  and _60921_ (_09714_, _09713_, _09693_);
  nor _60922_ (_09716_, _09714_, _09710_);
  not _60923_ (_09717_, _09716_);
  nor _60924_ (_09719_, _09657_, _09655_);
  nor _60925_ (_09720_, _09719_, _09658_);
  and _60926_ (_09722_, _09720_, _09717_);
  nor _60927_ (_09723_, _09665_, _09653_);
  nor _60928_ (_09725_, _09723_, _09666_);
  and _60929_ (_09726_, _09725_, _09722_);
  and _60930_ (_09728_, _09670_, _09667_);
  nor _60931_ (_09729_, _09728_, _09671_);
  and _60932_ (_09731_, _09729_, _09726_);
  nor _60933_ (_09732_, _09673_, _09671_);
  nor _60934_ (_09734_, _09732_, _09674_);
  and _60935_ (_09735_, _09734_, _09731_);
  nor _60936_ (_09736_, _09734_, _09731_);
  nor _60937_ (_09737_, _09736_, _09735_);
  and _60938_ (_09738_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and _60939_ (_09739_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and _60940_ (_09740_, _09739_, _09738_);
  and _60941_ (_09741_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor _60942_ (_09742_, _09739_, _09738_);
  nor _60943_ (_09743_, _09742_, _09740_);
  and _60944_ (_09744_, _09743_, _09741_);
  nor _60945_ (_09745_, _09744_, _09740_);
  not _60946_ (_09746_, _09745_);
  nor _60947_ (_09747_, _09685_, _09683_);
  nor _60948_ (_09748_, _09747_, _09686_);
  and _60949_ (_09749_, _09748_, _09746_);
  nor _60950_ (_09750_, _09748_, _09746_);
  nor _60951_ (_09751_, _09750_, _09749_);
  and _60952_ (_09752_, _09751_, _09692_);
  nor _60953_ (_09753_, _09752_, _09749_);
  not _60954_ (_09754_, _09753_);
  nor _60955_ (_09755_, _09701_, _09698_);
  nor _60956_ (_09756_, _09755_, _09702_);
  and _60957_ (_09757_, _09756_, _09754_);
  nor _60958_ (_09758_, _09713_, _09693_);
  nor _60959_ (_09759_, _09758_, _09714_);
  and _60960_ (_09760_, _09759_, _09757_);
  nor _60961_ (_09761_, _09720_, _09717_);
  nor _60962_ (_09762_, _09761_, _09722_);
  and _60963_ (_09763_, _09762_, _09760_);
  nor _60964_ (_09764_, _09725_, _09722_);
  nor _60965_ (_09765_, _09764_, _09726_);
  and _60966_ (_09766_, _09765_, _09763_);
  nor _60967_ (_09767_, _09729_, _09726_);
  nor _60968_ (_09768_, _09767_, _09731_);
  and _60969_ (_09769_, _09768_, _09766_);
  and _60970_ (_09770_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and _60971_ (_09771_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and _60972_ (_09772_, _09771_, _09770_);
  nor _60973_ (_09773_, _09743_, _09741_);
  nor _60974_ (_09774_, _09773_, _09744_);
  and _60975_ (_09775_, _09774_, _09772_);
  nor _60976_ (_09776_, _09751_, _09692_);
  nor _60977_ (_09777_, _09776_, _09752_);
  and _60978_ (_09778_, _09777_, _09775_);
  nor _60979_ (_09779_, _09756_, _09754_);
  nor _60980_ (_09780_, _09779_, _09757_);
  and _60981_ (_09781_, _09780_, _09778_);
  nor _60982_ (_09782_, _09759_, _09757_);
  nor _60983_ (_09783_, _09782_, _09760_);
  and _60984_ (_09784_, _09783_, _09781_);
  nor _60985_ (_09785_, _09762_, _09760_);
  nor _60986_ (_09786_, _09785_, _09763_);
  and _60987_ (_09787_, _09786_, _09784_);
  nor _60988_ (_09788_, _09765_, _09763_);
  nor _60989_ (_09789_, _09788_, _09766_);
  and _60990_ (_09790_, _09789_, _09787_);
  nor _60991_ (_09791_, _09768_, _09766_);
  nor _60992_ (_09793_, _09791_, _09769_);
  and _60993_ (_09795_, _09793_, _09790_);
  nor _60994_ (_09796_, _09795_, _09769_);
  not _60995_ (_09798_, _09796_);
  and _60996_ (_09799_, _09798_, _09737_);
  or _60997_ (_09801_, _09799_, _09735_);
  nand _60998_ (_09802_, _09801_, _09679_);
  and _60999_ (_09804_, _09802_, _09677_);
  not _61000_ (_09805_, _09804_);
  and _61001_ (_09807_, _09805_, _09621_);
  or _61002_ (_09808_, _09807_, _09619_);
  or _61003_ (_09810_, _09559_, _09557_);
  and _61004_ (_09811_, _09810_, _09560_);
  nand _61005_ (_09813_, _09811_, _09808_);
  and _61006_ (_09814_, _09813_, _09560_);
  nor _61007_ (_09816_, _09814_, _09493_);
  or _61008_ (_09817_, _09816_, _09492_);
  and _61009_ (_09819_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not _61010_ (_09820_, _09819_);
  nor _61011_ (_09822_, _09820_, _09444_);
  nor _61012_ (_09823_, _09822_, _09476_);
  nor _61013_ (_09825_, _09482_, _09479_);
  nor _61014_ (_09826_, _09825_, _09823_);
  and _61015_ (_09828_, _09825_, _09823_);
  nor _61016_ (_09829_, _09828_, _09826_);
  nor _61017_ (_09830_, _09489_, _09486_);
  not _61018_ (_09831_, _09830_);
  and _61019_ (_09832_, _09831_, _09829_);
  nor _61020_ (_09833_, _09831_, _09829_);
  nor _61021_ (_09834_, _09833_, _09832_);
  and _61022_ (_09835_, _09834_, _09817_);
  or _61023_ (_09836_, _09826_, _09473_);
  or _61024_ (_09837_, _09836_, _09832_);
  or _61025_ (_09838_, _09837_, _09835_);
  or _61026_ (_09839_, _09838_, _09301_);
  and _61027_ (_09840_, _09839_, _06140_);
  and _61028_ (_09841_, _09840_, _09300_);
  not _61029_ (_09842_, _06132_);
  and _61030_ (_09843_, _08587_, _08420_);
  or _61031_ (_09844_, _09843_, _09267_);
  and _61032_ (_09845_, _09844_, _06139_);
  or _61033_ (_09846_, _09845_, _09842_);
  or _61034_ (_09847_, _09846_, _09841_);
  and _61035_ (_09848_, _09847_, _09266_);
  or _61036_ (_09849_, _09848_, _06116_);
  and _61037_ (_09850_, _08535_, _07841_);
  or _61038_ (_09851_, _09263_, _06117_);
  or _61039_ (_09852_, _09851_, _09850_);
  and _61040_ (_09853_, _09852_, _06114_);
  and _61041_ (_09854_, _09853_, _09849_);
  and _61042_ (_09855_, _06294_, _05781_);
  and _61043_ (_09856_, _08782_, _07841_);
  or _61044_ (_09857_, _09856_, _09263_);
  and _61045_ (_09858_, _09857_, _05787_);
  or _61046_ (_09859_, _09858_, _09855_);
  or _61047_ (_09860_, _09859_, _09854_);
  not _61048_ (_09861_, _09855_);
  nor _61049_ (_09862_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor _61050_ (_09863_, _09862_, _09307_);
  not _61051_ (_09864_, \oc8051_golden_model_1.B [1]);
  nor _61052_ (_09865_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor _61053_ (_09866_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and _61054_ (_09867_, _09866_, _09865_);
  and _61055_ (_09868_, _09867_, _09864_);
  nor _61056_ (_09869_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not _61057_ (_09870_, _09869_);
  and _61058_ (_09871_, \oc8051_golden_model_1.B [0], _08430_);
  nor _61059_ (_09872_, _09871_, _09870_);
  and _61060_ (_09873_, _09872_, _09868_);
  and _61061_ (_09874_, _09873_, _09863_);
  or _61062_ (_09875_, _09873_, _08430_);
  not _61063_ (_09876_, \oc8051_golden_model_1.B [4]);
  not _61064_ (_09877_, \oc8051_golden_model_1.B [5]);
  nor _61065_ (_09878_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and _61066_ (_09879_, _09878_, _09877_);
  and _61067_ (_09880_, _09879_, _09876_);
  nor _61068_ (_09881_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.B [2]);
  and _61069_ (_09882_, _09881_, _09880_);
  not _61070_ (_09883_, \oc8051_golden_model_1.ACC [6]);
  and _61071_ (_09884_, \oc8051_golden_model_1.B [0], _09883_);
  nor _61072_ (_09885_, _09884_, _08430_);
  nor _61073_ (_09886_, _09885_, _09864_);
  not _61074_ (_09887_, _09886_);
  and _61075_ (_09888_, _09887_, _09882_);
  nor _61076_ (_09889_, _09888_, _09875_);
  nor _61077_ (_09890_, _09889_, _09874_);
  and _61078_ (_09891_, _09888_, \oc8051_golden_model_1.B [0]);
  nor _61079_ (_09892_, _09891_, _09883_);
  and _61080_ (_09893_, _09892_, _09864_);
  nor _61081_ (_09894_, _09892_, _09864_);
  nor _61082_ (_09895_, _09894_, _09893_);
  nor _61083_ (_09896_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor _61084_ (_09897_, _09896_, _09494_);
  nor _61085_ (_09898_, _09897_, \oc8051_golden_model_1.ACC [4]);
  not _61086_ (_09899_, \oc8051_golden_model_1.B [0]);
  and _61087_ (_09900_, \oc8051_golden_model_1.ACC [4], _09899_);
  nor _61088_ (_09901_, _09900_, \oc8051_golden_model_1.ACC [5]);
  not _61089_ (_09902_, \oc8051_golden_model_1.ACC [4]);
  and _61090_ (_09903_, _09902_, \oc8051_golden_model_1.B [0]);
  nor _61091_ (_09904_, _09903_, _09901_);
  nor _61092_ (_09905_, _09904_, _09898_);
  not _61093_ (_09906_, _09905_);
  and _61094_ (_09907_, _09906_, _09895_);
  nor _61095_ (_09908_, _09890_, \oc8051_golden_model_1.B [2]);
  nor _61096_ (_09909_, _09908_, _09893_);
  not _61097_ (_09910_, _09909_);
  nor _61098_ (_09911_, _09910_, _09907_);
  and _61099_ (_09912_, \oc8051_golden_model_1.B [2], _08430_);
  nor _61100_ (_09913_, _09912_, \oc8051_golden_model_1.B [7]);
  and _61101_ (_09914_, _09913_, _09867_);
  not _61102_ (_09915_, _09914_);
  nor _61103_ (_09916_, _09915_, _09911_);
  nor _61104_ (_09917_, _09916_, _09890_);
  nor _61105_ (_09918_, _09917_, _09874_);
  not _61106_ (_09919_, \oc8051_golden_model_1.B [2]);
  nor _61107_ (_09920_, _09906_, _09895_);
  nor _61108_ (_09921_, _09920_, _09907_);
  not _61109_ (_09922_, _09921_);
  and _61110_ (_09923_, _09922_, _09916_);
  nor _61111_ (_09924_, _09916_, _09892_);
  nor _61112_ (_09925_, _09924_, _09923_);
  and _61113_ (_09926_, _09925_, _09919_);
  nor _61114_ (_09927_, _09925_, _09919_);
  nor _61115_ (_09928_, _09927_, _09926_);
  not _61116_ (_09929_, _09928_);
  not _61117_ (_09930_, \oc8051_golden_model_1.ACC [5]);
  nor _61118_ (_09931_, _09916_, _09930_);
  and _61119_ (_09932_, _09916_, _09897_);
  or _61120_ (_09933_, _09932_, _09931_);
  and _61121_ (_09934_, _09933_, _09864_);
  nor _61122_ (_09935_, _09933_, _09864_);
  nor _61123_ (_09936_, _09935_, _09903_);
  nor _61124_ (_09937_, _09936_, _09934_);
  nor _61125_ (_09938_, _09937_, _09929_);
  nor _61126_ (_09939_, _09918_, \oc8051_golden_model_1.B [3]);
  nor _61127_ (_09940_, _09939_, _09926_);
  not _61128_ (_09941_, _09940_);
  nor _61129_ (_09942_, _09941_, _09938_);
  not _61130_ (_09943_, _09942_);
  and _61131_ (_09944_, \oc8051_golden_model_1.B [3], _08430_);
  not _61132_ (_09945_, _09944_);
  and _61133_ (_09946_, _09945_, _09880_);
  and _61134_ (_09947_, _09946_, _09943_);
  nor _61135_ (_09948_, _09947_, _09918_);
  nor _61136_ (_09949_, _09948_, _09874_);
  nor _61137_ (_09950_, _09949_, \oc8051_golden_model_1.B [4]);
  not _61138_ (_09951_, \oc8051_golden_model_1.B [3]);
  not _61139_ (_09952_, _09947_);
  and _61140_ (_09953_, _09937_, _09929_);
  nor _61141_ (_09954_, _09953_, _09938_);
  nor _61142_ (_09955_, _09954_, _09952_);
  nor _61143_ (_09956_, _09947_, _09925_);
  nor _61144_ (_09957_, _09956_, _09955_);
  and _61145_ (_09958_, _09957_, _09951_);
  nor _61146_ (_09959_, _09957_, _09951_);
  nor _61147_ (_09960_, _09959_, _09958_);
  not _61148_ (_09961_, _09960_);
  nor _61149_ (_09962_, _09947_, _09933_);
  nor _61150_ (_09963_, _09935_, _09934_);
  and _61151_ (_09964_, _09963_, _09903_);
  nor _61152_ (_09965_, _09963_, _09903_);
  nor _61153_ (_09966_, _09965_, _09964_);
  and _61154_ (_09967_, _09966_, _09947_);
  or _61155_ (_09968_, _09967_, _09962_);
  nor _61156_ (_09969_, _09968_, \oc8051_golden_model_1.B [2]);
  and _61157_ (_09970_, _09968_, \oc8051_golden_model_1.B [2]);
  nor _61158_ (_09971_, _09903_, _09900_);
  and _61159_ (_09972_, _09947_, _09971_);
  nor _61160_ (_09973_, _09947_, \oc8051_golden_model_1.ACC [4]);
  nor _61161_ (_09974_, _09973_, _09972_);
  and _61162_ (_09975_, _09974_, _09864_);
  nor _61163_ (_09976_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor _61164_ (_09977_, _09976_, _09680_);
  nor _61165_ (_09978_, _09977_, \oc8051_golden_model_1.ACC [2]);
  and _61166_ (_09979_, _09899_, \oc8051_golden_model_1.ACC [2]);
  nor _61167_ (_09980_, _09979_, \oc8051_golden_model_1.ACC [3]);
  not _61168_ (_09981_, \oc8051_golden_model_1.ACC [2]);
  and _61169_ (_09982_, \oc8051_golden_model_1.B [0], _09981_);
  nor _61170_ (_09983_, _09982_, _09980_);
  nor _61171_ (_09984_, _09983_, _09978_);
  not _61172_ (_09985_, _09984_);
  nor _61173_ (_09986_, _09974_, _09864_);
  nor _61174_ (_09987_, _09986_, _09975_);
  and _61175_ (_09988_, _09987_, _09985_);
  nor _61176_ (_09989_, _09988_, _09975_);
  nor _61177_ (_09990_, _09989_, _09970_);
  nor _61178_ (_09991_, _09990_, _09969_);
  nor _61179_ (_09992_, _09991_, _09961_);
  or _61180_ (_09993_, _09992_, _09958_);
  nor _61181_ (_09994_, _09993_, _09950_);
  and _61182_ (_09995_, _09879_, \oc8051_golden_model_1.ACC [7]);
  or _61183_ (_09996_, _09995_, _09880_);
  not _61184_ (_09997_, _09996_);
  nor _61185_ (_09998_, _09997_, _09994_);
  nor _61186_ (_09999_, _09998_, _09949_);
  nor _61187_ (_10000_, _09999_, _09874_);
  and _61188_ (_10001_, _09991_, _09961_);
  nor _61189_ (_10002_, _10001_, _09992_);
  not _61190_ (_10003_, _10002_);
  and _61191_ (_10004_, _10003_, _09998_);
  nor _61192_ (_10005_, _09998_, _09957_);
  nor _61193_ (_10006_, _10005_, _10004_);
  and _61194_ (_10007_, _10006_, _09876_);
  nor _61195_ (_10008_, _10006_, _09876_);
  nor _61196_ (_10009_, _10008_, _10007_);
  not _61197_ (_10010_, _10009_);
  nor _61198_ (_10011_, _09998_, _09968_);
  nor _61199_ (_10012_, _09970_, _09969_);
  and _61200_ (_10013_, _10012_, _09989_);
  nor _61201_ (_10014_, _10012_, _09989_);
  nor _61202_ (_10015_, _10014_, _10013_);
  not _61203_ (_10016_, _10015_);
  and _61204_ (_10017_, _10016_, _09998_);
  nor _61205_ (_10018_, _10017_, _10011_);
  nor _61206_ (_10019_, _10018_, \oc8051_golden_model_1.B [3]);
  and _61207_ (_10020_, _10018_, \oc8051_golden_model_1.B [3]);
  nor _61208_ (_10021_, _09987_, _09985_);
  nor _61209_ (_10022_, _10021_, _09988_);
  not _61210_ (_10023_, _10022_);
  and _61211_ (_10024_, _10023_, _09998_);
  nor _61212_ (_10025_, _09998_, _09974_);
  nor _61213_ (_10026_, _10025_, _10024_);
  and _61214_ (_10027_, _10026_, _09919_);
  not _61215_ (_10028_, \oc8051_golden_model_1.ACC [3]);
  nor _61216_ (_10029_, _09998_, _10028_);
  and _61217_ (_10030_, _09998_, _09977_);
  or _61218_ (_10031_, _10030_, _10029_);
  and _61219_ (_10032_, _10031_, _09864_);
  nor _61220_ (_10033_, _10031_, _09864_);
  nor _61221_ (_10034_, _10033_, _09982_);
  nor _61222_ (_10035_, _10034_, _10032_);
  nor _61223_ (_10036_, _10026_, _09919_);
  nor _61224_ (_10037_, _10036_, _10027_);
  not _61225_ (_10038_, _10037_);
  nor _61226_ (_10039_, _10038_, _10035_);
  nor _61227_ (_10040_, _10039_, _10027_);
  nor _61228_ (_10041_, _10040_, _10020_);
  nor _61229_ (_10042_, _10041_, _10019_);
  nor _61230_ (_10043_, _10042_, _10010_);
  nor _61231_ (_10044_, _10000_, \oc8051_golden_model_1.B [5]);
  nor _61232_ (_10045_, _10044_, _10007_);
  not _61233_ (_10046_, _10045_);
  nor _61234_ (_10047_, _10046_, _10043_);
  not _61235_ (_10048_, _10047_);
  not _61236_ (_10049_, _09878_);
  and _61237_ (_10050_, \oc8051_golden_model_1.B [5], _08430_);
  nor _61238_ (_10051_, _10050_, _10049_);
  and _61239_ (_10052_, _10051_, _10048_);
  nor _61240_ (_10053_, _10052_, _10000_);
  nor _61241_ (_10054_, _10053_, _09874_);
  not _61242_ (_10055_, _10052_);
  and _61243_ (_10056_, _10042_, _10010_);
  nor _61244_ (_10057_, _10056_, _10043_);
  nor _61245_ (_10058_, _10057_, _10055_);
  nor _61246_ (_10059_, _10052_, _10006_);
  nor _61247_ (_10060_, _10059_, _10058_);
  and _61248_ (_10061_, _10060_, _09877_);
  nor _61249_ (_10062_, _10060_, _09877_);
  nor _61250_ (_10063_, _10062_, _10061_);
  not _61251_ (_10064_, _10063_);
  nor _61252_ (_10065_, _10052_, _10018_);
  nor _61253_ (_10066_, _10020_, _10019_);
  nor _61254_ (_10067_, _10066_, _10040_);
  and _61255_ (_10068_, _10066_, _10040_);
  or _61256_ (_10069_, _10068_, _10067_);
  and _61257_ (_10070_, _10069_, _10052_);
  or _61258_ (_10071_, _10070_, _10065_);
  and _61259_ (_10072_, _10071_, _09876_);
  nor _61260_ (_10073_, _10071_, _09876_);
  and _61261_ (_10074_, _10038_, _10035_);
  nor _61262_ (_10075_, _10074_, _10039_);
  nor _61263_ (_10076_, _10075_, _10055_);
  nor _61264_ (_10077_, _10052_, _10026_);
  nor _61265_ (_10078_, _10077_, _10076_);
  and _61266_ (_10079_, _10078_, _09951_);
  nor _61267_ (_10080_, _10033_, _10032_);
  nor _61268_ (_10081_, _10080_, _09982_);
  and _61269_ (_10082_, _10080_, _09982_);
  or _61270_ (_10083_, _10082_, _10081_);
  nor _61271_ (_10084_, _10083_, _10055_);
  nor _61272_ (_10085_, _10052_, _10031_);
  nor _61273_ (_10086_, _10085_, _10084_);
  and _61274_ (_10087_, _10086_, _09919_);
  nor _61275_ (_10088_, _10086_, _09919_);
  nor _61276_ (_10089_, _09982_, _09979_);
  and _61277_ (_10090_, _10052_, _10089_);
  nor _61278_ (_10091_, _10052_, \oc8051_golden_model_1.ACC [2]);
  nor _61279_ (_10092_, _10091_, _10090_);
  and _61280_ (_10093_, _10092_, _09864_);
  and _61281_ (_10094_, _05887_, \oc8051_golden_model_1.B [0]);
  not _61282_ (_10095_, _10094_);
  nor _61283_ (_10096_, _10092_, _09864_);
  nor _61284_ (_10097_, _10096_, _10093_);
  and _61285_ (_10098_, _10097_, _10095_);
  nor _61286_ (_10099_, _10098_, _10093_);
  nor _61287_ (_10100_, _10099_, _10088_);
  nor _61288_ (_10101_, _10100_, _10087_);
  nor _61289_ (_10102_, _10078_, _09951_);
  nor _61290_ (_10103_, _10102_, _10079_);
  not _61291_ (_10104_, _10103_);
  nor _61292_ (_10105_, _10104_, _10101_);
  nor _61293_ (_10106_, _10105_, _10079_);
  nor _61294_ (_10107_, _10106_, _10073_);
  nor _61295_ (_10108_, _10107_, _10072_);
  nor _61296_ (_10109_, _10108_, _10064_);
  nor _61297_ (_10110_, _10054_, \oc8051_golden_model_1.B [6]);
  or _61298_ (_10111_, _10110_, _10061_);
  or _61299_ (_10112_, _10111_, _10109_);
  and _61300_ (_10113_, \oc8051_golden_model_1.B [6], _08430_);
  nor _61301_ (_10114_, _10113_, \oc8051_golden_model_1.B [7]);
  and _61302_ (_10115_, _10114_, _10112_);
  nor _61303_ (_10116_, _10115_, _10054_);
  or _61304_ (_10117_, _10116_, _09874_);
  nor _61305_ (_10118_, _10117_, \oc8051_golden_model_1.B [7]);
  nor _61306_ (_10119_, _10118_, _09819_);
  not _61307_ (_10120_, \oc8051_golden_model_1.B [6]);
  and _61308_ (_10121_, _10108_, _10064_);
  nor _61309_ (_10122_, _10121_, _10109_);
  not _61310_ (_10123_, _10122_);
  and _61311_ (_10124_, _10123_, _10115_);
  nor _61312_ (_10125_, _10115_, _10060_);
  nor _61313_ (_10126_, _10125_, _10124_);
  nor _61314_ (_10127_, _10126_, _10120_);
  not _61315_ (_10128_, _10127_);
  nor _61316_ (_10129_, _10128_, _10119_);
  nor _61317_ (_10130_, _10088_, _10087_);
  nor _61318_ (_10131_, _10130_, _10099_);
  and _61319_ (_10132_, _10130_, _10099_);
  or _61320_ (_10133_, _10132_, _10131_);
  not _61321_ (_10134_, _10133_);
  and _61322_ (_10135_, _10134_, _10115_);
  nor _61323_ (_10136_, _10115_, _10086_);
  nor _61324_ (_10137_, _10136_, _10135_);
  and _61325_ (_10138_, _10137_, _09951_);
  nor _61326_ (_10139_, _10137_, _09951_);
  nor _61327_ (_10140_, _10139_, _10138_);
  nor _61328_ (_10141_, _10097_, _10095_);
  nor _61329_ (_10142_, _10141_, _10098_);
  and _61330_ (_10143_, _10142_, _10115_);
  not _61331_ (_10144_, _10092_);
  nor _61332_ (_10145_, _10115_, _10144_);
  nor _61333_ (_10146_, _10145_, _10143_);
  and _61334_ (_10147_, _10146_, \oc8051_golden_model_1.B [2]);
  nor _61335_ (_10148_, _10146_, \oc8051_golden_model_1.B [2]);
  nor _61336_ (_10149_, _10148_, _10147_);
  and _61337_ (_10150_, _10149_, _10140_);
  nor _61338_ (_10151_, _10115_, \oc8051_golden_model_1.ACC [1]);
  nor _61339_ (_10152_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  or _61340_ (_10153_, _10152_, _09770_);
  and _61341_ (_10154_, _10115_, _10153_);
  nor _61342_ (_10155_, _10154_, _10151_);
  and _61343_ (_10156_, _10155_, _09864_);
  nor _61344_ (_10157_, _10155_, _09864_);
  and _61345_ (_10158_, _09899_, \oc8051_golden_model_1.ACC [0]);
  not _61346_ (_10159_, _10158_);
  nor _61347_ (_10160_, _10159_, _10157_);
  nor _61348_ (_10161_, _10160_, _10156_);
  and _61349_ (_10162_, _10161_, _10150_);
  not _61350_ (_10163_, _10162_);
  and _61351_ (_10164_, _10147_, _10140_);
  nor _61352_ (_10165_, _10164_, _10139_);
  and _61353_ (_10166_, _10165_, _10163_);
  and _61354_ (_10167_, _10126_, _10120_);
  nor _61355_ (_10168_, _10167_, _10127_);
  not _61356_ (_10169_, _10168_);
  nor _61357_ (_10170_, _10169_, _10119_);
  and _61358_ (_10171_, _10104_, _10101_);
  or _61359_ (_10172_, _10171_, _10105_);
  and _61360_ (_10173_, _10172_, _10115_);
  nor _61361_ (_10174_, _10115_, _10078_);
  nor _61362_ (_10175_, _10174_, _10173_);
  nor _61363_ (_10176_, _10175_, _09876_);
  and _61364_ (_10177_, _10175_, _09876_);
  nor _61365_ (_10178_, _10177_, _10176_);
  nor _61366_ (_10179_, _10073_, _10072_);
  nor _61367_ (_10180_, _10179_, _10106_);
  and _61368_ (_10181_, _10179_, _10106_);
  or _61369_ (_10182_, _10181_, _10180_);
  not _61370_ (_10183_, _10182_);
  and _61371_ (_10184_, _10183_, _10115_);
  nor _61372_ (_10185_, _10115_, _10071_);
  nor _61373_ (_10186_, _10185_, _10184_);
  nor _61374_ (_10187_, _10186_, _09877_);
  and _61375_ (_10188_, _10186_, _09877_);
  nor _61376_ (_10189_, _10188_, _10187_);
  and _61377_ (_10190_, _10189_, _10178_);
  and _61378_ (_10191_, _10190_, _10170_);
  not _61379_ (_10192_, _10191_);
  nor _61380_ (_10193_, _10192_, _10166_);
  and _61381_ (_10194_, _10054_, \oc8051_golden_model_1.B [7]);
  and _61382_ (_10195_, _10189_, _10176_);
  nor _61383_ (_10196_, _10195_, _10187_);
  not _61384_ (_10197_, _10196_);
  and _61385_ (_10198_, _10197_, _10170_);
  or _61386_ (_10199_, _10198_, _10194_);
  or _61387_ (_10200_, _10199_, _10193_);
  nor _61388_ (_10201_, _10200_, _10129_);
  and _61389_ (_10202_, \oc8051_golden_model_1.B [0], _05855_);
  not _61390_ (_10203_, _10202_);
  nor _61391_ (_10204_, _10157_, _10156_);
  and _61392_ (_10205_, _10204_, _10203_);
  and _61393_ (_10206_, _10205_, _10159_);
  and _61394_ (_10207_, _10206_, _10150_);
  and _61395_ (_10208_, _10207_, _10191_);
  nor _61396_ (_10209_, _10208_, _10201_);
  and _61397_ (_10210_, _10209_, _10117_);
  or _61398_ (_10211_, _10210_, _09874_);
  or _61399_ (_10212_, _10211_, _09861_);
  and _61400_ (_10213_, _10212_, _06298_);
  and _61401_ (_10214_, _10213_, _09860_);
  and _61402_ (_10215_, _08802_, _07841_);
  or _61403_ (_10216_, _10215_, _09263_);
  and _61404_ (_10217_, _10216_, _06297_);
  and _61405_ (_10218_, _08607_, _07841_);
  or _61406_ (_10219_, _10218_, _09263_);
  and _61407_ (_10220_, _10219_, _06110_);
  or _61408_ (_10221_, _10220_, _06402_);
  or _61409_ (_10222_, _10221_, _10217_);
  or _61410_ (_10223_, _10222_, _10214_);
  and _61411_ (_10224_, _08810_, _07841_);
  or _61412_ (_10225_, _09263_, _07125_);
  or _61413_ (_10226_, _10225_, _10224_);
  and _61414_ (_10227_, _10226_, _07132_);
  and _61415_ (_10228_, _10227_, _10223_);
  or _61416_ (_10229_, _09263_, _07926_);
  and _61417_ (_10230_, _10219_, _06306_);
  and _61418_ (_10231_, _10230_, _10229_);
  or _61419_ (_10232_, _10231_, _10228_);
  and _61420_ (_10233_, _10232_, _07130_);
  and _61421_ (_10234_, _09275_, _06411_);
  and _61422_ (_10235_, _10234_, _10229_);
  or _61423_ (_10236_, _10235_, _06303_);
  or _61424_ (_10237_, _10236_, _10233_);
  and _61425_ (_10238_, _08801_, _07841_);
  or _61426_ (_10239_, _09263_, _08819_);
  or _61427_ (_10240_, _10239_, _10238_);
  and _61428_ (_10241_, _10240_, _08824_);
  and _61429_ (_10242_, _10241_, _10237_);
  not _61430_ (_10243_, _07841_);
  nor _61431_ (_10244_, _08809_, _10243_);
  or _61432_ (_10245_, _10244_, _09263_);
  and _61433_ (_10246_, _10245_, _06396_);
  or _61434_ (_10247_, _10246_, _06433_);
  or _61435_ (_10248_, _10247_, _10242_);
  or _61436_ (_10249_, _09272_, _06829_);
  and _61437_ (_10250_, _10249_, _05749_);
  and _61438_ (_10251_, _10250_, _10248_);
  and _61439_ (_10252_, _09269_, _05748_);
  or _61440_ (_10253_, _10252_, _06440_);
  or _61441_ (_10254_, _10253_, _10251_);
  and _61442_ (_10255_, _08345_, _07841_);
  or _61443_ (_10256_, _09263_, _06444_);
  or _61444_ (_10257_, _10256_, _10255_);
  and _61445_ (_10258_, _10257_, _01317_);
  and _61446_ (_10259_, _10258_, _10254_);
  or _61447_ (_10260_, _10259_, _09262_);
  and _61448_ (_40980_, _10260_, _43100_);
  nor _61449_ (_10261_, _01317_, _08430_);
  and _61450_ (_10262_, _05825_, _06302_);
  nand _61451_ (_10263_, _10262_, _09883_);
  and _61452_ (_10264_, _06294_, _05825_);
  not _61453_ (_10265_, _10264_);
  nor _61454_ (_10266_, _08014_, _09883_);
  not _61455_ (_10267_, _10266_);
  nor _61456_ (_10268_, _08103_, _09930_);
  and _61457_ (_10269_, _08103_, _09930_);
  nor _61458_ (_10270_, _08338_, _09902_);
  not _61459_ (_10271_, _10270_);
  nor _61460_ (_10272_, _08139_, _10028_);
  and _61461_ (_10273_, _08139_, _10028_);
  nor _61462_ (_10274_, _08247_, _09981_);
  nor _61463_ (_10275_, _08175_, _05887_);
  and _61464_ (_10276_, _08211_, \oc8051_golden_model_1.ACC [0]);
  and _61465_ (_10277_, _08175_, _05887_);
  nor _61466_ (_10278_, _10277_, _10275_);
  and _61467_ (_10279_, _10278_, _10276_);
  nor _61468_ (_10280_, _10279_, _10275_);
  and _61469_ (_10281_, _08247_, _09981_);
  nor _61470_ (_10282_, _10281_, _10274_);
  not _61471_ (_10283_, _10282_);
  nor _61472_ (_10284_, _10283_, _10280_);
  nor _61473_ (_10285_, _10284_, _10274_);
  nor _61474_ (_10286_, _10285_, _10273_);
  or _61475_ (_10287_, _10286_, _10272_);
  and _61476_ (_10288_, _08338_, _09902_);
  nor _61477_ (_10289_, _10288_, _10270_);
  nand _61478_ (_10290_, _10289_, _10287_);
  and _61479_ (_10291_, _10290_, _10271_);
  nor _61480_ (_10292_, _10291_, _10269_);
  or _61481_ (_10293_, _10292_, _10268_);
  and _61482_ (_10294_, _08014_, _09883_);
  nor _61483_ (_10295_, _10294_, _10266_);
  nand _61484_ (_10296_, _10295_, _10293_);
  and _61485_ (_10297_, _10296_, _10267_);
  nor _61486_ (_10298_, _10297_, _08810_);
  and _61487_ (_10299_, _10297_, _08810_);
  or _61488_ (_10300_, _10299_, _10298_);
  and _61489_ (_10301_, _10300_, _06169_);
  and _61490_ (_10302_, _09200_, \oc8051_golden_model_1.PSW [7]);
  nor _61491_ (_10303_, _10302_, _09194_);
  and _61492_ (_10304_, _10302_, _09194_);
  nor _61493_ (_10305_, _10304_, _10303_);
  and _61494_ (_10306_, _10305_, \oc8051_golden_model_1.ACC [7]);
  nor _61495_ (_10307_, _10305_, \oc8051_golden_model_1.ACC [7]);
  nor _61496_ (_10308_, _10307_, _10306_);
  and _61497_ (_10309_, _09199_, \oc8051_golden_model_1.PSW [7]);
  nor _61498_ (_10310_, _10309_, _08012_);
  nor _61499_ (_10311_, _10310_, _10302_);
  nand _61500_ (_10312_, _10311_, \oc8051_golden_model_1.ACC [6]);
  nor _61501_ (_10313_, _10311_, _09883_);
  and _61502_ (_10314_, _10311_, _09883_);
  nor _61503_ (_10315_, _10314_, _10313_);
  not _61504_ (_10316_, _10315_);
  and _61505_ (_10317_, _09198_, \oc8051_golden_model_1.PSW [7]);
  nor _61506_ (_10318_, _10317_, _08101_);
  nor _61507_ (_10319_, _10318_, _10309_);
  and _61508_ (_10320_, _10319_, \oc8051_golden_model_1.ACC [5]);
  nor _61509_ (_10321_, _10319_, _09930_);
  and _61510_ (_10322_, _10319_, _09930_);
  nor _61511_ (_10323_, _10322_, _10321_);
  and _61512_ (_10324_, _09197_, \oc8051_golden_model_1.PSW [7]);
  nor _61513_ (_10325_, _10324_, _08336_);
  nor _61514_ (_10326_, _10325_, _10317_);
  nand _61515_ (_10327_, _10326_, \oc8051_golden_model_1.ACC [4]);
  nor _61516_ (_10328_, _10326_, _09902_);
  and _61517_ (_10329_, _10326_, _09902_);
  or _61518_ (_10330_, _10329_, _10328_);
  and _61519_ (_10331_, _09196_, \oc8051_golden_model_1.PSW [7]);
  nor _61520_ (_10332_, _10331_, _07544_);
  nor _61521_ (_10333_, _10332_, _10324_);
  and _61522_ (_10334_, _10333_, \oc8051_golden_model_1.ACC [3]);
  nor _61523_ (_10335_, _10333_, _10028_);
  and _61524_ (_10336_, _10333_, _10028_);
  nor _61525_ (_10337_, _10336_, _10335_);
  and _61526_ (_10338_, _09195_, \oc8051_golden_model_1.PSW [7]);
  nor _61527_ (_10339_, _10338_, _07708_);
  nor _61528_ (_10340_, _10339_, _10331_);
  and _61529_ (_10341_, _10340_, \oc8051_golden_model_1.ACC [2]);
  nor _61530_ (_10342_, _10340_, _09981_);
  and _61531_ (_10343_, _10340_, _09981_);
  nor _61532_ (_10344_, _10343_, _10342_);
  and _61533_ (_10345_, _07049_, \oc8051_golden_model_1.PSW [7]);
  nor _61534_ (_10346_, _10345_, _07306_);
  nor _61535_ (_10347_, _10346_, _10338_);
  and _61536_ (_10348_, _10347_, \oc8051_golden_model_1.ACC [1]);
  and _61537_ (_10349_, _10347_, _05887_);
  nor _61538_ (_10350_, _10347_, _05887_);
  nor _61539_ (_10351_, _10350_, _10349_);
  not _61540_ (_10352_, _10351_);
  nor _61541_ (_10353_, _07049_, \oc8051_golden_model_1.PSW [7]);
  nor _61542_ (_10354_, _10353_, _10345_);
  and _61543_ (_10355_, _10354_, \oc8051_golden_model_1.ACC [0]);
  and _61544_ (_10356_, _10355_, _10352_);
  nor _61545_ (_10357_, _10356_, _10348_);
  nor _61546_ (_10358_, _10357_, _10344_);
  nor _61547_ (_10359_, _10358_, _10341_);
  nor _61548_ (_10360_, _10359_, _10337_);
  or _61549_ (_10361_, _10360_, _10334_);
  nand _61550_ (_10362_, _10361_, _10330_);
  and _61551_ (_10363_, _10362_, _10327_);
  nor _61552_ (_10364_, _10363_, _10323_);
  or _61553_ (_10365_, _10364_, _10320_);
  nand _61554_ (_10366_, _10365_, _10316_);
  and _61555_ (_10367_, _10366_, _10312_);
  nor _61556_ (_10368_, _10367_, _10308_);
  and _61557_ (_10369_, _10367_, _10308_);
  nor _61558_ (_10370_, _10369_, _10368_);
  and _61559_ (_10371_, _06123_, _06300_);
  nor _61560_ (_10372_, _10371_, _06523_);
  and _61561_ (_10373_, _06119_, _06300_);
  not _61562_ (_10374_, _10373_);
  not _61563_ (_10375_, _06794_);
  and _61564_ (_10376_, _06957_, _06300_);
  nor _61565_ (_10377_, _10376_, _06795_);
  and _61566_ (_10378_, _10377_, _10375_);
  and _61567_ (_10379_, _10378_, _10374_);
  and _61568_ (_10380_, _10379_, _10372_);
  or _61569_ (_10381_, _10380_, _10370_);
  or _61570_ (_10382_, _06039_, _05802_);
  nor _61571_ (_10383_, _07809_, _08430_);
  and _61572_ (_10384_, _07923_, _07809_);
  or _61573_ (_10385_, _10384_, _10383_);
  or _61574_ (_10386_, _10385_, _06132_);
  and _61575_ (_10387_, _06294_, _05790_);
  not _61576_ (_10388_, _10387_);
  and _61577_ (_10389_, _08211_, \oc8051_golden_model_1.PSW [7]);
  and _61578_ (_10390_, _10389_, _08176_);
  and _61579_ (_10391_, _10390_, _08248_);
  and _61580_ (_10392_, _10391_, _08140_);
  and _61581_ (_10393_, _10392_, _08339_);
  and _61582_ (_10394_, _10393_, _08104_);
  and _61583_ (_10395_, _10394_, _08015_);
  nor _61584_ (_10396_, _10395_, _07925_);
  and _61585_ (_10397_, _10395_, _07925_);
  nor _61586_ (_10398_, _10397_, _10396_);
  and _61587_ (_10399_, _10398_, \oc8051_golden_model_1.ACC [7]);
  nor _61588_ (_10400_, _10398_, \oc8051_golden_model_1.ACC [7]);
  nor _61589_ (_10401_, _10400_, _10399_);
  not _61590_ (_10402_, _10401_);
  nor _61591_ (_10403_, _10394_, _08015_);
  nor _61592_ (_10404_, _10403_, _10395_);
  nor _61593_ (_10405_, _10404_, _09883_);
  nor _61594_ (_10406_, _10393_, _08104_);
  nor _61595_ (_10407_, _10406_, _10394_);
  nor _61596_ (_10408_, _10407_, _09930_);
  and _61597_ (_10409_, _10407_, _09930_);
  nor _61598_ (_10410_, _10409_, _10408_);
  not _61599_ (_10411_, _10410_);
  nor _61600_ (_10412_, _10392_, _08339_);
  nor _61601_ (_10413_, _10412_, _10393_);
  nor _61602_ (_10414_, _10413_, _09902_);
  and _61603_ (_10415_, _10413_, _09902_);
  or _61604_ (_10416_, _10415_, _10414_);
  or _61605_ (_10417_, _10416_, _10411_);
  nor _61606_ (_10418_, _10391_, _08140_);
  nor _61607_ (_10419_, _10418_, _10392_);
  nor _61608_ (_10420_, _10419_, _10028_);
  and _61609_ (_10421_, _10419_, _10028_);
  nor _61610_ (_10422_, _10421_, _10420_);
  nor _61611_ (_10423_, _10390_, _08248_);
  nor _61612_ (_10424_, _10423_, _10391_);
  nor _61613_ (_10425_, _10424_, _09981_);
  and _61614_ (_10426_, _10424_, _09981_);
  nor _61615_ (_10427_, _10426_, _10425_);
  and _61616_ (_10428_, _10427_, _10422_);
  nor _61617_ (_10429_, _10389_, _08176_);
  nor _61618_ (_10430_, _10429_, _10390_);
  nor _61619_ (_10431_, _10430_, _05887_);
  and _61620_ (_10432_, _10430_, _05887_);
  nor _61621_ (_10433_, _08211_, \oc8051_golden_model_1.PSW [7]);
  nor _61622_ (_10434_, _10433_, _10389_);
  and _61623_ (_10435_, _10434_, _05855_);
  nor _61624_ (_10436_, _10435_, _10432_);
  or _61625_ (_10437_, _10436_, _10431_);
  nand _61626_ (_10438_, _10437_, _10428_);
  nor _61627_ (_10439_, _10425_, _10420_);
  or _61628_ (_10440_, _10439_, _10421_);
  and _61629_ (_10441_, _10440_, _10438_);
  nor _61630_ (_10442_, _10441_, _10417_);
  nor _61631_ (_10443_, _10414_, _10408_);
  nor _61632_ (_10444_, _10443_, _10409_);
  nor _61633_ (_10445_, _10444_, _10442_);
  and _61634_ (_10446_, _10404_, _09883_);
  nor _61635_ (_10447_, _10405_, _10446_);
  not _61636_ (_10448_, _10447_);
  nor _61637_ (_10449_, _10448_, _10445_);
  or _61638_ (_10450_, _10449_, _10405_);
  and _61639_ (_10451_, _10450_, _10402_);
  nor _61640_ (_10452_, _10450_, _10402_);
  or _61641_ (_10453_, _10452_, _10451_);
  or _61642_ (_10454_, _10453_, _06265_);
  and _61643_ (_10455_, _10454_, _10388_);
  not _61644_ (_10456_, _06529_);
  nor _61645_ (_10457_, _07678_, _06538_);
  and _61646_ (_10458_, _10457_, _10456_);
  or _61647_ (_10459_, _10458_, _07923_);
  nor _61648_ (_10460_, _08409_, _08430_);
  and _61649_ (_10461_, _08552_, _08409_);
  or _61650_ (_10462_, _10461_, _10460_);
  or _61651_ (_10463_, _10462_, _06157_);
  and _61652_ (_10464_, _10463_, _07075_);
  not _61653_ (_10465_, _06658_);
  nor _61654_ (_10466_, _06119_, _06284_);
  nor _61655_ (_10467_, _10466_, _05771_);
  nor _61656_ (_10468_, _10467_, _10465_);
  nor _61657_ (_10469_, _06129_, _05771_);
  not _61658_ (_10470_, _10469_);
  and _61659_ (_10471_, _10470_, _10468_);
  or _61660_ (_10472_, _10471_, _07923_);
  and _61661_ (_10473_, _06294_, _06222_);
  not _61662_ (_10474_, _10473_);
  nor _61663_ (_10475_, _06653_, _08430_);
  and _61664_ (_10476_, _06653_, _08430_);
  nor _61665_ (_10477_, _10476_, _10475_);
  nand _61666_ (_10478_, _10477_, _10471_);
  and _61667_ (_10479_, _10478_, _10474_);
  and _61668_ (_10480_, _10479_, _10472_);
  and _61669_ (_10481_, _10473_, _08535_);
  or _61670_ (_10482_, _10481_, _10480_);
  not _61671_ (_10483_, _05772_);
  nor _61672_ (_10484_, _06160_, _10483_);
  and _61673_ (_10485_, _10484_, _10482_);
  and _61674_ (_10486_, _08548_, _07809_);
  or _61675_ (_10487_, _10486_, _10383_);
  and _61676_ (_10488_, _10487_, _06160_);
  or _61677_ (_10489_, _10488_, _10485_);
  and _61678_ (_10490_, _06294_, _06155_);
  not _61679_ (_10491_, _10490_);
  and _61680_ (_10492_, _10491_, _10489_);
  nor _61681_ (_10493_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor _61682_ (_10494_, _10493_, _10028_);
  and _61683_ (_10495_, _10494_, \oc8051_golden_model_1.ACC [4]);
  and _61684_ (_10496_, _10495_, \oc8051_golden_model_1.ACC [5]);
  and _61685_ (_10497_, _10496_, \oc8051_golden_model_1.ACC [6]);
  and _61686_ (_10498_, _10497_, \oc8051_golden_model_1.ACC [7]);
  nor _61687_ (_10499_, _10497_, \oc8051_golden_model_1.ACC [7]);
  nor _61688_ (_10500_, _10499_, _10498_);
  nor _61689_ (_10501_, _10495_, \oc8051_golden_model_1.ACC [5]);
  nor _61690_ (_10502_, _10501_, _10496_);
  nor _61691_ (_10503_, _10496_, \oc8051_golden_model_1.ACC [6]);
  nor _61692_ (_10504_, _10503_, _10497_);
  nor _61693_ (_10505_, _10504_, _10502_);
  not _61694_ (_10506_, _10505_);
  and _61695_ (_10507_, _10506_, _10500_);
  or _61696_ (_10508_, _10498_, \oc8051_golden_model_1.PSW [7]);
  and _61697_ (_10509_, _10508_, _10506_);
  nor _61698_ (_10510_, _10509_, _10500_);
  nor _61699_ (_10511_, _10510_, _10507_);
  and _61700_ (_10512_, _10511_, _10490_);
  or _61701_ (_10513_, _10512_, _06156_);
  or _61702_ (_10514_, _10513_, _10492_);
  and _61703_ (_10515_, _10514_, _10464_);
  not _61704_ (_10516_, _10458_);
  and _61705_ (_10517_, _10385_, _06217_);
  or _61706_ (_10518_, _10517_, _10516_);
  or _61707_ (_10519_, _10518_, _10515_);
  and _61708_ (_10520_, _10519_, _10459_);
  or _61709_ (_10521_, _10520_, _07081_);
  or _61710_ (_10522_, _08535_, _07082_);
  and _61711_ (_10523_, _10522_, _06229_);
  and _61712_ (_10524_, _10523_, _10521_);
  and _61713_ (_10525_, _06294_, _06150_);
  nor _61714_ (_10526_, _07925_, _06229_);
  or _61715_ (_10527_, _10526_, _10525_);
  or _61716_ (_10528_, _10527_, _10524_);
  nand _61717_ (_10529_, _10525_, _10028_);
  and _61718_ (_10530_, _10529_, _10528_);
  or _61719_ (_10531_, _10530_, _06152_);
  and _61720_ (_10532_, _08426_, _08409_);
  or _61721_ (_10533_, _10532_, _10460_);
  or _61722_ (_10534_, _10533_, _06153_);
  and _61723_ (_10535_, _10534_, _06146_);
  and _61724_ (_10536_, _10535_, _10531_);
  or _61725_ (_10537_, _10460_, _08568_);
  and _61726_ (_10538_, _10462_, _06145_);
  and _61727_ (_10539_, _10538_, _10537_);
  or _61728_ (_10540_, _10539_, _09295_);
  or _61729_ (_10541_, _10540_, _10536_);
  nor _61730_ (_10542_, _09789_, _09787_);
  nor _61731_ (_10543_, _10542_, _09790_);
  or _61732_ (_10544_, _10543_, _09301_);
  and _61733_ (_10545_, _06273_, _05790_);
  not _61734_ (_10546_, _10545_);
  and _61735_ (_10547_, _06125_, _05790_);
  nor _61736_ (_10548_, _10547_, _06536_);
  and _61737_ (_10549_, _06118_, _05790_);
  or _61738_ (_10550_, _06971_, _06276_);
  and _61739_ (_10551_, _10550_, _10549_);
  not _61740_ (_10552_, _10551_);
  and _61741_ (_10553_, _10552_, _10548_);
  and _61742_ (_10554_, _10553_, _10546_);
  and _61743_ (_10555_, _10554_, _10544_);
  and _61744_ (_10556_, _10555_, _10541_);
  not _61745_ (_10557_, _10554_);
  not _61746_ (_10558_, _10308_);
  not _61747_ (_10559_, _10323_);
  or _61748_ (_10560_, _10330_, _10559_);
  and _61749_ (_10561_, _10344_, _10337_);
  and _61750_ (_10562_, _10354_, _05855_);
  nor _61751_ (_10563_, _10562_, _10349_);
  or _61752_ (_10564_, _10563_, _10350_);
  nand _61753_ (_10565_, _10564_, _10561_);
  nor _61754_ (_10566_, _10342_, _10335_);
  or _61755_ (_10567_, _10566_, _10336_);
  and _61756_ (_10568_, _10567_, _10565_);
  nor _61757_ (_10569_, _10568_, _10560_);
  nor _61758_ (_10570_, _10328_, _10321_);
  nor _61759_ (_10571_, _10570_, _10322_);
  nor _61760_ (_10572_, _10571_, _10569_);
  nor _61761_ (_10573_, _10572_, _10316_);
  or _61762_ (_10574_, _10573_, _10313_);
  and _61763_ (_10575_, _10574_, _10558_);
  nor _61764_ (_10576_, _10574_, _10558_);
  or _61765_ (_10577_, _10576_, _10575_);
  and _61766_ (_10578_, _10577_, _10557_);
  or _61767_ (_10579_, _10578_, _10556_);
  and _61768_ (_10580_, _06284_, _05790_);
  not _61769_ (_10581_, _10580_);
  and _61770_ (_10582_, _10581_, _10579_);
  and _61771_ (_10583_, _09217_, \oc8051_golden_model_1.PSW [7]);
  nor _61772_ (_10584_, _10583_, _08838_);
  and _61773_ (_10585_, _10583_, _08838_);
  nor _61774_ (_10586_, _10585_, _10584_);
  and _61775_ (_10587_, _10586_, \oc8051_golden_model_1.ACC [7]);
  nor _61776_ (_10588_, _10586_, \oc8051_golden_model_1.ACC [7]);
  nor _61777_ (_10589_, _10588_, _10587_);
  and _61778_ (_10590_, _09216_, \oc8051_golden_model_1.PSW [7]);
  nor _61779_ (_10591_, _10590_, _09207_);
  nor _61780_ (_10592_, _10591_, _10583_);
  nor _61781_ (_10593_, _10592_, _09883_);
  and _61782_ (_10594_, _09215_, \oc8051_golden_model_1.PSW [7]);
  nor _61783_ (_10595_, _10594_, _09208_);
  nor _61784_ (_10596_, _10595_, _10590_);
  nor _61785_ (_10597_, _10596_, _09930_);
  and _61786_ (_10598_, _10596_, _09930_);
  nor _61787_ (_10599_, _10598_, _10597_);
  not _61788_ (_10600_, _10599_);
  and _61789_ (_10601_, _09214_, \oc8051_golden_model_1.PSW [7]);
  nor _61790_ (_10602_, _10601_, _09209_);
  nor _61791_ (_10603_, _10602_, _10594_);
  nor _61792_ (_10604_, _10603_, _09902_);
  and _61793_ (_10605_, _10603_, _09902_);
  or _61794_ (_10606_, _10605_, _10604_);
  or _61795_ (_10607_, _10606_, _10600_);
  and _61796_ (_10608_, _09213_, \oc8051_golden_model_1.PSW [7]);
  nor _61797_ (_10609_, _10608_, _09210_);
  nor _61798_ (_10610_, _10609_, _10601_);
  nor _61799_ (_10611_, _10610_, _10028_);
  and _61800_ (_10612_, _10610_, _10028_);
  nor _61801_ (_10613_, _10612_, _10611_);
  and _61802_ (_10614_, _09212_, \oc8051_golden_model_1.PSW [7]);
  nor _61803_ (_10615_, _10614_, _09211_);
  nor _61804_ (_10616_, _10615_, _10608_);
  nor _61805_ (_10617_, _10616_, _09981_);
  and _61806_ (_10618_, _10616_, _09981_);
  nor _61807_ (_10619_, _10618_, _10617_);
  and _61808_ (_10620_, _10619_, _10613_);
  and _61809_ (_10621_, _09160_, \oc8051_golden_model_1.PSW [7]);
  nor _61810_ (_10622_, _10621_, _09115_);
  nor _61811_ (_10623_, _10622_, _10614_);
  nor _61812_ (_10624_, _10623_, _05887_);
  and _61813_ (_10625_, _10623_, _05887_);
  nor _61814_ (_10626_, _09160_, \oc8051_golden_model_1.PSW [7]);
  nor _61815_ (_10627_, _10626_, _10621_);
  and _61816_ (_10628_, _10627_, _05855_);
  nor _61817_ (_10629_, _10628_, _10625_);
  or _61818_ (_10630_, _10629_, _10624_);
  nand _61819_ (_10631_, _10630_, _10620_);
  nor _61820_ (_10632_, _10617_, _10611_);
  or _61821_ (_10633_, _10632_, _10612_);
  and _61822_ (_10634_, _10633_, _10631_);
  nor _61823_ (_10635_, _10634_, _10607_);
  nor _61824_ (_10636_, _10604_, _10597_);
  nor _61825_ (_10637_, _10636_, _10598_);
  nor _61826_ (_10638_, _10637_, _10635_);
  and _61827_ (_10639_, _10592_, _09883_);
  nor _61828_ (_10640_, _10593_, _10639_);
  not _61829_ (_10641_, _10640_);
  nor _61830_ (_10642_, _10641_, _10638_);
  or _61831_ (_10643_, _10642_, _10593_);
  nor _61832_ (_10644_, _10643_, _10589_);
  and _61833_ (_10645_, _10643_, _10589_);
  or _61834_ (_10646_, _10645_, _10644_);
  nor _61835_ (_10647_, _10646_, _10581_);
  or _61836_ (_10648_, _10647_, _10582_);
  and _61837_ (_10649_, _10648_, _06710_);
  nor _61838_ (_10650_, _10646_, _06710_);
  or _61839_ (_10651_, _10650_, _10649_);
  or _61840_ (_10652_, _10651_, _06260_);
  and _61841_ (_10653_, _10652_, _10455_);
  and _61842_ (_10654_, _08586_, _06228_);
  and _61843_ (_10655_, _10654_, _07839_);
  and _61844_ (_10656_, _10654_, _07828_);
  and _61845_ (_10657_, _10656_, _07482_);
  nor _61846_ (_10658_, _10657_, _06039_);
  nor _61847_ (_10659_, _10658_, _10655_);
  nor _61848_ (_10660_, _10659_, _08430_);
  and _61849_ (_10661_, _10659_, _08430_);
  nor _61850_ (_10662_, _10661_, _10660_);
  nor _61851_ (_10663_, _10656_, _07482_);
  nor _61852_ (_10664_, _10663_, _10657_);
  nor _61853_ (_10665_, _10664_, _09883_);
  and _61854_ (_10666_, _10654_, _07775_);
  nor _61855_ (_10667_, _10666_, _07805_);
  nor _61856_ (_10668_, _10667_, _10656_);
  and _61857_ (_10669_, _10668_, _09930_);
  nor _61858_ (_10670_, _10668_, _09930_);
  nor _61859_ (_10671_, _10654_, _07775_);
  nor _61860_ (_10672_, _10671_, _10666_);
  nor _61861_ (_10673_, _10672_, _09902_);
  nor _61862_ (_10674_, _10673_, _10670_);
  nor _61863_ (_10675_, _10674_, _10669_);
  nor _61864_ (_10676_, _10670_, _10669_);
  not _61865_ (_10677_, _10676_);
  and _61866_ (_10678_, _10672_, _09902_);
  or _61867_ (_10679_, _10678_, _10673_);
  or _61868_ (_10680_, _10679_, _10677_);
  nor _61869_ (_10681_, _08586_, _06228_);
  nor _61870_ (_10682_, _10681_, _10654_);
  and _61871_ (_10683_, _10682_, _10028_);
  nor _61872_ (_10684_, _10682_, _10028_);
  nor _61873_ (_10685_, _10684_, _10683_);
  and _61874_ (_10686_, _07834_, \oc8051_golden_model_1.PSW [7]);
  nor _61875_ (_10687_, _10686_, _06626_);
  nor _61876_ (_10688_, _10687_, _08586_);
  and _61877_ (_10689_, _10688_, _09981_);
  nor _61878_ (_10690_, _10688_, _09981_);
  nor _61879_ (_10691_, _10690_, _10689_);
  and _61880_ (_10692_, _10691_, _10685_);
  not _61881_ (_10693_, \oc8051_golden_model_1.PSW [7]);
  nor _61882_ (_10694_, _06107_, _10693_);
  nor _61883_ (_10695_, _10694_, _06913_);
  nor _61884_ (_10696_, _10695_, _10686_);
  nor _61885_ (_10697_, _10696_, _05887_);
  and _61886_ (_10699_, _10696_, _05887_);
  and _61887_ (_10700_, _06107_, _10693_);
  nor _61888_ (_10701_, _10700_, _10694_);
  and _61889_ (_10702_, _10701_, _05855_);
  nor _61890_ (_10703_, _10702_, _10699_);
  or _61891_ (_10704_, _10703_, _10697_);
  nand _61892_ (_10705_, _10704_, _10692_);
  and _61893_ (_10706_, _10690_, _10685_);
  nor _61894_ (_10707_, _10706_, _10684_);
  and _61895_ (_10708_, _10707_, _10705_);
  nor _61896_ (_10710_, _10708_, _10680_);
  nor _61897_ (_10711_, _10710_, _10675_);
  and _61898_ (_10712_, _10664_, _09883_);
  nor _61899_ (_10713_, _10665_, _10712_);
  not _61900_ (_10714_, _10713_);
  nor _61901_ (_10715_, _10714_, _10711_);
  or _61902_ (_10716_, _10715_, _10665_);
  nor _61903_ (_10717_, _10716_, _10662_);
  and _61904_ (_10718_, _10716_, _10662_);
  or _61905_ (_10719_, _10718_, _10717_);
  nor _61906_ (_10721_, _10719_, _10388_);
  or _61907_ (_10722_, _10721_, _10653_);
  and _61908_ (_10723_, _10722_, _05805_);
  and _61909_ (_10724_, _06039_, _05870_);
  or _61910_ (_10725_, _10724_, _10723_);
  and _61911_ (_10726_, _10725_, _06140_);
  and _61912_ (_10727_, _08587_, _08409_);
  or _61913_ (_10728_, _10727_, _10460_);
  and _61914_ (_10729_, _10728_, _06139_);
  or _61915_ (_10730_, _10729_, _09842_);
  or _61916_ (_10732_, _10730_, _10726_);
  and _61917_ (_10733_, _10732_, _10386_);
  or _61918_ (_10734_, _10733_, _06116_);
  and _61919_ (_10735_, _08535_, _07809_);
  or _61920_ (_10736_, _10383_, _06117_);
  or _61921_ (_10737_, _10736_, _10735_);
  and _61922_ (_10738_, _10737_, _06114_);
  and _61923_ (_10739_, _10738_, _10734_);
  and _61924_ (_10740_, _08782_, _07809_);
  or _61925_ (_10741_, _10740_, _10383_);
  and _61926_ (_10743_, _10741_, _05787_);
  or _61927_ (_10744_, _10743_, _09855_);
  or _61928_ (_10745_, _10744_, _10739_);
  or _61929_ (_10746_, _09873_, _09861_);
  and _61930_ (_10747_, _10746_, _10745_);
  or _61931_ (_10748_, _10747_, _05801_);
  and _61932_ (_10749_, _10748_, _10382_);
  or _61933_ (_10750_, _10749_, _06110_);
  and _61934_ (_10751_, _06294_, _06109_);
  not _61935_ (_10752_, _10751_);
  and _61936_ (_10754_, _08607_, _07809_);
  or _61937_ (_10755_, _10754_, _10383_);
  or _61938_ (_10756_, _10755_, _06111_);
  and _61939_ (_10757_, _10756_, _10752_);
  and _61940_ (_10758_, _10757_, _10750_);
  and _61941_ (_10759_, _10751_, _06039_);
  or _61942_ (_10760_, _10759_, _06558_);
  or _61943_ (_10761_, _10760_, _10758_);
  not _61944_ (_10762_, _06558_);
  and _61945_ (_10763_, _09194_, _08430_);
  and _61946_ (_10765_, _07923_, \oc8051_golden_model_1.ACC [7]);
  nor _61947_ (_10766_, _10765_, _10763_);
  nor _61948_ (_10767_, _10766_, _10762_);
  nor _61949_ (_10768_, _06129_, _05833_);
  nor _61950_ (_10769_, _10768_, _10767_);
  and _61951_ (_10770_, _10769_, _10761_);
  and _61952_ (_10771_, _10768_, _10766_);
  and _61953_ (_10772_, _06119_, _06399_);
  or _61954_ (_10773_, _10772_, _10771_);
  or _61955_ (_10774_, _10773_, _10770_);
  and _61956_ (_10775_, _06115_, _06399_);
  not _61957_ (_10776_, _10775_);
  nand _61958_ (_10777_, _10776_, _10766_);
  nor _61959_ (_10778_, _07365_, _05833_);
  nand _61960_ (_10779_, _10778_, _10777_);
  and _61961_ (_10780_, _10779_, _10774_);
  and _61962_ (_10781_, _08838_, _08430_);
  and _61963_ (_10782_, _08535_, \oc8051_golden_model_1.ACC [7]);
  nor _61964_ (_10783_, _10782_, _10781_);
  and _61965_ (_10784_, _10775_, _10783_);
  or _61966_ (_10785_, _10784_, _06400_);
  or _61967_ (_10786_, _10785_, _10780_);
  and _61968_ (_10787_, _06294_, _06399_);
  not _61969_ (_10788_, _10787_);
  or _61970_ (_10789_, _08810_, _06401_);
  and _61971_ (_10790_, _10789_, _10788_);
  and _61972_ (_10791_, _10790_, _10786_);
  nor _61973_ (_10792_, _06039_, \oc8051_golden_model_1.ACC [7]);
  and _61974_ (_10793_, _06039_, \oc8051_golden_model_1.ACC [7]);
  nor _61975_ (_10794_, _10793_, _10792_);
  and _61976_ (_10795_, _10787_, _10794_);
  or _61977_ (_10796_, _10795_, _06297_);
  or _61978_ (_10797_, _10796_, _10791_);
  and _61979_ (_10798_, _08802_, _07809_);
  or _61980_ (_10799_, _10798_, _10383_);
  or _61981_ (_10800_, _10799_, _07127_);
  and _61982_ (_10801_, _10800_, _10797_);
  or _61983_ (_10802_, _10801_, _06402_);
  or _61984_ (_10803_, _10383_, _07125_);
  nor _61985_ (_10804_, _06129_, _05847_);
  and _61986_ (_10805_, _06125_, _06408_);
  or _61987_ (_10806_, _10805_, _10804_);
  and _61988_ (_10807_, _06119_, _06408_);
  nor _61989_ (_10808_, _10807_, _10806_);
  and _61990_ (_10809_, _10808_, _10803_);
  and _61991_ (_10810_, _10809_, _10802_);
  and _61992_ (_10811_, _06115_, _06408_);
  not _61993_ (_10812_, _10808_);
  and _61994_ (_10813_, _10812_, _10765_);
  or _61995_ (_10814_, _10813_, _10811_);
  or _61996_ (_10815_, _10814_, _10810_);
  not _61997_ (_10816_, _10811_);
  or _61998_ (_10817_, _10816_, _10782_);
  and _61999_ (_10818_, _10817_, _06410_);
  and _62000_ (_10819_, _10818_, _10815_);
  and _62001_ (_10820_, _06294_, _06408_);
  nor _62002_ (_10821_, _10820_, _06409_);
  not _62003_ (_10822_, _10821_);
  or _62004_ (_10823_, _10820_, _08808_);
  and _62005_ (_10824_, _10823_, _10822_);
  or _62006_ (_10825_, _10824_, _10819_);
  not _62007_ (_10826_, _10820_);
  or _62008_ (_10827_, _10826_, _10793_);
  and _62009_ (_10828_, _10827_, _07132_);
  and _62010_ (_10829_, _10828_, _10825_);
  nand _62011_ (_10830_, _10755_, _06306_);
  nor _62012_ (_10831_, _10830_, _08809_);
  or _62013_ (_10832_, _10831_, _06524_);
  or _62014_ (_10833_, _10832_, _10829_);
  not _62015_ (_10834_, _06555_);
  and _62016_ (_10835_, _06119_, _05840_);
  nor _62017_ (_10836_, _10835_, _06975_);
  and _62018_ (_10837_, _10836_, _10834_);
  nand _62019_ (_10838_, _10763_, _06524_);
  and _62020_ (_10839_, _10838_, _10837_);
  and _62021_ (_10840_, _10839_, _10833_);
  and _62022_ (_10841_, _06115_, _05840_);
  nor _62023_ (_10842_, _10837_, _10763_);
  or _62024_ (_10843_, _10842_, _10841_);
  or _62025_ (_10844_, _10843_, _10840_);
  nand _62026_ (_10845_, _10841_, _10781_);
  and _62027_ (_10846_, _10845_, _06395_);
  and _62028_ (_10847_, _10846_, _10844_);
  and _62029_ (_10848_, _06294_, _05840_);
  nor _62030_ (_10849_, _10848_, _06394_);
  not _62031_ (_10850_, _10849_);
  not _62032_ (_10851_, _10848_);
  nand _62033_ (_10852_, _10851_, _08809_);
  and _62034_ (_10853_, _10852_, _10850_);
  or _62035_ (_10854_, _10853_, _10847_);
  nand _62036_ (_10855_, _10848_, _10792_);
  and _62037_ (_10856_, _10855_, _08819_);
  and _62038_ (_10857_, _10856_, _10854_);
  not _62039_ (_10858_, _10380_);
  and _62040_ (_10859_, _08801_, _07809_);
  or _62041_ (_10860_, _10859_, _10383_);
  and _62042_ (_10861_, _10860_, _06303_);
  or _62043_ (_10862_, _10861_, _10858_);
  or _62044_ (_10863_, _10862_, _10857_);
  and _62045_ (_10864_, _10863_, _10381_);
  and _62046_ (_10865_, _06115_, _06300_);
  or _62047_ (_10866_, _10865_, _10864_);
  not _62048_ (_10867_, _10865_);
  nand _62049_ (_10868_, _10592_, \oc8051_golden_model_1.ACC [6]);
  and _62050_ (_10869_, _10596_, \oc8051_golden_model_1.ACC [5]);
  nand _62051_ (_10870_, _10603_, \oc8051_golden_model_1.ACC [4]);
  and _62052_ (_10871_, _10610_, \oc8051_golden_model_1.ACC [3]);
  and _62053_ (_10872_, _10616_, \oc8051_golden_model_1.ACC [2]);
  and _62054_ (_10873_, _10623_, \oc8051_golden_model_1.ACC [1]);
  nor _62055_ (_10874_, _10625_, _10624_);
  not _62056_ (_10875_, _10874_);
  and _62057_ (_10876_, _10627_, \oc8051_golden_model_1.ACC [0]);
  and _62058_ (_10877_, _10876_, _10875_);
  nor _62059_ (_10878_, _10877_, _10873_);
  nor _62060_ (_10879_, _10878_, _10619_);
  nor _62061_ (_10880_, _10879_, _10872_);
  nor _62062_ (_10881_, _10880_, _10613_);
  or _62063_ (_10882_, _10881_, _10871_);
  nand _62064_ (_10883_, _10882_, _10606_);
  and _62065_ (_10884_, _10883_, _10870_);
  nor _62066_ (_10885_, _10884_, _10599_);
  or _62067_ (_10886_, _10885_, _10869_);
  nand _62068_ (_10887_, _10886_, _10641_);
  and _62069_ (_10888_, _10887_, _10868_);
  nor _62070_ (_10889_, _10888_, _10589_);
  and _62071_ (_10890_, _10888_, _10589_);
  nor _62072_ (_10891_, _10890_, _10889_);
  or _62073_ (_10892_, _10891_, _10867_);
  and _62074_ (_10893_, _10892_, _06407_);
  and _62075_ (_10894_, _10893_, _10866_);
  and _62076_ (_10895_, _06294_, _06300_);
  nor _62077_ (_10896_, _10895_, _06406_);
  not _62078_ (_10897_, _10896_);
  and _62079_ (_10898_, _10404_, \oc8051_golden_model_1.ACC [6]);
  and _62080_ (_10899_, _10407_, \oc8051_golden_model_1.ACC [5]);
  nand _62081_ (_10900_, _10413_, \oc8051_golden_model_1.ACC [4]);
  and _62082_ (_10901_, _10419_, \oc8051_golden_model_1.ACC [3]);
  and _62083_ (_10902_, _10424_, \oc8051_golden_model_1.ACC [2]);
  and _62084_ (_10903_, _10430_, \oc8051_golden_model_1.ACC [1]);
  nor _62085_ (_10904_, _10432_, _10431_);
  not _62086_ (_10905_, _10904_);
  and _62087_ (_10906_, _10434_, \oc8051_golden_model_1.ACC [0]);
  and _62088_ (_10907_, _10906_, _10905_);
  nor _62089_ (_10908_, _10907_, _10903_);
  nor _62090_ (_10909_, _10908_, _10427_);
  nor _62091_ (_10910_, _10909_, _10902_);
  nor _62092_ (_10911_, _10910_, _10422_);
  or _62093_ (_10912_, _10911_, _10901_);
  nand _62094_ (_10913_, _10912_, _10416_);
  and _62095_ (_10914_, _10913_, _10900_);
  nor _62096_ (_10915_, _10914_, _10410_);
  or _62097_ (_10916_, _10915_, _10899_);
  and _62098_ (_10917_, _10916_, _10448_);
  nor _62099_ (_10918_, _10917_, _10898_);
  nor _62100_ (_10919_, _10918_, _10401_);
  and _62101_ (_10920_, _10918_, _10401_);
  nor _62102_ (_10921_, _10920_, _10919_);
  or _62103_ (_10922_, _10921_, _10895_);
  and _62104_ (_10923_, _10922_, _10897_);
  or _62105_ (_10924_, _10923_, _10894_);
  nor _62106_ (_10925_, _05844_, _05799_);
  not _62107_ (_10926_, _10925_);
  not _62108_ (_10927_, _10895_);
  and _62109_ (_10928_, _10664_, \oc8051_golden_model_1.ACC [6]);
  and _62110_ (_10929_, _10668_, \oc8051_golden_model_1.ACC [5]);
  nand _62111_ (_10930_, _10672_, \oc8051_golden_model_1.ACC [4]);
  and _62112_ (_10931_, _10682_, \oc8051_golden_model_1.ACC [3]);
  and _62113_ (_10932_, _10688_, \oc8051_golden_model_1.ACC [2]);
  and _62114_ (_10933_, _10696_, \oc8051_golden_model_1.ACC [1]);
  nor _62115_ (_10934_, _10699_, _10697_);
  not _62116_ (_10935_, _10934_);
  and _62117_ (_10936_, _10701_, \oc8051_golden_model_1.ACC [0]);
  and _62118_ (_10937_, _10936_, _10935_);
  nor _62119_ (_10938_, _10937_, _10933_);
  nor _62120_ (_10939_, _10938_, _10691_);
  nor _62121_ (_10940_, _10939_, _10932_);
  nor _62122_ (_10941_, _10940_, _10685_);
  or _62123_ (_10942_, _10941_, _10931_);
  nand _62124_ (_10943_, _10942_, _10679_);
  and _62125_ (_10944_, _10943_, _10930_);
  nor _62126_ (_10945_, _10944_, _10676_);
  or _62127_ (_10946_, _10945_, _10929_);
  and _62128_ (_10947_, _10946_, _10714_);
  nor _62129_ (_10948_, _10947_, _10928_);
  nor _62130_ (_10949_, _10948_, _10662_);
  and _62131_ (_10950_, _10948_, _10662_);
  nor _62132_ (_10951_, _10950_, _10949_);
  or _62133_ (_10952_, _10951_, _10927_);
  and _62134_ (_10953_, _10952_, _10926_);
  and _62135_ (_10954_, _10953_, _10924_);
  nand _62136_ (_10955_, _10925_, \oc8051_golden_model_1.ACC [6]);
  and _62137_ (_10956_, _06273_, _05825_);
  not _62138_ (_10957_, _10956_);
  and _62139_ (_10958_, _06288_, _05825_);
  nor _62140_ (_10959_, _10958_, _06952_);
  and _62141_ (_10960_, _06122_, _05825_);
  nor _62142_ (_10961_, _06958_, _10960_);
  and _62143_ (_10962_, _10961_, _10959_);
  and _62144_ (_10963_, _10962_, _10957_);
  nand _62145_ (_10964_, _10963_, _10955_);
  or _62146_ (_10965_, _10964_, _10954_);
  and _62147_ (_10966_, _08012_, \oc8051_golden_model_1.ACC [6]);
  or _62148_ (_10967_, _08012_, \oc8051_golden_model_1.ACC [6]);
  not _62149_ (_10968_, _10966_);
  and _62150_ (_10969_, _10968_, _10967_);
  and _62151_ (_10970_, _08101_, \oc8051_golden_model_1.ACC [5]);
  and _62152_ (_10971_, _08348_, _09930_);
  and _62153_ (_10972_, _08336_, \oc8051_golden_model_1.ACC [4]);
  or _62154_ (_10973_, _08336_, \oc8051_golden_model_1.ACC [4]);
  not _62155_ (_10974_, _10972_);
  and _62156_ (_10975_, _10974_, _10973_);
  and _62157_ (_10976_, _07544_, \oc8051_golden_model_1.ACC [3]);
  and _62158_ (_10977_, _07474_, _10028_);
  and _62159_ (_10978_, _07708_, \oc8051_golden_model_1.ACC [2]);
  and _62160_ (_10979_, _07657_, _09981_);
  nor _62161_ (_10980_, _10978_, _10979_);
  not _62162_ (_10981_, _10980_);
  and _62163_ (_10982_, _07306_, \oc8051_golden_model_1.ACC [1]);
  and _62164_ (_10983_, _07252_, _05887_);
  nor _62165_ (_10984_, _10982_, _10983_);
  and _62166_ (_10985_, _07049_, \oc8051_golden_model_1.ACC [0]);
  and _62167_ (_10986_, _10985_, _10984_);
  nor _62168_ (_10987_, _10986_, _10982_);
  nor _62169_ (_10988_, _10987_, _10981_);
  nor _62170_ (_10989_, _10988_, _10978_);
  nor _62171_ (_10990_, _10989_, _10977_);
  or _62172_ (_10991_, _10990_, _10976_);
  and _62173_ (_10992_, _10991_, _10975_);
  nor _62174_ (_10993_, _10992_, _10972_);
  nor _62175_ (_10994_, _10993_, _10971_);
  or _62176_ (_10995_, _10994_, _10970_);
  and _62177_ (_10996_, _10995_, _10969_);
  nor _62178_ (_10997_, _10996_, _10966_);
  and _62179_ (_10998_, _10997_, _10766_);
  nor _62180_ (_10999_, _10997_, _10766_);
  or _62181_ (_11000_, _10999_, _10998_);
  or _62182_ (_11001_, _11000_, _10963_);
  and _62183_ (_11002_, _11001_, _10965_);
  and _62184_ (_11003_, _06115_, _05825_);
  or _62185_ (_11004_, _11003_, _11002_);
  and _62186_ (_11005_, _09207_, \oc8051_golden_model_1.ACC [6]);
  or _62187_ (_11006_, _09207_, \oc8051_golden_model_1.ACC [6]);
  not _62188_ (_11007_, _11005_);
  and _62189_ (_11008_, _11007_, _11006_);
  and _62190_ (_11009_, _09208_, \oc8051_golden_model_1.ACC [5]);
  and _62191_ (_11010_, _08931_, _09930_);
  or _62192_ (_11011_, _11010_, _11009_);
  and _62193_ (_11012_, _09209_, \oc8051_golden_model_1.ACC [4]);
  not _62194_ (_11013_, _11012_);
  or _62195_ (_11014_, _09209_, \oc8051_golden_model_1.ACC [4]);
  and _62196_ (_11015_, _11013_, _11014_);
  and _62197_ (_11016_, _09210_, \oc8051_golden_model_1.ACC [3]);
  and _62198_ (_11017_, _09025_, _10028_);
  and _62199_ (_11018_, _09211_, \oc8051_golden_model_1.ACC [2]);
  or _62200_ (_11019_, _09211_, \oc8051_golden_model_1.ACC [2]);
  not _62201_ (_11020_, _11018_);
  and _62202_ (_11021_, _11020_, _11019_);
  not _62203_ (_11022_, _11021_);
  and _62204_ (_11023_, _09115_, \oc8051_golden_model_1.ACC [1]);
  or _62205_ (_11024_, _09115_, \oc8051_golden_model_1.ACC [1]);
  not _62206_ (_11025_, _11023_);
  and _62207_ (_11026_, _11025_, _11024_);
  and _62208_ (_11027_, _09160_, \oc8051_golden_model_1.ACC [0]);
  and _62209_ (_11028_, _11027_, _11026_);
  nor _62210_ (_11029_, _11028_, _11023_);
  nor _62211_ (_11030_, _11029_, _11022_);
  nor _62212_ (_11031_, _11030_, _11018_);
  nor _62213_ (_11032_, _11031_, _11017_);
  or _62214_ (_11033_, _11032_, _11016_);
  nand _62215_ (_11034_, _11033_, _11015_);
  and _62216_ (_11035_, _11034_, _11013_);
  nor _62217_ (_11036_, _11035_, _11011_);
  or _62218_ (_11037_, _11036_, _11009_);
  and _62219_ (_11038_, _11037_, _11008_);
  nor _62220_ (_11039_, _11038_, _11005_);
  and _62221_ (_11040_, _11039_, _10783_);
  not _62222_ (_11041_, _11003_);
  nor _62223_ (_11042_, _11039_, _10783_);
  or _62224_ (_11043_, _11042_, _11041_);
  or _62225_ (_11044_, _11043_, _11040_);
  and _62226_ (_11045_, _11044_, _06171_);
  and _62227_ (_11046_, _11045_, _11004_);
  or _62228_ (_11047_, _11046_, _10301_);
  and _62229_ (_11048_, _11047_, _10265_);
  nor _62230_ (_11049_, _06203_, _09883_);
  not _62231_ (_11050_, _11049_);
  and _62232_ (_11051_, _06203_, _09883_);
  nor _62233_ (_11052_, _11049_, _11051_);
  nor _62234_ (_11053_, _06477_, _09930_);
  and _62235_ (_11054_, _06477_, _09930_);
  nor _62236_ (_11055_, _06876_, _09902_);
  not _62237_ (_11056_, _11055_);
  and _62238_ (_11057_, _06876_, _09902_);
  nor _62239_ (_11058_, _11055_, _11057_);
  nor _62240_ (_11059_, _06070_, _10028_);
  and _62241_ (_11060_, _06070_, _10028_);
  nor _62242_ (_11061_, _06625_, _09981_);
  and _62243_ (_11062_, _06625_, _09981_);
  nor _62244_ (_11063_, _11061_, _11062_);
  nor _62245_ (_11064_, _06912_, _05887_);
  and _62246_ (_11065_, _06912_, _05887_);
  nor _62247_ (_11066_, _11064_, _11065_);
  nor _62248_ (_11067_, _06107_, _05855_);
  and _62249_ (_11068_, _11067_, _11066_);
  nor _62250_ (_11069_, _11068_, _11064_);
  not _62251_ (_11070_, _11069_);
  and _62252_ (_11071_, _11070_, _11063_);
  nor _62253_ (_11072_, _11071_, _11061_);
  nor _62254_ (_11073_, _11072_, _11060_);
  or _62255_ (_11074_, _11073_, _11059_);
  nand _62256_ (_11075_, _11074_, _11058_);
  and _62257_ (_11076_, _11075_, _11056_);
  nor _62258_ (_11077_, _11076_, _11054_);
  or _62259_ (_11078_, _11077_, _11053_);
  nand _62260_ (_11079_, _11078_, _11052_);
  and _62261_ (_11080_, _11079_, _11050_);
  nor _62262_ (_11081_, _11080_, _10794_);
  and _62263_ (_11082_, _11080_, _10794_);
  or _62264_ (_11083_, _11082_, _11081_);
  and _62265_ (_11084_, _11083_, _10264_);
  or _62266_ (_11085_, _11084_, _10262_);
  or _62267_ (_11086_, _11085_, _11048_);
  and _62268_ (_11087_, _11086_, _10263_);
  or _62269_ (_11088_, _11087_, _06433_);
  and _62270_ (_11089_, _06294_, _05591_);
  not _62271_ (_11090_, _11089_);
  or _62272_ (_11091_, _10487_, _06829_);
  and _62273_ (_11092_, _11091_, _11090_);
  and _62274_ (_11093_, _11092_, _11088_);
  and _62275_ (_11094_, _06302_, _05591_);
  and _62276_ (_11095_, _10493_, _05855_);
  and _62277_ (_11096_, _11095_, _10028_);
  and _62278_ (_11097_, _11096_, _09902_);
  and _62279_ (_11098_, _11097_, _09930_);
  and _62280_ (_11099_, _11098_, _09883_);
  nor _62281_ (_11100_, _11099_, _08430_);
  and _62282_ (_11101_, _11099_, _08430_);
  or _62283_ (_11102_, _11101_, _11100_);
  and _62284_ (_11103_, _11102_, _11089_);
  or _62285_ (_11104_, _11103_, _11094_);
  or _62286_ (_11105_, _11104_, _11093_);
  nand _62287_ (_11106_, _11094_, _10693_);
  and _62288_ (_11107_, _11106_, _05749_);
  and _62289_ (_11108_, _11107_, _11105_);
  and _62290_ (_11109_, _10533_, _05748_);
  or _62291_ (_11110_, _11109_, _06440_);
  or _62292_ (_11111_, _11110_, _11108_);
  and _62293_ (_11112_, _06294_, _05820_);
  not _62294_ (_11113_, _11112_);
  and _62295_ (_11114_, _08345_, _07809_);
  or _62296_ (_11115_, _10383_, _06444_);
  or _62297_ (_11116_, _11115_, _11114_);
  and _62298_ (_11117_, _11116_, _11113_);
  and _62299_ (_11118_, _11117_, _11111_);
  and _62300_ (_11119_, _05820_, _06302_);
  and _62301_ (_11120_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and _62302_ (_11121_, _11120_, \oc8051_golden_model_1.ACC [2]);
  and _62303_ (_11122_, _11121_, \oc8051_golden_model_1.ACC [3]);
  and _62304_ (_11123_, _11122_, \oc8051_golden_model_1.ACC [4]);
  and _62305_ (_11124_, _11123_, \oc8051_golden_model_1.ACC [5]);
  and _62306_ (_11125_, _11124_, \oc8051_golden_model_1.ACC [6]);
  nor _62307_ (_11126_, _11125_, _08430_);
  and _62308_ (_11127_, _11125_, _08430_);
  or _62309_ (_11128_, _11127_, _11126_);
  and _62310_ (_11129_, _11128_, _11112_);
  or _62311_ (_11130_, _11129_, _11119_);
  or _62312_ (_11131_, _11130_, _11118_);
  nand _62313_ (_11132_, _11119_, _05855_);
  and _62314_ (_11133_, _11132_, _01317_);
  and _62315_ (_11134_, _11133_, _11131_);
  or _62316_ (_11135_, _11134_, _10261_);
  and _62317_ (_40981_, _11135_, _43100_);
  not _62318_ (_11136_, _06298_);
  not _62319_ (_11137_, _07856_);
  and _62320_ (_11138_, _11137_, \oc8051_golden_model_1.PCON [7]);
  and _62321_ (_11139_, _07923_, _07856_);
  or _62322_ (_11140_, _11139_, _11138_);
  or _62323_ (_11141_, _11140_, _06132_);
  and _62324_ (_11142_, _08548_, _07856_);
  or _62325_ (_11143_, _11142_, _11138_);
  or _62326_ (_11144_, _11143_, _06161_);
  and _62327_ (_11145_, _07856_, \oc8051_golden_model_1.ACC [7]);
  or _62328_ (_11146_, _11145_, _11138_);
  and _62329_ (_11147_, _11146_, _07056_);
  and _62330_ (_11148_, _07057_, \oc8051_golden_model_1.PCON [7]);
  or _62331_ (_11149_, _11148_, _06160_);
  or _62332_ (_11150_, _11149_, _11147_);
  and _62333_ (_11151_, _11150_, _07075_);
  and _62334_ (_11152_, _11151_, _11144_);
  and _62335_ (_11153_, _11140_, _06217_);
  or _62336_ (_11154_, _11153_, _11152_);
  and _62337_ (_11155_, _11154_, _06229_);
  and _62338_ (_11156_, _11146_, _06220_);
  or _62339_ (_11157_, _11156_, _09842_);
  or _62340_ (_11158_, _11157_, _11155_);
  and _62341_ (_11159_, _11158_, _11141_);
  or _62342_ (_11160_, _11159_, _06116_);
  and _62343_ (_11161_, _08535_, _07856_);
  or _62344_ (_11162_, _11138_, _06117_);
  or _62345_ (_11163_, _11162_, _11161_);
  and _62346_ (_11164_, _11163_, _06114_);
  and _62347_ (_11165_, _11164_, _11160_);
  and _62348_ (_11166_, _08782_, _07856_);
  or _62349_ (_11167_, _11166_, _11138_);
  and _62350_ (_11168_, _11167_, _05787_);
  or _62351_ (_11169_, _11168_, _11165_);
  or _62352_ (_11170_, _11169_, _11136_);
  and _62353_ (_11171_, _08802_, _07856_);
  or _62354_ (_11172_, _11138_, _07127_);
  or _62355_ (_11173_, _11172_, _11171_);
  and _62356_ (_11174_, _08607_, _07856_);
  or _62357_ (_11175_, _11174_, _11138_);
  or _62358_ (_11176_, _11175_, _06111_);
  and _62359_ (_11177_, _11176_, _07125_);
  and _62360_ (_11178_, _11177_, _11173_);
  and _62361_ (_11179_, _11178_, _11170_);
  and _62362_ (_11180_, _08810_, _07856_);
  or _62363_ (_11181_, _11180_, _11138_);
  and _62364_ (_11182_, _11181_, _06402_);
  or _62365_ (_11183_, _11182_, _11179_);
  and _62366_ (_11184_, _11183_, _07132_);
  or _62367_ (_11185_, _11138_, _07926_);
  and _62368_ (_11186_, _11175_, _06306_);
  and _62369_ (_11187_, _11186_, _11185_);
  or _62370_ (_11188_, _11187_, _11184_);
  and _62371_ (_11189_, _11188_, _07130_);
  and _62372_ (_11190_, _11146_, _06411_);
  and _62373_ (_11191_, _11190_, _11185_);
  or _62374_ (_11192_, _11191_, _06303_);
  or _62375_ (_11193_, _11192_, _11189_);
  and _62376_ (_11194_, _08801_, _07856_);
  or _62377_ (_11195_, _11138_, _08819_);
  or _62378_ (_11196_, _11195_, _11194_);
  and _62379_ (_11197_, _11196_, _08824_);
  and _62380_ (_11198_, _11197_, _11193_);
  nor _62381_ (_11199_, _08809_, _11137_);
  or _62382_ (_11200_, _11199_, _11138_);
  and _62383_ (_11201_, _11200_, _06396_);
  or _62384_ (_11202_, _11201_, _06433_);
  or _62385_ (_11203_, _11202_, _11198_);
  or _62386_ (_11204_, _11143_, _06829_);
  and _62387_ (_11205_, _11204_, _06444_);
  and _62388_ (_11206_, _11205_, _11203_);
  and _62389_ (_11207_, _08345_, _07856_);
  or _62390_ (_11208_, _11207_, _11138_);
  and _62391_ (_11209_, _11208_, _06440_);
  or _62392_ (_11210_, _11209_, _01321_);
  or _62393_ (_11211_, _11210_, _11206_);
  or _62394_ (_11212_, _01317_, \oc8051_golden_model_1.PCON [7]);
  and _62395_ (_11213_, _11212_, _43100_);
  and _62396_ (_40982_, _11213_, _11211_);
  not _62397_ (_11214_, _07812_);
  and _62398_ (_11215_, _11214_, \oc8051_golden_model_1.TMOD [7]);
  and _62399_ (_11216_, _07923_, _07812_);
  or _62400_ (_11217_, _11216_, _11215_);
  or _62401_ (_11218_, _11217_, _06132_);
  and _62402_ (_11219_, _08548_, _07812_);
  or _62403_ (_11220_, _11219_, _11215_);
  or _62404_ (_11221_, _11220_, _06161_);
  and _62405_ (_11222_, _07812_, \oc8051_golden_model_1.ACC [7]);
  or _62406_ (_11223_, _11222_, _11215_);
  and _62407_ (_11224_, _11223_, _07056_);
  and _62408_ (_11225_, _07057_, \oc8051_golden_model_1.TMOD [7]);
  or _62409_ (_11226_, _11225_, _06160_);
  or _62410_ (_11227_, _11226_, _11224_);
  and _62411_ (_11228_, _11227_, _07075_);
  and _62412_ (_11229_, _11228_, _11221_);
  and _62413_ (_11230_, _11217_, _06217_);
  or _62414_ (_11231_, _11230_, _11229_);
  and _62415_ (_11232_, _11231_, _06229_);
  and _62416_ (_11233_, _11223_, _06220_);
  or _62417_ (_11234_, _11233_, _09842_);
  or _62418_ (_11235_, _11234_, _11232_);
  and _62419_ (_11236_, _11235_, _11218_);
  or _62420_ (_11237_, _11236_, _06116_);
  and _62421_ (_11238_, _08535_, _07812_);
  or _62422_ (_11239_, _11215_, _06117_);
  or _62423_ (_11240_, _11239_, _11238_);
  and _62424_ (_11241_, _11240_, _06114_);
  and _62425_ (_11242_, _11241_, _11237_);
  and _62426_ (_11243_, _08782_, _07812_);
  or _62427_ (_11244_, _11243_, _11215_);
  and _62428_ (_11245_, _11244_, _05787_);
  or _62429_ (_11246_, _11245_, _11242_);
  or _62430_ (_11247_, _11246_, _11136_);
  and _62431_ (_11248_, _08802_, _07812_);
  or _62432_ (_11249_, _11215_, _07127_);
  or _62433_ (_11250_, _11249_, _11248_);
  and _62434_ (_11251_, _08607_, _07812_);
  or _62435_ (_11252_, _11251_, _11215_);
  or _62436_ (_11253_, _11252_, _06111_);
  and _62437_ (_11254_, _11253_, _07125_);
  and _62438_ (_11255_, _11254_, _11250_);
  and _62439_ (_11256_, _11255_, _11247_);
  and _62440_ (_11257_, _08810_, _07812_);
  or _62441_ (_11258_, _11257_, _11215_);
  and _62442_ (_11259_, _11258_, _06402_);
  or _62443_ (_11260_, _11259_, _11256_);
  and _62444_ (_11261_, _11260_, _07132_);
  or _62445_ (_11262_, _11215_, _07926_);
  and _62446_ (_11263_, _11252_, _06306_);
  and _62447_ (_11264_, _11263_, _11262_);
  or _62448_ (_11265_, _11264_, _11261_);
  and _62449_ (_11266_, _11265_, _07130_);
  and _62450_ (_11267_, _11223_, _06411_);
  and _62451_ (_11268_, _11267_, _11262_);
  or _62452_ (_11269_, _11268_, _06303_);
  or _62453_ (_11270_, _11269_, _11266_);
  and _62454_ (_11271_, _08801_, _07812_);
  or _62455_ (_11272_, _11215_, _08819_);
  or _62456_ (_11273_, _11272_, _11271_);
  and _62457_ (_11274_, _11273_, _08824_);
  and _62458_ (_11275_, _11274_, _11270_);
  nor _62459_ (_11276_, _08809_, _11214_);
  or _62460_ (_11277_, _11276_, _11215_);
  and _62461_ (_11278_, _11277_, _06396_);
  or _62462_ (_11279_, _11278_, _06433_);
  or _62463_ (_11280_, _11279_, _11275_);
  or _62464_ (_11281_, _11220_, _06829_);
  and _62465_ (_11282_, _11281_, _06444_);
  and _62466_ (_11283_, _11282_, _11280_);
  and _62467_ (_11284_, _08345_, _07812_);
  or _62468_ (_11285_, _11284_, _11215_);
  and _62469_ (_11286_, _11285_, _06440_);
  or _62470_ (_11287_, _11286_, _01321_);
  or _62471_ (_11288_, _11287_, _11283_);
  or _62472_ (_11289_, _01317_, \oc8051_golden_model_1.TMOD [7]);
  and _62473_ (_11290_, _11289_, _43100_);
  and _62474_ (_40983_, _11290_, _11288_);
  not _62475_ (_11291_, \oc8051_golden_model_1.DPL [7]);
  nor _62476_ (_11292_, _07849_, _11291_);
  and _62477_ (_11293_, _07923_, _07849_);
  or _62478_ (_11294_, _11293_, _11292_);
  or _62479_ (_11295_, _11294_, _06132_);
  not _62480_ (_11296_, _06293_);
  and _62481_ (_11297_, _08548_, _07849_);
  or _62482_ (_11298_, _11297_, _11292_);
  or _62483_ (_11299_, _11298_, _06161_);
  and _62484_ (_11300_, _07849_, \oc8051_golden_model_1.ACC [7]);
  or _62485_ (_11301_, _11300_, _11292_);
  and _62486_ (_11302_, _11301_, _07056_);
  nor _62487_ (_11303_, _07056_, _11291_);
  or _62488_ (_11304_, _11303_, _06160_);
  or _62489_ (_11305_, _11304_, _11302_);
  and _62490_ (_11306_, _11305_, _07075_);
  and _62491_ (_11307_, _11306_, _11299_);
  and _62492_ (_11308_, _11294_, _06217_);
  or _62493_ (_11309_, _11308_, _06220_);
  or _62494_ (_11310_, _11309_, _11307_);
  nor _62495_ (_11311_, _05799_, _05774_);
  not _62496_ (_11312_, _11311_);
  or _62497_ (_11313_, _11301_, _06229_);
  and _62498_ (_11314_, _11313_, _11312_);
  and _62499_ (_11315_, _11314_, _11310_);
  and _62500_ (_11316_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and _62501_ (_11317_, _11316_, \oc8051_golden_model_1.DPL [2]);
  and _62502_ (_11318_, _11317_, \oc8051_golden_model_1.DPL [3]);
  and _62503_ (_11319_, _11318_, \oc8051_golden_model_1.DPL [4]);
  and _62504_ (_11320_, _11319_, \oc8051_golden_model_1.DPL [5]);
  and _62505_ (_11321_, _11320_, \oc8051_golden_model_1.DPL [6]);
  nor _62506_ (_11322_, _11321_, \oc8051_golden_model_1.DPL [7]);
  and _62507_ (_11323_, _11321_, \oc8051_golden_model_1.DPL [7]);
  nor _62508_ (_11324_, _11323_, _11322_);
  and _62509_ (_11325_, _11324_, _11311_);
  or _62510_ (_11326_, _11325_, _11315_);
  and _62511_ (_11327_, _11326_, _11296_);
  nor _62512_ (_11328_, _08395_, _11296_);
  or _62513_ (_11329_, _11328_, _09842_);
  or _62514_ (_11330_, _11329_, _11327_);
  and _62515_ (_11331_, _11330_, _11295_);
  or _62516_ (_11332_, _11331_, _06116_);
  and _62517_ (_11333_, _08535_, _07849_);
  or _62518_ (_11334_, _11292_, _06117_);
  or _62519_ (_11335_, _11334_, _11333_);
  and _62520_ (_11336_, _11335_, _06114_);
  and _62521_ (_11337_, _11336_, _11332_);
  and _62522_ (_11338_, _08782_, _07849_);
  or _62523_ (_11339_, _11338_, _11292_);
  and _62524_ (_11340_, _11339_, _05787_);
  or _62525_ (_11341_, _11340_, _11337_);
  or _62526_ (_11342_, _11341_, _11136_);
  and _62527_ (_11343_, _08802_, _07849_);
  or _62528_ (_11344_, _11292_, _07127_);
  or _62529_ (_11345_, _11344_, _11343_);
  and _62530_ (_11346_, _08607_, _07849_);
  or _62531_ (_11347_, _11346_, _11292_);
  or _62532_ (_11348_, _11347_, _06111_);
  and _62533_ (_11349_, _11348_, _07125_);
  and _62534_ (_11350_, _11349_, _11345_);
  and _62535_ (_11351_, _11350_, _11342_);
  and _62536_ (_11352_, _08810_, _07849_);
  or _62537_ (_11353_, _11352_, _11292_);
  and _62538_ (_11354_, _11353_, _06402_);
  or _62539_ (_11355_, _11354_, _11351_);
  and _62540_ (_11356_, _11355_, _07132_);
  or _62541_ (_11357_, _11292_, _07926_);
  and _62542_ (_11358_, _11347_, _06306_);
  and _62543_ (_11359_, _11358_, _11357_);
  or _62544_ (_11360_, _11359_, _11356_);
  and _62545_ (_11361_, _11360_, _07130_);
  and _62546_ (_11362_, _11301_, _06411_);
  and _62547_ (_11363_, _11362_, _11357_);
  or _62548_ (_11364_, _11363_, _06303_);
  or _62549_ (_11365_, _11364_, _11361_);
  and _62550_ (_11366_, _08801_, _07849_);
  or _62551_ (_11367_, _11292_, _08819_);
  or _62552_ (_11368_, _11367_, _11366_);
  and _62553_ (_11369_, _11368_, _08824_);
  and _62554_ (_11370_, _11369_, _11365_);
  not _62555_ (_11371_, _07849_);
  nor _62556_ (_11372_, _08809_, _11371_);
  or _62557_ (_11373_, _11372_, _11292_);
  and _62558_ (_11374_, _11373_, _06396_);
  or _62559_ (_11375_, _11374_, _06433_);
  or _62560_ (_11376_, _11375_, _11370_);
  or _62561_ (_11377_, _11298_, _06829_);
  and _62562_ (_11378_, _11377_, _06444_);
  and _62563_ (_11379_, _11378_, _11376_);
  and _62564_ (_11380_, _08345_, _07849_);
  or _62565_ (_11381_, _11380_, _11292_);
  and _62566_ (_11382_, _11381_, _06440_);
  or _62567_ (_11383_, _11382_, _01321_);
  or _62568_ (_11384_, _11383_, _11379_);
  or _62569_ (_11385_, _01317_, \oc8051_golden_model_1.DPL [7]);
  and _62570_ (_11386_, _11385_, _43100_);
  and _62571_ (_40985_, _11386_, _11384_);
  not _62572_ (_11387_, \oc8051_golden_model_1.DPH [7]);
  nand _62573_ (_11388_, _06625_, _06070_);
  nor _62574_ (_11389_, _07835_, _11388_);
  and _62575_ (_11390_, _11389_, _07787_);
  nor _62576_ (_11391_, _11390_, _11387_);
  and _62577_ (_11392_, _07923_, _07852_);
  or _62578_ (_11393_, _11392_, _11391_);
  or _62579_ (_11394_, _11393_, _06132_);
  and _62580_ (_11395_, _08548_, _07852_);
  or _62581_ (_11396_, _11395_, _11391_);
  or _62582_ (_11397_, _11396_, _06161_);
  and _62583_ (_11398_, _11390_, \oc8051_golden_model_1.ACC [7]);
  or _62584_ (_11399_, _11398_, _11391_);
  and _62585_ (_11400_, _11399_, _07056_);
  nor _62586_ (_11401_, _07056_, _11387_);
  or _62587_ (_11402_, _11401_, _06160_);
  or _62588_ (_11403_, _11402_, _11400_);
  and _62589_ (_11404_, _11403_, _07075_);
  and _62590_ (_11405_, _11404_, _11397_);
  and _62591_ (_11406_, _11393_, _06217_);
  or _62592_ (_11407_, _11406_, _06220_);
  or _62593_ (_11408_, _11407_, _11405_);
  or _62594_ (_11409_, _11399_, _06229_);
  and _62595_ (_11410_, _11409_, _11312_);
  and _62596_ (_11411_, _11410_, _11408_);
  and _62597_ (_11412_, _11323_, \oc8051_golden_model_1.DPH [0]);
  and _62598_ (_11413_, _11412_, \oc8051_golden_model_1.DPH [1]);
  and _62599_ (_11414_, _11413_, \oc8051_golden_model_1.DPH [2]);
  and _62600_ (_11415_, _11414_, \oc8051_golden_model_1.DPH [3]);
  and _62601_ (_11416_, _11415_, \oc8051_golden_model_1.DPH [4]);
  and _62602_ (_11417_, _11416_, \oc8051_golden_model_1.DPH [5]);
  and _62603_ (_11418_, _11417_, \oc8051_golden_model_1.DPH [6]);
  nand _62604_ (_11419_, _11418_, \oc8051_golden_model_1.DPH [7]);
  or _62605_ (_11420_, _11418_, \oc8051_golden_model_1.DPH [7]);
  and _62606_ (_11421_, _11420_, _11311_);
  and _62607_ (_11422_, _11421_, _11419_);
  or _62608_ (_11423_, _11422_, _11411_);
  and _62609_ (_11424_, _11423_, _11296_);
  and _62610_ (_11425_, _06293_, _06039_);
  or _62611_ (_11426_, _11425_, _09842_);
  or _62612_ (_11427_, _11426_, _11424_);
  and _62613_ (_11428_, _11427_, _11394_);
  or _62614_ (_11429_, _11428_, _06116_);
  or _62615_ (_11430_, _11391_, _06117_);
  and _62616_ (_11431_, _08535_, _11390_);
  or _62617_ (_11432_, _11431_, _11430_);
  and _62618_ (_11433_, _11432_, _06114_);
  and _62619_ (_11434_, _11433_, _11429_);
  and _62620_ (_11435_, _08782_, _11390_);
  or _62621_ (_11436_, _11435_, _11391_);
  and _62622_ (_11437_, _11436_, _05787_);
  or _62623_ (_11438_, _11437_, _11434_);
  or _62624_ (_11439_, _11438_, _11136_);
  and _62625_ (_11440_, _08802_, _07852_);
  or _62626_ (_11441_, _11391_, _07127_);
  or _62627_ (_11442_, _11441_, _11440_);
  and _62628_ (_11443_, _08607_, _11390_);
  or _62629_ (_11444_, _11443_, _11391_);
  or _62630_ (_11445_, _11444_, _06111_);
  and _62631_ (_11446_, _11445_, _07125_);
  and _62632_ (_11447_, _11446_, _11442_);
  and _62633_ (_11448_, _11447_, _11439_);
  and _62634_ (_11449_, _08810_, _07852_);
  or _62635_ (_11450_, _11449_, _11391_);
  and _62636_ (_11451_, _11450_, _06402_);
  or _62637_ (_11452_, _11451_, _11448_);
  and _62638_ (_11453_, _11452_, _07132_);
  or _62639_ (_11454_, _11391_, _07926_);
  and _62640_ (_11455_, _11444_, _06306_);
  and _62641_ (_11456_, _11455_, _11454_);
  or _62642_ (_11457_, _11456_, _11453_);
  and _62643_ (_11458_, _11457_, _07130_);
  and _62644_ (_11459_, _11399_, _06411_);
  and _62645_ (_11460_, _11459_, _11454_);
  or _62646_ (_11461_, _11460_, _06303_);
  or _62647_ (_11462_, _11461_, _11458_);
  and _62648_ (_11463_, _08801_, _07852_);
  or _62649_ (_11464_, _11391_, _08819_);
  or _62650_ (_11465_, _11464_, _11463_);
  and _62651_ (_11466_, _11465_, _08824_);
  and _62652_ (_11467_, _11466_, _11462_);
  not _62653_ (_11468_, _07852_);
  nor _62654_ (_11469_, _08809_, _11468_);
  or _62655_ (_11470_, _11469_, _11391_);
  and _62656_ (_11471_, _11470_, _06396_);
  or _62657_ (_11472_, _11471_, _06433_);
  or _62658_ (_11473_, _11472_, _11467_);
  or _62659_ (_11474_, _11396_, _06829_);
  and _62660_ (_11475_, _11474_, _06444_);
  and _62661_ (_11476_, _11475_, _11473_);
  and _62662_ (_11477_, _08345_, _07852_);
  or _62663_ (_11478_, _11477_, _11391_);
  and _62664_ (_11479_, _11478_, _06440_);
  or _62665_ (_11480_, _11479_, _01321_);
  or _62666_ (_11481_, _11480_, _11476_);
  or _62667_ (_11482_, _01317_, \oc8051_golden_model_1.DPH [7]);
  and _62668_ (_11483_, _11482_, _43100_);
  and _62669_ (_40986_, _11483_, _11481_);
  not _62670_ (_11484_, _07837_);
  and _62671_ (_11485_, _11484_, \oc8051_golden_model_1.TL1 [7]);
  and _62672_ (_11486_, _07923_, _07837_);
  or _62673_ (_11487_, _11486_, _11485_);
  or _62674_ (_11488_, _11487_, _06132_);
  and _62675_ (_11489_, _08548_, _07837_);
  or _62676_ (_11490_, _11489_, _11485_);
  or _62677_ (_11491_, _11490_, _06161_);
  and _62678_ (_11492_, _07837_, \oc8051_golden_model_1.ACC [7]);
  or _62679_ (_11493_, _11492_, _11485_);
  and _62680_ (_11494_, _11493_, _07056_);
  and _62681_ (_11495_, _07057_, \oc8051_golden_model_1.TL1 [7]);
  or _62682_ (_11496_, _11495_, _06160_);
  or _62683_ (_11497_, _11496_, _11494_);
  and _62684_ (_11498_, _11497_, _07075_);
  and _62685_ (_11499_, _11498_, _11491_);
  and _62686_ (_11500_, _11487_, _06217_);
  or _62687_ (_11501_, _11500_, _11499_);
  and _62688_ (_11502_, _11501_, _06229_);
  and _62689_ (_11503_, _11493_, _06220_);
  or _62690_ (_11504_, _11503_, _09842_);
  or _62691_ (_11505_, _11504_, _11502_);
  and _62692_ (_11506_, _11505_, _11488_);
  or _62693_ (_11507_, _11506_, _06116_);
  and _62694_ (_11508_, _08535_, _07837_);
  or _62695_ (_11509_, _11485_, _06117_);
  or _62696_ (_11510_, _11509_, _11508_);
  and _62697_ (_11511_, _11510_, _06114_);
  and _62698_ (_11512_, _11511_, _11507_);
  and _62699_ (_11513_, _08782_, _07837_);
  or _62700_ (_11514_, _11513_, _11485_);
  and _62701_ (_11515_, _11514_, _05787_);
  or _62702_ (_11516_, _11515_, _11512_);
  or _62703_ (_11517_, _11516_, _11136_);
  and _62704_ (_11518_, _08802_, _07837_);
  or _62705_ (_11519_, _11485_, _07127_);
  or _62706_ (_11520_, _11519_, _11518_);
  and _62707_ (_11521_, _08607_, _07837_);
  or _62708_ (_11522_, _11521_, _11485_);
  or _62709_ (_11523_, _11522_, _06111_);
  and _62710_ (_11524_, _11523_, _07125_);
  and _62711_ (_11525_, _11524_, _11520_);
  and _62712_ (_11526_, _11525_, _11517_);
  and _62713_ (_11527_, _08810_, _07837_);
  or _62714_ (_11528_, _11527_, _11485_);
  and _62715_ (_11529_, _11528_, _06402_);
  or _62716_ (_11530_, _11529_, _11526_);
  and _62717_ (_11531_, _11530_, _07132_);
  or _62718_ (_11532_, _11485_, _07926_);
  and _62719_ (_11533_, _11522_, _06306_);
  and _62720_ (_11534_, _11533_, _11532_);
  or _62721_ (_11535_, _11534_, _11531_);
  and _62722_ (_11536_, _11535_, _07130_);
  and _62723_ (_11537_, _11493_, _06411_);
  and _62724_ (_11538_, _11537_, _11532_);
  or _62725_ (_11539_, _11538_, _06303_);
  or _62726_ (_11540_, _11539_, _11536_);
  and _62727_ (_11541_, _08801_, _07837_);
  or _62728_ (_11542_, _11485_, _08819_);
  or _62729_ (_11543_, _11542_, _11541_);
  and _62730_ (_11544_, _11543_, _08824_);
  and _62731_ (_11545_, _11544_, _11540_);
  nor _62732_ (_11546_, _08809_, _11484_);
  or _62733_ (_11547_, _11546_, _11485_);
  and _62734_ (_11548_, _11547_, _06396_);
  or _62735_ (_11549_, _11548_, _06433_);
  or _62736_ (_11550_, _11549_, _11545_);
  or _62737_ (_11551_, _11490_, _06829_);
  and _62738_ (_11552_, _11551_, _06444_);
  and _62739_ (_11553_, _11552_, _11550_);
  and _62740_ (_11554_, _08345_, _07837_);
  or _62741_ (_11555_, _11554_, _11485_);
  and _62742_ (_11556_, _11555_, _06440_);
  or _62743_ (_11557_, _11556_, _01321_);
  or _62744_ (_11558_, _11557_, _11553_);
  or _62745_ (_11559_, _01317_, \oc8051_golden_model_1.TL1 [7]);
  and _62746_ (_11560_, _11559_, _43100_);
  and _62747_ (_40987_, _11560_, _11558_);
  not _62748_ (_11561_, _07803_);
  and _62749_ (_11562_, _11561_, \oc8051_golden_model_1.TL0 [7]);
  and _62750_ (_11563_, _07923_, _07803_);
  or _62751_ (_11564_, _11563_, _11562_);
  or _62752_ (_11565_, _11564_, _06132_);
  and _62753_ (_11566_, _08548_, _07803_);
  or _62754_ (_11567_, _11566_, _11562_);
  or _62755_ (_11568_, _11567_, _06161_);
  and _62756_ (_11569_, _07803_, \oc8051_golden_model_1.ACC [7]);
  or _62757_ (_11570_, _11569_, _11562_);
  and _62758_ (_11571_, _11570_, _07056_);
  and _62759_ (_11572_, _07057_, \oc8051_golden_model_1.TL0 [7]);
  or _62760_ (_11573_, _11572_, _06160_);
  or _62761_ (_11574_, _11573_, _11571_);
  and _62762_ (_11575_, _11574_, _07075_);
  and _62763_ (_11576_, _11575_, _11568_);
  and _62764_ (_11577_, _11564_, _06217_);
  or _62765_ (_11578_, _11577_, _11576_);
  and _62766_ (_11579_, _11578_, _06229_);
  and _62767_ (_11580_, _11570_, _06220_);
  or _62768_ (_11581_, _11580_, _09842_);
  or _62769_ (_11582_, _11581_, _11579_);
  and _62770_ (_11583_, _11582_, _11565_);
  or _62771_ (_11584_, _11583_, _06116_);
  and _62772_ (_11585_, _08535_, _07803_);
  or _62773_ (_11586_, _11562_, _06117_);
  or _62774_ (_11587_, _11586_, _11585_);
  and _62775_ (_11588_, _11587_, _06114_);
  and _62776_ (_11589_, _11588_, _11584_);
  and _62777_ (_11590_, _08782_, _07803_);
  or _62778_ (_11591_, _11590_, _11562_);
  and _62779_ (_11592_, _11591_, _05787_);
  or _62780_ (_11593_, _11592_, _11589_);
  or _62781_ (_11594_, _11593_, _11136_);
  and _62782_ (_11595_, _08802_, _07803_);
  or _62783_ (_11596_, _11562_, _07127_);
  or _62784_ (_11597_, _11596_, _11595_);
  and _62785_ (_11598_, _08607_, _07803_);
  or _62786_ (_11599_, _11598_, _11562_);
  or _62787_ (_11600_, _11599_, _06111_);
  and _62788_ (_11601_, _11600_, _07125_);
  and _62789_ (_11602_, _11601_, _11597_);
  and _62790_ (_11603_, _11602_, _11594_);
  and _62791_ (_11604_, _08810_, _07803_);
  or _62792_ (_11605_, _11604_, _11562_);
  and _62793_ (_11606_, _11605_, _06402_);
  or _62794_ (_11607_, _11606_, _11603_);
  and _62795_ (_11608_, _11607_, _07132_);
  or _62796_ (_11609_, _11562_, _07926_);
  and _62797_ (_11610_, _11599_, _06306_);
  and _62798_ (_11611_, _11610_, _11609_);
  or _62799_ (_11612_, _11611_, _11608_);
  and _62800_ (_11613_, _11612_, _07130_);
  and _62801_ (_11614_, _11570_, _06411_);
  and _62802_ (_11615_, _11614_, _11609_);
  or _62803_ (_11616_, _11615_, _06303_);
  or _62804_ (_11617_, _11616_, _11613_);
  and _62805_ (_11618_, _08801_, _07803_);
  or _62806_ (_11619_, _11562_, _08819_);
  or _62807_ (_11620_, _11619_, _11618_);
  and _62808_ (_11621_, _11620_, _08824_);
  and _62809_ (_11622_, _11621_, _11617_);
  nor _62810_ (_11623_, _08809_, _11561_);
  or _62811_ (_11624_, _11623_, _11562_);
  and _62812_ (_11625_, _11624_, _06396_);
  or _62813_ (_11626_, _11625_, _06433_);
  or _62814_ (_11627_, _11626_, _11622_);
  or _62815_ (_11628_, _11567_, _06829_);
  and _62816_ (_11629_, _11628_, _06444_);
  and _62817_ (_11630_, _11629_, _11627_);
  and _62818_ (_11631_, _08345_, _07803_);
  or _62819_ (_11632_, _11631_, _11562_);
  and _62820_ (_11633_, _11632_, _06440_);
  or _62821_ (_11634_, _11633_, _01321_);
  or _62822_ (_11635_, _11634_, _11630_);
  or _62823_ (_11636_, _01317_, \oc8051_golden_model_1.TL0 [7]);
  and _62824_ (_11637_, _11636_, _43100_);
  and _62825_ (_40988_, _11637_, _11635_);
  and _62826_ (_11638_, _01321_, \oc8051_golden_model_1.TCON [7]);
  not _62827_ (_11639_, _07788_);
  and _62828_ (_11640_, _11639_, \oc8051_golden_model_1.TCON [7]);
  and _62829_ (_11641_, _07923_, _07788_);
  or _62830_ (_11642_, _11641_, _11640_);
  or _62831_ (_11643_, _11642_, _06132_);
  not _62832_ (_11644_, _08407_);
  and _62833_ (_11645_, _11644_, \oc8051_golden_model_1.TCON [7]);
  and _62834_ (_11646_, _08426_, _08407_);
  or _62835_ (_11647_, _11646_, _11645_);
  and _62836_ (_11648_, _11647_, _06152_);
  and _62837_ (_11649_, _08548_, _07788_);
  or _62838_ (_11650_, _11649_, _11640_);
  or _62839_ (_11651_, _11650_, _06161_);
  and _62840_ (_11652_, _07788_, \oc8051_golden_model_1.ACC [7]);
  or _62841_ (_11653_, _11652_, _11640_);
  and _62842_ (_11654_, _11653_, _07056_);
  and _62843_ (_11655_, _07057_, \oc8051_golden_model_1.TCON [7]);
  or _62844_ (_11656_, _11655_, _06160_);
  or _62845_ (_11657_, _11656_, _11654_);
  and _62846_ (_11658_, _11657_, _06157_);
  and _62847_ (_11659_, _11658_, _11651_);
  and _62848_ (_11660_, _08552_, _08407_);
  or _62849_ (_11661_, _11660_, _11645_);
  and _62850_ (_11662_, _11661_, _06156_);
  or _62851_ (_11663_, _11662_, _06217_);
  or _62852_ (_11664_, _11663_, _11659_);
  or _62853_ (_11665_, _11642_, _07075_);
  and _62854_ (_11666_, _11665_, _11664_);
  or _62855_ (_11667_, _11666_, _06220_);
  or _62856_ (_11668_, _11653_, _06229_);
  and _62857_ (_11669_, _11668_, _06153_);
  and _62858_ (_11670_, _11669_, _11667_);
  or _62859_ (_11671_, _11670_, _11648_);
  and _62860_ (_11672_, _11671_, _06146_);
  and _62861_ (_11673_, _08569_, _08407_);
  or _62862_ (_11674_, _11673_, _11645_);
  and _62863_ (_11675_, _11674_, _06145_);
  or _62864_ (_11676_, _11675_, _11672_);
  and _62865_ (_11677_, _11676_, _06140_);
  and _62866_ (_11678_, _08587_, _08407_);
  or _62867_ (_11679_, _11678_, _11645_);
  and _62868_ (_11680_, _11679_, _06139_);
  or _62869_ (_11681_, _11680_, _09842_);
  or _62870_ (_11682_, _11681_, _11677_);
  and _62871_ (_11683_, _11682_, _11643_);
  or _62872_ (_11684_, _11683_, _06116_);
  and _62873_ (_11685_, _08535_, _07788_);
  or _62874_ (_11686_, _11640_, _06117_);
  or _62875_ (_11687_, _11686_, _11685_);
  and _62876_ (_11688_, _11687_, _06114_);
  and _62877_ (_11689_, _11688_, _11684_);
  and _62878_ (_11690_, _08782_, _07788_);
  or _62879_ (_11691_, _11690_, _11640_);
  and _62880_ (_11692_, _11691_, _05787_);
  or _62881_ (_11693_, _11692_, _11136_);
  or _62882_ (_11694_, _11693_, _11689_);
  and _62883_ (_11695_, _08802_, _07788_);
  or _62884_ (_11696_, _11640_, _07127_);
  or _62885_ (_11697_, _11696_, _11695_);
  and _62886_ (_11698_, _08607_, _07788_);
  or _62887_ (_11699_, _11698_, _11640_);
  or _62888_ (_11700_, _11699_, _06111_);
  and _62889_ (_11701_, _11700_, _07125_);
  and _62890_ (_11702_, _11701_, _11697_);
  and _62891_ (_11703_, _11702_, _11694_);
  and _62892_ (_11704_, _08810_, _07788_);
  or _62893_ (_11705_, _11704_, _11640_);
  and _62894_ (_11706_, _11705_, _06402_);
  or _62895_ (_11707_, _11706_, _11703_);
  and _62896_ (_11708_, _11707_, _07132_);
  or _62897_ (_11709_, _11640_, _07926_);
  and _62898_ (_11710_, _11699_, _06306_);
  and _62899_ (_11711_, _11710_, _11709_);
  or _62900_ (_11712_, _11711_, _11708_);
  and _62901_ (_11713_, _11712_, _07130_);
  and _62902_ (_11714_, _11653_, _06411_);
  and _62903_ (_11715_, _11714_, _11709_);
  or _62904_ (_11716_, _11715_, _06303_);
  or _62905_ (_11717_, _11716_, _11713_);
  and _62906_ (_11718_, _08801_, _07788_);
  or _62907_ (_11719_, _11640_, _08819_);
  or _62908_ (_11720_, _11719_, _11718_);
  and _62909_ (_11721_, _11720_, _08824_);
  and _62910_ (_11722_, _11721_, _11717_);
  nor _62911_ (_11723_, _08809_, _11639_);
  or _62912_ (_11724_, _11723_, _11640_);
  and _62913_ (_11725_, _11724_, _06396_);
  or _62914_ (_11726_, _11725_, _06433_);
  or _62915_ (_11727_, _11726_, _11722_);
  or _62916_ (_11728_, _11650_, _06829_);
  and _62917_ (_11729_, _11728_, _05749_);
  and _62918_ (_11730_, _11729_, _11727_);
  and _62919_ (_11731_, _11647_, _05748_);
  or _62920_ (_11732_, _11731_, _06440_);
  or _62921_ (_11733_, _11732_, _11730_);
  and _62922_ (_11734_, _08345_, _07788_);
  or _62923_ (_11735_, _11640_, _06444_);
  or _62924_ (_11736_, _11735_, _11734_);
  and _62925_ (_11737_, _11736_, _01317_);
  and _62926_ (_11738_, _11737_, _11733_);
  or _62927_ (_11739_, _11738_, _11638_);
  and _62928_ (_40989_, _11739_, _43100_);
  not _62929_ (_11740_, _07817_);
  and _62930_ (_11741_, _11740_, \oc8051_golden_model_1.TH1 [7]);
  and _62931_ (_11742_, _08548_, _07817_);
  or _62932_ (_11743_, _11742_, _11741_);
  or _62933_ (_11744_, _11743_, _06161_);
  and _62934_ (_11745_, _07817_, \oc8051_golden_model_1.ACC [7]);
  or _62935_ (_11746_, _11745_, _11741_);
  and _62936_ (_11747_, _11746_, _07056_);
  and _62937_ (_11748_, _07057_, \oc8051_golden_model_1.TH1 [7]);
  or _62938_ (_11749_, _11748_, _06160_);
  or _62939_ (_11750_, _11749_, _11747_);
  and _62940_ (_11751_, _11750_, _07075_);
  and _62941_ (_11752_, _11751_, _11744_);
  and _62942_ (_11753_, _07923_, _07817_);
  or _62943_ (_11754_, _11753_, _11741_);
  and _62944_ (_11755_, _11754_, _06217_);
  or _62945_ (_11756_, _11755_, _11752_);
  and _62946_ (_11757_, _11756_, _06229_);
  and _62947_ (_11758_, _11746_, _06220_);
  or _62948_ (_11759_, _11758_, _09842_);
  or _62949_ (_11760_, _11759_, _11757_);
  or _62950_ (_11761_, _11754_, _06132_);
  and _62951_ (_11762_, _11761_, _11760_);
  or _62952_ (_11763_, _11762_, _06116_);
  and _62953_ (_11764_, _08535_, _07817_);
  or _62954_ (_11765_, _11741_, _06117_);
  or _62955_ (_11766_, _11765_, _11764_);
  and _62956_ (_11767_, _11766_, _06114_);
  and _62957_ (_11768_, _11767_, _11763_);
  and _62958_ (_11769_, _08782_, _07817_);
  or _62959_ (_11770_, _11769_, _11741_);
  and _62960_ (_11771_, _11770_, _05787_);
  or _62961_ (_11772_, _11771_, _11768_);
  or _62962_ (_11773_, _11772_, _11136_);
  and _62963_ (_11774_, _08802_, _07817_);
  or _62964_ (_11775_, _11741_, _07127_);
  or _62965_ (_11776_, _11775_, _11774_);
  and _62966_ (_11777_, _08607_, _07817_);
  or _62967_ (_11778_, _11777_, _11741_);
  or _62968_ (_11779_, _11778_, _06111_);
  and _62969_ (_11780_, _11779_, _07125_);
  and _62970_ (_11781_, _11780_, _11776_);
  and _62971_ (_11782_, _11781_, _11773_);
  and _62972_ (_11783_, _08810_, _07817_);
  or _62973_ (_11784_, _11783_, _11741_);
  and _62974_ (_11785_, _11784_, _06402_);
  or _62975_ (_11786_, _11785_, _11782_);
  and _62976_ (_11787_, _11786_, _07132_);
  or _62977_ (_11788_, _11741_, _07926_);
  and _62978_ (_11789_, _11778_, _06306_);
  and _62979_ (_11790_, _11789_, _11788_);
  or _62980_ (_11791_, _11790_, _11787_);
  and _62981_ (_11792_, _11791_, _07130_);
  and _62982_ (_11793_, _11746_, _06411_);
  and _62983_ (_11794_, _11793_, _11788_);
  or _62984_ (_11795_, _11794_, _06303_);
  or _62985_ (_11796_, _11795_, _11792_);
  and _62986_ (_11797_, _08801_, _07817_);
  or _62987_ (_11798_, _11741_, _08819_);
  or _62988_ (_11799_, _11798_, _11797_);
  and _62989_ (_11800_, _11799_, _08824_);
  and _62990_ (_11801_, _11800_, _11796_);
  nor _62991_ (_11802_, _08809_, _11740_);
  or _62992_ (_11803_, _11802_, _11741_);
  and _62993_ (_11804_, _11803_, _06396_);
  or _62994_ (_11805_, _11804_, _06433_);
  or _62995_ (_11806_, _11805_, _11801_);
  or _62996_ (_11807_, _11743_, _06829_);
  and _62997_ (_11808_, _11807_, _06444_);
  and _62998_ (_11809_, _11808_, _11806_);
  and _62999_ (_11810_, _08345_, _07817_);
  or _63000_ (_11811_, _11810_, _11741_);
  and _63001_ (_11812_, _11811_, _06440_);
  or _63002_ (_11813_, _11812_, _01321_);
  or _63003_ (_11814_, _11813_, _11809_);
  or _63004_ (_11815_, _01317_, \oc8051_golden_model_1.TH1 [7]);
  and _63005_ (_11816_, _11815_, _43100_);
  and _63006_ (_40991_, _11816_, _11814_);
  not _63007_ (_11817_, _07823_);
  and _63008_ (_11818_, _11817_, \oc8051_golden_model_1.TH0 [7]);
  and _63009_ (_11819_, _08548_, _07823_);
  or _63010_ (_11820_, _11819_, _11818_);
  or _63011_ (_11821_, _11820_, _06161_);
  and _63012_ (_11822_, _07823_, \oc8051_golden_model_1.ACC [7]);
  or _63013_ (_11823_, _11822_, _11818_);
  and _63014_ (_11824_, _11823_, _07056_);
  and _63015_ (_11825_, _07057_, \oc8051_golden_model_1.TH0 [7]);
  or _63016_ (_11826_, _11825_, _06160_);
  or _63017_ (_11827_, _11826_, _11824_);
  and _63018_ (_11828_, _11827_, _07075_);
  and _63019_ (_11829_, _11828_, _11821_);
  and _63020_ (_11830_, _07923_, _07823_);
  or _63021_ (_11831_, _11830_, _11818_);
  and _63022_ (_11832_, _11831_, _06217_);
  or _63023_ (_11833_, _11832_, _11829_);
  and _63024_ (_11834_, _11833_, _06229_);
  and _63025_ (_11835_, _11823_, _06220_);
  or _63026_ (_11836_, _11835_, _09842_);
  or _63027_ (_11837_, _11836_, _11834_);
  or _63028_ (_11838_, _11831_, _06132_);
  and _63029_ (_11839_, _11838_, _11837_);
  or _63030_ (_11840_, _11839_, _06116_);
  and _63031_ (_11841_, _08535_, _07823_);
  or _63032_ (_11842_, _11818_, _06117_);
  or _63033_ (_11843_, _11842_, _11841_);
  and _63034_ (_11844_, _11843_, _06114_);
  and _63035_ (_11845_, _11844_, _11840_);
  and _63036_ (_11846_, _08782_, _07823_);
  or _63037_ (_11847_, _11846_, _11818_);
  and _63038_ (_11848_, _11847_, _05787_);
  or _63039_ (_11849_, _11848_, _11845_);
  or _63040_ (_11850_, _11849_, _11136_);
  and _63041_ (_11851_, _08802_, _07823_);
  or _63042_ (_11852_, _11818_, _07127_);
  or _63043_ (_11853_, _11852_, _11851_);
  and _63044_ (_11854_, _08607_, _07823_);
  or _63045_ (_11855_, _11854_, _11818_);
  or _63046_ (_11856_, _11855_, _06111_);
  and _63047_ (_11857_, _11856_, _07125_);
  and _63048_ (_11858_, _11857_, _11853_);
  and _63049_ (_11859_, _11858_, _11850_);
  and _63050_ (_11860_, _08810_, _07823_);
  or _63051_ (_11861_, _11860_, _11818_);
  and _63052_ (_11862_, _11861_, _06402_);
  or _63053_ (_11863_, _11862_, _11859_);
  and _63054_ (_11864_, _11863_, _07132_);
  or _63055_ (_11865_, _11818_, _07926_);
  and _63056_ (_11866_, _11855_, _06306_);
  and _63057_ (_11867_, _11866_, _11865_);
  or _63058_ (_11868_, _11867_, _11864_);
  and _63059_ (_11869_, _11868_, _07130_);
  and _63060_ (_11870_, _11823_, _06411_);
  and _63061_ (_11871_, _11870_, _11865_);
  or _63062_ (_11872_, _11871_, _06303_);
  or _63063_ (_11873_, _11872_, _11869_);
  and _63064_ (_11874_, _08801_, _07823_);
  or _63065_ (_11875_, _11818_, _08819_);
  or _63066_ (_11876_, _11875_, _11874_);
  and _63067_ (_11877_, _11876_, _08824_);
  and _63068_ (_11878_, _11877_, _11873_);
  nor _63069_ (_11879_, _08809_, _11817_);
  or _63070_ (_11880_, _11879_, _11818_);
  and _63071_ (_11881_, _11880_, _06396_);
  or _63072_ (_11882_, _11881_, _06433_);
  or _63073_ (_11883_, _11882_, _11878_);
  or _63074_ (_11884_, _11820_, _06829_);
  and _63075_ (_11885_, _11884_, _06444_);
  and _63076_ (_11886_, _11885_, _11883_);
  and _63077_ (_11887_, _08345_, _07823_);
  or _63078_ (_11888_, _11887_, _11818_);
  and _63079_ (_11889_, _11888_, _06440_);
  or _63080_ (_11890_, _11889_, _01321_);
  or _63081_ (_11891_, _11890_, _11886_);
  or _63082_ (_11892_, _01317_, \oc8051_golden_model_1.TH0 [7]);
  and _63083_ (_11893_, _11892_, _43100_);
  and _63084_ (_40992_, _11893_, _11891_);
  and _63085_ (_11894_, _08433_, _05426_);
  and _63086_ (_11895_, _11894_, \oc8051_golden_model_1.PC [7]);
  and _63087_ (_11896_, _11895_, _09231_);
  and _63088_ (_11897_, _11896_, \oc8051_golden_model_1.PC [10]);
  and _63089_ (_11898_, _11897_, \oc8051_golden_model_1.PC [11]);
  and _63090_ (_11899_, _11898_, \oc8051_golden_model_1.PC [12]);
  and _63091_ (_11900_, _11899_, \oc8051_golden_model_1.PC [13]);
  and _63092_ (_11901_, _11900_, \oc8051_golden_model_1.PC [14]);
  or _63093_ (_11902_, _11901_, \oc8051_golden_model_1.PC [15]);
  nand _63094_ (_11903_, _11901_, \oc8051_golden_model_1.PC [15]);
  and _63095_ (_11904_, _11903_, _11902_);
  and _63096_ (_11905_, _11041_, _10963_);
  or _63097_ (_11906_, _11905_, _11904_);
  and _63098_ (_11907_, _10867_, _10380_);
  or _63099_ (_11908_, _11907_, _11904_);
  nor _63100_ (_11909_, _08441_, _06783_);
  not _63101_ (_11910_, _11909_);
  nor _63102_ (_11911_, _10841_, _10835_);
  and _63103_ (_11912_, _11911_, _11910_);
  or _63104_ (_11913_, _11912_, _11904_);
  and _63105_ (_11914_, _10816_, _10808_);
  or _63106_ (_11915_, _11914_, _11904_);
  nor _63107_ (_11916_, _10787_, _06400_);
  not _63108_ (_11917_, _11916_);
  nor _63109_ (_11918_, _10778_, _10768_);
  and _63110_ (_11919_, _11918_, _10762_);
  or _63111_ (_11920_, _11919_, _11904_);
  or _63112_ (_11921_, _09256_, _08787_);
  nor _63113_ (_11922_, _09855_, _05801_);
  and _63114_ (_11923_, _09239_, _05787_);
  nor _63115_ (_11924_, _05799_, _05758_);
  not _63116_ (_11925_, _11924_);
  or _63117_ (_11926_, _09210_, _06070_);
  or _63118_ (_11927_, _09025_, _06228_);
  and _63119_ (_11928_, _11927_, _11926_);
  or _63120_ (_11929_, _09211_, _06625_);
  or _63121_ (_11930_, _09070_, _06626_);
  and _63122_ (_11931_, _11930_, _11929_);
  and _63123_ (_11932_, _11931_, _11928_);
  nand _63124_ (_11933_, _09160_, _06107_);
  or _63125_ (_11934_, _09115_, _06912_);
  nor _63126_ (_11935_, _09114_, _09092_);
  or _63127_ (_11936_, _11935_, _06913_);
  and _63128_ (_11937_, _11936_, _11934_);
  and _63129_ (_11938_, _11937_, _11933_);
  and _63130_ (_11939_, _11938_, _11932_);
  or _63131_ (_11940_, _09160_, _06107_);
  and _63132_ (_11941_, _08838_, _06039_);
  nor _63133_ (_11942_, _11941_, _08581_);
  or _63134_ (_11943_, _09207_, _06203_);
  or _63135_ (_11944_, _08883_, _07482_);
  and _63136_ (_11945_, _11944_, _11943_);
  and _63137_ (_11946_, _11945_, _11942_);
  or _63138_ (_11947_, _08931_, _07805_);
  or _63139_ (_11948_, _09208_, _06477_);
  and _63140_ (_11949_, _11948_, _11947_);
  or _63141_ (_11950_, _08980_, _07775_);
  or _63142_ (_11951_, _09209_, _06876_);
  and _63143_ (_11952_, _11951_, _11950_);
  and _63144_ (_11953_, _11952_, _11949_);
  and _63145_ (_11954_, _11953_, _11946_);
  and _63146_ (_11955_, _11954_, _11940_);
  nand _63147_ (_11956_, _11955_, _11939_);
  or _63148_ (_11957_, _11956_, _09239_);
  and _63149_ (_11958_, _11955_, _11939_);
  and _63150_ (_11959_, _09242_, _09178_);
  and _63151_ (_11960_, _11959_, \oc8051_golden_model_1.PC [11]);
  and _63152_ (_11961_, _11960_, \oc8051_golden_model_1.PC [12]);
  and _63153_ (_11962_, _11961_, \oc8051_golden_model_1.PC [13]);
  and _63154_ (_11963_, _11962_, \oc8051_golden_model_1.PC [14]);
  nor _63155_ (_11964_, _11962_, \oc8051_golden_model_1.PC [14]);
  nor _63156_ (_11965_, _11964_, _11963_);
  not _63157_ (_11966_, _11965_);
  nor _63158_ (_11967_, _11966_, _08395_);
  and _63159_ (_11968_, _11966_, _08395_);
  nor _63160_ (_11969_, _11968_, _11967_);
  not _63161_ (_11970_, _11969_);
  nor _63162_ (_11971_, _11961_, \oc8051_golden_model_1.PC [13]);
  nor _63163_ (_11972_, _11971_, _11962_);
  not _63164_ (_11973_, _11972_);
  nor _63165_ (_11974_, _11973_, _08395_);
  and _63166_ (_11975_, _11973_, _08395_);
  nor _63167_ (_11976_, _11960_, \oc8051_golden_model_1.PC [12]);
  nor _63168_ (_11977_, _11976_, _11961_);
  not _63169_ (_11978_, _11977_);
  nor _63170_ (_11979_, _11978_, _08395_);
  nor _63171_ (_11980_, _11959_, \oc8051_golden_model_1.PC [11]);
  nor _63172_ (_11981_, _11980_, _11960_);
  not _63173_ (_11982_, _11981_);
  nor _63174_ (_11983_, _11982_, _08395_);
  and _63175_ (_11984_, _11982_, _08395_);
  nor _63176_ (_11985_, _11984_, _11983_);
  and _63177_ (_11986_, _09231_, _09178_);
  nor _63178_ (_11987_, _11986_, \oc8051_golden_model_1.PC [10]);
  nor _63179_ (_11988_, _11987_, _11959_);
  not _63180_ (_11989_, _11988_);
  nor _63181_ (_11990_, _11989_, _08395_);
  and _63182_ (_11991_, _11989_, _08395_);
  nor _63183_ (_11992_, _11991_, _11990_);
  and _63184_ (_11993_, _11992_, _11985_);
  and _63185_ (_11994_, _09178_, \oc8051_golden_model_1.PC [8]);
  nor _63186_ (_11995_, _11994_, \oc8051_golden_model_1.PC [9]);
  nor _63187_ (_11996_, _11995_, _11986_);
  not _63188_ (_11997_, _11996_);
  nor _63189_ (_11998_, _11997_, _08395_);
  and _63190_ (_11999_, _11997_, _08395_);
  nor _63191_ (_12000_, _11999_, _11998_);
  nor _63192_ (_12001_, _09181_, _08395_);
  and _63193_ (_12002_, _09181_, _08395_);
  and _63194_ (_12003_, _09176_, _08432_);
  nor _63195_ (_12004_, _12003_, \oc8051_golden_model_1.PC [6]);
  nor _63196_ (_12005_, _12004_, _09177_);
  not _63197_ (_12006_, _12005_);
  nor _63198_ (_12007_, _12006_, _08638_);
  and _63199_ (_12008_, _12006_, _08638_);
  nor _63200_ (_12009_, _12008_, _12007_);
  not _63201_ (_12010_, _12009_);
  and _63202_ (_12011_, _09176_, \oc8051_golden_model_1.PC [4]);
  nor _63203_ (_12012_, _12011_, \oc8051_golden_model_1.PC [5]);
  nor _63204_ (_12013_, _12012_, _12003_);
  not _63205_ (_12014_, _12013_);
  nor _63206_ (_12015_, _12014_, _08701_);
  and _63207_ (_12016_, _12014_, _08701_);
  nor _63208_ (_12017_, _09176_, \oc8051_golden_model_1.PC [4]);
  nor _63209_ (_12018_, _12017_, _12011_);
  not _63210_ (_12019_, _12018_);
  nor _63211_ (_12020_, _12019_, _08670_);
  and _63212_ (_12021_, _05449_, \oc8051_golden_model_1.PC [2]);
  nor _63213_ (_12022_, _12021_, \oc8051_golden_model_1.PC [3]);
  nor _63214_ (_12023_, _12022_, _09176_);
  not _63215_ (_12024_, _12023_);
  nor _63216_ (_12025_, _12024_, _06389_);
  and _63217_ (_12026_, _12024_, _06389_);
  nor _63218_ (_12027_, _05449_, \oc8051_golden_model_1.PC [2]);
  nor _63219_ (_12028_, _12027_, _12021_);
  not _63220_ (_12029_, _12028_);
  nor _63221_ (_12030_, _12029_, _06521_);
  nor _63222_ (_12031_, _06945_, _05879_);
  nor _63223_ (_12032_, _06758_, \oc8051_golden_model_1.PC [0]);
  and _63224_ (_12033_, _06945_, _05879_);
  nor _63225_ (_12034_, _12033_, _12031_);
  and _63226_ (_12035_, _12034_, _12032_);
  nor _63227_ (_12036_, _12035_, _12031_);
  and _63228_ (_12037_, _12029_, _06521_);
  nor _63229_ (_12038_, _12037_, _12030_);
  not _63230_ (_12039_, _12038_);
  nor _63231_ (_12040_, _12039_, _12036_);
  nor _63232_ (_12041_, _12040_, _12030_);
  nor _63233_ (_12042_, _12041_, _12026_);
  nor _63234_ (_12043_, _12042_, _12025_);
  and _63235_ (_12044_, _12019_, _08670_);
  nor _63236_ (_12045_, _12044_, _12020_);
  not _63237_ (_12046_, _12045_);
  nor _63238_ (_12047_, _12046_, _12043_);
  nor _63239_ (_12048_, _12047_, _12020_);
  nor _63240_ (_12049_, _12048_, _12016_);
  nor _63241_ (_12050_, _12049_, _12015_);
  nor _63242_ (_12051_, _12050_, _12010_);
  nor _63243_ (_12052_, _12051_, _12007_);
  nor _63244_ (_12053_, _12052_, _12002_);
  or _63245_ (_12054_, _12053_, _12001_);
  nor _63246_ (_12055_, _09178_, \oc8051_golden_model_1.PC [8]);
  nor _63247_ (_12056_, _12055_, _11994_);
  not _63248_ (_12057_, _12056_);
  nor _63249_ (_12058_, _12057_, _08395_);
  and _63250_ (_12059_, _12057_, _08395_);
  nor _63251_ (_12060_, _12059_, _12058_);
  and _63252_ (_12061_, _12060_, _12054_);
  and _63253_ (_12062_, _12061_, _12000_);
  and _63254_ (_12063_, _12062_, _11993_);
  nor _63255_ (_12064_, _12058_, _11998_);
  not _63256_ (_12065_, _12064_);
  and _63257_ (_12066_, _12065_, _11993_);
  or _63258_ (_12067_, _12066_, _11990_);
  or _63259_ (_12068_, _12067_, _12063_);
  nor _63260_ (_12069_, _12068_, _11983_);
  and _63261_ (_12070_, _11978_, _08395_);
  nor _63262_ (_12071_, _12070_, _11979_);
  not _63263_ (_12072_, _12071_);
  nor _63264_ (_12073_, _12072_, _12069_);
  nor _63265_ (_12074_, _12073_, _11979_);
  nor _63266_ (_12075_, _12074_, _11975_);
  nor _63267_ (_12076_, _12075_, _11974_);
  nor _63268_ (_12077_, _12076_, _11970_);
  nor _63269_ (_12078_, _12077_, _11967_);
  and _63270_ (_12079_, _09240_, _08395_);
  nor _63271_ (_12080_, _09240_, _08395_);
  nor _63272_ (_12081_, _12080_, _12079_);
  and _63273_ (_12082_, _12081_, _12078_);
  nor _63274_ (_12083_, _12081_, _12078_);
  nor _63275_ (_12084_, _12083_, _12082_);
  not _63276_ (_12085_, _12084_);
  or _63277_ (_12086_, _12085_, _11958_);
  and _63278_ (_12087_, _12086_, _06687_);
  and _63279_ (_12088_, _12087_, _11957_);
  not _63280_ (_12089_, _06687_);
  nor _63281_ (_12090_, _07049_, _06107_);
  not _63282_ (_12091_, _12090_);
  and _63283_ (_12092_, _09194_, _06039_);
  and _63284_ (_12093_, _08347_, _07482_);
  nor _63285_ (_12094_, _12093_, _12092_);
  and _63286_ (_12095_, _08012_, _06203_);
  and _63287_ (_12096_, _08101_, _06477_);
  nor _63288_ (_12097_, _12096_, _12095_);
  and _63289_ (_12098_, _12097_, _12094_);
  and _63290_ (_12099_, _08348_, _07805_);
  and _63291_ (_12100_, _08349_, _07775_);
  nor _63292_ (_12101_, _12100_, _12099_);
  and _63293_ (_12102_, _08336_, _06876_);
  nor _63294_ (_12103_, _12102_, _07924_);
  and _63295_ (_12104_, _12103_, _12101_);
  and _63296_ (_12105_, _12104_, _12098_);
  and _63297_ (_12106_, _07474_, _06228_);
  and _63298_ (_12107_, _07544_, _06070_);
  nor _63299_ (_12108_, _12107_, _12106_);
  and _63300_ (_12109_, _07657_, _06626_);
  and _63301_ (_12110_, _07708_, _06625_);
  nor _63302_ (_12111_, _12110_, _12109_);
  and _63303_ (_12112_, _12111_, _12108_);
  and _63304_ (_12113_, _07252_, _06913_);
  and _63305_ (_12114_, _07306_, _06912_);
  and _63306_ (_12115_, _07049_, _06107_);
  or _63307_ (_12116_, _12115_, _12114_);
  nor _63308_ (_12117_, _12116_, _12113_);
  and _63309_ (_12118_, _12117_, _12112_);
  and _63310_ (_12119_, _12118_, _12105_);
  and _63311_ (_12120_, _12119_, _12091_);
  nand _63312_ (_12121_, _12120_, _09240_);
  nand _63313_ (_12122_, _06125_, _06144_);
  and _63314_ (_12123_, _06119_, _06144_);
  nor _63315_ (_12124_, _12123_, _06290_);
  and _63316_ (_12125_, _12124_, _12122_);
  not _63317_ (_12126_, _12125_);
  or _63318_ (_12127_, _12120_, _12085_);
  and _63319_ (_12128_, _12127_, _12126_);
  and _63320_ (_12129_, _12128_, _12121_);
  and _63321_ (_12130_, _09256_, _06220_);
  and _63322_ (_12131_, _06221_, _05764_);
  or _63323_ (_12132_, _12131_, _09256_);
  nor _63324_ (_12133_, _05799_, _05762_);
  nor _63325_ (_12134_, _12133_, _10490_);
  and _63326_ (_12135_, _08211_, _08175_);
  and _63327_ (_12136_, _08542_, _12135_);
  and _63328_ (_12137_, _08014_, _07925_);
  and _63329_ (_12138_, _12137_, _08539_);
  nand _63330_ (_12139_, _12138_, _12136_);
  or _63331_ (_12140_, _12139_, _09239_);
  and _63332_ (_12141_, _12138_, _12136_);
  or _63333_ (_12142_, _12141_, _12085_);
  and _63334_ (_12143_, _12142_, _06160_);
  and _63335_ (_12144_, _12143_, _12140_);
  nor _63336_ (_12145_, _09246_, \oc8051_golden_model_1.PC [14]);
  nor _63337_ (_12146_, _12145_, _09247_);
  and _63338_ (_12147_, _12146_, _06039_);
  nor _63339_ (_12148_, _12146_, _06039_);
  nor _63340_ (_12149_, _12148_, _12147_);
  not _63341_ (_12150_, _12149_);
  nor _63342_ (_12151_, _09245_, \oc8051_golden_model_1.PC [13]);
  nor _63343_ (_12152_, _12151_, _09246_);
  and _63344_ (_12153_, _12152_, _06039_);
  nor _63345_ (_12154_, _12152_, _06039_);
  nor _63346_ (_12155_, _09244_, \oc8051_golden_model_1.PC [12]);
  nor _63347_ (_12156_, _12155_, _09245_);
  and _63348_ (_12157_, _12156_, _06039_);
  nor _63349_ (_12158_, _09249_, \oc8051_golden_model_1.PC [10]);
  nor _63350_ (_12159_, _12158_, _09250_);
  and _63351_ (_12160_, _12159_, _06039_);
  not _63352_ (_12161_, _12160_);
  nor _63353_ (_12162_, _09250_, \oc8051_golden_model_1.PC [11]);
  nor _63354_ (_12163_, _12162_, _09251_);
  and _63355_ (_12164_, _12163_, _06039_);
  nor _63356_ (_12165_, _12163_, _06039_);
  nor _63357_ (_12166_, _12165_, _12164_);
  nor _63358_ (_12167_, _12159_, _06039_);
  nor _63359_ (_12168_, _12167_, _12160_);
  and _63360_ (_12169_, _12168_, _12166_);
  and _63361_ (_12170_, _08435_, \oc8051_golden_model_1.PC [8]);
  nor _63362_ (_12171_, _12170_, \oc8051_golden_model_1.PC [9]);
  nor _63363_ (_12172_, _12171_, _09249_);
  and _63364_ (_12173_, _12172_, _06039_);
  nor _63365_ (_12174_, _12172_, _06039_);
  nor _63366_ (_12175_, _12174_, _12173_);
  and _63367_ (_12176_, _08437_, _06039_);
  nor _63368_ (_12177_, _08437_, _06039_);
  and _63369_ (_12178_, _08432_, _05972_);
  nor _63370_ (_12179_, _12178_, \oc8051_golden_model_1.PC [6]);
  nor _63371_ (_12180_, _12179_, _08434_);
  not _63372_ (_12181_, _12180_);
  nor _63373_ (_12182_, _12181_, _06203_);
  and _63374_ (_12183_, _12181_, _06203_);
  nor _63375_ (_12184_, _12183_, _12182_);
  not _63376_ (_12185_, _12184_);
  and _63377_ (_12186_, _05972_, \oc8051_golden_model_1.PC [4]);
  nor _63378_ (_12187_, _12186_, \oc8051_golden_model_1.PC [5]);
  nor _63379_ (_12188_, _12187_, _12178_);
  not _63380_ (_12189_, _12188_);
  nor _63381_ (_12190_, _12189_, _06477_);
  and _63382_ (_12191_, _12189_, _06477_);
  nor _63383_ (_12192_, _05972_, \oc8051_golden_model_1.PC [4]);
  nor _63384_ (_12193_, _12192_, _12186_);
  not _63385_ (_12194_, _12193_);
  nor _63386_ (_12195_, _12194_, _06876_);
  nor _63387_ (_12196_, _06070_, _06322_);
  and _63388_ (_12197_, _06070_, _06322_);
  nor _63389_ (_12198_, _06625_, _05923_);
  nor _63390_ (_12199_, _06912_, \oc8051_golden_model_1.PC [1]);
  nor _63391_ (_12200_, _06107_, _05444_);
  and _63392_ (_12201_, _06912_, \oc8051_golden_model_1.PC [1]);
  nor _63393_ (_12202_, _12201_, _12199_);
  and _63394_ (_12203_, _12202_, _12200_);
  nor _63395_ (_12204_, _12203_, _12199_);
  and _63396_ (_12205_, _06625_, _05923_);
  nor _63397_ (_12206_, _12205_, _12198_);
  not _63398_ (_12207_, _12206_);
  nor _63399_ (_12208_, _12207_, _12204_);
  nor _63400_ (_12209_, _12208_, _12198_);
  nor _63401_ (_12210_, _12209_, _12197_);
  nor _63402_ (_12211_, _12210_, _12196_);
  and _63403_ (_12212_, _12194_, _06876_);
  nor _63404_ (_12213_, _12212_, _12195_);
  not _63405_ (_12214_, _12213_);
  nor _63406_ (_12215_, _12214_, _12211_);
  nor _63407_ (_12216_, _12215_, _12195_);
  nor _63408_ (_12217_, _12216_, _12191_);
  nor _63409_ (_12218_, _12217_, _12190_);
  nor _63410_ (_12219_, _12218_, _12185_);
  nor _63411_ (_12220_, _12219_, _12182_);
  nor _63412_ (_12221_, _12220_, _12177_);
  or _63413_ (_12222_, _12221_, _12176_);
  nor _63414_ (_12223_, _08435_, \oc8051_golden_model_1.PC [8]);
  nor _63415_ (_12224_, _12223_, _12170_);
  and _63416_ (_12225_, _12224_, _06039_);
  nor _63417_ (_12226_, _12224_, _06039_);
  nor _63418_ (_12227_, _12226_, _12225_);
  and _63419_ (_12228_, _12227_, _12222_);
  and _63420_ (_12229_, _12228_, _12175_);
  and _63421_ (_12230_, _12229_, _12169_);
  nor _63422_ (_12231_, _12225_, _12173_);
  not _63423_ (_12232_, _12231_);
  and _63424_ (_12233_, _12232_, _12169_);
  or _63425_ (_12234_, _12233_, _12164_);
  nor _63426_ (_12235_, _12234_, _12230_);
  and _63427_ (_12236_, _12235_, _12161_);
  nor _63428_ (_12237_, _12156_, _06039_);
  nor _63429_ (_12238_, _12237_, _12157_);
  not _63430_ (_12239_, _12238_);
  nor _63431_ (_12240_, _12239_, _12236_);
  nor _63432_ (_12241_, _12240_, _12157_);
  nor _63433_ (_12242_, _12241_, _12154_);
  nor _63434_ (_12243_, _12242_, _12153_);
  nor _63435_ (_12244_, _12243_, _12150_);
  nor _63436_ (_12245_, _12244_, _12147_);
  nor _63437_ (_12246_, _09256_, _06039_);
  and _63438_ (_12247_, _09256_, _06039_);
  nor _63439_ (_12248_, _12247_, _12246_);
  and _63440_ (_12249_, _12248_, _12245_);
  nor _63441_ (_12250_, _12248_, _12245_);
  or _63442_ (_12251_, _12250_, _12249_);
  and _63443_ (_12252_, _07252_, _07049_);
  and _63444_ (_12253_, _08347_, _09194_);
  and _63445_ (_12254_, _12253_, _12252_);
  and _63446_ (_12255_, _08351_, _08350_);
  nand _63447_ (_12256_, _12255_, _12254_);
  and _63448_ (_12257_, _12256_, _12251_);
  and _63449_ (_12258_, _12255_, _12254_);
  and _63450_ (_12259_, _12258_, _09256_);
  or _63451_ (_12260_, _12259_, _08443_);
  or _63452_ (_12261_, _12260_, _12257_);
  nor _63453_ (_12262_, _10473_, _10483_);
  and _63454_ (_12263_, _12262_, _10471_);
  not _63455_ (_12264_, _06653_);
  nor _63456_ (_12265_, _07382_, _07372_);
  and _63457_ (_12266_, _12265_, _12264_);
  and _63458_ (_12267_, _12266_, _12263_);
  not _63459_ (_12268_, _12267_);
  and _63460_ (_12269_, _12268_, _11904_);
  and _63461_ (_12270_, _09256_, _06581_);
  and _63462_ (_12271_, _09256_, _07056_);
  nor _63463_ (_12272_, _06581_, _09229_);
  and _63464_ (_12273_, _12272_, _07057_);
  and _63465_ (_12274_, _12273_, _12265_);
  or _63466_ (_12275_, _12274_, _12271_);
  and _63467_ (_12276_, _12275_, _12264_);
  or _63468_ (_12277_, _12276_, _12270_);
  and _63469_ (_12278_, _12277_, _12263_);
  or _63470_ (_12279_, _12278_, _08445_);
  or _63471_ (_12280_, _12279_, _12269_);
  nor _63472_ (_12281_, _07064_, _06160_);
  and _63473_ (_12282_, _12281_, _12280_);
  and _63474_ (_12283_, _12282_, _12261_);
  or _63475_ (_12284_, _12283_, _12144_);
  and _63476_ (_12285_, _12284_, _12134_);
  not _63477_ (_12286_, _12131_);
  nand _63478_ (_12287_, _12134_, _07065_);
  and _63479_ (_12288_, _12287_, _11904_);
  or _63480_ (_12289_, _12288_, _12286_);
  or _63481_ (_12290_, _12289_, _12285_);
  and _63482_ (_12291_, _12290_, _12132_);
  and _63483_ (_12292_, _10458_, _07082_);
  not _63484_ (_12293_, _12292_);
  or _63485_ (_12294_, _12293_, _12291_);
  or _63486_ (_12295_, _12292_, _11904_);
  and _63487_ (_12296_, _12295_, _06229_);
  and _63488_ (_12297_, _12296_, _12294_);
  or _63489_ (_12298_, _12297_, _12130_);
  nor _63490_ (_12299_, _05799_, _05768_);
  nor _63491_ (_12300_, _12299_, _10525_);
  and _63492_ (_12301_, _12300_, _12298_);
  not _63493_ (_12302_, _12300_);
  and _63494_ (_12303_, _12302_, _11904_);
  not _63495_ (_12304_, _05769_);
  nor _63496_ (_12305_, _06151_, _12304_);
  and _63497_ (_12306_, _12305_, _06153_);
  not _63498_ (_12307_, _12306_);
  or _63499_ (_12308_, _12307_, _12303_);
  or _63500_ (_12309_, _12308_, _12301_);
  or _63501_ (_12310_, _12306_, _09256_);
  and _63502_ (_12311_, _12310_, _12125_);
  and _63503_ (_12312_, _12311_, _12309_);
  or _63504_ (_12313_, _12312_, _12129_);
  and _63505_ (_12314_, _12313_, _12089_);
  or _63506_ (_12315_, _12314_, _06236_);
  or _63507_ (_12316_, _12315_, _12088_);
  not _63508_ (_12317_, _06295_);
  nor _63509_ (_12318_, _10273_, _10272_);
  nor _63510_ (_12319_, _12318_, _10282_);
  not _63511_ (_12320_, _10278_);
  nor _63512_ (_12321_, _08211_, \oc8051_golden_model_1.ACC [0]);
  or _63513_ (_12322_, _12321_, _10276_);
  and _63514_ (_12323_, _12322_, _12320_);
  and _63515_ (_12324_, _12323_, _12319_);
  nor _63516_ (_12325_, _10268_, _10269_);
  nor _63517_ (_12326_, _12325_, _10289_);
  nor _63518_ (_12327_, _10295_, _08810_);
  and _63519_ (_12328_, _12327_, _12326_);
  and _63520_ (_12329_, _12328_, _12324_);
  and _63521_ (_12330_, _12329_, _09239_);
  nor _63522_ (_12331_, _12329_, _12084_);
  or _63523_ (_12332_, _12331_, _06643_);
  or _63524_ (_12333_, _12332_, _12330_);
  and _63525_ (_12334_, _12333_, _12317_);
  and _63526_ (_12335_, _12334_, _12316_);
  nor _63527_ (_12336_, _11059_, _11060_);
  nor _63528_ (_12337_, _12336_, _11063_);
  and _63529_ (_12338_, _06107_, _05855_);
  nor _63530_ (_12339_, _12338_, _11067_);
  nor _63531_ (_12340_, _12339_, _11066_);
  and _63532_ (_12341_, _12340_, _12337_);
  nor _63533_ (_12342_, _11053_, _11054_);
  nor _63534_ (_12343_, _12342_, _11058_);
  nor _63535_ (_12344_, _11052_, _10794_);
  and _63536_ (_12345_, _12344_, _12343_);
  and _63537_ (_12346_, _12345_, _12341_);
  not _63538_ (_12347_, _12346_);
  nand _63539_ (_12348_, _12347_, _12084_);
  nand _63540_ (_12349_, _12346_, _09240_);
  and _63541_ (_12350_, _12349_, _06295_);
  and _63542_ (_12351_, _12350_, _12348_);
  or _63543_ (_12352_, _12351_, _12335_);
  and _63544_ (_12353_, _12352_, _11925_);
  nand _63545_ (_12354_, _11924_, _11904_);
  and _63546_ (_12355_, _06124_, _06245_);
  nor _63547_ (_12356_, _12355_, _06212_);
  nor _63548_ (_12357_, _06701_, _07388_);
  and _63549_ (_12358_, _06128_, _06245_);
  not _63550_ (_12359_, _12358_);
  nor _63551_ (_12360_, _07292_, _06145_);
  and _63552_ (_12361_, _12360_, _12359_);
  and _63553_ (_12362_, _12361_, _12357_);
  and _63554_ (_12363_, _12362_, _12356_);
  nand _63555_ (_12364_, _12363_, _12354_);
  or _63556_ (_12365_, _12364_, _12353_);
  and _63557_ (_12366_, _05786_, _06245_);
  not _63558_ (_12367_, _12366_);
  nor _63559_ (_12368_, _11311_, _09295_);
  and _63560_ (_12369_, _12368_, _12367_);
  or _63561_ (_12370_, _12363_, _09256_);
  and _63562_ (_12371_, _12370_, _12369_);
  and _63563_ (_12372_, _12371_, _12365_);
  not _63564_ (_12373_, _12369_);
  and _63565_ (_12374_, _12373_, _11904_);
  and _63566_ (_12375_, _06256_, _05775_);
  not _63567_ (_12376_, _12375_);
  or _63568_ (_12377_, _12376_, _12374_);
  or _63569_ (_12378_, _12377_, _12372_);
  and _63570_ (_12379_, _06115_, _05790_);
  not _63571_ (_12380_, _12379_);
  and _63572_ (_12381_, _10554_, _12380_);
  or _63573_ (_12382_, _12375_, _09256_);
  and _63574_ (_12383_, _12382_, _12381_);
  and _63575_ (_12384_, _12383_, _12378_);
  nor _63576_ (_12385_, _10387_, _06260_);
  not _63577_ (_12386_, _12385_);
  not _63578_ (_12387_, _12381_);
  and _63579_ (_12388_, _12387_, _11904_);
  or _63580_ (_12389_, _12388_, _12386_);
  or _63581_ (_12390_, _12389_, _12384_);
  or _63582_ (_12391_, _12385_, _09256_);
  and _63583_ (_12392_, _12391_, _05805_);
  and _63584_ (_12393_, _12392_, _12390_);
  and _63585_ (_12394_, _11904_, _05870_);
  nor _63586_ (_12395_, _06139_, _05791_);
  not _63587_ (_12396_, _12395_);
  or _63588_ (_12397_, _12396_, _12394_);
  or _63589_ (_12398_, _12397_, _12393_);
  or _63590_ (_12399_, _12395_, _09256_);
  and _63591_ (_12400_, _12399_, _11296_);
  and _63592_ (_12401_, _12400_, _12398_);
  nand _63593_ (_12402_, _09239_, _06293_);
  nand _63594_ (_12403_, _12402_, _06133_);
  or _63595_ (_12404_, _12403_, _12401_);
  or _63596_ (_12405_, _09256_, _06133_);
  and _63597_ (_12406_, _12405_, _06114_);
  and _63598_ (_12407_, _12406_, _12404_);
  or _63599_ (_12408_, _12407_, _11923_);
  and _63600_ (_12409_, _12408_, _11922_);
  nor _63601_ (_12410_, _06209_, _05829_);
  not _63602_ (_12411_, _12410_);
  not _63603_ (_12412_, _11922_);
  and _63604_ (_12413_, _12412_, _11904_);
  or _63605_ (_12414_, _12413_, _12411_);
  or _63606_ (_12415_, _12414_, _12409_);
  and _63607_ (_12416_, _05781_, _05746_);
  not _63608_ (_12417_, _12416_);
  or _63609_ (_12418_, _12410_, _09256_);
  and _63610_ (_12419_, _12418_, _12417_);
  and _63611_ (_12420_, _12419_, _12415_);
  and _63612_ (_12421_, _12416_, _12251_);
  or _63613_ (_12422_, _12421_, _08788_);
  or _63614_ (_12423_, _12422_, _12420_);
  and _63615_ (_12424_, _12423_, _11921_);
  or _63616_ (_12425_, _12424_, _06110_);
  nand _63617_ (_12426_, _09240_, _06110_);
  and _63618_ (_12427_, _12426_, _10752_);
  and _63619_ (_12428_, _12427_, _12425_);
  and _63620_ (_12429_, _10751_, _09256_);
  or _63621_ (_12430_, _12429_, _12428_);
  nor _63622_ (_12431_, _05835_, _05799_);
  not _63623_ (_12432_, _12431_);
  and _63624_ (_12433_, _12432_, _12430_);
  not _63625_ (_12434_, \oc8051_golden_model_1.DPH [0]);
  and _63626_ (_12435_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor _63627_ (_12436_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and _63628_ (_12437_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _63629_ (_12438_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _63630_ (_12439_, _12438_, _12437_);
  not _63631_ (_12440_, _12439_);
  and _63632_ (_12441_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _63633_ (_12442_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _63634_ (_12443_, _12442_, _12441_);
  not _63635_ (_12444_, _12443_);
  and _63636_ (_12445_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _63637_ (_12446_, _05966_, _05962_);
  nor _63638_ (_12447_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _63639_ (_12448_, _12447_, _12445_);
  not _63640_ (_12449_, _12448_);
  nor _63641_ (_12450_, _12449_, _12446_);
  nor _63642_ (_12451_, _12450_, _12445_);
  nor _63643_ (_12452_, _12451_, _12444_);
  nor _63644_ (_12453_, _12452_, _12441_);
  nor _63645_ (_12454_, _12453_, _12440_);
  nor _63646_ (_12455_, _12454_, _12437_);
  nor _63647_ (_12456_, _12455_, _12436_);
  nor _63648_ (_12457_, _12456_, _12435_);
  nor _63649_ (_12458_, _12457_, _12434_);
  and _63650_ (_12459_, _12458_, \oc8051_golden_model_1.DPH [1]);
  and _63651_ (_12460_, _12459_, \oc8051_golden_model_1.DPH [2]);
  and _63652_ (_12461_, _12460_, \oc8051_golden_model_1.DPH [3]);
  and _63653_ (_12462_, _12461_, \oc8051_golden_model_1.DPH [4]);
  and _63654_ (_12463_, _12462_, \oc8051_golden_model_1.DPH [5]);
  and _63655_ (_12464_, _12463_, \oc8051_golden_model_1.DPH [6]);
  nand _63656_ (_12465_, _12464_, \oc8051_golden_model_1.DPH [7]);
  or _63657_ (_12466_, _12464_, \oc8051_golden_model_1.DPH [7]);
  and _63658_ (_12467_, _12466_, _12431_);
  and _63659_ (_12468_, _12467_, _12465_);
  nor _63660_ (_12469_, _06208_, _06076_);
  not _63661_ (_12470_, _12469_);
  or _63662_ (_12471_, _12470_, _12468_);
  or _63663_ (_12472_, _12471_, _12433_);
  and _63664_ (_12473_, _06109_, _05746_);
  not _63665_ (_12474_, _12473_);
  or _63666_ (_12475_, _12469_, _09256_);
  and _63667_ (_12476_, _12475_, _12474_);
  and _63668_ (_12477_, _12476_, _12472_);
  not _63669_ (_12478_, _11919_);
  or _63670_ (_12479_, _12251_, _11101_);
  not _63671_ (_12480_, _11101_);
  or _63672_ (_12481_, _12480_, _09256_);
  and _63673_ (_12482_, _12481_, _12473_);
  and _63674_ (_12483_, _12482_, _12479_);
  or _63675_ (_12484_, _12483_, _12478_);
  or _63676_ (_12485_, _12484_, _12477_);
  and _63677_ (_12486_, _12485_, _11920_);
  or _63678_ (_12487_, _12486_, _11917_);
  or _63679_ (_12488_, _11916_, _09256_);
  and _63680_ (_12489_, _12488_, _07127_);
  and _63681_ (_12490_, _12489_, _12487_);
  nand _63682_ (_12491_, _09239_, _06297_);
  not _63683_ (_12492_, _05834_);
  nor _63684_ (_12493_, _06402_, _12492_);
  nand _63685_ (_12494_, _12493_, _12491_);
  or _63686_ (_12495_, _12494_, _12490_);
  and _63687_ (_12496_, _06399_, _05746_);
  not _63688_ (_12497_, _12496_);
  or _63689_ (_12498_, _12493_, _09256_);
  and _63690_ (_12499_, _12498_, _12497_);
  and _63691_ (_12500_, _12499_, _12495_);
  or _63692_ (_12501_, _12251_, _12480_);
  or _63693_ (_12502_, _11101_, _09256_);
  and _63694_ (_12503_, _12502_, _12496_);
  and _63695_ (_12504_, _12503_, _12501_);
  not _63696_ (_12505_, _11914_);
  or _63697_ (_12506_, _12505_, _12504_);
  or _63698_ (_12507_, _12506_, _12500_);
  and _63699_ (_12508_, _12507_, _11915_);
  or _63700_ (_12509_, _12508_, _10822_);
  or _63701_ (_12510_, _10821_, _09256_);
  and _63702_ (_12511_, _12510_, _07132_);
  and _63703_ (_12512_, _12511_, _12509_);
  nand _63704_ (_12513_, _09239_, _06306_);
  nor _63705_ (_12514_, _06411_, _07124_);
  nand _63706_ (_12515_, _12514_, _12513_);
  or _63707_ (_12516_, _12515_, _12512_);
  and _63708_ (_12517_, _06408_, _05746_);
  not _63709_ (_12518_, _12517_);
  or _63710_ (_12519_, _12514_, _09256_);
  and _63711_ (_12520_, _12519_, _12518_);
  and _63712_ (_12521_, _12520_, _12516_);
  not _63713_ (_12522_, _11912_);
  or _63714_ (_12523_, _12251_, \oc8051_golden_model_1.PSW [7]);
  or _63715_ (_12524_, _09256_, _10693_);
  and _63716_ (_12525_, _12524_, _12517_);
  and _63717_ (_12526_, _12525_, _12523_);
  or _63718_ (_12527_, _12526_, _12522_);
  or _63719_ (_12528_, _12527_, _12521_);
  and _63720_ (_12529_, _12528_, _11913_);
  or _63721_ (_12530_, _12529_, _10850_);
  or _63722_ (_12531_, _10849_, _09256_);
  and _63723_ (_12532_, _12531_, _08819_);
  and _63724_ (_12533_, _12532_, _12530_);
  nand _63725_ (_12534_, _09239_, _06303_);
  nor _63726_ (_12535_, _06396_, _05842_);
  nand _63727_ (_12536_, _12535_, _12534_);
  or _63728_ (_12537_, _12536_, _12533_);
  and _63729_ (_12538_, _05840_, _05746_);
  not _63730_ (_12539_, _12538_);
  or _63731_ (_12540_, _12535_, _09256_);
  and _63732_ (_12541_, _12540_, _12539_);
  and _63733_ (_12542_, _12541_, _12537_);
  or _63734_ (_12543_, _12251_, _10693_);
  or _63735_ (_12544_, _09256_, \oc8051_golden_model_1.PSW [7]);
  and _63736_ (_12545_, _12544_, _12538_);
  and _63737_ (_12546_, _12545_, _12543_);
  not _63738_ (_12547_, _11907_);
  or _63739_ (_12548_, _12547_, _12546_);
  or _63740_ (_12549_, _12548_, _12542_);
  and _63741_ (_12550_, _12549_, _11908_);
  or _63742_ (_12551_, _12550_, _10897_);
  or _63743_ (_12552_, _10896_, _09256_);
  and _63744_ (_12553_, _12552_, _10926_);
  and _63745_ (_12554_, _12553_, _12551_);
  and _63746_ (_12555_, _11904_, _10925_);
  or _63747_ (_12556_, _12555_, _06417_);
  or _63748_ (_12557_, _12556_, _12554_);
  not _63749_ (_12558_, _06417_);
  or _63750_ (_12559_, _07923_, _12558_);
  and _63751_ (_12560_, _12559_, _12557_);
  or _63752_ (_12561_, _12560_, _07142_);
  nor _63753_ (_12562_, _09256_, _05846_);
  nor _63754_ (_12563_, _12562_, _06301_);
  and _63755_ (_12564_, _12563_, _12561_);
  not _63756_ (_12565_, _11905_);
  and _63757_ (_12566_, _08415_, \oc8051_golden_model_1.IP [6]);
  and _63758_ (_12567_, _08418_, \oc8051_golden_model_1.IE [6]);
  and _63759_ (_12568_, _08409_, \oc8051_golden_model_1.ACC [6]);
  or _63760_ (_12569_, _12568_, _12567_);
  or _63761_ (_12570_, _12569_, _12566_);
  and _63762_ (_12571_, _08413_, \oc8051_golden_model_1.SCON [6]);
  and _63763_ (_12572_, _08404_, \oc8051_golden_model_1.PSW [6]);
  or _63764_ (_12573_, _12572_, _12571_);
  and _63765_ (_12574_, _08407_, \oc8051_golden_model_1.TCON [6]);
  and _63766_ (_12575_, _08420_, \oc8051_golden_model_1.B [6]);
  or _63767_ (_12576_, _12575_, _12574_);
  or _63768_ (_12577_, _12576_, _12573_);
  or _63769_ (_12578_, _12577_, _12570_);
  or _63770_ (_12579_, _12578_, _08013_);
  and _63771_ (_12580_, _07800_, _06626_);
  and _63772_ (_12581_, _12580_, _12579_);
  and _63773_ (_12582_, _08415_, \oc8051_golden_model_1.IP [3]);
  and _63774_ (_12583_, _08420_, \oc8051_golden_model_1.B [3]);
  and _63775_ (_12584_, _08409_, \oc8051_golden_model_1.ACC [3]);
  or _63776_ (_12585_, _12584_, _12583_);
  or _63777_ (_12586_, _12585_, _12582_);
  and _63778_ (_12587_, _08407_, \oc8051_golden_model_1.TCON [3]);
  and _63779_ (_12588_, _08413_, \oc8051_golden_model_1.SCON [3]);
  or _63780_ (_12589_, _12588_, _12587_);
  and _63781_ (_12590_, _08418_, \oc8051_golden_model_1.IE [3]);
  and _63782_ (_12591_, _08404_, \oc8051_golden_model_1.PSW [3]);
  or _63783_ (_12592_, _12591_, _12590_);
  or _63784_ (_12593_, _12592_, _12589_);
  or _63785_ (_12594_, _12593_, _12586_);
  or _63786_ (_12595_, _12594_, _08138_);
  and _63787_ (_12596_, _12595_, _07851_);
  nor _63788_ (_12597_, _12596_, _12581_);
  and _63789_ (_12598_, _08413_, \oc8051_golden_model_1.SCON [5]);
  and _63790_ (_12599_, _08418_, \oc8051_golden_model_1.IE [5]);
  and _63791_ (_12600_, _08409_, \oc8051_golden_model_1.ACC [5]);
  or _63792_ (_12601_, _12600_, _12599_);
  or _63793_ (_12602_, _12601_, _12598_);
  and _63794_ (_12603_, _08404_, \oc8051_golden_model_1.PSW [5]);
  and _63795_ (_12604_, _08420_, \oc8051_golden_model_1.B [5]);
  or _63796_ (_12605_, _12604_, _12603_);
  and _63797_ (_12606_, _08407_, \oc8051_golden_model_1.TCON [5]);
  and _63798_ (_12607_, _08415_, \oc8051_golden_model_1.IP [5]);
  or _63799_ (_12608_, _12607_, _12606_);
  or _63800_ (_12609_, _12608_, _12605_);
  or _63801_ (_12610_, _12609_, _12602_);
  or _63802_ (_12611_, _12610_, _08102_);
  and _63803_ (_12612_, _07780_, _06626_);
  and _63804_ (_12613_, _12612_, _12611_);
  and _63805_ (_12614_, _08409_, \oc8051_golden_model_1.ACC [1]);
  and _63806_ (_12615_, _08415_, \oc8051_golden_model_1.IP [1]);
  and _63807_ (_12616_, _08420_, \oc8051_golden_model_1.B [1]);
  or _63808_ (_12617_, _12616_, _12615_);
  or _63809_ (_12618_, _12617_, _12614_);
  and _63810_ (_12619_, _08407_, \oc8051_golden_model_1.TCON [1]);
  and _63811_ (_12620_, _08413_, \oc8051_golden_model_1.SCON [1]);
  or _63812_ (_12621_, _12620_, _12619_);
  and _63813_ (_12622_, _08418_, \oc8051_golden_model_1.IE [1]);
  and _63814_ (_12623_, _08404_, \oc8051_golden_model_1.PSW [1]);
  or _63815_ (_12624_, _12623_, _12622_);
  or _63816_ (_12625_, _12624_, _12621_);
  or _63817_ (_12626_, _12625_, _12618_);
  or _63818_ (_12627_, _12626_, _08174_);
  and _63819_ (_12628_, _12627_, _07781_);
  nor _63820_ (_12629_, _12628_, _12613_);
  and _63821_ (_12630_, _12629_, _12597_);
  and _63822_ (_12631_, _08413_, \oc8051_golden_model_1.SCON [2]);
  and _63823_ (_12632_, _08407_, \oc8051_golden_model_1.TCON [2]);
  and _63824_ (_12633_, _08409_, \oc8051_golden_model_1.ACC [2]);
  or _63825_ (_12634_, _12633_, _12632_);
  or _63826_ (_12635_, _12634_, _12631_);
  and _63827_ (_12636_, _08404_, \oc8051_golden_model_1.PSW [2]);
  and _63828_ (_12637_, _08420_, \oc8051_golden_model_1.B [2]);
  or _63829_ (_12638_, _12637_, _12636_);
  and _63830_ (_12639_, _08418_, \oc8051_golden_model_1.IE [2]);
  and _63831_ (_12640_, _08415_, \oc8051_golden_model_1.IP [2]);
  or _63832_ (_12641_, _12640_, _12639_);
  or _63833_ (_12642_, _12641_, _12638_);
  or _63834_ (_12643_, _12642_, _12635_);
  or _63835_ (_12644_, _12643_, _08246_);
  and _63836_ (_12645_, _12644_, _07848_);
  nor _63837_ (_12646_, _12645_, _08567_);
  and _63838_ (_12647_, _08413_, \oc8051_golden_model_1.SCON [0]);
  and _63839_ (_12648_, _08407_, \oc8051_golden_model_1.TCON [0]);
  and _63840_ (_12649_, _08409_, \oc8051_golden_model_1.ACC [0]);
  or _63841_ (_12650_, _12649_, _12648_);
  or _63842_ (_12651_, _12650_, _12647_);
  and _63843_ (_12652_, _08415_, \oc8051_golden_model_1.IP [0]);
  and _63844_ (_12653_, _08420_, \oc8051_golden_model_1.B [0]);
  or _63845_ (_12654_, _12653_, _12652_);
  and _63846_ (_12655_, _08418_, \oc8051_golden_model_1.IE [0]);
  and _63847_ (_12656_, _08404_, \oc8051_golden_model_1.PSW [0]);
  or _63848_ (_12657_, _12656_, _12655_);
  or _63849_ (_12658_, _12657_, _12654_);
  or _63850_ (_12659_, _12658_, _12651_);
  or _63851_ (_12660_, _12659_, _08210_);
  and _63852_ (_12661_, _12660_, _07772_);
  and _63853_ (_12662_, _08420_, \oc8051_golden_model_1.B [4]);
  and _63854_ (_12663_, _08413_, \oc8051_golden_model_1.SCON [4]);
  and _63855_ (_12664_, _08418_, \oc8051_golden_model_1.IE [4]);
  or _63856_ (_12665_, _12664_, _12663_);
  or _63857_ (_12666_, _12665_, _12662_);
  and _63858_ (_12667_, _08415_, \oc8051_golden_model_1.IP [4]);
  and _63859_ (_12668_, _08404_, \oc8051_golden_model_1.PSW [4]);
  or _63860_ (_12669_, _12668_, _12667_);
  and _63861_ (_12670_, _08407_, \oc8051_golden_model_1.TCON [4]);
  and _63862_ (_12671_, _08409_, \oc8051_golden_model_1.ACC [4]);
  or _63863_ (_12672_, _12671_, _12670_);
  or _63864_ (_12673_, _12672_, _12669_);
  nor _63865_ (_12674_, _12673_, _12666_);
  not _63866_ (_12675_, _12674_);
  nor _63867_ (_12676_, _12675_, _08337_);
  and _63868_ (_12677_, _07771_, _06626_);
  not _63869_ (_12678_, _12677_);
  nor _63870_ (_12679_, _12678_, _12676_);
  nor _63871_ (_12680_, _12679_, _12661_);
  and _63872_ (_12681_, _12680_, _12646_);
  and _63873_ (_12682_, _12681_, _12630_);
  nand _63874_ (_12683_, _12084_, _12682_);
  or _63875_ (_12684_, _09239_, _12682_);
  and _63876_ (_12685_, _12684_, _06301_);
  and _63877_ (_12686_, _12685_, _12683_);
  or _63878_ (_12687_, _12686_, _12565_);
  or _63879_ (_12688_, _12687_, _12564_);
  and _63880_ (_12689_, _12688_, _11906_);
  nor _63881_ (_12690_, _10264_, _06169_);
  not _63882_ (_12691_, _12690_);
  or _63883_ (_12692_, _12691_, _12689_);
  not _63884_ (_12693_, _10262_);
  or _63885_ (_12694_, _12690_, _09256_);
  and _63886_ (_12695_, _12694_, _12693_);
  and _63887_ (_12696_, _12695_, _12692_);
  and _63888_ (_12697_, _11904_, _10262_);
  or _63889_ (_12698_, _12697_, _06167_);
  or _63890_ (_12699_, _12698_, _12696_);
  or _63891_ (_12700_, _07923_, _06168_);
  and _63892_ (_12701_, _12700_, _12699_);
  or _63893_ (_12702_, _12701_, _05826_);
  not _63894_ (_12703_, _05826_);
  or _63895_ (_12704_, _09256_, _12703_);
  and _63896_ (_12705_, _12704_, _06166_);
  and _63897_ (_12706_, _12705_, _12702_);
  or _63898_ (_12707_, _12085_, _12682_);
  nand _63899_ (_12708_, _09240_, _12682_);
  and _63900_ (_12709_, _12708_, _12707_);
  and _63901_ (_12710_, _12709_, _06165_);
  and _63902_ (_12711_, _08362_, _07154_);
  not _63903_ (_12712_, _12711_);
  or _63904_ (_12713_, _12712_, _12710_);
  or _63905_ (_12714_, _12713_, _12706_);
  or _63906_ (_12716_, _12711_, _11904_);
  and _63907_ (_12717_, _12716_, _06829_);
  and _63908_ (_12718_, _12717_, _12714_);
  nor _63909_ (_12719_, _11094_, _11089_);
  nand _63910_ (_12720_, _09256_, _06433_);
  nand _63911_ (_12721_, _12720_, _12719_);
  or _63912_ (_12722_, _12721_, _12718_);
  not _63913_ (_12723_, _06310_);
  or _63914_ (_12724_, _11904_, _12719_);
  and _63915_ (_12725_, _12724_, _12723_);
  and _63916_ (_12726_, _12725_, _12722_);
  and _63917_ (_12727_, _06310_, _06039_);
  or _63918_ (_12728_, _12727_, _05823_);
  or _63919_ (_12729_, _12728_, _12726_);
  not _63920_ (_12730_, _05823_);
  or _63921_ (_12731_, _09256_, _12730_);
  and _63922_ (_12732_, _12731_, _05749_);
  and _63923_ (_12733_, _12732_, _12729_);
  and _63924_ (_12734_, _12709_, _05748_);
  nor _63925_ (_12735_, _09189_, _07168_);
  not _63926_ (_12737_, _12735_);
  or _63927_ (_12738_, _12737_, _12734_);
  or _63928_ (_12739_, _12738_, _12733_);
  or _63929_ (_12740_, _12735_, _11904_);
  and _63930_ (_12741_, _12740_, _06444_);
  and _63931_ (_12742_, _12741_, _12739_);
  nand _63932_ (_12743_, _09256_, _06440_);
  nor _63933_ (_12744_, _11119_, _11112_);
  nand _63934_ (_12745_, _12744_, _12743_);
  or _63935_ (_12746_, _12745_, _12742_);
  not _63936_ (_12747_, _06305_);
  or _63937_ (_12748_, _12744_, _11904_);
  and _63938_ (_12749_, _12748_, _12747_);
  and _63939_ (_12750_, _12749_, _12746_);
  and _63940_ (_12751_, _06305_, _06039_);
  or _63941_ (_12752_, _12751_, _05821_);
  or _63942_ (_12753_, _12752_, _12750_);
  and _63943_ (_12754_, _05820_, _05746_);
  not _63944_ (_12755_, _12754_);
  or _63945_ (_12756_, _09256_, _05822_);
  and _63946_ (_12757_, _12756_, _12755_);
  and _63947_ (_12758_, _12757_, _12753_);
  and _63948_ (_12759_, _12754_, _11904_);
  or _63949_ (_12760_, _12759_, _12758_);
  or _63950_ (_12761_, _12760_, _01321_);
  or _63951_ (_12762_, _01317_, \oc8051_golden_model_1.PC [15]);
  and _63952_ (_12763_, _12762_, _43100_);
  and _63953_ (_40993_, _12763_, _12761_);
  nor _63954_ (_12764_, \oc8051_golden_model_1.P2 [7], rst);
  nor _63955_ (_12765_, _12764_, _00000_);
  not _63956_ (_12766_, \oc8051_golden_model_1.P2 [7]);
  not _63957_ (_12767_, _07825_);
  nor _63958_ (_12768_, _12767_, _07790_);
  nor _63959_ (_12769_, _12768_, _12766_);
  and _63960_ (_12770_, _12768_, _07923_);
  or _63961_ (_12771_, _12770_, _12769_);
  or _63962_ (_12772_, _12771_, _06132_);
  and _63963_ (_12773_, _08403_, _07825_);
  nor _63964_ (_12774_, _12773_, _12766_);
  and _63965_ (_12775_, _07847_, \oc8051_golden_model_1.P0 [7]);
  and _63966_ (_12776_, _12773_, \oc8051_golden_model_1.P2 [7]);
  or _63967_ (_12777_, _12776_, _12775_);
  and _63968_ (_12778_, _08403_, _07777_);
  and _63969_ (_12779_, _12778_, \oc8051_golden_model_1.P1 [7]);
  and _63970_ (_12780_, _08403_, _07829_);
  and _63971_ (_12781_, _12780_, \oc8051_golden_model_1.P3 [7]);
  or _63972_ (_12782_, _12781_, _12779_);
  or _63973_ (_12783_, _12782_, _12777_);
  or _63974_ (_12784_, _12783_, _08425_);
  and _63975_ (_12785_, _12784_, _08399_);
  and _63976_ (_12786_, _12785_, _12773_);
  or _63977_ (_12787_, _12786_, _12774_);
  and _63978_ (_12788_, _12787_, _06152_);
  and _63979_ (_12789_, _07847_, _07772_);
  and _63980_ (_12790_, _12789_, \oc8051_golden_model_1.P0 [7]);
  not _63981_ (_12791_, _07777_);
  nor _63982_ (_12792_, _07790_, _12791_);
  and _63983_ (_12793_, _12792_, \oc8051_golden_model_1.P1 [7]);
  nor _63984_ (_12794_, _12793_, _12790_);
  and _63985_ (_12795_, _12768_, \oc8051_golden_model_1.P2 [7]);
  not _63986_ (_12796_, _07829_);
  nor _63987_ (_12797_, _12796_, _07790_);
  and _63988_ (_12798_, _12797_, \oc8051_golden_model_1.P3 [7]);
  nor _63989_ (_12799_, _12798_, _12795_);
  and _63990_ (_12800_, _12799_, _12794_);
  and _63991_ (_12801_, _12800_, _07925_);
  not _63992_ (_12802_, _12801_);
  and _63993_ (_12803_, _12797_, \oc8051_golden_model_1.P3 [6]);
  and _63994_ (_12804_, _12792_, \oc8051_golden_model_1.P1 [6]);
  or _63995_ (_12805_, _12804_, _12803_);
  and _63996_ (_12806_, _12789_, \oc8051_golden_model_1.P0 [6]);
  and _63997_ (_12807_, _12768_, \oc8051_golden_model_1.P2 [6]);
  or _63998_ (_12808_, _12807_, _12806_);
  nor _63999_ (_12809_, _12808_, _12805_);
  nand _64000_ (_12810_, _12809_, _08014_);
  and _64001_ (_12811_, _12797_, \oc8051_golden_model_1.P3 [5]);
  and _64002_ (_12812_, _12792_, \oc8051_golden_model_1.P1 [5]);
  or _64003_ (_12813_, _12812_, _12811_);
  and _64004_ (_12814_, _12789_, \oc8051_golden_model_1.P0 [5]);
  and _64005_ (_12815_, _12768_, \oc8051_golden_model_1.P2 [5]);
  or _64006_ (_12816_, _12815_, _12814_);
  nor _64007_ (_12817_, _12816_, _12813_);
  nand _64008_ (_12818_, _12817_, _08103_);
  and _64009_ (_12819_, _12797_, \oc8051_golden_model_1.P3 [4]);
  and _64010_ (_12820_, _12792_, \oc8051_golden_model_1.P1 [4]);
  or _64011_ (_12821_, _12820_, _12819_);
  and _64012_ (_12822_, _12789_, \oc8051_golden_model_1.P0 [4]);
  and _64013_ (_12823_, _12768_, \oc8051_golden_model_1.P2 [4]);
  or _64014_ (_12824_, _12823_, _12822_);
  nor _64015_ (_12825_, _12824_, _12821_);
  nand _64016_ (_12826_, _12825_, _08338_);
  and _64017_ (_12827_, _12797_, \oc8051_golden_model_1.P3 [3]);
  and _64018_ (_12828_, _12792_, \oc8051_golden_model_1.P1 [3]);
  or _64019_ (_12829_, _12828_, _12827_);
  and _64020_ (_12830_, _12789_, \oc8051_golden_model_1.P0 [3]);
  and _64021_ (_12831_, _12768_, \oc8051_golden_model_1.P2 [3]);
  or _64022_ (_12832_, _12831_, _12830_);
  nor _64023_ (_12833_, _12832_, _12829_);
  nand _64024_ (_12834_, _12833_, _08139_);
  and _64025_ (_12835_, _12797_, \oc8051_golden_model_1.P3 [2]);
  and _64026_ (_12836_, _12792_, \oc8051_golden_model_1.P1 [2]);
  or _64027_ (_12837_, _12836_, _12835_);
  and _64028_ (_12838_, _12789_, \oc8051_golden_model_1.P0 [2]);
  and _64029_ (_12839_, _12768_, \oc8051_golden_model_1.P2 [2]);
  or _64030_ (_12840_, _12839_, _12838_);
  nor _64031_ (_12841_, _12840_, _12837_);
  nand _64032_ (_12842_, _12841_, _08247_);
  and _64033_ (_12843_, _12789_, \oc8051_golden_model_1.P0 [1]);
  and _64034_ (_12844_, _12792_, \oc8051_golden_model_1.P1 [1]);
  or _64035_ (_12845_, _12844_, _12843_);
  and _64036_ (_12846_, _12768_, \oc8051_golden_model_1.P2 [1]);
  and _64037_ (_12847_, _12797_, \oc8051_golden_model_1.P3 [1]);
  or _64038_ (_12848_, _12847_, _12846_);
  nor _64039_ (_12849_, _12848_, _12845_);
  nand _64040_ (_12850_, _12849_, _08175_);
  and _64041_ (_12851_, _12789_, \oc8051_golden_model_1.P0 [0]);
  and _64042_ (_12852_, _12792_, \oc8051_golden_model_1.P1 [0]);
  or _64043_ (_12853_, _12852_, _12851_);
  and _64044_ (_12854_, _12768_, \oc8051_golden_model_1.P2 [0]);
  and _64045_ (_12855_, _12797_, \oc8051_golden_model_1.P3 [0]);
  or _64046_ (_12856_, _12855_, _12854_);
  or _64047_ (_12857_, _12856_, _12853_);
  or _64048_ (_12858_, _12857_, _08211_);
  or _64049_ (_12859_, _12858_, _12850_);
  nor _64050_ (_12860_, _12859_, _12842_);
  not _64051_ (_12861_, _12860_);
  nor _64052_ (_12862_, _12861_, _12834_);
  not _64053_ (_12863_, _12862_);
  nor _64054_ (_12864_, _12863_, _12826_);
  not _64055_ (_12865_, _12864_);
  nor _64056_ (_12866_, _12865_, _12818_);
  not _64057_ (_12867_, _12866_);
  nor _64058_ (_12868_, _12867_, _12810_);
  or _64059_ (_12869_, _12868_, _12802_);
  nand _64060_ (_12870_, _12868_, _12802_);
  and _64061_ (_12871_, _12870_, _12869_);
  and _64062_ (_12872_, _12871_, _12768_);
  or _64063_ (_12873_, _12872_, _12769_);
  or _64064_ (_12874_, _12873_, _06161_);
  and _64065_ (_12875_, _12768_, \oc8051_golden_model_1.ACC [7]);
  or _64066_ (_12876_, _12875_, _12769_);
  and _64067_ (_12877_, _12876_, _07056_);
  nor _64068_ (_12878_, _07056_, _12766_);
  or _64069_ (_12879_, _12878_, _06160_);
  or _64070_ (_12880_, _12879_, _12877_);
  and _64071_ (_12881_, _12880_, _06157_);
  and _64072_ (_12882_, _12881_, _12874_);
  or _64073_ (_12883_, _12783_, _08552_);
  and _64074_ (_12884_, _12883_, _12773_);
  or _64075_ (_12885_, _12884_, _12774_);
  and _64076_ (_12886_, _12885_, _06156_);
  or _64077_ (_12887_, _12886_, _06217_);
  or _64078_ (_12888_, _12887_, _12882_);
  or _64079_ (_12889_, _12771_, _07075_);
  and _64080_ (_12890_, _12889_, _12888_);
  or _64081_ (_12891_, _12890_, _06220_);
  or _64082_ (_12892_, _12876_, _06229_);
  and _64083_ (_12893_, _12892_, _06153_);
  and _64084_ (_12894_, _12893_, _12891_);
  or _64085_ (_12895_, _12894_, _12788_);
  and _64086_ (_12896_, _12895_, _06146_);
  nand _64087_ (_12897_, _12784_, _07855_);
  or _64088_ (_12898_, _12897_, _12774_);
  and _64089_ (_12899_, _12885_, _06145_);
  and _64090_ (_12900_, _12899_, _12898_);
  or _64091_ (_12901_, _12900_, _12896_);
  and _64092_ (_12902_, _12901_, _06140_);
  or _64093_ (_12903_, _12785_, _08586_);
  and _64094_ (_12904_, _12903_, _12773_);
  or _64095_ (_12905_, _12904_, _12774_);
  and _64096_ (_12906_, _12905_, _06139_);
  or _64097_ (_12907_, _12906_, _09842_);
  or _64098_ (_12908_, _12907_, _12902_);
  and _64099_ (_12909_, _12908_, _12772_);
  or _64100_ (_12910_, _12909_, _06116_);
  and _64101_ (_12911_, _12768_, _08535_);
  or _64102_ (_12912_, _12769_, _06117_);
  or _64103_ (_12913_, _12912_, _12911_);
  and _64104_ (_12914_, _12913_, _06114_);
  and _64105_ (_12915_, _12914_, _12910_);
  and _64106_ (_12916_, _08731_, _08703_);
  and _64107_ (_12917_, _12916_, \oc8051_golden_model_1.P0 [7]);
  and _64108_ (_12918_, _08717_, _08731_);
  and _64109_ (_12919_, _12918_, \oc8051_golden_model_1.P1 [7]);
  and _64110_ (_12920_, _08748_, _08731_);
  and _64111_ (_12921_, _12920_, \oc8051_golden_model_1.P2 [7]);
  and _64112_ (_12922_, _08731_, _08745_);
  and _64113_ (_12923_, _12922_, \oc8051_golden_model_1.P3 [7]);
  or _64114_ (_12924_, _12923_, _12921_);
  or _64115_ (_12925_, _12924_, _12919_);
  or _64116_ (_12926_, _12925_, _12917_);
  or _64117_ (_12927_, _12926_, _08782_);
  and _64118_ (_12928_, _12927_, _12768_);
  or _64119_ (_12929_, _12928_, _12769_);
  and _64120_ (_12930_, _12929_, _05787_);
  or _64121_ (_12931_, _12930_, _06110_);
  or _64122_ (_12932_, _12931_, _12915_);
  and _64123_ (_12933_, _12768_, _08607_);
  or _64124_ (_12934_, _12933_, _12769_);
  or _64125_ (_12935_, _12934_, _06111_);
  and _64126_ (_12936_, _12935_, _07127_);
  and _64127_ (_12937_, _12936_, _12932_);
  nand _64128_ (_12938_, _12801_, _08395_);
  and _64129_ (_12939_, _12938_, _12768_);
  or _64130_ (_12940_, _12939_, _12769_);
  or _64131_ (_12941_, _12801_, _08395_);
  or _64132_ (_12942_, _12941_, _12769_);
  and _64133_ (_12943_, _12942_, _06297_);
  and _64134_ (_12944_, _12943_, _12940_);
  or _64135_ (_12945_, _12944_, _12937_);
  and _64136_ (_12946_, _12945_, _07125_);
  nand _64137_ (_12947_, _12801_, _08430_);
  and _64138_ (_12948_, _12947_, _12768_);
  or _64139_ (_12949_, _12948_, _12769_);
  or _64140_ (_12950_, _12801_, _08430_);
  or _64141_ (_12951_, _12950_, _12769_);
  and _64142_ (_12952_, _12951_, _06402_);
  and _64143_ (_12953_, _12952_, _12949_);
  or _64144_ (_12954_, _12953_, _12946_);
  and _64145_ (_12955_, _12954_, _07132_);
  or _64146_ (_12956_, _12802_, _12769_);
  and _64147_ (_12957_, _12934_, _06306_);
  and _64148_ (_12958_, _12957_, _12956_);
  or _64149_ (_12959_, _12958_, _12955_);
  and _64150_ (_12960_, _12959_, _07130_);
  and _64151_ (_12961_, _12876_, _06411_);
  and _64152_ (_12962_, _12961_, _12956_);
  or _64153_ (_12963_, _12962_, _06303_);
  or _64154_ (_12964_, _12963_, _12960_);
  or _64155_ (_12965_, _12940_, _08819_);
  and _64156_ (_12966_, _12965_, _08824_);
  and _64157_ (_12967_, _12966_, _12964_);
  and _64158_ (_12968_, _12949_, _06396_);
  or _64159_ (_12969_, _12968_, _06433_);
  or _64160_ (_12970_, _12969_, _12967_);
  or _64161_ (_12971_, _12873_, _06829_);
  and _64162_ (_12972_, _12971_, _05749_);
  and _64163_ (_12973_, _12972_, _12970_);
  and _64164_ (_12974_, _12787_, _05748_);
  or _64165_ (_12975_, _12974_, _06440_);
  or _64166_ (_12976_, _12975_, _12973_);
  and _64167_ (_12977_, _12858_, _12850_);
  and _64168_ (_12978_, _12977_, _12842_);
  and _64169_ (_12979_, _12978_, _12834_);
  and _64170_ (_12980_, _12979_, _12826_);
  and _64171_ (_12981_, _12980_, _12818_);
  nand _64172_ (_12982_, _12981_, _12810_);
  nand _64173_ (_12983_, _12982_, _12801_);
  or _64174_ (_12984_, _12982_, _12801_);
  and _64175_ (_12985_, _12984_, _12983_);
  and _64176_ (_12986_, _12985_, _12768_);
  or _64177_ (_12987_, _12769_, _06444_);
  or _64178_ (_12988_, _12987_, _12986_);
  and _64179_ (_12989_, _12988_, _01317_);
  and _64180_ (_12990_, _12989_, _12976_);
  or _64181_ (_40994_, _12990_, _12765_);
  not _64182_ (_12991_, _12797_);
  and _64183_ (_12992_, _12991_, \oc8051_golden_model_1.P3 [7]);
  and _64184_ (_12993_, _12797_, _07923_);
  or _64185_ (_12994_, _12993_, _12992_);
  or _64186_ (_12995_, _12994_, _06132_);
  not _64187_ (_12996_, _12780_);
  and _64188_ (_12997_, _12996_, \oc8051_golden_model_1.P3 [7]);
  and _64189_ (_12998_, _12785_, _12780_);
  or _64190_ (_12999_, _12998_, _12997_);
  and _64191_ (_13000_, _12999_, _06152_);
  and _64192_ (_13001_, _12871_, _12797_);
  or _64193_ (_13002_, _13001_, _12992_);
  or _64194_ (_13003_, _13002_, _06161_);
  and _64195_ (_13004_, _12797_, \oc8051_golden_model_1.ACC [7]);
  or _64196_ (_13005_, _13004_, _12992_);
  and _64197_ (_13006_, _13005_, _07056_);
  and _64198_ (_13007_, _07057_, \oc8051_golden_model_1.P3 [7]);
  or _64199_ (_13008_, _13007_, _06160_);
  or _64200_ (_13009_, _13008_, _13006_);
  and _64201_ (_13010_, _13009_, _06157_);
  and _64202_ (_13011_, _13010_, _13003_);
  and _64203_ (_13012_, _12883_, _12780_);
  or _64204_ (_13013_, _13012_, _12997_);
  and _64205_ (_13014_, _13013_, _06156_);
  or _64206_ (_13015_, _13014_, _06217_);
  or _64207_ (_13016_, _13015_, _13011_);
  or _64208_ (_13017_, _12994_, _07075_);
  and _64209_ (_13018_, _13017_, _13016_);
  or _64210_ (_13019_, _13018_, _06220_);
  or _64211_ (_13020_, _13005_, _06229_);
  and _64212_ (_13021_, _13020_, _06153_);
  and _64213_ (_13022_, _13021_, _13019_);
  or _64214_ (_13023_, _13022_, _13000_);
  and _64215_ (_13024_, _13023_, _06146_);
  or _64216_ (_13025_, _12997_, _12897_);
  and _64217_ (_13026_, _13013_, _06145_);
  and _64218_ (_13027_, _13026_, _13025_);
  or _64219_ (_13028_, _13027_, _13024_);
  and _64220_ (_13029_, _13028_, _06140_);
  and _64221_ (_13030_, _12903_, _12780_);
  or _64222_ (_13031_, _13030_, _12997_);
  and _64223_ (_13032_, _13031_, _06139_);
  or _64224_ (_13033_, _13032_, _09842_);
  or _64225_ (_13034_, _13033_, _13029_);
  and _64226_ (_13035_, _13034_, _12995_);
  or _64227_ (_13036_, _13035_, _06116_);
  and _64228_ (_13037_, _12797_, _08535_);
  or _64229_ (_13038_, _12992_, _06117_);
  or _64230_ (_13039_, _13038_, _13037_);
  and _64231_ (_13040_, _13039_, _06114_);
  and _64232_ (_13041_, _13040_, _13036_);
  and _64233_ (_13042_, _12927_, _12797_);
  or _64234_ (_13043_, _13042_, _12992_);
  and _64235_ (_13044_, _13043_, _05787_);
  or _64236_ (_13045_, _13044_, _06110_);
  or _64237_ (_13046_, _13045_, _13041_);
  and _64238_ (_13047_, _12797_, _08607_);
  or _64239_ (_13048_, _13047_, _12992_);
  or _64240_ (_13049_, _13048_, _06111_);
  and _64241_ (_13050_, _13049_, _07127_);
  and _64242_ (_13051_, _13050_, _13046_);
  and _64243_ (_13052_, _12938_, _12797_);
  or _64244_ (_13053_, _13052_, _12992_);
  or _64245_ (_13054_, _12992_, _12941_);
  and _64246_ (_13055_, _13054_, _06297_);
  and _64247_ (_13056_, _13055_, _13053_);
  or _64248_ (_13057_, _13056_, _13051_);
  and _64249_ (_13058_, _13057_, _07125_);
  and _64250_ (_13059_, _12947_, _12797_);
  or _64251_ (_13060_, _13059_, _12992_);
  or _64252_ (_13061_, _12992_, _12950_);
  and _64253_ (_13062_, _13061_, _06402_);
  and _64254_ (_13063_, _13062_, _13060_);
  or _64255_ (_13064_, _13063_, _13058_);
  and _64256_ (_13065_, _13064_, _07132_);
  or _64257_ (_13066_, _12992_, _12802_);
  and _64258_ (_13067_, _13048_, _06306_);
  and _64259_ (_13068_, _13067_, _13066_);
  or _64260_ (_13069_, _13068_, _13065_);
  and _64261_ (_13070_, _13069_, _07130_);
  and _64262_ (_13071_, _13005_, _06411_);
  and _64263_ (_13072_, _13071_, _13066_);
  or _64264_ (_13073_, _13072_, _06303_);
  or _64265_ (_13074_, _13073_, _13070_);
  or _64266_ (_13075_, _13053_, _08819_);
  and _64267_ (_13076_, _13075_, _08824_);
  and _64268_ (_13077_, _13076_, _13074_);
  and _64269_ (_13078_, _13060_, _06396_);
  or _64270_ (_13079_, _13078_, _06433_);
  or _64271_ (_13080_, _13079_, _13077_);
  or _64272_ (_13081_, _13002_, _06829_);
  and _64273_ (_13082_, _13081_, _05749_);
  and _64274_ (_13083_, _13082_, _13080_);
  and _64275_ (_13084_, _12999_, _05748_);
  or _64276_ (_13085_, _13084_, _06440_);
  or _64277_ (_13086_, _13085_, _13083_);
  and _64278_ (_13087_, _12985_, _12797_);
  or _64279_ (_13088_, _12992_, _06444_);
  or _64280_ (_13089_, _13088_, _13087_);
  and _64281_ (_13090_, _13089_, _01317_);
  and _64282_ (_13091_, _13090_, _13086_);
  nor _64283_ (_13092_, \oc8051_golden_model_1.P3 [7], rst);
  nor _64284_ (_13093_, _13092_, _00000_);
  or _64285_ (_40995_, _13093_, _13091_);
  nor _64286_ (_13094_, \oc8051_golden_model_1.P0 [7], rst);
  nor _64287_ (_13095_, _13094_, _00000_);
  not _64288_ (_13096_, _12789_);
  and _64289_ (_13097_, _13096_, \oc8051_golden_model_1.P0 [7]);
  and _64290_ (_13098_, _12789_, _07923_);
  or _64291_ (_13099_, _13098_, _13097_);
  or _64292_ (_13100_, _13099_, _06132_);
  not _64293_ (_13101_, _07847_);
  and _64294_ (_13102_, _13101_, \oc8051_golden_model_1.P0 [7]);
  and _64295_ (_13103_, _12785_, _07847_);
  or _64296_ (_13104_, _13103_, _13102_);
  and _64297_ (_13105_, _13104_, _06152_);
  and _64298_ (_13106_, _12871_, _12789_);
  or _64299_ (_13107_, _13106_, _13097_);
  or _64300_ (_13108_, _13107_, _06161_);
  and _64301_ (_13109_, _12789_, \oc8051_golden_model_1.ACC [7]);
  or _64302_ (_13110_, _13109_, _13097_);
  and _64303_ (_13111_, _13110_, _07056_);
  and _64304_ (_13112_, _07057_, \oc8051_golden_model_1.P0 [7]);
  or _64305_ (_13113_, _13112_, _06160_);
  or _64306_ (_13114_, _13113_, _13111_);
  and _64307_ (_13115_, _13114_, _06157_);
  and _64308_ (_13116_, _13115_, _13108_);
  and _64309_ (_13117_, _12883_, _07847_);
  or _64310_ (_13118_, _13117_, _13102_);
  and _64311_ (_13119_, _13118_, _06156_);
  or _64312_ (_13120_, _13119_, _06217_);
  or _64313_ (_13121_, _13120_, _13116_);
  or _64314_ (_13122_, _13099_, _07075_);
  and _64315_ (_13123_, _13122_, _13121_);
  or _64316_ (_13124_, _13123_, _06220_);
  or _64317_ (_13125_, _13110_, _06229_);
  and _64318_ (_13126_, _13125_, _06153_);
  and _64319_ (_13127_, _13126_, _13124_);
  or _64320_ (_13128_, _13127_, _13105_);
  and _64321_ (_13129_, _13128_, _06146_);
  or _64322_ (_13130_, _13102_, _12897_);
  and _64323_ (_13131_, _13118_, _06145_);
  and _64324_ (_13132_, _13131_, _13130_);
  or _64325_ (_13133_, _13132_, _13129_);
  and _64326_ (_13134_, _13133_, _06140_);
  and _64327_ (_13135_, _12903_, _07847_);
  or _64328_ (_13136_, _13135_, _13102_);
  and _64329_ (_13137_, _13136_, _06139_);
  or _64330_ (_13138_, _13137_, _09842_);
  or _64331_ (_13139_, _13138_, _13134_);
  and _64332_ (_13140_, _13139_, _13100_);
  or _64333_ (_13141_, _13140_, _06116_);
  and _64334_ (_13142_, _12789_, _08535_);
  or _64335_ (_13143_, _13097_, _06117_);
  or _64336_ (_13144_, _13143_, _13142_);
  and _64337_ (_13145_, _13144_, _06114_);
  and _64338_ (_13146_, _13145_, _13141_);
  and _64339_ (_13147_, _12927_, _12789_);
  or _64340_ (_13148_, _13147_, _13097_);
  and _64341_ (_13149_, _13148_, _05787_);
  or _64342_ (_13150_, _13149_, _11136_);
  or _64343_ (_13151_, _13150_, _13146_);
  and _64344_ (_13152_, _12938_, _12789_);
  and _64345_ (_13153_, _13152_, _12941_);
  or _64346_ (_13154_, _13097_, _07127_);
  or _64347_ (_13155_, _13154_, _13153_);
  and _64348_ (_13156_, _12789_, _08607_);
  or _64349_ (_13157_, _13156_, _13097_);
  or _64350_ (_13158_, _13157_, _06111_);
  and _64351_ (_13159_, _13158_, _07125_);
  and _64352_ (_13160_, _13159_, _13155_);
  and _64353_ (_13161_, _13160_, _13151_);
  and _64354_ (_13162_, _12947_, _12789_);
  and _64355_ (_13163_, _13162_, _12950_);
  or _64356_ (_13164_, _13163_, _13097_);
  and _64357_ (_13165_, _13164_, _06402_);
  or _64358_ (_13166_, _13165_, _13161_);
  and _64359_ (_13167_, _13166_, _07132_);
  or _64360_ (_13168_, _13097_, _12802_);
  and _64361_ (_13169_, _13157_, _06306_);
  and _64362_ (_13170_, _13169_, _13168_);
  or _64363_ (_13171_, _13170_, _13167_);
  and _64364_ (_13172_, _13171_, _07130_);
  and _64365_ (_13173_, _13110_, _06411_);
  and _64366_ (_13174_, _13173_, _13168_);
  or _64367_ (_13175_, _13174_, _06303_);
  or _64368_ (_13176_, _13175_, _13172_);
  or _64369_ (_13177_, _13097_, _08819_);
  or _64370_ (_13178_, _13177_, _13152_);
  and _64371_ (_13179_, _13178_, _08824_);
  and _64372_ (_13180_, _13179_, _13176_);
  or _64373_ (_13181_, _13162_, _13097_);
  and _64374_ (_13182_, _13181_, _06396_);
  or _64375_ (_13183_, _13182_, _06433_);
  or _64376_ (_13184_, _13183_, _13180_);
  or _64377_ (_13185_, _13107_, _06829_);
  and _64378_ (_13186_, _13185_, _05749_);
  and _64379_ (_13187_, _13186_, _13184_);
  and _64380_ (_13188_, _13104_, _05748_);
  or _64381_ (_13189_, _13188_, _06440_);
  or _64382_ (_13190_, _13189_, _13187_);
  and _64383_ (_13191_, _12985_, _12789_);
  or _64384_ (_13192_, _13097_, _06444_);
  or _64385_ (_13193_, _13192_, _13191_);
  and _64386_ (_13194_, _13193_, _01317_);
  and _64387_ (_13195_, _13194_, _13190_);
  or _64388_ (_40997_, _13195_, _13095_);
  not _64389_ (_13196_, _12792_);
  and _64390_ (_13197_, _13196_, \oc8051_golden_model_1.P1 [7]);
  and _64391_ (_13198_, _12792_, _07923_);
  or _64392_ (_13199_, _13198_, _13197_);
  or _64393_ (_13200_, _13199_, _06132_);
  not _64394_ (_13201_, _12778_);
  and _64395_ (_13202_, _13201_, \oc8051_golden_model_1.P1 [7]);
  and _64396_ (_13203_, _12785_, _12778_);
  or _64397_ (_13204_, _13203_, _13202_);
  and _64398_ (_13205_, _13204_, _06152_);
  and _64399_ (_13206_, _12871_, _12792_);
  or _64400_ (_13207_, _13206_, _13197_);
  or _64401_ (_13208_, _13207_, _06161_);
  and _64402_ (_13209_, _12792_, \oc8051_golden_model_1.ACC [7]);
  or _64403_ (_13210_, _13209_, _13197_);
  and _64404_ (_13211_, _13210_, _07056_);
  and _64405_ (_13212_, _07057_, \oc8051_golden_model_1.P1 [7]);
  or _64406_ (_13213_, _13212_, _06160_);
  or _64407_ (_13214_, _13213_, _13211_);
  and _64408_ (_13215_, _13214_, _06157_);
  and _64409_ (_13216_, _13215_, _13208_);
  and _64410_ (_13217_, _12883_, _12778_);
  or _64411_ (_13218_, _13217_, _13202_);
  and _64412_ (_13219_, _13218_, _06156_);
  or _64413_ (_13220_, _13219_, _06217_);
  or _64414_ (_13221_, _13220_, _13216_);
  or _64415_ (_13222_, _13199_, _07075_);
  and _64416_ (_13223_, _13222_, _13221_);
  or _64417_ (_13224_, _13223_, _06220_);
  or _64418_ (_13225_, _13210_, _06229_);
  and _64419_ (_13226_, _13225_, _06153_);
  and _64420_ (_13227_, _13226_, _13224_);
  or _64421_ (_13228_, _13227_, _13205_);
  and _64422_ (_13229_, _13228_, _06146_);
  or _64423_ (_13230_, _13202_, _12897_);
  and _64424_ (_13231_, _13218_, _06145_);
  and _64425_ (_13232_, _13231_, _13230_);
  or _64426_ (_13233_, _13232_, _13229_);
  and _64427_ (_13234_, _13233_, _06140_);
  and _64428_ (_13235_, _12903_, _12778_);
  or _64429_ (_13236_, _13235_, _13202_);
  and _64430_ (_13237_, _13236_, _06139_);
  or _64431_ (_13238_, _13237_, _09842_);
  or _64432_ (_13239_, _13238_, _13234_);
  and _64433_ (_13240_, _13239_, _13200_);
  or _64434_ (_13241_, _13240_, _06116_);
  and _64435_ (_13242_, _12792_, _08535_);
  or _64436_ (_13243_, _13197_, _06117_);
  or _64437_ (_13244_, _13243_, _13242_);
  and _64438_ (_13245_, _13244_, _06114_);
  and _64439_ (_13246_, _13245_, _13241_);
  and _64440_ (_13247_, _12927_, _12792_);
  or _64441_ (_13248_, _13247_, _13197_);
  and _64442_ (_13249_, _13248_, _05787_);
  or _64443_ (_13250_, _13249_, _06110_);
  or _64444_ (_13251_, _13250_, _13246_);
  and _64445_ (_13252_, _12792_, _08607_);
  or _64446_ (_13253_, _13252_, _13197_);
  or _64447_ (_13254_, _13253_, _06111_);
  and _64448_ (_13255_, _13254_, _07127_);
  and _64449_ (_13256_, _13255_, _13251_);
  and _64450_ (_13257_, _12938_, _12792_);
  or _64451_ (_13258_, _13257_, _13197_);
  or _64452_ (_13259_, _13197_, _12941_);
  and _64453_ (_13260_, _13259_, _06297_);
  and _64454_ (_13261_, _13260_, _13258_);
  or _64455_ (_13262_, _13261_, _13256_);
  and _64456_ (_13263_, _13262_, _07125_);
  and _64457_ (_13264_, _12947_, _12792_);
  or _64458_ (_13265_, _13264_, _13197_);
  or _64459_ (_13266_, _13197_, _12950_);
  and _64460_ (_13267_, _13266_, _06402_);
  and _64461_ (_13268_, _13267_, _13265_);
  or _64462_ (_13269_, _13268_, _13263_);
  and _64463_ (_13270_, _13269_, _07132_);
  or _64464_ (_13271_, _13197_, _12802_);
  and _64465_ (_13272_, _13253_, _06306_);
  and _64466_ (_13273_, _13272_, _13271_);
  or _64467_ (_13274_, _13273_, _13270_);
  and _64468_ (_13275_, _13274_, _07130_);
  and _64469_ (_13276_, _13210_, _06411_);
  and _64470_ (_13277_, _13276_, _13271_);
  or _64471_ (_13278_, _13277_, _06303_);
  or _64472_ (_13279_, _13278_, _13275_);
  or _64473_ (_13280_, _13258_, _08819_);
  and _64474_ (_13281_, _13280_, _08824_);
  and _64475_ (_13282_, _13281_, _13279_);
  and _64476_ (_13283_, _13265_, _06396_);
  or _64477_ (_13284_, _13283_, _06433_);
  or _64478_ (_13285_, _13284_, _13282_);
  or _64479_ (_13286_, _13207_, _06829_);
  and _64480_ (_13287_, _13286_, _05749_);
  and _64481_ (_13288_, _13287_, _13285_);
  and _64482_ (_13289_, _13204_, _05748_);
  or _64483_ (_13290_, _13289_, _06440_);
  or _64484_ (_13291_, _13290_, _13288_);
  and _64485_ (_13292_, _12985_, _12792_);
  or _64486_ (_13293_, _13197_, _06444_);
  or _64487_ (_13294_, _13293_, _13292_);
  and _64488_ (_13295_, _13294_, _01317_);
  and _64489_ (_13296_, _13295_, _13291_);
  nor _64490_ (_13297_, \oc8051_golden_model_1.P1 [7], rst);
  nor _64491_ (_13298_, _13297_, _00000_);
  or _64492_ (_40998_, _13298_, _13296_);
  and _64493_ (_13299_, _01321_, \oc8051_golden_model_1.IP [7]);
  not _64494_ (_13300_, _07830_);
  and _64495_ (_13301_, _13300_, \oc8051_golden_model_1.IP [7]);
  and _64496_ (_13302_, _07923_, _07830_);
  or _64497_ (_13303_, _13302_, _13301_);
  or _64498_ (_13304_, _13303_, _06132_);
  not _64499_ (_13305_, _08415_);
  and _64500_ (_13306_, _13305_, \oc8051_golden_model_1.IP [7]);
  and _64501_ (_13307_, _08426_, _08415_);
  or _64502_ (_13308_, _13307_, _13306_);
  and _64503_ (_13309_, _13308_, _06152_);
  and _64504_ (_13310_, _08548_, _07830_);
  or _64505_ (_13311_, _13310_, _13301_);
  or _64506_ (_13312_, _13311_, _06161_);
  and _64507_ (_13313_, _07830_, \oc8051_golden_model_1.ACC [7]);
  or _64508_ (_13314_, _13313_, _13301_);
  and _64509_ (_13315_, _13314_, _07056_);
  and _64510_ (_13316_, _07057_, \oc8051_golden_model_1.IP [7]);
  or _64511_ (_13317_, _13316_, _06160_);
  or _64512_ (_13318_, _13317_, _13315_);
  and _64513_ (_13319_, _13318_, _06157_);
  and _64514_ (_13320_, _13319_, _13312_);
  and _64515_ (_13321_, _08552_, _08415_);
  or _64516_ (_13322_, _13321_, _13306_);
  and _64517_ (_13323_, _13322_, _06156_);
  or _64518_ (_13324_, _13323_, _06217_);
  or _64519_ (_13325_, _13324_, _13320_);
  or _64520_ (_13326_, _13303_, _07075_);
  and _64521_ (_13327_, _13326_, _13325_);
  or _64522_ (_13328_, _13327_, _06220_);
  or _64523_ (_13329_, _13314_, _06229_);
  and _64524_ (_13330_, _13329_, _06153_);
  and _64525_ (_13331_, _13330_, _13328_);
  or _64526_ (_13332_, _13331_, _13309_);
  and _64527_ (_13333_, _13332_, _06146_);
  and _64528_ (_13334_, _08569_, _08415_);
  or _64529_ (_13335_, _13334_, _13306_);
  and _64530_ (_13336_, _13335_, _06145_);
  or _64531_ (_13337_, _13336_, _13333_);
  and _64532_ (_13338_, _13337_, _06140_);
  and _64533_ (_13339_, _08587_, _08415_);
  or _64534_ (_13340_, _13339_, _13306_);
  and _64535_ (_13341_, _13340_, _06139_);
  or _64536_ (_13342_, _13341_, _09842_);
  or _64537_ (_13343_, _13342_, _13338_);
  and _64538_ (_13344_, _13343_, _13304_);
  or _64539_ (_13345_, _13344_, _06116_);
  and _64540_ (_13346_, _08535_, _07830_);
  or _64541_ (_13347_, _13301_, _06117_);
  or _64542_ (_13348_, _13347_, _13346_);
  and _64543_ (_13349_, _13348_, _06114_);
  and _64544_ (_13350_, _13349_, _13345_);
  and _64545_ (_13351_, _08782_, _07830_);
  or _64546_ (_13352_, _13351_, _13301_);
  and _64547_ (_13353_, _13352_, _05787_);
  or _64548_ (_13354_, _13353_, _11136_);
  or _64549_ (_13355_, _13354_, _13350_);
  and _64550_ (_13356_, _08802_, _07830_);
  or _64551_ (_13357_, _13301_, _07127_);
  or _64552_ (_13358_, _13357_, _13356_);
  and _64553_ (_13359_, _08607_, _07830_);
  or _64554_ (_13360_, _13359_, _13301_);
  or _64555_ (_13361_, _13360_, _06111_);
  and _64556_ (_13362_, _13361_, _07125_);
  and _64557_ (_13363_, _13362_, _13358_);
  and _64558_ (_13364_, _13363_, _13355_);
  and _64559_ (_13365_, _08810_, _07830_);
  or _64560_ (_13366_, _13365_, _13301_);
  and _64561_ (_13367_, _13366_, _06402_);
  or _64562_ (_13368_, _13367_, _13364_);
  and _64563_ (_13369_, _13368_, _07132_);
  or _64564_ (_13370_, _13301_, _07926_);
  and _64565_ (_13371_, _13360_, _06306_);
  and _64566_ (_13372_, _13371_, _13370_);
  or _64567_ (_13373_, _13372_, _13369_);
  and _64568_ (_13374_, _13373_, _07130_);
  and _64569_ (_13375_, _13314_, _06411_);
  and _64570_ (_13376_, _13375_, _13370_);
  or _64571_ (_13377_, _13376_, _06303_);
  or _64572_ (_13378_, _13377_, _13374_);
  and _64573_ (_13379_, _08801_, _07830_);
  or _64574_ (_13380_, _13301_, _08819_);
  or _64575_ (_13381_, _13380_, _13379_);
  and _64576_ (_13382_, _13381_, _08824_);
  and _64577_ (_13383_, _13382_, _13378_);
  nor _64578_ (_13384_, _08809_, _13300_);
  or _64579_ (_13385_, _13384_, _13301_);
  and _64580_ (_13386_, _13385_, _06396_);
  or _64581_ (_13387_, _13386_, _06433_);
  or _64582_ (_13388_, _13387_, _13383_);
  or _64583_ (_13389_, _13311_, _06829_);
  and _64584_ (_13390_, _13389_, _05749_);
  and _64585_ (_13391_, _13390_, _13388_);
  and _64586_ (_13392_, _13308_, _05748_);
  or _64587_ (_13393_, _13392_, _06440_);
  or _64588_ (_13394_, _13393_, _13391_);
  and _64589_ (_13395_, _08345_, _07830_);
  or _64590_ (_13396_, _13301_, _06444_);
  or _64591_ (_13397_, _13396_, _13395_);
  and _64592_ (_13398_, _13397_, _01317_);
  and _64593_ (_13399_, _13398_, _13394_);
  or _64594_ (_13400_, _13399_, _13299_);
  and _64595_ (_40999_, _13400_, _43100_);
  and _64596_ (_13401_, _01321_, \oc8051_golden_model_1.IE [7]);
  not _64597_ (_13402_, _07826_);
  and _64598_ (_13403_, _13402_, \oc8051_golden_model_1.IE [7]);
  and _64599_ (_13404_, _07923_, _07826_);
  or _64600_ (_13405_, _13404_, _13403_);
  or _64601_ (_13406_, _13405_, _06132_);
  not _64602_ (_13407_, _08418_);
  and _64603_ (_13408_, _13407_, \oc8051_golden_model_1.IE [7]);
  and _64604_ (_13409_, _08426_, _08418_);
  or _64605_ (_13410_, _13409_, _13408_);
  and _64606_ (_13411_, _13410_, _06152_);
  and _64607_ (_13412_, _08548_, _07826_);
  or _64608_ (_13413_, _13412_, _13403_);
  or _64609_ (_13414_, _13413_, _06161_);
  and _64610_ (_13415_, _07826_, \oc8051_golden_model_1.ACC [7]);
  or _64611_ (_13416_, _13415_, _13403_);
  and _64612_ (_13417_, _13416_, _07056_);
  and _64613_ (_13418_, _07057_, \oc8051_golden_model_1.IE [7]);
  or _64614_ (_13419_, _13418_, _06160_);
  or _64615_ (_13420_, _13419_, _13417_);
  and _64616_ (_13421_, _13420_, _06157_);
  and _64617_ (_13422_, _13421_, _13414_);
  and _64618_ (_13423_, _08552_, _08418_);
  or _64619_ (_13424_, _13423_, _13408_);
  and _64620_ (_13425_, _13424_, _06156_);
  or _64621_ (_13426_, _13425_, _06217_);
  or _64622_ (_13427_, _13426_, _13422_);
  or _64623_ (_13428_, _13405_, _07075_);
  and _64624_ (_13429_, _13428_, _13427_);
  or _64625_ (_13430_, _13429_, _06220_);
  or _64626_ (_13431_, _13416_, _06229_);
  and _64627_ (_13432_, _13431_, _06153_);
  and _64628_ (_13433_, _13432_, _13430_);
  or _64629_ (_13434_, _13433_, _13411_);
  and _64630_ (_13435_, _13434_, _06146_);
  and _64631_ (_13436_, _08569_, _08418_);
  or _64632_ (_13437_, _13436_, _13408_);
  and _64633_ (_13438_, _13437_, _06145_);
  or _64634_ (_13439_, _13438_, _13435_);
  and _64635_ (_13440_, _13439_, _06140_);
  and _64636_ (_13441_, _08587_, _08418_);
  or _64637_ (_13442_, _13441_, _13408_);
  and _64638_ (_13443_, _13442_, _06139_);
  or _64639_ (_13444_, _13443_, _09842_);
  or _64640_ (_13445_, _13444_, _13440_);
  and _64641_ (_13446_, _13445_, _13406_);
  or _64642_ (_13447_, _13446_, _06116_);
  and _64643_ (_13448_, _08535_, _07826_);
  or _64644_ (_13449_, _13403_, _06117_);
  or _64645_ (_13450_, _13449_, _13448_);
  and _64646_ (_13451_, _13450_, _06114_);
  and _64647_ (_13452_, _13451_, _13447_);
  and _64648_ (_13453_, _08782_, _07826_);
  or _64649_ (_13454_, _13453_, _13403_);
  and _64650_ (_13455_, _13454_, _05787_);
  or _64651_ (_13456_, _13455_, _11136_);
  or _64652_ (_13457_, _13456_, _13452_);
  and _64653_ (_13458_, _08802_, _07826_);
  or _64654_ (_13459_, _13403_, _07127_);
  or _64655_ (_13460_, _13459_, _13458_);
  and _64656_ (_13461_, _08607_, _07826_);
  or _64657_ (_13462_, _13461_, _13403_);
  or _64658_ (_13463_, _13462_, _06111_);
  and _64659_ (_13464_, _13463_, _07125_);
  and _64660_ (_13465_, _13464_, _13460_);
  and _64661_ (_13466_, _13465_, _13457_);
  and _64662_ (_13467_, _08810_, _07826_);
  or _64663_ (_13468_, _13467_, _13403_);
  and _64664_ (_13469_, _13468_, _06402_);
  or _64665_ (_13470_, _13469_, _13466_);
  and _64666_ (_13471_, _13470_, _07132_);
  or _64667_ (_13472_, _13403_, _07926_);
  and _64668_ (_13473_, _13462_, _06306_);
  and _64669_ (_13474_, _13473_, _13472_);
  or _64670_ (_13475_, _13474_, _13471_);
  and _64671_ (_13476_, _13475_, _07130_);
  and _64672_ (_13477_, _13416_, _06411_);
  and _64673_ (_13478_, _13477_, _13472_);
  or _64674_ (_13479_, _13478_, _06303_);
  or _64675_ (_13480_, _13479_, _13476_);
  and _64676_ (_13481_, _08801_, _07826_);
  or _64677_ (_13482_, _13403_, _08819_);
  or _64678_ (_13483_, _13482_, _13481_);
  and _64679_ (_13484_, _13483_, _08824_);
  and _64680_ (_13485_, _13484_, _13480_);
  nor _64681_ (_13486_, _08809_, _13402_);
  or _64682_ (_13487_, _13486_, _13403_);
  and _64683_ (_13488_, _13487_, _06396_);
  or _64684_ (_13489_, _13488_, _06433_);
  or _64685_ (_13490_, _13489_, _13485_);
  or _64686_ (_13491_, _13413_, _06829_);
  and _64687_ (_13492_, _13491_, _05749_);
  and _64688_ (_13493_, _13492_, _13490_);
  and _64689_ (_13494_, _13410_, _05748_);
  or _64690_ (_13495_, _13494_, _06440_);
  or _64691_ (_13496_, _13495_, _13493_);
  and _64692_ (_13497_, _08345_, _07826_);
  or _64693_ (_13498_, _13403_, _06444_);
  or _64694_ (_13499_, _13498_, _13497_);
  and _64695_ (_13500_, _13499_, _01317_);
  and _64696_ (_13501_, _13500_, _13496_);
  or _64697_ (_13502_, _13501_, _13401_);
  and _64698_ (_41000_, _13502_, _43100_);
  and _64699_ (_13503_, _01321_, \oc8051_golden_model_1.SCON [7]);
  not _64700_ (_13504_, _07778_);
  and _64701_ (_13505_, _13504_, \oc8051_golden_model_1.SCON [7]);
  and _64702_ (_13506_, _07923_, _07778_);
  or _64703_ (_13507_, _13506_, _13505_);
  or _64704_ (_13508_, _13507_, _06132_);
  not _64705_ (_13509_, _08413_);
  and _64706_ (_13510_, _13509_, \oc8051_golden_model_1.SCON [7]);
  and _64707_ (_13511_, _08426_, _08413_);
  or _64708_ (_13512_, _13511_, _13510_);
  and _64709_ (_13513_, _13512_, _06152_);
  and _64710_ (_13514_, _08548_, _07778_);
  or _64711_ (_13515_, _13514_, _13505_);
  or _64712_ (_13516_, _13515_, _06161_);
  and _64713_ (_13517_, _07778_, \oc8051_golden_model_1.ACC [7]);
  or _64714_ (_13518_, _13517_, _13505_);
  and _64715_ (_13519_, _13518_, _07056_);
  and _64716_ (_13520_, _07057_, \oc8051_golden_model_1.SCON [7]);
  or _64717_ (_13521_, _13520_, _06160_);
  or _64718_ (_13522_, _13521_, _13519_);
  and _64719_ (_13523_, _13522_, _06157_);
  and _64720_ (_13524_, _13523_, _13516_);
  and _64721_ (_13525_, _08552_, _08413_);
  or _64722_ (_13526_, _13525_, _13510_);
  and _64723_ (_13527_, _13526_, _06156_);
  or _64724_ (_13528_, _13527_, _06217_);
  or _64725_ (_13529_, _13528_, _13524_);
  or _64726_ (_13530_, _13507_, _07075_);
  and _64727_ (_13531_, _13530_, _13529_);
  or _64728_ (_13532_, _13531_, _06220_);
  or _64729_ (_13533_, _13518_, _06229_);
  and _64730_ (_13534_, _13533_, _06153_);
  and _64731_ (_13535_, _13534_, _13532_);
  or _64732_ (_13536_, _13535_, _13513_);
  and _64733_ (_13537_, _13536_, _06146_);
  and _64734_ (_13538_, _08569_, _08413_);
  or _64735_ (_13539_, _13538_, _13510_);
  and _64736_ (_13540_, _13539_, _06145_);
  or _64737_ (_13541_, _13540_, _13537_);
  and _64738_ (_13542_, _13541_, _06140_);
  and _64739_ (_13543_, _08587_, _08413_);
  or _64740_ (_13544_, _13543_, _13510_);
  and _64741_ (_13545_, _13544_, _06139_);
  or _64742_ (_13546_, _13545_, _09842_);
  or _64743_ (_13547_, _13546_, _13542_);
  and _64744_ (_13548_, _13547_, _13508_);
  or _64745_ (_13549_, _13548_, _06116_);
  and _64746_ (_13550_, _08535_, _07778_);
  or _64747_ (_13551_, _13505_, _06117_);
  or _64748_ (_13552_, _13551_, _13550_);
  and _64749_ (_13553_, _13552_, _06114_);
  and _64750_ (_13554_, _13553_, _13549_);
  and _64751_ (_13555_, _08782_, _07778_);
  or _64752_ (_13556_, _13555_, _13505_);
  and _64753_ (_13557_, _13556_, _05787_);
  or _64754_ (_13558_, _13557_, _11136_);
  or _64755_ (_13559_, _13558_, _13554_);
  and _64756_ (_13560_, _08802_, _07778_);
  or _64757_ (_13561_, _13505_, _07127_);
  or _64758_ (_13562_, _13561_, _13560_);
  and _64759_ (_13563_, _08607_, _07778_);
  or _64760_ (_13564_, _13563_, _13505_);
  or _64761_ (_13565_, _13564_, _06111_);
  and _64762_ (_13566_, _13565_, _07125_);
  and _64763_ (_13567_, _13566_, _13562_);
  and _64764_ (_13568_, _13567_, _13559_);
  and _64765_ (_13569_, _08810_, _07778_);
  or _64766_ (_13570_, _13569_, _13505_);
  and _64767_ (_13571_, _13570_, _06402_);
  or _64768_ (_13572_, _13571_, _13568_);
  and _64769_ (_13573_, _13572_, _07132_);
  or _64770_ (_13574_, _13505_, _07926_);
  and _64771_ (_13575_, _13564_, _06306_);
  and _64772_ (_13576_, _13575_, _13574_);
  or _64773_ (_13577_, _13576_, _13573_);
  and _64774_ (_13578_, _13577_, _07130_);
  and _64775_ (_13579_, _13518_, _06411_);
  and _64776_ (_13580_, _13579_, _13574_);
  or _64777_ (_13581_, _13580_, _06303_);
  or _64778_ (_13582_, _13581_, _13578_);
  and _64779_ (_13583_, _08801_, _07778_);
  or _64780_ (_13584_, _13505_, _08819_);
  or _64781_ (_13585_, _13584_, _13583_);
  and _64782_ (_13586_, _13585_, _08824_);
  and _64783_ (_13587_, _13586_, _13582_);
  nor _64784_ (_13588_, _08809_, _13504_);
  or _64785_ (_13589_, _13588_, _13505_);
  and _64786_ (_13590_, _13589_, _06396_);
  or _64787_ (_13591_, _13590_, _06433_);
  or _64788_ (_13592_, _13591_, _13587_);
  or _64789_ (_13593_, _13515_, _06829_);
  and _64790_ (_13594_, _13593_, _05749_);
  and _64791_ (_13595_, _13594_, _13592_);
  and _64792_ (_13596_, _13512_, _05748_);
  or _64793_ (_13597_, _13596_, _06440_);
  or _64794_ (_13598_, _13597_, _13595_);
  and _64795_ (_13599_, _08345_, _07778_);
  or _64796_ (_13600_, _13505_, _06444_);
  or _64797_ (_13601_, _13600_, _13599_);
  and _64798_ (_13602_, _13601_, _01317_);
  and _64799_ (_13603_, _13602_, _13598_);
  or _64800_ (_13604_, _13603_, _13503_);
  and _64801_ (_41001_, _13604_, _43100_);
  not _64802_ (_13605_, \oc8051_golden_model_1.SP [7]);
  nor _64803_ (_13606_, _01317_, _13605_);
  and _64804_ (_13607_, _07756_, \oc8051_golden_model_1.SP [4]);
  and _64805_ (_13608_, _13607_, \oc8051_golden_model_1.SP [5]);
  and _64806_ (_13609_, _13608_, \oc8051_golden_model_1.SP [6]);
  or _64807_ (_13610_, _13609_, \oc8051_golden_model_1.SP [7]);
  nand _64808_ (_13611_, _13609_, \oc8051_golden_model_1.SP [7]);
  and _64809_ (_13612_, _13611_, _13610_);
  or _64810_ (_13613_, _13612_, _07160_);
  nor _64811_ (_13614_, _11388_, _07814_);
  and _64812_ (_13615_, _13614_, _07787_);
  nor _64813_ (_13616_, _13615_, _13605_);
  and _64814_ (_13617_, _08810_, _07858_);
  or _64815_ (_13618_, _13617_, _13616_);
  and _64816_ (_13619_, _13618_, _06402_);
  not _64817_ (_13620_, _06133_);
  and _64818_ (_13621_, _07923_, _07858_);
  or _64819_ (_13622_, _13616_, _06116_);
  or _64820_ (_13623_, _13622_, _13621_);
  and _64821_ (_13624_, _13623_, _13620_);
  and _64822_ (_13625_, _08548_, _07858_);
  or _64823_ (_13626_, _13625_, _13616_);
  or _64824_ (_13627_, _13626_, _06161_);
  and _64825_ (_13628_, _13615_, \oc8051_golden_model_1.ACC [7]);
  or _64826_ (_13629_, _13628_, _13616_);
  or _64827_ (_13630_, _13629_, _07057_);
  or _64828_ (_13631_, _07056_, \oc8051_golden_model_1.SP [7]);
  and _64829_ (_13632_, _13631_, _06582_);
  and _64830_ (_13633_, _13632_, _13630_);
  and _64831_ (_13634_, _13612_, _06581_);
  or _64832_ (_13635_, _13634_, _06160_);
  or _64833_ (_13636_, _13635_, _13633_);
  and _64834_ (_13637_, _13636_, _05764_);
  and _64835_ (_13638_, _13637_, _13627_);
  and _64836_ (_13639_, _13612_, _07485_);
  or _64837_ (_13640_, _13639_, _06217_);
  or _64838_ (_13641_, _13640_, _13638_);
  not _64839_ (_13642_, \oc8051_golden_model_1.SP [6]);
  not _64840_ (_13643_, \oc8051_golden_model_1.SP [5]);
  not _64841_ (_13644_, \oc8051_golden_model_1.SP [4]);
  and _64842_ (_13645_, _08453_, _13644_);
  and _64843_ (_13646_, _13645_, _13643_);
  and _64844_ (_13647_, _13646_, _13642_);
  and _64845_ (_13648_, _13647_, _06142_);
  nor _64846_ (_13650_, _13648_, _13605_);
  and _64847_ (_13651_, _13648_, _13605_);
  nor _64848_ (_13652_, _13651_, _13650_);
  nand _64849_ (_13653_, _13652_, _06217_);
  and _64850_ (_13654_, _13653_, _13641_);
  or _64851_ (_13655_, _13654_, _06220_);
  or _64852_ (_13656_, _13629_, _06229_);
  and _64853_ (_13657_, _13656_, _07191_);
  and _64854_ (_13658_, _13657_, _13655_);
  and _64855_ (_13659_, _13608_, \oc8051_golden_model_1.SP [0]);
  and _64856_ (_13661_, _13659_, \oc8051_golden_model_1.SP [6]);
  nor _64857_ (_13662_, _13661_, _13605_);
  and _64858_ (_13663_, _13661_, _13605_);
  or _64859_ (_13664_, _13663_, _13662_);
  nand _64860_ (_13665_, _13664_, _06151_);
  nand _64861_ (_13666_, _13665_, _07389_);
  or _64862_ (_13667_, _13666_, _13658_);
  or _64863_ (_13668_, _13612_, _07389_);
  and _64864_ (_13669_, _13668_, _06132_);
  and _64865_ (_13670_, _13669_, _13667_);
  or _64866_ (_13672_, _13670_, _13624_);
  or _64867_ (_13673_, _13616_, _06117_);
  and _64868_ (_13674_, _08535_, _13615_);
  or _64869_ (_13675_, _13674_, _13673_);
  and _64870_ (_13676_, _13675_, _06114_);
  and _64871_ (_13677_, _13676_, _13672_);
  and _64872_ (_13678_, _08782_, _07858_);
  or _64873_ (_13679_, _13678_, _13616_);
  and _64874_ (_13680_, _13679_, _05787_);
  or _64875_ (_13681_, _13680_, _06110_);
  or _64876_ (_13683_, _13681_, _13677_);
  and _64877_ (_13684_, _08607_, _13615_);
  or _64878_ (_13685_, _13684_, _13616_);
  or _64879_ (_13686_, _13685_, _06111_);
  and _64880_ (_13687_, _13686_, _13683_);
  or _64881_ (_13688_, _13687_, _06076_);
  or _64882_ (_13689_, _13612_, _05836_);
  and _64883_ (_13690_, _13689_, _13688_);
  or _64884_ (_13691_, _13690_, _06297_);
  and _64885_ (_13692_, _08802_, _13615_);
  or _64886_ (_13694_, _13692_, _13616_);
  or _64887_ (_13695_, _13694_, _07127_);
  and _64888_ (_13696_, _13695_, _07125_);
  and _64889_ (_13697_, _13696_, _13691_);
  or _64890_ (_13698_, _13697_, _13619_);
  and _64891_ (_13699_, _13698_, _07132_);
  or _64892_ (_13700_, _13616_, _07926_);
  and _64893_ (_13701_, _13685_, _06306_);
  and _64894_ (_13702_, _13701_, _13700_);
  or _64895_ (_13703_, _13702_, _13699_);
  and _64896_ (_13705_, _13703_, _12514_);
  and _64897_ (_13706_, _13629_, _06411_);
  and _64898_ (_13707_, _13706_, _13700_);
  and _64899_ (_13708_, _13612_, _07124_);
  or _64900_ (_13709_, _13708_, _06303_);
  or _64901_ (_13710_, _13709_, _13707_);
  or _64902_ (_13711_, _13710_, _13705_);
  and _64903_ (_13712_, _08801_, _07858_);
  or _64904_ (_13713_, _13616_, _08819_);
  or _64905_ (_13714_, _13713_, _13712_);
  and _64906_ (_13716_, _13714_, _13711_);
  or _64907_ (_13717_, _13716_, _06396_);
  not _64908_ (_13718_, _07858_);
  nor _64909_ (_13719_, _08809_, _13718_);
  or _64910_ (_13720_, _13616_, _08824_);
  or _64911_ (_13721_, _13720_, _13719_);
  and _64912_ (_13722_, _13721_, _12558_);
  and _64913_ (_13723_, _13722_, _13717_);
  or _64914_ (_13724_, _13647_, \oc8051_golden_model_1.SP [7]);
  nand _64915_ (_13725_, _13647_, \oc8051_golden_model_1.SP [7]);
  and _64916_ (_13727_, _13725_, _13724_);
  and _64917_ (_13728_, _13727_, _06417_);
  or _64918_ (_13729_, _13728_, _07142_);
  or _64919_ (_13730_, _13729_, _13723_);
  or _64920_ (_13731_, _13612_, _05846_);
  and _64921_ (_13732_, _13731_, _13730_);
  or _64922_ (_13733_, _13732_, _06167_);
  or _64923_ (_13734_, _13727_, _06168_);
  and _64924_ (_13735_, _13734_, _06829_);
  and _64925_ (_13736_, _13735_, _13733_);
  and _64926_ (_13738_, _13626_, _06433_);
  or _64927_ (_13739_, _13738_, _07577_);
  or _64928_ (_13740_, _13739_, _13736_);
  and _64929_ (_13741_, _13740_, _13613_);
  or _64930_ (_13742_, _13741_, _06440_);
  and _64931_ (_13743_, _08345_, _07858_);
  or _64932_ (_13744_, _13616_, _06444_);
  or _64933_ (_13745_, _13744_, _13743_);
  and _64934_ (_13746_, _13745_, _01317_);
  and _64935_ (_13747_, _13746_, _13742_);
  or _64936_ (_13749_, _13747_, _13606_);
  and _64937_ (_41003_, _13749_, _43100_);
  not _64938_ (_13750_, _07783_);
  and _64939_ (_13751_, _13750_, \oc8051_golden_model_1.SBUF [7]);
  and _64940_ (_13752_, _08548_, _07783_);
  or _64941_ (_13753_, _13752_, _13751_);
  or _64942_ (_13754_, _13753_, _06161_);
  and _64943_ (_13755_, _07783_, \oc8051_golden_model_1.ACC [7]);
  or _64944_ (_13756_, _13755_, _13751_);
  and _64945_ (_13757_, _13756_, _07056_);
  and _64946_ (_13759_, _07057_, \oc8051_golden_model_1.SBUF [7]);
  or _64947_ (_13760_, _13759_, _06160_);
  or _64948_ (_13761_, _13760_, _13757_);
  and _64949_ (_13762_, _13761_, _07075_);
  and _64950_ (_13763_, _13762_, _13754_);
  and _64951_ (_13764_, _07923_, _07783_);
  or _64952_ (_13765_, _13764_, _13751_);
  and _64953_ (_13766_, _13765_, _06217_);
  or _64954_ (_13767_, _13766_, _13763_);
  and _64955_ (_13768_, _13767_, _06229_);
  and _64956_ (_13770_, _13756_, _06220_);
  or _64957_ (_13771_, _13770_, _09842_);
  or _64958_ (_13772_, _13771_, _13768_);
  or _64959_ (_13773_, _13765_, _06132_);
  and _64960_ (_13774_, _13773_, _13772_);
  or _64961_ (_13775_, _13774_, _06116_);
  and _64962_ (_13776_, _08535_, _07783_);
  or _64963_ (_13777_, _13751_, _06117_);
  or _64964_ (_13778_, _13777_, _13776_);
  and _64965_ (_13779_, _13778_, _06114_);
  and _64966_ (_13781_, _13779_, _13775_);
  and _64967_ (_13782_, _08782_, _07783_);
  or _64968_ (_13783_, _13782_, _13751_);
  and _64969_ (_13784_, _13783_, _05787_);
  or _64970_ (_13785_, _13784_, _13781_);
  or _64971_ (_13786_, _13785_, _11136_);
  and _64972_ (_13787_, _08802_, _07783_);
  or _64973_ (_13788_, _13751_, _07127_);
  or _64974_ (_13789_, _13788_, _13787_);
  and _64975_ (_13790_, _08607_, _07783_);
  or _64976_ (_13792_, _13790_, _13751_);
  or _64977_ (_13793_, _13792_, _06111_);
  and _64978_ (_13794_, _13793_, _07125_);
  and _64979_ (_13795_, _13794_, _13789_);
  and _64980_ (_13796_, _13795_, _13786_);
  and _64981_ (_13797_, _08810_, _07783_);
  or _64982_ (_13798_, _13797_, _13751_);
  and _64983_ (_13799_, _13798_, _06402_);
  or _64984_ (_13800_, _13799_, _13796_);
  and _64985_ (_13801_, _13800_, _07132_);
  or _64986_ (_13802_, _13751_, _07926_);
  and _64987_ (_13803_, _13792_, _06306_);
  and _64988_ (_13804_, _13803_, _13802_);
  or _64989_ (_13805_, _13804_, _13801_);
  and _64990_ (_13806_, _13805_, _07130_);
  and _64991_ (_13807_, _13756_, _06411_);
  and _64992_ (_13808_, _13807_, _13802_);
  or _64993_ (_13809_, _13808_, _06303_);
  or _64994_ (_13810_, _13809_, _13806_);
  and _64995_ (_13811_, _08801_, _07783_);
  or _64996_ (_13812_, _13751_, _08819_);
  or _64997_ (_13813_, _13812_, _13811_);
  and _64998_ (_13814_, _13813_, _08824_);
  and _64999_ (_13815_, _13814_, _13810_);
  nor _65000_ (_13816_, _08809_, _13750_);
  or _65001_ (_13817_, _13816_, _13751_);
  and _65002_ (_13818_, _13817_, _06396_);
  or _65003_ (_13819_, _13818_, _06433_);
  or _65004_ (_13820_, _13819_, _13815_);
  or _65005_ (_13821_, _13753_, _06829_);
  and _65006_ (_13822_, _13821_, _06444_);
  and _65007_ (_13823_, _13822_, _13820_);
  and _65008_ (_13824_, _08345_, _07783_);
  or _65009_ (_13825_, _13824_, _13751_);
  and _65010_ (_13826_, _13825_, _06440_);
  or _65011_ (_13827_, _13826_, _01321_);
  or _65012_ (_13828_, _13827_, _13823_);
  or _65013_ (_13829_, _01317_, \oc8051_golden_model_1.SBUF [7]);
  and _65014_ (_13830_, _13829_, _43100_);
  and _65015_ (_41004_, _13830_, _13828_);
  nor _65016_ (_13831_, _01317_, _10693_);
  and _65017_ (_13832_, _11094_, \oc8051_golden_model_1.ACC [0]);
  nor _65018_ (_13833_, _07794_, _10693_);
  and _65019_ (_13834_, _08810_, _07794_);
  or _65020_ (_13835_, _13834_, _13833_);
  and _65021_ (_13836_, _13835_, _06402_);
  and _65022_ (_13837_, _08782_, _07794_);
  or _65023_ (_13838_, _13837_, _13833_);
  and _65024_ (_13839_, _13838_, _05787_);
  and _65025_ (_13840_, _07923_, _07794_);
  or _65026_ (_13841_, _13840_, _13833_);
  or _65027_ (_13842_, _13841_, _06132_);
  not _65028_ (_13843_, _06254_);
  not _65029_ (_13844_, _06255_);
  nor _65030_ (_13845_, _12682_, _13844_);
  nor _65031_ (_13846_, _09295_, _06255_);
  and _65032_ (_13847_, _08548_, _07794_);
  or _65033_ (_13848_, _13847_, _13833_);
  or _65034_ (_13849_, _13848_, _06161_);
  and _65035_ (_13850_, _07794_, \oc8051_golden_model_1.ACC [7]);
  or _65036_ (_13851_, _13850_, _13833_);
  and _65037_ (_13852_, _13851_, _07056_);
  nor _65038_ (_13853_, _07056_, _10693_);
  or _65039_ (_13854_, _13853_, _06160_);
  or _65040_ (_13855_, _13854_, _13852_);
  and _65041_ (_13856_, _13855_, _10491_);
  and _65042_ (_13857_, _13856_, _13849_);
  nor _65043_ (_13858_, _10508_, _10507_);
  nor _65044_ (_13859_, _13858_, _10491_);
  not _65045_ (_13860_, _06221_);
  or _65046_ (_13861_, _12133_, _13860_);
  or _65047_ (_13862_, _13861_, _13859_);
  or _65048_ (_13863_, _13862_, _13857_);
  nor _65049_ (_13864_, _08404_, _10693_);
  and _65050_ (_13865_, _08552_, _08404_);
  or _65051_ (_13866_, _13865_, _13864_);
  or _65052_ (_13867_, _13866_, _06157_);
  or _65053_ (_13868_, _13841_, _07075_);
  and _65054_ (_13869_, _13868_, _13867_);
  and _65055_ (_13870_, _13869_, _13863_);
  or _65056_ (_13871_, _13870_, _06220_);
  or _65057_ (_13872_, _13851_, _06229_);
  nor _65058_ (_13873_, _12299_, _06152_);
  and _65059_ (_13874_, _13873_, _13872_);
  and _65060_ (_13875_, _13874_, _13871_);
  and _65061_ (_13876_, _08426_, _08404_);
  or _65062_ (_13877_, _13876_, _13864_);
  and _65063_ (_13878_, _13877_, _06152_);
  or _65064_ (_13879_, _13878_, _12126_);
  or _65065_ (_13880_, _13879_, _13875_);
  and _65066_ (_13881_, _12108_, _12109_);
  or _65067_ (_13882_, _13881_, _12106_);
  and _65068_ (_13883_, _12113_, _12112_);
  or _65069_ (_13884_, _13883_, _13882_);
  and _65070_ (_13885_, _13884_, _12105_);
  not _65071_ (_13886_, _12101_);
  nand _65072_ (_13887_, _13886_, _12098_);
  and _65073_ (_13888_, _13887_, _12094_);
  nor _65074_ (_13889_, _13888_, _07924_);
  or _65075_ (_13890_, _13889_, _12119_);
  nor _65076_ (_13891_, _13890_, _13885_);
  nor _65077_ (_13892_, _13891_, _12120_);
  or _65078_ (_13893_, _13892_, _12125_);
  and _65079_ (_13894_, _13893_, _12089_);
  and _65080_ (_13895_, _13894_, _13880_);
  not _65081_ (_13896_, _11929_);
  nand _65082_ (_13897_, _11927_, _13896_);
  nand _65083_ (_13898_, _13897_, _11926_);
  not _65084_ (_13899_, _11934_);
  or _65085_ (_13900_, _11938_, _13899_);
  and _65086_ (_13901_, _13900_, _11932_);
  or _65087_ (_13902_, _13901_, _13898_);
  and _65088_ (_13903_, _13902_, _11954_);
  nor _65089_ (_13904_, _11943_, _08581_);
  nand _65090_ (_13905_, _11951_, _11948_);
  and _65091_ (_13906_, _11946_, _13905_);
  and _65092_ (_13907_, _13906_, _11947_);
  or _65093_ (_13908_, _13907_, _11941_);
  or _65094_ (_13909_, _13908_, _13904_);
  or _65095_ (_13910_, _13909_, _13903_);
  and _65096_ (_13911_, _11956_, _06687_);
  and _65097_ (_13912_, _13911_, _13910_);
  or _65098_ (_13913_, _13912_, _13895_);
  and _65099_ (_13914_, _13913_, _06643_);
  nand _65100_ (_13915_, _08139_, \oc8051_golden_model_1.ACC [3]);
  nor _65101_ (_13916_, _08247_, \oc8051_golden_model_1.ACC [2]);
  nor _65102_ (_13917_, _08139_, \oc8051_golden_model_1.ACC [3]);
  or _65103_ (_13918_, _13917_, _13916_);
  and _65104_ (_13919_, _13918_, _13915_);
  nor _65105_ (_13920_, _08175_, \oc8051_golden_model_1.ACC [1]);
  nor _65106_ (_13921_, _08211_, _05855_);
  nor _65107_ (_13922_, _13921_, _10278_);
  or _65108_ (_13923_, _13922_, _13920_);
  and _65109_ (_13924_, _13923_, _12319_);
  or _65110_ (_13925_, _13924_, _13919_);
  and _65111_ (_13926_, _13925_, _12328_);
  nand _65112_ (_13927_, _08103_, \oc8051_golden_model_1.ACC [5]);
  nor _65113_ (_13928_, _08338_, \oc8051_golden_model_1.ACC [4]);
  nor _65114_ (_13929_, _08103_, \oc8051_golden_model_1.ACC [5]);
  or _65115_ (_13930_, _13929_, _13928_);
  and _65116_ (_13931_, _13930_, _13927_);
  and _65117_ (_13932_, _13931_, _12327_);
  nor _65118_ (_13933_, _07925_, \oc8051_golden_model_1.ACC [7]);
  or _65119_ (_13934_, _08014_, \oc8051_golden_model_1.ACC [6]);
  nor _65120_ (_13935_, _13934_, _08810_);
  or _65121_ (_13936_, _13935_, _13933_);
  or _65122_ (_13937_, _13936_, _13932_);
  or _65123_ (_13938_, _13937_, _13926_);
  nor _65124_ (_13939_, _12329_, _06643_);
  and _65125_ (_13940_, _13939_, _13938_);
  or _65126_ (_13941_, _13940_, _13914_);
  and _65127_ (_13942_, _13941_, _12317_);
  nor _65128_ (_13943_, _06912_, \oc8051_golden_model_1.ACC [1]);
  and _65129_ (_13944_, _06912_, \oc8051_golden_model_1.ACC [1]);
  and _65130_ (_13945_, _06107_, \oc8051_golden_model_1.ACC [0]);
  nor _65131_ (_13946_, _13945_, _13944_);
  or _65132_ (_13947_, _13946_, _13943_);
  and _65133_ (_13948_, _13947_, _12337_);
  nand _65134_ (_13949_, _06070_, \oc8051_golden_model_1.ACC [3]);
  nor _65135_ (_13950_, _06070_, \oc8051_golden_model_1.ACC [3]);
  nor _65136_ (_13951_, _06625_, \oc8051_golden_model_1.ACC [2]);
  or _65137_ (_13952_, _13951_, _13950_);
  and _65138_ (_13953_, _13952_, _13949_);
  or _65139_ (_13954_, _13953_, _13948_);
  and _65140_ (_13955_, _13954_, _12345_);
  nand _65141_ (_13956_, _06477_, \oc8051_golden_model_1.ACC [5]);
  nor _65142_ (_13957_, _06477_, \oc8051_golden_model_1.ACC [5]);
  nor _65143_ (_13958_, _06876_, \oc8051_golden_model_1.ACC [4]);
  or _65144_ (_13959_, _13958_, _13957_);
  and _65145_ (_13960_, _13959_, _13956_);
  and _65146_ (_13961_, _13960_, _12344_);
  and _65147_ (_13962_, _06039_, _08430_);
  or _65148_ (_13963_, _06203_, \oc8051_golden_model_1.ACC [6]);
  nor _65149_ (_13964_, _13963_, _10794_);
  or _65150_ (_13965_, _13964_, _13962_);
  or _65151_ (_13966_, _13965_, _13961_);
  or _65152_ (_13967_, _13966_, _13955_);
  nor _65153_ (_13968_, _12346_, _12317_);
  and _65154_ (_13969_, _13968_, _13967_);
  or _65155_ (_13970_, _13969_, _11924_);
  or _65156_ (_13971_, _13970_, _13942_);
  nand _65157_ (_13972_, _11924_, \oc8051_golden_model_1.PSW [7]);
  and _65158_ (_13973_, _13972_, _06146_);
  and _65159_ (_13974_, _13973_, _13971_);
  or _65160_ (_13975_, _13864_, _08568_);
  and _65161_ (_13976_, _13975_, _06145_);
  and _65162_ (_13977_, _13976_, _13866_);
  nor _65163_ (_13978_, _13977_, _13974_);
  nor _65164_ (_13979_, _13978_, _06212_);
  and _65165_ (_13980_, _12682_, \oc8051_golden_model_1.PSW [7]);
  and _65166_ (_13981_, _13980_, _06212_);
  or _65167_ (_13982_, _13981_, _13979_);
  and _65168_ (_13983_, _13982_, _13846_);
  or _65169_ (_13984_, _13983_, _13845_);
  and _65170_ (_13985_, _13984_, _13843_);
  or _65171_ (_13986_, _12682_, \oc8051_golden_model_1.PSW [7]);
  nand _65172_ (_13987_, _13986_, _06254_);
  nand _65173_ (_13988_, _13987_, _10553_);
  or _65174_ (_13989_, _13988_, _13985_);
  and _65175_ (_13990_, _10302_, _07923_);
  and _65176_ (_13991_, _10313_, _10308_);
  nor _65177_ (_13992_, _13991_, _10306_);
  nand _65178_ (_13993_, _10315_, _10308_);
  or _65179_ (_13994_, _13993_, _10572_);
  and _65180_ (_13995_, _13994_, _13992_);
  or _65181_ (_13996_, _13995_, _13990_);
  and _65182_ (_13997_, _13996_, _10546_);
  or _65183_ (_13998_, _13997_, _10554_);
  and _65184_ (_13999_, _13998_, _13989_);
  and _65185_ (_14000_, _13996_, _10545_);
  or _65186_ (_14001_, _14000_, _12379_);
  or _65187_ (_14002_, _14001_, _13999_);
  and _65188_ (_14003_, _10593_, _10589_);
  nor _65189_ (_14004_, _14003_, _10587_);
  nand _65190_ (_14005_, _10640_, _10589_);
  or _65191_ (_14006_, _14005_, _10638_);
  and _65192_ (_14007_, _14006_, _14004_);
  and _65193_ (_14008_, _10583_, _08535_);
  or _65194_ (_14009_, _14008_, _12380_);
  or _65195_ (_14010_, _14009_, _14007_);
  and _65196_ (_14011_, _14010_, _14002_);
  or _65197_ (_14012_, _14011_, _06260_);
  and _65198_ (_14013_, _10405_, _10401_);
  nor _65199_ (_14014_, _14013_, _10399_);
  nand _65200_ (_14015_, _10447_, _10401_);
  or _65201_ (_14016_, _14015_, _10445_);
  and _65202_ (_14017_, _14016_, _14014_);
  and _65203_ (_14018_, _10395_, _07926_);
  or _65204_ (_14019_, _14018_, _06265_);
  or _65205_ (_14020_, _14019_, _14017_);
  and _65206_ (_14021_, _14020_, _10388_);
  and _65207_ (_14022_, _14021_, _14012_);
  and _65208_ (_14023_, _10665_, _10662_);
  nor _65209_ (_14024_, _14023_, _10660_);
  nand _65210_ (_14025_, _10713_, _10662_);
  or _65211_ (_14026_, _14025_, _10711_);
  and _65212_ (_14027_, _14026_, _14024_);
  or _65213_ (_14028_, _14027_, _10655_);
  and _65214_ (_14029_, _14028_, _10387_);
  or _65215_ (_14030_, _14029_, _09842_);
  or _65216_ (_14031_, _14030_, _14022_);
  and _65217_ (_14032_, _14031_, _13842_);
  or _65218_ (_14033_, _14032_, _06116_);
  and _65219_ (_14034_, _08535_, _07794_);
  or _65220_ (_14035_, _13833_, _06117_);
  or _65221_ (_14036_, _14035_, _14034_);
  and _65222_ (_14037_, _14036_, _06114_);
  and _65223_ (_14038_, _14037_, _14033_);
  or _65224_ (_14039_, _14038_, _13839_);
  nor _65225_ (_14040_, _09855_, _06209_);
  and _65226_ (_14041_, _14040_, _14039_);
  nor _65227_ (_14042_, _12682_, _10693_);
  and _65228_ (_14043_, _14042_, _06209_);
  or _65229_ (_14044_, _14043_, _06110_);
  or _65230_ (_14045_, _14044_, _14041_);
  and _65231_ (_14046_, _08607_, _07794_);
  or _65232_ (_14047_, _14046_, _13833_);
  or _65233_ (_14048_, _14047_, _06111_);
  and _65234_ (_14049_, _14048_, _14045_);
  or _65235_ (_14050_, _14049_, _06208_);
  nand _65236_ (_14051_, _12682_, _10693_);
  or _65237_ (_14052_, _14051_, _06768_);
  and _65238_ (_14053_, _14052_, _14050_);
  or _65239_ (_14054_, _14053_, _06297_);
  and _65240_ (_14055_, _08802_, _07794_);
  or _65241_ (_14056_, _14055_, _13833_);
  or _65242_ (_14057_, _14056_, _07127_);
  and _65243_ (_14058_, _14057_, _07125_);
  and _65244_ (_14059_, _14058_, _14054_);
  or _65245_ (_14060_, _14059_, _13836_);
  and _65246_ (_14061_, _14060_, _07132_);
  or _65247_ (_14062_, _13833_, _07926_);
  and _65248_ (_14063_, _14047_, _06306_);
  and _65249_ (_14064_, _14063_, _14062_);
  or _65250_ (_14065_, _14064_, _14061_);
  and _65251_ (_14066_, _14065_, _07130_);
  and _65252_ (_14067_, _13851_, _06411_);
  and _65253_ (_14068_, _14067_, _14062_);
  or _65254_ (_14069_, _14068_, _06303_);
  or _65255_ (_14070_, _14069_, _14066_);
  and _65256_ (_14071_, _08801_, _07794_);
  or _65257_ (_14072_, _13833_, _08819_);
  or _65258_ (_14073_, _14072_, _14071_);
  and _65259_ (_14074_, _14073_, _08824_);
  and _65260_ (_14075_, _14074_, _14070_);
  not _65261_ (_14076_, _07794_);
  nor _65262_ (_14077_, _08809_, _14076_);
  or _65263_ (_14078_, _14077_, _13833_);
  and _65264_ (_14079_, _14078_, _06396_);
  or _65265_ (_14080_, _14079_, _12547_);
  or _65266_ (_14081_, _14080_, _14075_);
  nor _65267_ (_14082_, _10586_, _08430_);
  or _65268_ (_14083_, _14082_, _10889_);
  or _65269_ (_14084_, _10867_, _14008_);
  or _65270_ (_14085_, _14084_, _14083_);
  nor _65271_ (_14086_, _10305_, _08430_);
  or _65272_ (_14087_, _14086_, _10368_);
  or _65273_ (_14088_, _10380_, _13990_);
  or _65274_ (_14089_, _14088_, _14087_);
  and _65275_ (_14090_, _14089_, _06407_);
  and _65276_ (_14091_, _14090_, _14085_);
  and _65277_ (_14092_, _14091_, _14081_);
  nor _65278_ (_14093_, _10398_, _08430_);
  or _65279_ (_14094_, _14093_, _10919_);
  or _65280_ (_14095_, _10895_, _14018_);
  or _65281_ (_14096_, _14095_, _14094_);
  and _65282_ (_14097_, _14096_, _10897_);
  or _65283_ (_14098_, _14097_, _14092_);
  and _65284_ (_14099_, _10659_, \oc8051_golden_model_1.ACC [7]);
  or _65285_ (_14100_, _14099_, _10949_);
  or _65286_ (_14101_, _10927_, _10655_);
  or _65287_ (_14102_, _14101_, _14100_);
  and _65288_ (_14103_, _14102_, _10926_);
  and _65289_ (_14104_, _14103_, _14098_);
  nand _65290_ (_14105_, _10925_, \oc8051_golden_model_1.ACC [7]);
  nand _65291_ (_14106_, _14105_, _10962_);
  or _65292_ (_14107_, _14106_, _14104_);
  nor _65293_ (_14108_, _10997_, _10763_);
  or _65294_ (_14109_, _14108_, _10765_);
  and _65295_ (_14110_, _14109_, _10957_);
  or _65296_ (_14111_, _14110_, _10963_);
  and _65297_ (_14112_, _14111_, _14107_);
  and _65298_ (_14113_, _14109_, _10956_);
  or _65299_ (_14114_, _14113_, _11003_);
  or _65300_ (_14115_, _14114_, _14112_);
  and _65301_ (_14116_, _11038_, _10783_);
  not _65302_ (_14117_, _10781_);
  or _65303_ (_14118_, _11005_, _10782_);
  and _65304_ (_14119_, _14118_, _14117_);
  or _65305_ (_14120_, _14119_, _11041_);
  or _65306_ (_14121_, _14120_, _14116_);
  and _65307_ (_14122_, _14121_, _06171_);
  and _65308_ (_14123_, _14122_, _14115_);
  not _65309_ (_14124_, _08809_);
  not _65310_ (_14125_, _08808_);
  nand _65311_ (_14126_, _10297_, _14125_);
  and _65312_ (_14127_, _14126_, _06169_);
  and _65313_ (_14128_, _14127_, _14124_);
  or _65314_ (_14129_, _14128_, _10264_);
  or _65315_ (_14130_, _14129_, _14123_);
  not _65316_ (_14131_, _10793_);
  or _65317_ (_14132_, _11080_, _10792_);
  and _65318_ (_14133_, _14132_, _10264_);
  nand _65319_ (_14134_, _14133_, _14131_);
  and _65320_ (_14135_, _14134_, _06829_);
  and _65321_ (_14136_, _14135_, _14130_);
  and _65322_ (_14137_, _13848_, _06433_);
  nor _65323_ (_14138_, _14137_, _14136_);
  nor _65324_ (_14139_, _14138_, _11094_);
  or _65325_ (_14140_, _14139_, _13832_);
  and _65326_ (_14141_, _14140_, _05749_);
  and _65327_ (_14142_, _13877_, _05748_);
  or _65328_ (_14143_, _14142_, _06440_);
  or _65329_ (_14144_, _14143_, _14141_);
  and _65330_ (_14145_, _08345_, _07794_);
  or _65331_ (_14146_, _13833_, _06444_);
  or _65332_ (_14147_, _14146_, _14145_);
  and _65333_ (_14148_, _14147_, _01317_);
  and _65334_ (_14149_, _14148_, _14144_);
  or _65335_ (_14150_, _14149_, _13831_);
  and _65336_ (_41005_, _14150_, _43100_);
  nor _65337_ (_14151_, _07593_, _07418_);
  nor _65338_ (_14152_, _14151_, _07747_);
  nor _65339_ (_14153_, _07418_, _07174_);
  nor _65340_ (_14154_, _14153_, _07419_);
  and _65341_ (_14155_, _14154_, _07417_);
  and _65342_ (_14156_, _14155_, _14152_);
  or _65343_ (_14157_, _14156_, \oc8051_golden_model_1.IRAM[0] [0]);
  and _65344_ (_14158_, _07764_, _07755_);
  nor _65345_ (_14159_, _07765_, _14158_);
  and _65346_ (_14160_, _14159_, _07178_);
  and _65347_ (_14161_, _14160_, _07764_);
  not _65348_ (_14162_, _14161_);
  and _65349_ (_14163_, _14162_, _14157_);
  not _65350_ (_14164_, _14156_);
  nand _65351_ (_14165_, _05823_, _05444_);
  not _65352_ (_14166_, _08825_);
  or _65353_ (_14167_, _08211_, _08708_);
  and _65354_ (_14168_, _14167_, _08820_);
  or _65355_ (_14169_, _12660_, _07772_);
  nand _65356_ (_14170_, _07772_, _10693_);
  and _65357_ (_14171_, _14170_, _14169_);
  and _65358_ (_14172_, _14171_, _07103_);
  or _65359_ (_14173_, _08211_, _06251_);
  not _65360_ (_14174_, _07772_);
  and _65361_ (_14175_, _12660_, _14174_);
  or _65362_ (_14176_, _14175_, _08398_);
  nor _65363_ (_14177_, _08443_, _07049_);
  and _65364_ (_14178_, _06581_, \oc8051_golden_model_1.PC [0]);
  nor _65365_ (_14179_, _06581_, _05855_);
  or _65366_ (_14180_, _14179_, _14178_);
  and _65367_ (_14181_, _14180_, _08443_);
  or _65368_ (_14182_, _14181_, _14177_);
  and _65369_ (_14183_, _14182_, _08429_);
  nor _65370_ (_14184_, _08211_, _08429_);
  or _65371_ (_14185_, _14184_, _14183_);
  and _65372_ (_14186_, _14185_, _08428_);
  and _65373_ (_14187_, _14169_, _06159_);
  or _65374_ (_14188_, _14187_, _07485_);
  or _65375_ (_14189_, _14188_, _14186_);
  nor _65376_ (_14190_, _05764_, \oc8051_golden_model_1.PC [0]);
  nor _65377_ (_14191_, _14190_, _07076_);
  and _65378_ (_14192_, _14191_, _14189_);
  and _65379_ (_14193_, _07076_, _07049_);
  or _65380_ (_14194_, _14193_, _07086_);
  or _65381_ (_14195_, _14194_, _14192_);
  and _65382_ (_14196_, _14195_, _14176_);
  or _65383_ (_14197_, _14196_, _06151_);
  or _65384_ (_14198_, _08211_, _07191_);
  and _65385_ (_14199_, _14198_, _06149_);
  and _65386_ (_14200_, _14199_, _14197_);
  nor _65387_ (_14201_, _12661_, _06149_);
  and _65388_ (_14202_, _14201_, _14169_);
  or _65389_ (_14203_, _14202_, _14200_);
  and _65390_ (_14204_, _14203_, _05760_);
  or _65391_ (_14205_, _05760_, _05444_);
  nand _65392_ (_14206_, _06251_, _14205_);
  or _65393_ (_14207_, _14206_, _14204_);
  and _65394_ (_14208_, _14207_, _14173_);
  or _65395_ (_14209_, _14208_, _06701_);
  and _65396_ (_14210_, _09160_, _06172_);
  or _65397_ (_14211_, _08209_, _07104_);
  or _65398_ (_14212_, _14211_, _14210_);
  and _65399_ (_14213_, _14212_, _08580_);
  and _65400_ (_14214_, _14213_, _14209_);
  or _65401_ (_14215_, _14214_, _14172_);
  or _65402_ (_14216_, _14215_, _05791_);
  and _65403_ (_14217_, _05791_, _05444_);
  nor _65404_ (_14218_, _14217_, _08591_);
  and _65405_ (_14219_, _14218_, _14216_);
  and _65406_ (_14220_, _08591_, _07049_);
  or _65407_ (_14221_, _14220_, _08595_);
  or _65408_ (_14222_, _14221_, _14219_);
  or _65409_ (_14223_, _09160_, _08601_);
  and _65410_ (_14224_, _14223_, _08600_);
  and _65411_ (_14225_, _14224_, _14222_);
  and _65412_ (_14226_, _08395_, _07049_);
  and _65413_ (_14227_, _08765_, \oc8051_golden_model_1.DPL [0]);
  and _65414_ (_14228_, _08760_, \oc8051_golden_model_1.DPH [0]);
  and _65415_ (_14229_, _08758_, \oc8051_golden_model_1.SP [0]);
  or _65416_ (_14230_, _14229_, _14228_);
  or _65417_ (_14231_, _14230_, _14227_);
  and _65418_ (_14232_, _08726_, \oc8051_golden_model_1.TCON [0]);
  and _65419_ (_14233_, _08775_, \oc8051_golden_model_1.TMOD [0]);
  and _65420_ (_14234_, _08773_, \oc8051_golden_model_1.TL0 [0]);
  or _65421_ (_14235_, _14234_, _14233_);
  or _65422_ (_14236_, _14235_, _14232_);
  or _65423_ (_14237_, _14236_, _14231_);
  and _65424_ (_14238_, _08734_, \oc8051_golden_model_1.PSW [0]);
  and _65425_ (_14239_, _08738_, \oc8051_golden_model_1.ACC [0]);
  and _65426_ (_14240_, _08741_, \oc8051_golden_model_1.B [0]);
  or _65427_ (_14241_, _14240_, _14239_);
  or _65428_ (_14242_, _14241_, _14238_);
  and _65429_ (_14243_, _08746_, \oc8051_golden_model_1.IP [0]);
  and _65430_ (_14244_, _08749_, \oc8051_golden_model_1.IE [0]);
  and _65431_ (_14245_, _08752_, \oc8051_golden_model_1.SBUF [0]);
  or _65432_ (_14246_, _14245_, _14244_);
  or _65433_ (_14247_, _14246_, _14243_);
  or _65434_ (_14248_, _14247_, _14242_);
  and _65435_ (_14249_, _08724_, \oc8051_golden_model_1.TL1 [0]);
  and _65436_ (_14250_, _08710_, \oc8051_golden_model_1.TH1 [0]);
  and _65437_ (_14251_, _08718_, \oc8051_golden_model_1.SCON [0]);
  or _65438_ (_14252_, _14251_, _14250_);
  or _65439_ (_14253_, _14252_, _14249_);
  and _65440_ (_14254_, _08706_, \oc8051_golden_model_1.TH0 [0]);
  and _65441_ (_14255_, _08770_, \oc8051_golden_model_1.PCON [0]);
  or _65442_ (_14256_, _14255_, _14254_);
  or _65443_ (_14257_, _14256_, _14253_);
  or _65444_ (_14258_, _14257_, _14248_);
  or _65445_ (_14259_, _14258_, _14237_);
  or _65446_ (_14260_, _14259_, _14226_);
  and _65447_ (_14261_, _14260_, _08599_);
  or _65448_ (_14262_, _14261_, _08788_);
  or _65449_ (_14263_, _14262_, _14225_);
  and _65450_ (_14264_, _08788_, _06107_);
  nor _65451_ (_14265_, _14264_, _06112_);
  and _65452_ (_14266_, _14265_, _14263_);
  and _65453_ (_14267_, _08708_, _06112_);
  or _65454_ (_14268_, _14267_, _06076_);
  or _65455_ (_14269_, _14268_, _14266_);
  nor _65456_ (_14270_, _05836_, \oc8051_golden_model_1.PC [0]);
  nor _65457_ (_14271_, _14270_, _07128_);
  and _65458_ (_14272_, _14271_, _14269_);
  and _65459_ (_14273_, _08211_, _08708_);
  not _65460_ (_14274_, _14273_);
  and _65461_ (_14275_, _14274_, _14167_);
  and _65462_ (_14276_, _14275_, _07128_);
  or _65463_ (_14277_, _14276_, _14272_);
  and _65464_ (_14278_, _14277_, _08807_);
  nor _65465_ (_14279_, _12322_, _08807_);
  or _65466_ (_14280_, _14279_, _07133_);
  or _65467_ (_14281_, _14280_, _14278_);
  or _65468_ (_14282_, _14273_, _08806_);
  and _65469_ (_14283_, _14282_, _08364_);
  and _65470_ (_14284_, _14283_, _14281_);
  and _65471_ (_14285_, _10276_, _07131_);
  or _65472_ (_14286_, _14285_, _07124_);
  or _65473_ (_14287_, _14286_, _14284_);
  nor _65474_ (_14288_, _05848_, \oc8051_golden_model_1.PC [0]);
  nor _65475_ (_14289_, _14288_, _08820_);
  and _65476_ (_14290_, _14289_, _14287_);
  or _65477_ (_14291_, _14290_, _14168_);
  and _65478_ (_14292_, _14291_, _14166_);
  nor _65479_ (_14293_, _12321_, _14166_);
  or _65480_ (_14294_, _14293_, _07142_);
  or _65481_ (_14295_, _14294_, _14292_);
  or _65482_ (_14296_, _05846_, \oc8051_golden_model_1.PC [0]);
  and _65483_ (_14297_, _14296_, _08362_);
  and _65484_ (_14298_, _14297_, _14295_);
  nor _65485_ (_14299_, _08362_, _07049_);
  or _65486_ (_14300_, _14299_, _14298_);
  and _65487_ (_14301_, _14300_, _07154_);
  nor _65488_ (_14302_, _09160_, _07154_);
  or _65489_ (_14303_, _14302_, _07152_);
  or _65490_ (_14304_, _14303_, _14301_);
  nand _65491_ (_14305_, _08211_, _07152_);
  and _65492_ (_14306_, _14305_, _12723_);
  and _65493_ (_14307_, _14306_, _14304_);
  and _65494_ (_14308_, _06310_, _05444_);
  or _65495_ (_14309_, _14308_, _05823_);
  or _65496_ (_14310_, _14309_, _14307_);
  and _65497_ (_14311_, _14310_, _14165_);
  or _65498_ (_14312_, _14311_, _06073_);
  or _65499_ (_14313_, _14175_, _06074_);
  and _65500_ (_14314_, _14313_, _09193_);
  and _65501_ (_14315_, _14314_, _14312_);
  nor _65502_ (_14316_, _09193_, _07049_);
  or _65503_ (_14317_, _14316_, _14315_);
  and _65504_ (_14318_, _14317_, _07169_);
  nor _65505_ (_14319_, _09160_, _07169_);
  or _65506_ (_14320_, _14319_, _07167_);
  or _65507_ (_14321_, _14320_, _14318_);
  nand _65508_ (_14322_, _08211_, _07167_);
  and _65509_ (_14323_, _14322_, _07417_);
  and _65510_ (_14324_, _14323_, _14321_);
  or _65511_ (_14325_, _14324_, _14164_);
  and _65512_ (_14326_, _14325_, _14163_);
  and _65513_ (_14327_, _07764_, _07178_);
  and _65514_ (_14328_, _14327_, _14159_);
  nand _65515_ (_14329_, _12057_, _06310_);
  or _65516_ (_14330_, _12224_, _06310_);
  and _65517_ (_14331_, _14330_, _14329_);
  and _65518_ (_14332_, _14331_, _07764_);
  and _65519_ (_14333_, _14332_, _14328_);
  or _65520_ (_41013_, _14333_, _14326_);
  or _65521_ (_14334_, _14156_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _65522_ (_14335_, _14334_, _14162_);
  and _65523_ (_14336_, _06284_, _05820_);
  nor _65524_ (_14337_, _09212_, _09161_);
  and _65525_ (_14338_, _14337_, _14336_);
  not _65526_ (_14339_, _14336_);
  or _65527_ (_14340_, _09195_, _08352_);
  nor _65528_ (_14341_, _14340_, _09193_);
  nor _65529_ (_14342_, _05846_, \oc8051_golden_model_1.PC [1]);
  nand _65530_ (_14343_, _08175_, _06945_);
  nor _65531_ (_14344_, _08175_, _06945_);
  not _65532_ (_14345_, _14344_);
  and _65533_ (_14346_, _14345_, _14343_);
  and _65534_ (_14347_, _14346_, _07128_);
  not _65535_ (_14348_, _07781_);
  and _65536_ (_14349_, _12627_, _14348_);
  and _65537_ (_14350_, _07781_, \oc8051_golden_model_1.PSW [7]);
  or _65538_ (_14351_, _14350_, _14349_);
  and _65539_ (_14352_, _14351_, _07103_);
  nand _65540_ (_14353_, _08175_, _06252_);
  or _65541_ (_14354_, _14349_, _08398_);
  or _65542_ (_14355_, _14340_, _08443_);
  nor _65543_ (_14356_, _06581_, _05887_);
  and _65544_ (_14357_, _06581_, _05407_);
  or _65545_ (_14358_, _14357_, _14356_);
  nor _65546_ (_14359_, _14358_, _07377_);
  nand _65547_ (_14360_, _14359_, _07667_);
  and _65548_ (_14361_, _14360_, _14355_);
  and _65549_ (_14362_, _14361_, _08429_);
  nor _65550_ (_14363_, _08541_, _08212_);
  nor _65551_ (_14364_, _14363_, _08429_);
  or _65552_ (_14365_, _14364_, _14362_);
  or _65553_ (_14366_, _14365_, _06159_);
  or _65554_ (_14367_, _12627_, _07781_);
  or _65555_ (_14368_, _14367_, _08428_);
  and _65556_ (_14369_, _14368_, _14366_);
  or _65557_ (_14370_, _14369_, _07485_);
  nor _65558_ (_14371_, _05764_, _05407_);
  nor _65559_ (_14372_, _14371_, _07076_);
  and _65560_ (_14373_, _14372_, _14370_);
  and _65561_ (_14374_, _07306_, _07076_);
  or _65562_ (_14375_, _14374_, _07086_);
  or _65563_ (_14376_, _14375_, _14373_);
  and _65564_ (_14377_, _14376_, _14354_);
  or _65565_ (_14378_, _14377_, _06151_);
  nand _65566_ (_14379_, _08175_, _06151_);
  and _65567_ (_14380_, _14379_, _06149_);
  and _65568_ (_14381_, _14380_, _14378_);
  not _65569_ (_14382_, _12628_);
  and _65570_ (_14383_, _14367_, _14382_);
  and _65571_ (_14384_, _14383_, _06148_);
  or _65572_ (_14385_, _14384_, _14381_);
  and _65573_ (_14386_, _14385_, _05760_);
  or _65574_ (_14387_, _05760_, \oc8051_golden_model_1.PC [1]);
  nand _65575_ (_14388_, _06251_, _14387_);
  or _65576_ (_14389_, _14388_, _14386_);
  and _65577_ (_14390_, _14389_, _14353_);
  or _65578_ (_14391_, _14390_, _06701_);
  and _65579_ (_14392_, _09115_, _06172_);
  or _65580_ (_14393_, _08173_, _07104_);
  or _65581_ (_14394_, _14393_, _14392_);
  and _65582_ (_14395_, _14394_, _08580_);
  and _65583_ (_14396_, _14395_, _14391_);
  or _65584_ (_14397_, _14396_, _14352_);
  or _65585_ (_14398_, _14397_, _05791_);
  and _65586_ (_14399_, _05791_, \oc8051_golden_model_1.PC [1]);
  nor _65587_ (_14400_, _14399_, _08591_);
  and _65588_ (_14401_, _14400_, _14398_);
  and _65589_ (_14402_, _07306_, _08591_);
  or _65590_ (_14403_, _14402_, _08595_);
  or _65591_ (_14404_, _14403_, _14401_);
  or _65592_ (_14405_, _09115_, _08601_);
  and _65593_ (_14406_, _14405_, _08600_);
  and _65594_ (_14407_, _14406_, _14404_);
  and _65595_ (_14408_, _08395_, _07306_);
  and _65596_ (_14409_, _08773_, \oc8051_golden_model_1.TL0 [1]);
  and _65597_ (_14410_, _08775_, \oc8051_golden_model_1.TMOD [1]);
  and _65598_ (_14411_, _08710_, \oc8051_golden_model_1.TH1 [1]);
  or _65599_ (_14412_, _14411_, _14410_);
  or _65600_ (_14413_, _14412_, _14409_);
  and _65601_ (_14414_, _08724_, \oc8051_golden_model_1.TL1 [1]);
  and _65602_ (_14415_, _08770_, \oc8051_golden_model_1.PCON [1]);
  and _65603_ (_14416_, _08760_, \oc8051_golden_model_1.DPH [1]);
  or _65604_ (_14417_, _14416_, _14415_);
  or _65605_ (_14418_, _14417_, _14414_);
  and _65606_ (_14419_, _08738_, \oc8051_golden_model_1.ACC [1]);
  and _65607_ (_14420_, _08741_, \oc8051_golden_model_1.B [1]);
  or _65608_ (_14421_, _14420_, _14419_);
  and _65609_ (_14422_, _08749_, \oc8051_golden_model_1.IE [1]);
  and _65610_ (_14423_, _08746_, \oc8051_golden_model_1.IP [1]);
  or _65611_ (_14424_, _14423_, _14422_);
  or _65612_ (_14425_, _14424_, _14421_);
  and _65613_ (_14426_, _08765_, \oc8051_golden_model_1.DPL [1]);
  and _65614_ (_14427_, _08758_, \oc8051_golden_model_1.SP [1]);
  or _65615_ (_14428_, _14427_, _14426_);
  or _65616_ (_14429_, _14428_, _14425_);
  and _65617_ (_14430_, _08706_, \oc8051_golden_model_1.TH0 [1]);
  and _65618_ (_14431_, _08726_, \oc8051_golden_model_1.TCON [1]);
  and _65619_ (_14432_, _08734_, \oc8051_golden_model_1.PSW [1]);
  or _65620_ (_14433_, _14432_, _14431_);
  and _65621_ (_14434_, _08718_, \oc8051_golden_model_1.SCON [1]);
  and _65622_ (_14435_, _08752_, \oc8051_golden_model_1.SBUF [1]);
  or _65623_ (_14436_, _14435_, _14434_);
  or _65624_ (_14437_, _14436_, _14433_);
  or _65625_ (_14438_, _14437_, _14430_);
  or _65626_ (_14439_, _14438_, _14429_);
  or _65627_ (_14440_, _14439_, _14418_);
  or _65628_ (_14441_, _14440_, _14413_);
  or _65629_ (_14442_, _14441_, _14408_);
  and _65630_ (_14443_, _14442_, _08599_);
  or _65631_ (_14444_, _14443_, _08788_);
  or _65632_ (_14445_, _14444_, _14407_);
  and _65633_ (_14446_, _08788_, _06912_);
  nor _65634_ (_14447_, _14446_, _06112_);
  and _65635_ (_14448_, _14447_, _14445_);
  and _65636_ (_14449_, _08763_, _06112_);
  or _65637_ (_14450_, _14449_, _06076_);
  or _65638_ (_14451_, _14450_, _14448_);
  nor _65639_ (_14452_, _05836_, _05407_);
  nor _65640_ (_14453_, _14452_, _07128_);
  and _65641_ (_14454_, _14453_, _14451_);
  or _65642_ (_14455_, _14454_, _14347_);
  and _65643_ (_14456_, _14455_, _08807_);
  and _65644_ (_14457_, _10278_, _07126_);
  or _65645_ (_14458_, _14457_, _07133_);
  or _65646_ (_14459_, _14458_, _14456_);
  or _65647_ (_14460_, _14344_, _08806_);
  and _65648_ (_14461_, _14460_, _08364_);
  and _65649_ (_14462_, _14461_, _14459_);
  and _65650_ (_14463_, _10275_, _07131_);
  or _65651_ (_14464_, _14463_, _07124_);
  or _65652_ (_14465_, _14464_, _14462_);
  nor _65653_ (_14466_, _05848_, _05407_);
  nor _65654_ (_14467_, _14466_, _08820_);
  and _65655_ (_14468_, _14467_, _14465_);
  and _65656_ (_14469_, _14343_, _08820_);
  or _65657_ (_14470_, _14469_, _08825_);
  or _65658_ (_14471_, _14470_, _14468_);
  nand _65659_ (_14472_, _10277_, _08825_);
  and _65660_ (_14473_, _14472_, _05846_);
  and _65661_ (_14474_, _14473_, _14471_);
  nor _65662_ (_14475_, _14474_, _14342_);
  nor _65663_ (_14476_, _14475_, _06530_);
  and _65664_ (_14477_, _14340_, _06530_);
  or _65665_ (_14478_, _14477_, _06565_);
  or _65666_ (_14479_, _14478_, _14476_);
  not _65667_ (_14480_, _06972_);
  or _65668_ (_14481_, _14340_, _06564_);
  and _65669_ (_14482_, _14481_, _14480_);
  and _65670_ (_14483_, _14482_, _14479_);
  and _65671_ (_14484_, _14340_, _06972_);
  or _65672_ (_14485_, _14484_, _07325_);
  or _65673_ (_14486_, _14485_, _14483_);
  and _65674_ (_14487_, _06284_, _05591_);
  not _65675_ (_14488_, _14487_);
  or _65676_ (_14489_, _14340_, _07326_);
  and _65677_ (_14490_, _14489_, _14488_);
  and _65678_ (_14491_, _14490_, _14486_);
  nand _65679_ (_14492_, _14337_, _06276_);
  and _65680_ (_14493_, _14492_, _07153_);
  or _65681_ (_14494_, _14493_, _14491_);
  and _65682_ (_14495_, _06281_, _05591_);
  nand _65683_ (_14496_, _14337_, _14495_);
  and _65684_ (_14497_, _14496_, _08837_);
  and _65685_ (_14498_, _14497_, _14494_);
  nor _65686_ (_14499_, _14363_, _08837_);
  or _65687_ (_14500_, _14499_, _06310_);
  or _65688_ (_14501_, _14500_, _14498_);
  nand _65689_ (_14502_, _06310_, _05879_);
  and _65690_ (_14503_, _14502_, _12730_);
  and _65691_ (_14504_, _14503_, _14501_);
  and _65692_ (_14505_, _05823_, _05407_);
  or _65693_ (_14506_, _06073_, _14505_);
  or _65694_ (_14507_, _14506_, _14504_);
  or _65695_ (_14508_, _14349_, _06074_);
  and _65696_ (_14509_, _14508_, _09193_);
  and _65697_ (_14510_, _14509_, _14507_);
  or _65698_ (_14511_, _14510_, _14341_);
  and _65699_ (_14512_, _14511_, _14339_);
  or _65700_ (_14513_, _14512_, _14338_);
  and _65701_ (_14514_, _14513_, _06835_);
  and _65702_ (_14515_, _14337_, _06834_);
  or _65703_ (_14516_, _14515_, _07167_);
  or _65704_ (_14517_, _14516_, _14514_);
  not _65705_ (_14518_, _07167_);
  or _65706_ (_14519_, _14363_, _14518_);
  and _65707_ (_14520_, _14519_, _07417_);
  and _65708_ (_14521_, _14520_, _14517_);
  or _65709_ (_14522_, _14521_, _14164_);
  and _65710_ (_14523_, _14522_, _14335_);
  nand _65711_ (_14524_, _11997_, _06310_);
  or _65712_ (_14525_, _12172_, _06310_);
  and _65713_ (_14526_, _14525_, _14524_);
  and _65714_ (_14527_, _14526_, _07764_);
  and _65715_ (_14528_, _14527_, _14328_);
  or _65716_ (_41014_, _14528_, _14523_);
  or _65717_ (_14529_, _14156_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _65718_ (_14530_, _14529_, _14162_);
  nor _65719_ (_14531_, _05923_, _05846_);
  and _65720_ (_14532_, _09211_, _06172_);
  or _65721_ (_14533_, _14532_, _08245_);
  and _65722_ (_14534_, _14533_, _06701_);
  not _65723_ (_14535_, _07848_);
  and _65724_ (_14536_, _12644_, _14535_);
  or _65725_ (_14537_, _14536_, _08398_);
  or _65726_ (_14538_, _12644_, _07848_);
  or _65727_ (_14539_, _14538_, _08428_);
  nand _65728_ (_14540_, _08541_, _08247_);
  or _65729_ (_14541_, _08541_, _08247_);
  nand _65730_ (_14542_, _14541_, _14540_);
  and _65731_ (_14543_, _14542_, _06162_);
  and _65732_ (_14544_, _08352_, _07657_);
  nor _65733_ (_14545_, _08352_, _07657_);
  nor _65734_ (_14546_, _14545_, _14544_);
  nand _65735_ (_14547_, _14546_, _08445_);
  and _65736_ (_14548_, _06581_, _05921_);
  nor _65737_ (_14549_, _06581_, _09981_);
  nor _65738_ (_14550_, _14549_, _14548_);
  and _65739_ (_14551_, _14550_, _08443_);
  nor _65740_ (_14552_, _14551_, _06162_);
  and _65741_ (_14553_, _14552_, _14547_);
  or _65742_ (_14554_, _14553_, _06159_);
  or _65743_ (_14555_, _14554_, _14543_);
  and _65744_ (_14556_, _14555_, _14539_);
  or _65745_ (_14557_, _14556_, _07485_);
  nor _65746_ (_14558_, _05921_, _05764_);
  nor _65747_ (_14559_, _14558_, _07076_);
  and _65748_ (_14560_, _14559_, _14557_);
  and _65749_ (_14561_, _07708_, _07076_);
  or _65750_ (_14562_, _14561_, _07086_);
  or _65751_ (_14563_, _14562_, _14560_);
  and _65752_ (_14564_, _14563_, _14537_);
  or _65753_ (_14565_, _14564_, _06151_);
  nand _65754_ (_14566_, _08247_, _06151_);
  and _65755_ (_14567_, _14566_, _06149_);
  and _65756_ (_14568_, _14567_, _14565_);
  not _65757_ (_14569_, _12645_);
  and _65758_ (_14570_, _14538_, _14569_);
  and _65759_ (_14571_, _14570_, _06148_);
  or _65760_ (_14572_, _14571_, _14568_);
  and _65761_ (_14573_, _14572_, _05760_);
  or _65762_ (_14574_, _05923_, _05760_);
  nand _65763_ (_14575_, _06251_, _14574_);
  or _65764_ (_14576_, _14575_, _14573_);
  nand _65765_ (_14577_, _08247_, _06252_);
  and _65766_ (_14578_, _14577_, _07104_);
  and _65767_ (_14579_, _14578_, _14576_);
  or _65768_ (_14580_, _14579_, _14534_);
  and _65769_ (_14581_, _14580_, _08580_);
  and _65770_ (_14582_, _07848_, \oc8051_golden_model_1.PSW [7]);
  or _65771_ (_14583_, _14582_, _14536_);
  and _65772_ (_14584_, _14583_, _07103_);
  or _65773_ (_14585_, _14584_, _05791_);
  or _65774_ (_14586_, _14585_, _14581_);
  and _65775_ (_14587_, _05923_, _05791_);
  nor _65776_ (_14588_, _14587_, _08591_);
  and _65777_ (_14589_, _14588_, _14586_);
  and _65778_ (_14590_, _07708_, _08591_);
  or _65779_ (_14591_, _14590_, _08595_);
  or _65780_ (_14592_, _14591_, _14589_);
  or _65781_ (_14593_, _09211_, _08601_);
  and _65782_ (_14594_, _14593_, _08600_);
  and _65783_ (_14595_, _14594_, _14592_);
  and _65784_ (_14596_, _08395_, _07708_);
  and _65785_ (_14597_, _08724_, \oc8051_golden_model_1.TL1 [2]);
  and _65786_ (_14598_, _08710_, \oc8051_golden_model_1.TH1 [2]);
  and _65787_ (_14599_, _08718_, \oc8051_golden_model_1.SCON [2]);
  or _65788_ (_14600_, _14599_, _14598_);
  or _65789_ (_14601_, _14600_, _14597_);
  and _65790_ (_14602_, _08706_, \oc8051_golden_model_1.TH0 [2]);
  and _65791_ (_14603_, _08726_, \oc8051_golden_model_1.TCON [2]);
  or _65792_ (_14604_, _14603_, _14602_);
  or _65793_ (_14605_, _14604_, _14601_);
  and _65794_ (_14606_, _08734_, \oc8051_golden_model_1.PSW [2]);
  and _65795_ (_14607_, _08741_, \oc8051_golden_model_1.B [2]);
  and _65796_ (_14608_, _08738_, \oc8051_golden_model_1.ACC [2]);
  or _65797_ (_14609_, _14608_, _14607_);
  or _65798_ (_14610_, _14609_, _14606_);
  and _65799_ (_14611_, _08746_, \oc8051_golden_model_1.IP [2]);
  and _65800_ (_14612_, _08749_, \oc8051_golden_model_1.IE [2]);
  and _65801_ (_14613_, _08752_, \oc8051_golden_model_1.SBUF [2]);
  or _65802_ (_14614_, _14613_, _14612_);
  or _65803_ (_14615_, _14614_, _14611_);
  or _65804_ (_14616_, _14615_, _14610_);
  and _65805_ (_14617_, _08760_, \oc8051_golden_model_1.DPH [2]);
  and _65806_ (_14618_, _08758_, \oc8051_golden_model_1.SP [2]);
  or _65807_ (_14619_, _14618_, _14617_);
  and _65808_ (_14620_, _08765_, \oc8051_golden_model_1.DPL [2]);
  or _65809_ (_14621_, _14620_, _14619_);
  and _65810_ (_14622_, _08770_, \oc8051_golden_model_1.PCON [2]);
  and _65811_ (_14623_, _08775_, \oc8051_golden_model_1.TMOD [2]);
  and _65812_ (_14624_, _08773_, \oc8051_golden_model_1.TL0 [2]);
  or _65813_ (_14625_, _14624_, _14623_);
  or _65814_ (_14626_, _14625_, _14622_);
  or _65815_ (_14627_, _14626_, _14621_);
  or _65816_ (_14628_, _14627_, _14616_);
  or _65817_ (_14629_, _14628_, _14605_);
  or _65818_ (_14630_, _14629_, _14596_);
  and _65819_ (_14631_, _14630_, _08599_);
  or _65820_ (_14632_, _14631_, _08788_);
  or _65821_ (_14633_, _14632_, _14595_);
  and _65822_ (_14634_, _08788_, _06625_);
  nor _65823_ (_14635_, _14634_, _06112_);
  and _65824_ (_14636_, _14635_, _14633_);
  and _65825_ (_14637_, _08768_, _06112_);
  or _65826_ (_14638_, _14637_, _06076_);
  or _65827_ (_14639_, _14638_, _14636_);
  nor _65828_ (_14640_, _05921_, _05836_);
  nor _65829_ (_14641_, _14640_, _07128_);
  and _65830_ (_14642_, _14641_, _14639_);
  nand _65831_ (_14643_, _08247_, _06521_);
  nor _65832_ (_14644_, _08247_, _06521_);
  not _65833_ (_14645_, _14644_);
  and _65834_ (_14646_, _14645_, _14643_);
  and _65835_ (_14647_, _14646_, _07128_);
  or _65836_ (_14648_, _14647_, _14642_);
  and _65837_ (_14649_, _14648_, _08807_);
  and _65838_ (_14650_, _10282_, _07126_);
  or _65839_ (_14651_, _14650_, _14649_);
  and _65840_ (_14652_, _14651_, _08806_);
  and _65841_ (_14653_, _14644_, _07133_);
  or _65842_ (_14654_, _14653_, _14652_);
  and _65843_ (_14655_, _14654_, _08364_);
  and _65844_ (_14656_, _10274_, _07131_);
  or _65845_ (_14657_, _14656_, _07124_);
  or _65846_ (_14658_, _14657_, _14655_);
  nor _65847_ (_14659_, _05921_, _05848_);
  nor _65848_ (_14660_, _14659_, _08820_);
  and _65849_ (_14661_, _14660_, _14658_);
  and _65850_ (_14662_, _14643_, _08820_);
  or _65851_ (_14663_, _14662_, _08825_);
  or _65852_ (_14664_, _14663_, _14661_);
  nand _65853_ (_14665_, _10281_, _08825_);
  and _65854_ (_14666_, _14665_, _05846_);
  and _65855_ (_14667_, _14666_, _14664_);
  or _65856_ (_14668_, _14667_, _14531_);
  and _65857_ (_14669_, _14668_, _08361_);
  nor _65858_ (_14670_, _14546_, _08361_);
  or _65859_ (_14671_, _14670_, _07325_);
  nor _65860_ (_14672_, _14671_, _14669_);
  and _65861_ (_14673_, _14546_, _07325_);
  or _65862_ (_14674_, _14673_, _14487_);
  nor _65863_ (_14675_, _14674_, _14672_);
  nor _65864_ (_14676_, _09161_, _09070_);
  nor _65865_ (_14677_, _14676_, _09162_);
  nand _65866_ (_14678_, _14677_, _06276_);
  and _65867_ (_14679_, _14678_, _07153_);
  or _65868_ (_14680_, _14679_, _14675_);
  nand _65869_ (_14681_, _14677_, _14495_);
  and _65870_ (_14682_, _14681_, _08837_);
  and _65871_ (_14683_, _14682_, _14680_);
  and _65872_ (_14684_, _14542_, _07152_);
  or _65873_ (_14685_, _14684_, _06310_);
  or _65874_ (_14686_, _14685_, _14683_);
  nand _65875_ (_14687_, _12029_, _06310_);
  and _65876_ (_14688_, _14687_, _12730_);
  and _65877_ (_14689_, _14688_, _14686_);
  and _65878_ (_14690_, _05921_, _05823_);
  or _65879_ (_14691_, _06073_, _14690_);
  or _65880_ (_14692_, _14691_, _14689_);
  or _65881_ (_14693_, _14536_, _06074_);
  and _65882_ (_14694_, _14693_, _09193_);
  and _65883_ (_14695_, _14694_, _14692_);
  nor _65884_ (_14696_, _09195_, _07708_);
  nor _65885_ (_14697_, _14696_, _09196_);
  and _65886_ (_14698_, _14697_, _09189_);
  or _65887_ (_14699_, _14698_, _14336_);
  or _65888_ (_14700_, _14699_, _14695_);
  nor _65889_ (_14701_, _09212_, _09211_);
  nor _65890_ (_14702_, _14701_, _09213_);
  or _65891_ (_14703_, _14702_, _14339_);
  and _65892_ (_14704_, _14703_, _14700_);
  and _65893_ (_14705_, _14704_, _06835_);
  and _65894_ (_14706_, _14702_, _06834_);
  or _65895_ (_14707_, _14706_, _07167_);
  or _65896_ (_14708_, _14707_, _14705_);
  nor _65897_ (_14709_, _08248_, _08212_);
  nor _65898_ (_14710_, _14709_, _08249_);
  or _65899_ (_14711_, _14710_, _14518_);
  and _65900_ (_14712_, _14711_, _07417_);
  and _65901_ (_14713_, _14712_, _14708_);
  or _65902_ (_14714_, _14713_, _14164_);
  and _65903_ (_14715_, _14714_, _14530_);
  nand _65904_ (_14716_, _11989_, _06310_);
  or _65905_ (_14717_, _12159_, _06310_);
  and _65906_ (_14718_, _14717_, _14716_);
  and _65907_ (_14719_, _14718_, _07764_);
  and _65908_ (_14720_, _14719_, _14328_);
  or _65909_ (_41016_, _14720_, _14715_);
  or _65910_ (_14721_, _14156_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _65911_ (_14722_, _14721_, _14162_);
  nor _65912_ (_14723_, _06322_, _05846_);
  nand _65913_ (_14724_, _08139_, _06389_);
  nor _65914_ (_14725_, _08139_, _06389_);
  not _65915_ (_14726_, _14725_);
  and _65916_ (_14727_, _14726_, _14724_);
  and _65917_ (_14728_, _14727_, _07128_);
  and _65918_ (_14729_, _07851_, \oc8051_golden_model_1.PSW [7]);
  not _65919_ (_14730_, _07851_);
  and _65920_ (_14731_, _12595_, _14730_);
  or _65921_ (_14732_, _14731_, _14729_);
  and _65922_ (_14733_, _14732_, _07103_);
  or _65923_ (_14734_, _14731_, _08398_);
  or _65924_ (_14735_, _12595_, _07851_);
  or _65925_ (_14736_, _14735_, _08428_);
  and _65926_ (_14737_, _14540_, _08140_);
  or _65927_ (_14738_, _14737_, _08543_);
  and _65928_ (_14739_, _14738_, _06162_);
  nor _65929_ (_14740_, _14544_, _07474_);
  nor _65930_ (_14741_, _14740_, _08353_);
  nand _65931_ (_14742_, _14741_, _08445_);
  and _65932_ (_14743_, _06581_, _05974_);
  nor _65933_ (_14744_, _06581_, _10028_);
  nor _65934_ (_14745_, _14744_, _14743_);
  and _65935_ (_14746_, _14745_, _08443_);
  nor _65936_ (_14747_, _14746_, _06162_);
  and _65937_ (_14748_, _14747_, _14742_);
  or _65938_ (_14749_, _14748_, _06159_);
  or _65939_ (_14750_, _14749_, _14739_);
  and _65940_ (_14751_, _14750_, _14736_);
  or _65941_ (_14752_, _14751_, _07485_);
  nor _65942_ (_14753_, _05974_, _05764_);
  nor _65943_ (_14754_, _14753_, _07076_);
  and _65944_ (_14755_, _14754_, _14752_);
  and _65945_ (_14756_, _07544_, _07076_);
  or _65946_ (_14757_, _14756_, _07086_);
  or _65947_ (_14758_, _14757_, _14755_);
  and _65948_ (_14759_, _14758_, _14734_);
  or _65949_ (_14760_, _14759_, _06151_);
  nand _65950_ (_14761_, _08139_, _06151_);
  and _65951_ (_14762_, _14761_, _06149_);
  and _65952_ (_14763_, _14762_, _14760_);
  not _65953_ (_14764_, _12596_);
  and _65954_ (_14765_, _14735_, _14764_);
  and _65955_ (_14766_, _14765_, _06148_);
  or _65956_ (_14767_, _14766_, _14763_);
  and _65957_ (_14768_, _14767_, _05760_);
  or _65958_ (_14769_, _06322_, _05760_);
  nand _65959_ (_14770_, _06251_, _14769_);
  or _65960_ (_14771_, _14770_, _14768_);
  nand _65961_ (_14772_, _08139_, _06252_);
  and _65962_ (_14773_, _14772_, _14771_);
  or _65963_ (_14774_, _14773_, _06701_);
  and _65964_ (_14775_, _09210_, _06172_);
  or _65965_ (_14776_, _08137_, _07104_);
  or _65966_ (_14777_, _14776_, _14775_);
  and _65967_ (_14778_, _14777_, _08580_);
  and _65968_ (_14779_, _14778_, _14774_);
  or _65969_ (_14780_, _14779_, _14733_);
  or _65970_ (_14781_, _14780_, _05791_);
  and _65971_ (_14782_, _06322_, _05791_);
  nor _65972_ (_14783_, _14782_, _08591_);
  and _65973_ (_14784_, _14783_, _14781_);
  and _65974_ (_14785_, _07544_, _08591_);
  or _65975_ (_14786_, _14785_, _08595_);
  or _65976_ (_14787_, _14786_, _14784_);
  or _65977_ (_14788_, _09210_, _08601_);
  and _65978_ (_14789_, _14788_, _08600_);
  and _65979_ (_14790_, _14789_, _14787_);
  and _65980_ (_14791_, _08395_, _07544_);
  and _65981_ (_14792_, _08724_, \oc8051_golden_model_1.TL1 [3]);
  and _65982_ (_14793_, _08710_, \oc8051_golden_model_1.TH1 [3]);
  and _65983_ (_14794_, _08718_, \oc8051_golden_model_1.SCON [3]);
  or _65984_ (_14795_, _14794_, _14793_);
  or _65985_ (_14796_, _14795_, _14792_);
  and _65986_ (_14797_, _08770_, \oc8051_golden_model_1.PCON [3]);
  and _65987_ (_14798_, _08706_, \oc8051_golden_model_1.TH0 [3]);
  or _65988_ (_14799_, _14798_, _14797_);
  or _65989_ (_14800_, _14799_, _14796_);
  and _65990_ (_14801_, _08734_, \oc8051_golden_model_1.PSW [3]);
  and _65991_ (_14802_, _08741_, \oc8051_golden_model_1.B [3]);
  and _65992_ (_14803_, _08738_, \oc8051_golden_model_1.ACC [3]);
  or _65993_ (_14804_, _14803_, _14802_);
  or _65994_ (_14805_, _14804_, _14801_);
  and _65995_ (_14806_, _08746_, \oc8051_golden_model_1.IP [3]);
  and _65996_ (_14807_, _08749_, \oc8051_golden_model_1.IE [3]);
  and _65997_ (_14808_, _08752_, \oc8051_golden_model_1.SBUF [3]);
  or _65998_ (_14809_, _14808_, _14807_);
  or _65999_ (_14810_, _14809_, _14806_);
  or _66000_ (_14811_, _14810_, _14805_);
  and _66001_ (_14812_, _08765_, \oc8051_golden_model_1.DPL [3]);
  and _66002_ (_14813_, _08758_, \oc8051_golden_model_1.SP [3]);
  and _66003_ (_14814_, _08760_, \oc8051_golden_model_1.DPH [3]);
  or _66004_ (_14815_, _14814_, _14813_);
  or _66005_ (_14816_, _14815_, _14812_);
  and _66006_ (_14817_, _08775_, \oc8051_golden_model_1.TMOD [3]);
  and _66007_ (_14818_, _08773_, \oc8051_golden_model_1.TL0 [3]);
  or _66008_ (_14819_, _14818_, _14817_);
  and _66009_ (_14820_, _08726_, \oc8051_golden_model_1.TCON [3]);
  or _66010_ (_14821_, _14820_, _14819_);
  or _66011_ (_14822_, _14821_, _14816_);
  or _66012_ (_14823_, _14822_, _14811_);
  or _66013_ (_14824_, _14823_, _14800_);
  or _66014_ (_14825_, _14824_, _14791_);
  and _66015_ (_14826_, _14825_, _08599_);
  or _66016_ (_14827_, _14826_, _08788_);
  or _66017_ (_14828_, _14827_, _14790_);
  and _66018_ (_14829_, _08788_, _06070_);
  nor _66019_ (_14830_, _14829_, _06112_);
  and _66020_ (_14831_, _14830_, _14828_);
  and _66021_ (_14832_, _08712_, _06112_);
  or _66022_ (_14833_, _14832_, _06076_);
  or _66023_ (_14834_, _14833_, _14831_);
  nor _66024_ (_14835_, _05974_, _05836_);
  nor _66025_ (_14836_, _14835_, _07128_);
  and _66026_ (_14837_, _14836_, _14834_);
  or _66027_ (_14838_, _14837_, _14728_);
  and _66028_ (_14839_, _14838_, _08807_);
  and _66029_ (_14840_, _12318_, _07126_);
  or _66030_ (_14841_, _14840_, _07133_);
  or _66031_ (_14842_, _14841_, _14839_);
  or _66032_ (_14843_, _14725_, _08806_);
  and _66033_ (_14844_, _14843_, _08364_);
  and _66034_ (_14845_, _14844_, _14842_);
  and _66035_ (_14846_, _10272_, _07131_);
  or _66036_ (_14847_, _14846_, _07124_);
  or _66037_ (_14848_, _14847_, _14845_);
  nor _66038_ (_14849_, _05974_, _05848_);
  nor _66039_ (_14850_, _14849_, _08820_);
  and _66040_ (_14851_, _14850_, _14848_);
  and _66041_ (_14852_, _14724_, _08820_);
  or _66042_ (_14853_, _14852_, _08825_);
  or _66043_ (_14854_, _14853_, _14851_);
  nand _66044_ (_14855_, _10273_, _08825_);
  and _66045_ (_14856_, _14855_, _05846_);
  and _66046_ (_14857_, _14856_, _14854_);
  or _66047_ (_14858_, _14857_, _14723_);
  and _66048_ (_14859_, _14858_, _08361_);
  nor _66049_ (_14860_, _14741_, _08361_);
  or _66050_ (_14861_, _14860_, _07325_);
  nor _66051_ (_14862_, _14861_, _14859_);
  and _66052_ (_14863_, _14741_, _07325_);
  or _66053_ (_14864_, _14863_, _14487_);
  nor _66054_ (_14865_, _14864_, _14862_);
  nor _66055_ (_14866_, _09162_, _09025_);
  nor _66056_ (_14867_, _14866_, _09163_);
  nand _66057_ (_14868_, _14867_, _06276_);
  and _66058_ (_14869_, _14868_, _07153_);
  or _66059_ (_14870_, _14869_, _14865_);
  nand _66060_ (_14871_, _14867_, _14495_);
  and _66061_ (_14872_, _14871_, _08837_);
  and _66062_ (_14873_, _14872_, _14870_);
  and _66063_ (_14874_, _14738_, _07152_);
  or _66064_ (_14875_, _14874_, _06310_);
  or _66065_ (_14876_, _14875_, _14873_);
  nand _66066_ (_14877_, _12024_, _06310_);
  and _66067_ (_14878_, _14877_, _12730_);
  and _66068_ (_14879_, _14878_, _14876_);
  and _66069_ (_14880_, _05974_, _05823_);
  or _66070_ (_14881_, _06073_, _14880_);
  or _66071_ (_14882_, _14881_, _14879_);
  or _66072_ (_14883_, _14731_, _06074_);
  and _66073_ (_14884_, _14883_, _09193_);
  and _66074_ (_14885_, _14884_, _14882_);
  nor _66075_ (_14886_, _09196_, _07544_);
  nor _66076_ (_14887_, _14886_, _09197_);
  or _66077_ (_14888_, _14887_, _07168_);
  and _66078_ (_14889_, _14888_, _12737_);
  or _66079_ (_14890_, _14889_, _14885_);
  nor _66080_ (_14891_, _09213_, _09210_);
  nor _66081_ (_14892_, _14891_, _09214_);
  or _66082_ (_14893_, _14892_, _07169_);
  and _66083_ (_14894_, _14893_, _14890_);
  or _66084_ (_14895_, _14894_, _07167_);
  nor _66085_ (_14896_, _08249_, _08140_);
  nor _66086_ (_14897_, _14896_, _08250_);
  or _66087_ (_14898_, _14897_, _14518_);
  and _66088_ (_14899_, _14898_, _07417_);
  and _66089_ (_14900_, _14899_, _14895_);
  or _66090_ (_14901_, _14900_, _14164_);
  and _66091_ (_14902_, _14901_, _14722_);
  nand _66092_ (_14903_, _11982_, _06310_);
  or _66093_ (_14904_, _12163_, _06310_);
  and _66094_ (_14905_, _14904_, _14903_);
  and _66095_ (_14906_, _14905_, _07764_);
  and _66096_ (_14907_, _14906_, _14328_);
  or _66097_ (_41017_, _14907_, _14902_);
  nor _66098_ (_14908_, _14156_, _08284_);
  nor _66099_ (_14909_, _09214_, _09209_);
  nor _66100_ (_14910_, _14909_, _09215_);
  or _66101_ (_14911_, _14910_, _07169_);
  nor _66102_ (_14912_, _12194_, _05846_);
  and _66103_ (_14913_, _08353_, _08349_);
  nor _66104_ (_14914_, _08353_, _08349_);
  nor _66105_ (_14915_, _14914_, _14913_);
  nand _66106_ (_14916_, _14915_, _08445_);
  nor _66107_ (_14917_, _06581_, _09902_);
  and _66108_ (_14918_, _12193_, _06581_);
  nor _66109_ (_14919_, _14918_, _14917_);
  nand _66110_ (_14920_, _14919_, _08443_);
  and _66111_ (_14921_, _14920_, _14916_);
  or _66112_ (_14922_, _14921_, _07064_);
  or _66113_ (_14923_, _09209_, _07065_);
  and _66114_ (_14924_, _14923_, _14922_);
  and _66115_ (_14925_, _14924_, _08429_);
  nand _66116_ (_14926_, _08543_, _08338_);
  or _66117_ (_14927_, _08543_, _08338_);
  nand _66118_ (_14928_, _14927_, _14926_);
  and _66119_ (_14929_, _14928_, _06162_);
  or _66120_ (_14930_, _14929_, _14925_);
  and _66121_ (_14931_, _14930_, _08428_);
  nand _66122_ (_14932_, _12678_, _12676_);
  and _66123_ (_14933_, _14932_, _06159_);
  or _66124_ (_14934_, _14933_, _07485_);
  or _66125_ (_14935_, _14934_, _14931_);
  nor _66126_ (_14936_, _12193_, _05764_);
  nor _66127_ (_14937_, _14936_, _07076_);
  and _66128_ (_14938_, _14937_, _14935_);
  and _66129_ (_14939_, _08336_, _07076_);
  or _66130_ (_14940_, _14939_, _07086_);
  or _66131_ (_14941_, _14940_, _14938_);
  nor _66132_ (_14942_, _12677_, _12676_);
  or _66133_ (_14943_, _14942_, _08398_);
  and _66134_ (_14944_, _14943_, _14941_);
  or _66135_ (_14945_, _14944_, _06151_);
  nand _66136_ (_14946_, _08338_, _06151_);
  and _66137_ (_14947_, _14946_, _06149_);
  and _66138_ (_14948_, _14947_, _14945_);
  not _66139_ (_14949_, _12679_);
  and _66140_ (_14950_, _14932_, _14949_);
  and _66141_ (_14951_, _14950_, _06148_);
  or _66142_ (_14952_, _14951_, _14948_);
  and _66143_ (_14953_, _14952_, _05760_);
  or _66144_ (_14954_, _12194_, _05760_);
  nand _66145_ (_14955_, _14954_, _06251_);
  or _66146_ (_14956_, _14955_, _14953_);
  nand _66147_ (_14957_, _08338_, _06252_);
  and _66148_ (_14958_, _14957_, _14956_);
  or _66149_ (_14959_, _14958_, _06701_);
  and _66150_ (_14960_, _09209_, _06172_);
  or _66151_ (_14961_, _08283_, _07104_);
  or _66152_ (_14962_, _14961_, _14960_);
  and _66153_ (_14963_, _14962_, _08580_);
  and _66154_ (_14964_, _14963_, _14959_);
  and _66155_ (_14965_, _12677_, \oc8051_golden_model_1.PSW [7]);
  or _66156_ (_14966_, _14965_, _14942_);
  and _66157_ (_14967_, _14966_, _07103_);
  or _66158_ (_14968_, _14967_, _05791_);
  or _66159_ (_14969_, _14968_, _14964_);
  and _66160_ (_14970_, _12194_, _05791_);
  nor _66161_ (_14971_, _14970_, _08591_);
  and _66162_ (_14972_, _14971_, _14969_);
  and _66163_ (_14973_, _08336_, _08591_);
  or _66164_ (_14974_, _14973_, _08595_);
  or _66165_ (_14975_, _14974_, _14972_);
  or _66166_ (_14976_, _09209_, _08601_);
  and _66167_ (_14977_, _14976_, _08600_);
  and _66168_ (_14978_, _14977_, _14975_);
  and _66169_ (_14979_, _08395_, _08336_);
  and _66170_ (_14980_, _08710_, \oc8051_golden_model_1.TH1 [4]);
  and _66171_ (_14981_, _08775_, \oc8051_golden_model_1.TMOD [4]);
  and _66172_ (_14982_, _08706_, \oc8051_golden_model_1.TH0 [4]);
  or _66173_ (_14983_, _14982_, _14981_);
  or _66174_ (_14984_, _14983_, _14980_);
  and _66175_ (_14985_, _08760_, \oc8051_golden_model_1.DPH [4]);
  and _66176_ (_14986_, _08724_, \oc8051_golden_model_1.TL1 [4]);
  and _66177_ (_14987_, _08758_, \oc8051_golden_model_1.SP [4]);
  or _66178_ (_14988_, _14987_, _14986_);
  or _66179_ (_14989_, _14988_, _14985_);
  and _66180_ (_14990_, _08752_, \oc8051_golden_model_1.SBUF [4]);
  and _66181_ (_14991_, _08746_, \oc8051_golden_model_1.IP [4]);
  or _66182_ (_14992_, _14991_, _14990_);
  and _66183_ (_14993_, _08718_, \oc8051_golden_model_1.SCON [4]);
  and _66184_ (_14994_, _08741_, \oc8051_golden_model_1.B [4]);
  or _66185_ (_14995_, _14994_, _14993_);
  or _66186_ (_14996_, _14995_, _14992_);
  and _66187_ (_14997_, _08765_, \oc8051_golden_model_1.DPL [4]);
  and _66188_ (_14998_, _08770_, \oc8051_golden_model_1.PCON [4]);
  or _66189_ (_14999_, _14998_, _14997_);
  or _66190_ (_15000_, _14999_, _14996_);
  and _66191_ (_15001_, _08773_, \oc8051_golden_model_1.TL0 [4]);
  and _66192_ (_15002_, _08726_, \oc8051_golden_model_1.TCON [4]);
  and _66193_ (_15003_, _08749_, \oc8051_golden_model_1.IE [4]);
  or _66194_ (_15004_, _15003_, _15002_);
  and _66195_ (_15005_, _08738_, \oc8051_golden_model_1.ACC [4]);
  and _66196_ (_15006_, _08734_, \oc8051_golden_model_1.PSW [4]);
  or _66197_ (_15007_, _15006_, _15005_);
  or _66198_ (_15008_, _15007_, _15004_);
  or _66199_ (_15009_, _15008_, _15001_);
  or _66200_ (_15010_, _15009_, _15000_);
  or _66201_ (_15011_, _15010_, _14989_);
  or _66202_ (_15012_, _15011_, _14984_);
  or _66203_ (_15013_, _15012_, _14979_);
  and _66204_ (_15014_, _15013_, _08599_);
  or _66205_ (_15015_, _15014_, _08788_);
  or _66206_ (_15016_, _15015_, _14978_);
  and _66207_ (_15017_, _08788_, _06876_);
  nor _66208_ (_15018_, _15017_, _06112_);
  and _66209_ (_15019_, _15018_, _15016_);
  and _66210_ (_15020_, _08715_, _06112_);
  or _66211_ (_15021_, _15020_, _06076_);
  or _66212_ (_15022_, _15021_, _15019_);
  nor _66213_ (_15023_, _12193_, _05836_);
  nor _66214_ (_15024_, _15023_, _07128_);
  and _66215_ (_15025_, _15024_, _15022_);
  nand _66216_ (_15026_, _08670_, _08338_);
  nor _66217_ (_15027_, _08670_, _08338_);
  not _66218_ (_15028_, _15027_);
  and _66219_ (_15029_, _15028_, _15026_);
  and _66220_ (_15030_, _15029_, _07128_);
  or _66221_ (_15031_, _15030_, _15025_);
  and _66222_ (_15032_, _15031_, _08807_);
  and _66223_ (_15033_, _10289_, _07126_);
  or _66224_ (_15034_, _15033_, _07133_);
  or _66225_ (_15035_, _15034_, _15032_);
  or _66226_ (_15036_, _15027_, _08806_);
  and _66227_ (_15037_, _15036_, _08364_);
  and _66228_ (_15038_, _15037_, _15035_);
  and _66229_ (_15039_, _10270_, _07131_);
  or _66230_ (_15040_, _15039_, _07124_);
  or _66231_ (_15041_, _15040_, _15038_);
  nor _66232_ (_15042_, _12193_, _05848_);
  nor _66233_ (_15043_, _15042_, _08820_);
  and _66234_ (_15044_, _15043_, _15041_);
  and _66235_ (_15045_, _15026_, _08820_);
  or _66236_ (_15046_, _15045_, _08825_);
  or _66237_ (_15047_, _15046_, _15044_);
  nand _66238_ (_15048_, _10288_, _08825_);
  and _66239_ (_15049_, _15048_, _05846_);
  and _66240_ (_15050_, _15049_, _15047_);
  or _66241_ (_15051_, _15050_, _14912_);
  and _66242_ (_15052_, _15051_, _08361_);
  nor _66243_ (_15053_, _14915_, _08361_);
  or _66244_ (_15054_, _15053_, _07325_);
  nor _66245_ (_15055_, _15054_, _15052_);
  and _66246_ (_15056_, _14915_, _07325_);
  or _66247_ (_15057_, _15056_, _14487_);
  nor _66248_ (_15058_, _15057_, _15055_);
  nor _66249_ (_15059_, _09163_, _08980_);
  nor _66250_ (_15060_, _15059_, _09164_);
  nand _66251_ (_15061_, _15060_, _06276_);
  and _66252_ (_15062_, _15061_, _07153_);
  or _66253_ (_15063_, _15062_, _15058_);
  nand _66254_ (_15064_, _15060_, _14495_);
  and _66255_ (_15065_, _15064_, _08837_);
  and _66256_ (_15066_, _15065_, _15063_);
  and _66257_ (_15067_, _14928_, _07152_);
  or _66258_ (_15068_, _15067_, _06310_);
  or _66259_ (_15069_, _15068_, _15066_);
  nand _66260_ (_15070_, _12019_, _06310_);
  and _66261_ (_15071_, _15070_, _12730_);
  and _66262_ (_15072_, _15071_, _15069_);
  and _66263_ (_15073_, _12193_, _05823_);
  or _66264_ (_15074_, _15073_, _06073_);
  or _66265_ (_15075_, _15074_, _15072_);
  or _66266_ (_15076_, _14942_, _06074_);
  and _66267_ (_15077_, _15076_, _09193_);
  and _66268_ (_15078_, _15077_, _15075_);
  nor _66269_ (_15079_, _09197_, _08336_);
  nor _66270_ (_15080_, _15079_, _09198_);
  and _66271_ (_15081_, _15080_, _09189_);
  or _66272_ (_15082_, _15081_, _07168_);
  or _66273_ (_15083_, _15082_, _15078_);
  and _66274_ (_15084_, _15083_, _14911_);
  or _66275_ (_15085_, _15084_, _07167_);
  nor _66276_ (_15086_, _08339_, _08250_);
  nor _66277_ (_15087_, _15086_, _08340_);
  or _66278_ (_15088_, _15087_, _14518_);
  and _66279_ (_15089_, _15088_, _07417_);
  and _66280_ (_15090_, _15089_, _15085_);
  and _66281_ (_15091_, _15090_, _14156_);
  or _66282_ (_15092_, _15091_, _14908_);
  and _66283_ (_15093_, _15092_, _14162_);
  nand _66284_ (_15094_, _11978_, _06310_);
  or _66285_ (_15095_, _12156_, _06310_);
  and _66286_ (_15096_, _15095_, _15094_);
  and _66287_ (_15097_, _15096_, _07764_);
  and _66288_ (_15098_, _15097_, _14328_);
  or _66289_ (_41018_, _15098_, _15093_);
  nor _66290_ (_15099_, _14156_, _08049_);
  nor _66291_ (_15100_, _09164_, _08931_);
  or _66292_ (_15101_, _15100_, _09165_);
  and _66293_ (_15102_, _15101_, _14495_);
  not _66294_ (_15103_, _12612_);
  and _66295_ (_15104_, _15103_, _12611_);
  or _66296_ (_15105_, _15104_, _08398_);
  nor _66297_ (_15106_, _06581_, _09930_);
  and _66298_ (_15107_, _12188_, _06581_);
  or _66299_ (_15108_, _15107_, _15106_);
  and _66300_ (_15109_, _15108_, _08443_);
  nor _66301_ (_15110_, _14913_, _08348_);
  or _66302_ (_15111_, _15110_, _08354_);
  and _66303_ (_15112_, _15111_, _08445_);
  or _66304_ (_15113_, _15112_, _15109_);
  and _66305_ (_15114_, _15113_, _07065_);
  and _66306_ (_15115_, _09208_, _07064_);
  or _66307_ (_15116_, _15115_, _15114_);
  and _66308_ (_15117_, _15116_, _08429_);
  and _66309_ (_15118_, _14926_, _08104_);
  or _66310_ (_15119_, _15118_, _08544_);
  and _66311_ (_15120_, _15119_, _06162_);
  or _66312_ (_15121_, _15120_, _15117_);
  and _66313_ (_15122_, _15121_, _08428_);
  or _66314_ (_15123_, _12612_, _12611_);
  and _66315_ (_15124_, _15123_, _06159_);
  or _66316_ (_15125_, _15124_, _07485_);
  or _66317_ (_15126_, _15125_, _15122_);
  nor _66318_ (_15127_, _12188_, _05764_);
  nor _66319_ (_15128_, _15127_, _07076_);
  and _66320_ (_15129_, _15128_, _15126_);
  and _66321_ (_15130_, _08101_, _07076_);
  or _66322_ (_15131_, _15130_, _07086_);
  or _66323_ (_15132_, _15131_, _15129_);
  and _66324_ (_15133_, _15132_, _15105_);
  or _66325_ (_15134_, _15133_, _06151_);
  nand _66326_ (_15135_, _08103_, _06151_);
  and _66327_ (_15136_, _15135_, _06149_);
  and _66328_ (_15137_, _15136_, _15134_);
  not _66329_ (_15138_, _12613_);
  and _66330_ (_15139_, _15123_, _15138_);
  and _66331_ (_15140_, _15139_, _06148_);
  or _66332_ (_15141_, _15140_, _15137_);
  and _66333_ (_15142_, _15141_, _05760_);
  or _66334_ (_15143_, _12189_, _05760_);
  nand _66335_ (_15144_, _15143_, _06251_);
  or _66336_ (_15145_, _15144_, _15142_);
  nand _66337_ (_15146_, _08103_, _06252_);
  and _66338_ (_15147_, _15146_, _15145_);
  or _66339_ (_15148_, _15147_, _06701_);
  and _66340_ (_15149_, _09208_, _06172_);
  or _66341_ (_15150_, _08048_, _07104_);
  or _66342_ (_15151_, _15150_, _15149_);
  and _66343_ (_15152_, _15151_, _08580_);
  and _66344_ (_15153_, _15152_, _15148_);
  and _66345_ (_15154_, _12612_, \oc8051_golden_model_1.PSW [7]);
  or _66346_ (_15155_, _15154_, _15104_);
  and _66347_ (_15156_, _15155_, _07103_);
  or _66348_ (_15157_, _15156_, _05791_);
  or _66349_ (_15158_, _15157_, _15153_);
  and _66350_ (_15159_, _12189_, _05791_);
  nor _66351_ (_15160_, _15159_, _08591_);
  and _66352_ (_15161_, _15160_, _15158_);
  and _66353_ (_15162_, _08101_, _08591_);
  or _66354_ (_15163_, _15162_, _08595_);
  or _66355_ (_15164_, _15163_, _15161_);
  or _66356_ (_15165_, _09208_, _08601_);
  and _66357_ (_15166_, _15165_, _08600_);
  and _66358_ (_15167_, _15166_, _15164_);
  and _66359_ (_15168_, _08395_, _08101_);
  and _66360_ (_15169_, _08775_, \oc8051_golden_model_1.TMOD [5]);
  and _66361_ (_15170_, _08706_, \oc8051_golden_model_1.TH0 [5]);
  and _66362_ (_15171_, _08710_, \oc8051_golden_model_1.TH1 [5]);
  or _66363_ (_15172_, _15171_, _15170_);
  or _66364_ (_15173_, _15172_, _15169_);
  and _66365_ (_15174_, _08770_, \oc8051_golden_model_1.PCON [5]);
  and _66366_ (_15175_, _08724_, \oc8051_golden_model_1.TL1 [5]);
  and _66367_ (_15176_, _08758_, \oc8051_golden_model_1.SP [5]);
  or _66368_ (_15177_, _15176_, _15175_);
  or _66369_ (_15178_, _15177_, _15174_);
  and _66370_ (_15179_, _08741_, \oc8051_golden_model_1.B [5]);
  and _66371_ (_15180_, _08738_, \oc8051_golden_model_1.ACC [5]);
  or _66372_ (_15181_, _15180_, _15179_);
  and _66373_ (_15182_, _08718_, \oc8051_golden_model_1.SCON [5]);
  and _66374_ (_15183_, _08734_, \oc8051_golden_model_1.PSW [5]);
  or _66375_ (_15184_, _15183_, _15182_);
  or _66376_ (_15185_, _15184_, _15181_);
  and _66377_ (_15186_, _08765_, \oc8051_golden_model_1.DPL [5]);
  and _66378_ (_15187_, _08760_, \oc8051_golden_model_1.DPH [5]);
  or _66379_ (_15188_, _15187_, _15186_);
  or _66380_ (_15189_, _15188_, _15185_);
  and _66381_ (_15190_, _08773_, \oc8051_golden_model_1.TL0 [5]);
  and _66382_ (_15191_, _08752_, \oc8051_golden_model_1.SBUF [5]);
  and _66383_ (_15192_, _08749_, \oc8051_golden_model_1.IE [5]);
  or _66384_ (_15193_, _15192_, _15191_);
  and _66385_ (_15194_, _08726_, \oc8051_golden_model_1.TCON [5]);
  and _66386_ (_15196_, _08746_, \oc8051_golden_model_1.IP [5]);
  or _66387_ (_15197_, _15196_, _15194_);
  or _66388_ (_15198_, _15197_, _15193_);
  or _66389_ (_15199_, _15198_, _15190_);
  or _66390_ (_15200_, _15199_, _15189_);
  or _66391_ (_15201_, _15200_, _15178_);
  or _66392_ (_15202_, _15201_, _15173_);
  or _66393_ (_15203_, _15202_, _15168_);
  and _66394_ (_15204_, _15203_, _08599_);
  or _66395_ (_15205_, _15204_, _08788_);
  or _66396_ (_15206_, _15205_, _15167_);
  and _66397_ (_15207_, _08788_, _06477_);
  nor _66398_ (_15208_, _15207_, _06112_);
  and _66399_ (_15209_, _15208_, _15206_);
  and _66400_ (_15210_, _08736_, _06112_);
  or _66401_ (_15211_, _15210_, _06076_);
  or _66402_ (_15212_, _15211_, _15209_);
  nor _66403_ (_15213_, _12188_, _05836_);
  nor _66404_ (_15214_, _15213_, _07128_);
  and _66405_ (_15215_, _15214_, _15212_);
  nand _66406_ (_15216_, _08701_, _08103_);
  nor _66407_ (_15217_, _08701_, _08103_);
  not _66408_ (_15218_, _15217_);
  and _66409_ (_15219_, _15218_, _15216_);
  and _66410_ (_15220_, _15219_, _07128_);
  or _66411_ (_15221_, _15220_, _15215_);
  and _66412_ (_15222_, _15221_, _08807_);
  and _66413_ (_15223_, _12325_, _07126_);
  or _66414_ (_15224_, _15223_, _07133_);
  or _66415_ (_15225_, _15224_, _15222_);
  or _66416_ (_15226_, _15217_, _08806_);
  and _66417_ (_15227_, _15226_, _08364_);
  and _66418_ (_15228_, _15227_, _15225_);
  and _66419_ (_15229_, _10268_, _07131_);
  or _66420_ (_15230_, _15229_, _07124_);
  or _66421_ (_15231_, _15230_, _15228_);
  nor _66422_ (_15232_, _12188_, _05848_);
  nor _66423_ (_15233_, _15232_, _08820_);
  and _66424_ (_15234_, _15233_, _15231_);
  and _66425_ (_15235_, _15216_, _08820_);
  or _66426_ (_15236_, _15235_, _08825_);
  or _66427_ (_15237_, _15236_, _15234_);
  nand _66428_ (_15238_, _10269_, _08825_);
  and _66429_ (_15239_, _15238_, _05846_);
  and _66430_ (_15240_, _15239_, _15237_);
  or _66431_ (_15241_, _12189_, _05846_);
  nand _66432_ (_15242_, _15241_, _08362_);
  or _66433_ (_15243_, _15242_, _15240_);
  or _66434_ (_15244_, _15111_, _08362_);
  and _66435_ (_15245_, _15244_, _14488_);
  and _66436_ (_15246_, _15245_, _15243_);
  and _66437_ (_15247_, _15101_, _14487_);
  nor _66438_ (_15248_, _15247_, _15246_);
  nor _66439_ (_15249_, _15248_, _14495_);
  or _66440_ (_15250_, _15249_, _15102_);
  and _66441_ (_15251_, _15250_, _08837_);
  and _66442_ (_15252_, _15119_, _07152_);
  or _66443_ (_15253_, _15252_, _06310_);
  or _66444_ (_15254_, _15253_, _15251_);
  nand _66445_ (_15255_, _12014_, _06310_);
  and _66446_ (_15256_, _15255_, _12730_);
  and _66447_ (_15257_, _15256_, _15254_);
  and _66448_ (_15258_, _12188_, _05823_);
  or _66449_ (_15259_, _15258_, _06073_);
  or _66450_ (_15260_, _15259_, _15257_);
  or _66451_ (_15261_, _15104_, _06074_);
  and _66452_ (_15262_, _15261_, _09193_);
  and _66453_ (_15263_, _15262_, _15260_);
  nor _66454_ (_15264_, _09198_, _08101_);
  nor _66455_ (_15265_, _15264_, _09199_);
  or _66456_ (_15266_, _15265_, _07168_);
  and _66457_ (_15267_, _15266_, _12737_);
  or _66458_ (_15268_, _15267_, _15263_);
  nor _66459_ (_15269_, _09215_, _09208_);
  nor _66460_ (_15270_, _15269_, _09216_);
  or _66461_ (_15271_, _15270_, _07169_);
  and _66462_ (_15272_, _15271_, _15268_);
  or _66463_ (_15273_, _15272_, _07167_);
  nor _66464_ (_15274_, _08340_, _08104_);
  nor _66465_ (_15275_, _15274_, _08341_);
  or _66466_ (_15276_, _15275_, _14518_);
  and _66467_ (_15277_, _15276_, _07417_);
  and _66468_ (_15278_, _15277_, _15273_);
  and _66469_ (_15279_, _15278_, _14156_);
  or _66470_ (_15280_, _15279_, _15099_);
  and _66471_ (_15281_, _15280_, _14162_);
  nand _66472_ (_15282_, _11973_, _06310_);
  or _66473_ (_15283_, _12152_, _06310_);
  and _66474_ (_15284_, _15283_, _15282_);
  and _66475_ (_15285_, _15284_, _07764_);
  and _66476_ (_15286_, _15285_, _14328_);
  or _66477_ (_41020_, _15286_, _15281_);
  or _66478_ (_15287_, _14156_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _66479_ (_15288_, _15287_, _14162_);
  nor _66480_ (_15289_, _09216_, _09207_);
  nor _66481_ (_15290_, _15289_, _09217_);
  or _66482_ (_15291_, _15290_, _07169_);
  not _66483_ (_15292_, _05820_);
  nor _66484_ (_15293_, _06129_, _15292_);
  nor _66485_ (_15294_, _12181_, _05846_);
  and _66486_ (_15295_, _10295_, _07126_);
  not _66487_ (_15296_, _12580_);
  and _66488_ (_15297_, _15296_, _12579_);
  or _66489_ (_15298_, _15297_, _08398_);
  nor _66490_ (_15299_, _08544_, _08014_);
  or _66491_ (_15300_, _15299_, _08545_);
  and _66492_ (_15301_, _15300_, _06162_);
  or _66493_ (_15302_, _09207_, _07065_);
  nor _66494_ (_15303_, _08354_, _08347_);
  nor _66495_ (_15304_, _15303_, _08355_);
  nor _66496_ (_15305_, _15304_, _08443_);
  nand _66497_ (_15306_, _12181_, _06581_);
  or _66498_ (_15307_, _06581_, \oc8051_golden_model_1.ACC [6]);
  and _66499_ (_15308_, _15307_, _15306_);
  and _66500_ (_15309_, _15308_, _08443_);
  or _66501_ (_15310_, _15309_, _07064_);
  or _66502_ (_15311_, _15310_, _15305_);
  and _66503_ (_15312_, _15311_, _08429_);
  and _66504_ (_15313_, _15312_, _15302_);
  or _66505_ (_15314_, _15313_, _15301_);
  and _66506_ (_15315_, _15314_, _08428_);
  or _66507_ (_15316_, _12580_, _12579_);
  and _66508_ (_15317_, _15316_, _06159_);
  or _66509_ (_15318_, _15317_, _07485_);
  or _66510_ (_15319_, _15318_, _15315_);
  nor _66511_ (_15320_, _12180_, _05764_);
  nor _66512_ (_15321_, _15320_, _07076_);
  and _66513_ (_15322_, _15321_, _15319_);
  and _66514_ (_15323_, _08012_, _07076_);
  or _66515_ (_15324_, _15323_, _07086_);
  or _66516_ (_15325_, _15324_, _15322_);
  and _66517_ (_15326_, _15325_, _15298_);
  or _66518_ (_15327_, _15326_, _06151_);
  nand _66519_ (_15328_, _08014_, _06151_);
  and _66520_ (_15329_, _15328_, _06149_);
  and _66521_ (_15330_, _15329_, _15327_);
  not _66522_ (_15331_, _12581_);
  and _66523_ (_15332_, _15316_, _15331_);
  and _66524_ (_15333_, _15332_, _06148_);
  or _66525_ (_15334_, _15333_, _15330_);
  and _66526_ (_15335_, _15334_, _05760_);
  or _66527_ (_15336_, _12181_, _05760_);
  nand _66528_ (_15337_, _15336_, _06251_);
  or _66529_ (_15338_, _15337_, _15335_);
  nand _66530_ (_15339_, _08014_, _06252_);
  and _66531_ (_15340_, _15339_, _15338_);
  or _66532_ (_15341_, _15340_, _06701_);
  and _66533_ (_15342_, _09207_, _06172_);
  or _66534_ (_15343_, _07959_, _07104_);
  or _66535_ (_15344_, _15343_, _15342_);
  and _66536_ (_15345_, _15344_, _08580_);
  and _66537_ (_15346_, _15345_, _15341_);
  and _66538_ (_15347_, _12580_, \oc8051_golden_model_1.PSW [7]);
  or _66539_ (_15348_, _15347_, _15297_);
  and _66540_ (_15349_, _15348_, _07103_);
  or _66541_ (_15350_, _15349_, _05791_);
  or _66542_ (_15351_, _15350_, _15346_);
  and _66543_ (_15352_, _12181_, _05791_);
  nor _66544_ (_15353_, _15352_, _08591_);
  and _66545_ (_15354_, _15353_, _15351_);
  and _66546_ (_15355_, _08012_, _08591_);
  or _66547_ (_15356_, _15355_, _08595_);
  or _66548_ (_15357_, _15356_, _15354_);
  or _66549_ (_15358_, _09207_, _08601_);
  and _66550_ (_15359_, _15358_, _08600_);
  and _66551_ (_15360_, _15359_, _15357_);
  and _66552_ (_15361_, _08395_, _08012_);
  and _66553_ (_15362_, _08738_, \oc8051_golden_model_1.ACC [6]);
  and _66554_ (_15363_, _08741_, \oc8051_golden_model_1.B [6]);
  or _66555_ (_15364_, _15363_, _15362_);
  and _66556_ (_15365_, _08734_, \oc8051_golden_model_1.PSW [6]);
  or _66557_ (_15366_, _15365_, _15364_);
  and _66558_ (_15367_, _08752_, \oc8051_golden_model_1.SBUF [6]);
  and _66559_ (_15368_, _08749_, \oc8051_golden_model_1.IE [6]);
  or _66560_ (_15369_, _15368_, _15367_);
  and _66561_ (_15370_, _08746_, \oc8051_golden_model_1.IP [6]);
  or _66562_ (_15371_, _15370_, _15369_);
  or _66563_ (_15372_, _15371_, _15366_);
  and _66564_ (_15373_, _08724_, \oc8051_golden_model_1.TL1 [6]);
  and _66565_ (_15374_, _08706_, \oc8051_golden_model_1.TH0 [6]);
  and _66566_ (_15375_, _08710_, \oc8051_golden_model_1.TH1 [6]);
  and _66567_ (_15376_, _08718_, \oc8051_golden_model_1.SCON [6]);
  or _66568_ (_15377_, _15376_, _15375_);
  or _66569_ (_15378_, _15377_, _15374_);
  or _66570_ (_15379_, _15378_, _15373_);
  or _66571_ (_15380_, _15379_, _15372_);
  and _66572_ (_15381_, _08765_, \oc8051_golden_model_1.DPL [6]);
  and _66573_ (_15382_, _08758_, \oc8051_golden_model_1.SP [6]);
  and _66574_ (_15383_, _08760_, \oc8051_golden_model_1.DPH [6]);
  or _66575_ (_15384_, _15383_, _15382_);
  or _66576_ (_15385_, _15384_, _15381_);
  and _66577_ (_15386_, _08773_, \oc8051_golden_model_1.TL0 [6]);
  and _66578_ (_15387_, _08775_, \oc8051_golden_model_1.TMOD [6]);
  or _66579_ (_15388_, _15387_, _15386_);
  and _66580_ (_15389_, _08770_, \oc8051_golden_model_1.PCON [6]);
  and _66581_ (_15390_, _08726_, \oc8051_golden_model_1.TCON [6]);
  or _66582_ (_15391_, _15390_, _15389_);
  or _66583_ (_15392_, _15391_, _15388_);
  or _66584_ (_15393_, _15392_, _15385_);
  or _66585_ (_15394_, _15393_, _15380_);
  or _66586_ (_15395_, _15394_, _15361_);
  and _66587_ (_15396_, _15395_, _08599_);
  or _66588_ (_15397_, _15396_, _08788_);
  or _66589_ (_15398_, _15397_, _15360_);
  and _66590_ (_15399_, _08788_, _06203_);
  nor _66591_ (_15400_, _15399_, _06112_);
  and _66592_ (_15401_, _15400_, _15398_);
  not _66593_ (_15402_, _08638_);
  and _66594_ (_15403_, _15402_, _06112_);
  or _66595_ (_15404_, _15403_, _06076_);
  or _66596_ (_15405_, _15404_, _15401_);
  or _66597_ (_15406_, _12180_, _05836_);
  and _66598_ (_15407_, _15406_, _15405_);
  or _66599_ (_15408_, _15407_, _07128_);
  not _66600_ (_15409_, _07128_);
  nand _66601_ (_15410_, _08638_, _08014_);
  nor _66602_ (_15411_, _08638_, _08014_);
  not _66603_ (_15412_, _15411_);
  and _66604_ (_15413_, _15412_, _15410_);
  or _66605_ (_15414_, _15413_, _15409_);
  and _66606_ (_15415_, _15414_, _08807_);
  and _66607_ (_15416_, _15415_, _15408_);
  or _66608_ (_15417_, _15416_, _15295_);
  and _66609_ (_15418_, _15417_, _08806_);
  and _66610_ (_15419_, _15411_, _07133_);
  or _66611_ (_15420_, _15419_, _15418_);
  and _66612_ (_15421_, _15420_, _08364_);
  and _66613_ (_15422_, _10266_, _07131_);
  or _66614_ (_15423_, _15422_, _07124_);
  or _66615_ (_15424_, _15423_, _15421_);
  nor _66616_ (_15425_, _12180_, _05848_);
  nor _66617_ (_15426_, _15425_, _08820_);
  and _66618_ (_15427_, _15426_, _15424_);
  and _66619_ (_15428_, _15410_, _08820_);
  or _66620_ (_15429_, _15428_, _08825_);
  or _66621_ (_15430_, _15429_, _15427_);
  nand _66622_ (_15431_, _10294_, _08825_);
  and _66623_ (_15432_, _15431_, _05846_);
  and _66624_ (_15433_, _15432_, _15430_);
  or _66625_ (_15434_, _15433_, _15294_);
  and _66626_ (_15435_, _15434_, _08361_);
  nor _66627_ (_15436_, _15304_, _08361_);
  or _66628_ (_15437_, _15436_, _07325_);
  nor _66629_ (_15438_, _15437_, _15435_);
  and _66630_ (_15439_, _15304_, _07325_);
  or _66631_ (_15440_, _15439_, _14487_);
  nor _66632_ (_15441_, _15440_, _15438_);
  nor _66633_ (_15442_, _09165_, _08883_);
  nor _66634_ (_15443_, _15442_, _09166_);
  nand _66635_ (_15444_, _15443_, _06276_);
  and _66636_ (_15445_, _15444_, _07153_);
  or _66637_ (_15446_, _15445_, _15441_);
  nand _66638_ (_15447_, _15443_, _14495_);
  and _66639_ (_15448_, _15447_, _08837_);
  and _66640_ (_15449_, _15448_, _15446_);
  and _66641_ (_15450_, _15300_, _07152_);
  or _66642_ (_15451_, _15450_, _06310_);
  or _66643_ (_15452_, _15451_, _15449_);
  nand _66644_ (_15453_, _12006_, _06310_);
  and _66645_ (_15454_, _15453_, _12730_);
  and _66646_ (_15455_, _15454_, _15452_);
  and _66647_ (_15456_, _12180_, _05823_);
  or _66648_ (_15457_, _15456_, _06073_);
  or _66649_ (_15458_, _15457_, _15455_);
  and _66650_ (_15459_, _06539_, _07369_);
  nor _66651_ (_15460_, _15297_, _06074_);
  nor _66652_ (_15461_, _15460_, _15459_);
  and _66653_ (_15462_, _15461_, _15458_);
  nor _66654_ (_15463_, _09199_, _08012_);
  nor _66655_ (_15464_, _15463_, _09200_);
  and _66656_ (_15465_, _15464_, _15459_);
  or _66657_ (_15466_, _15465_, _15462_);
  or _66658_ (_15467_, _15466_, _15293_);
  not _66659_ (_15468_, _15293_);
  nor _66660_ (_15469_, _15464_, _15468_);
  nor _66661_ (_15470_, _15469_, _07394_);
  and _66662_ (_15471_, _15470_, _15467_);
  and _66663_ (_15472_, _15464_, _07394_);
  or _66664_ (_15473_, _15472_, _07168_);
  or _66665_ (_15474_, _15473_, _15471_);
  and _66666_ (_15475_, _15474_, _15291_);
  or _66667_ (_15476_, _15475_, _07167_);
  nor _66668_ (_15477_, _08341_, _08015_);
  nor _66669_ (_15478_, _15477_, _08342_);
  or _66670_ (_15479_, _15478_, _14518_);
  and _66671_ (_15480_, _15479_, _07417_);
  and _66672_ (_15481_, _15480_, _15476_);
  or _66673_ (_15482_, _15481_, _14164_);
  and _66674_ (_15483_, _15482_, _15288_);
  nand _66675_ (_15484_, _11966_, _06310_);
  or _66676_ (_15485_, _12146_, _06310_);
  and _66677_ (_15486_, _15485_, _15484_);
  and _66678_ (_15487_, _15486_, _07764_);
  and _66679_ (_15488_, _15487_, _14328_);
  or _66680_ (_41021_, _15488_, _15483_);
  or _66681_ (_15489_, _14156_, \oc8051_golden_model_1.IRAM[0] [7]);
  nand _66682_ (_15490_, _14156_, _09225_);
  and _66683_ (_15491_, _15490_, _15489_);
  or _66684_ (_15492_, _15491_, _14161_);
  or _66685_ (_15493_, _14162_, _09258_);
  and _66686_ (_41022_, _15493_, _15492_);
  and _66687_ (_15494_, _14153_, _07345_);
  and _66688_ (_15495_, _15494_, _14152_);
  not _66689_ (_15496_, _15495_);
  or _66690_ (_15497_, _15496_, _14324_);
  or _66691_ (_15498_, _15495_, \oc8051_golden_model_1.IRAM[1] [0]);
  not _66692_ (_15499_, _07764_);
  nand _66693_ (_15500_, _14159_, _07476_);
  or _66694_ (_15501_, _15500_, _15499_);
  and _66695_ (_15502_, _15501_, _15498_);
  and _66696_ (_15503_, _15502_, _15497_);
  and _66697_ (_15504_, _07764_, _07476_);
  and _66698_ (_15505_, _15504_, _14159_);
  and _66699_ (_15506_, _15505_, _14332_);
  or _66700_ (_41027_, _15506_, _15503_);
  or _66701_ (_15507_, _15496_, _14521_);
  or _66702_ (_15508_, _15495_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _66703_ (_15509_, _15508_, _15501_);
  and _66704_ (_15510_, _15509_, _15507_);
  and _66705_ (_15511_, _15505_, _14527_);
  or _66706_ (_41028_, _15511_, _15510_);
  or _66707_ (_15512_, _15496_, _14713_);
  or _66708_ (_15513_, _15495_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _66709_ (_15514_, _15513_, _15501_);
  and _66710_ (_15515_, _15514_, _15512_);
  and _66711_ (_15516_, _15505_, _14719_);
  or _66712_ (_41029_, _15516_, _15515_);
  or _66713_ (_15517_, _15496_, _14900_);
  or _66714_ (_15518_, _15495_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _66715_ (_15519_, _15518_, _15501_);
  and _66716_ (_15520_, _15519_, _15517_);
  and _66717_ (_15521_, _15505_, _14906_);
  or _66718_ (_41030_, _15521_, _15520_);
  or _66719_ (_15522_, _15496_, _15090_);
  or _66720_ (_15523_, _15495_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _66721_ (_15524_, _15523_, _15501_);
  and _66722_ (_15525_, _15524_, _15522_);
  and _66723_ (_15526_, _15505_, _15097_);
  or _66724_ (_41031_, _15526_, _15525_);
  or _66725_ (_15527_, _15496_, _15278_);
  or _66726_ (_15528_, _15495_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _66727_ (_15529_, _15528_, _15501_);
  and _66728_ (_15530_, _15529_, _15527_);
  and _66729_ (_15531_, _15505_, _15285_);
  or _66730_ (_41033_, _15531_, _15530_);
  or _66731_ (_15532_, _15496_, _15481_);
  or _66732_ (_15533_, _15495_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _66733_ (_15534_, _15533_, _15501_);
  and _66734_ (_15535_, _15534_, _15532_);
  and _66735_ (_15536_, _15505_, _15487_);
  or _66736_ (_41034_, _15536_, _15535_);
  or _66737_ (_15537_, _15496_, _09226_);
  or _66738_ (_15538_, _15495_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _66739_ (_15539_, _15538_, _15501_);
  and _66740_ (_15540_, _15539_, _15537_);
  and _66741_ (_15541_, _15505_, _09259_);
  or _66742_ (_41035_, _15541_, _15540_);
  and _66743_ (_15542_, _07419_, _07174_);
  and _66744_ (_15543_, _15542_, _14152_);
  not _66745_ (_15544_, _15543_);
  or _66746_ (_15545_, _15544_, _14324_);
  or _66747_ (_15546_, _15543_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand _66748_ (_15547_, _14159_, _08449_);
  or _66749_ (_15548_, _15547_, _15499_);
  and _66750_ (_15549_, _15548_, _15546_);
  and _66751_ (_15550_, _15549_, _15545_);
  and _66752_ (_15551_, _08449_, _07764_);
  and _66753_ (_15552_, _15551_, _14159_);
  and _66754_ (_15553_, _15552_, _14332_);
  or _66755_ (_41038_, _15553_, _15550_);
  or _66756_ (_15554_, _15544_, _14521_);
  or _66757_ (_15555_, _15543_, \oc8051_golden_model_1.IRAM[2] [1]);
  and _66758_ (_15556_, _15555_, _15548_);
  and _66759_ (_15557_, _15556_, _15554_);
  and _66760_ (_15558_, _15552_, _14527_);
  or _66761_ (_41041_, _15558_, _15557_);
  or _66762_ (_15559_, _15544_, _14713_);
  or _66763_ (_15560_, _15543_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _66764_ (_15561_, _15560_, _15548_);
  and _66765_ (_15562_, _15561_, _15559_);
  and _66766_ (_15563_, _15552_, _14719_);
  or _66767_ (_41042_, _15563_, _15562_);
  or _66768_ (_15564_, _15544_, _14900_);
  or _66769_ (_15565_, _15543_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _66770_ (_15566_, _15565_, _15548_);
  and _66771_ (_15567_, _15566_, _15564_);
  and _66772_ (_15568_, _15552_, _14906_);
  or _66773_ (_41043_, _15568_, _15567_);
  or _66774_ (_15569_, _15544_, _15090_);
  or _66775_ (_15570_, _15543_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _66776_ (_15571_, _15570_, _15548_);
  and _66777_ (_15572_, _15571_, _15569_);
  and _66778_ (_15573_, _15552_, _15097_);
  or _66779_ (_41044_, _15573_, _15572_);
  or _66780_ (_15574_, _15544_, _15278_);
  or _66781_ (_15575_, _15543_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _66782_ (_15576_, _15575_, _15548_);
  and _66783_ (_15577_, _15576_, _15574_);
  and _66784_ (_15578_, _15552_, _15285_);
  or _66785_ (_41045_, _15578_, _15577_);
  or _66786_ (_15579_, _15544_, _15481_);
  or _66787_ (_15580_, _15543_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _66788_ (_15581_, _15580_, _15548_);
  and _66789_ (_15582_, _15581_, _15579_);
  and _66790_ (_15583_, _15552_, _15487_);
  or _66791_ (_41047_, _15583_, _15582_);
  and _66792_ (_15584_, _15543_, _09226_);
  or _66793_ (_15585_, _15543_, _07871_);
  nand _66794_ (_15586_, _15585_, _15548_);
  or _66795_ (_15587_, _15586_, _15584_);
  or _66796_ (_15588_, _15548_, _09258_);
  and _66797_ (_41048_, _15588_, _15587_);
  and _66798_ (_15589_, _14152_, _07421_);
  or _66799_ (_15590_, _15589_, \oc8051_golden_model_1.IRAM[3] [0]);
  nand _66800_ (_15591_, _14159_, _07177_);
  or _66801_ (_15592_, _15591_, _15499_);
  and _66802_ (_15593_, _15592_, _15590_);
  not _66803_ (_15594_, _15589_);
  or _66804_ (_15595_, _15594_, _14324_);
  and _66805_ (_15596_, _15595_, _15593_);
  and _66806_ (_15597_, _07764_, _07177_);
  and _66807_ (_15598_, _15597_, _14159_);
  and _66808_ (_15599_, _15598_, _14332_);
  or _66809_ (_41052_, _15599_, _15596_);
  or _66810_ (_15600_, _15589_, \oc8051_golden_model_1.IRAM[3] [1]);
  and _66811_ (_15601_, _15600_, _15592_);
  or _66812_ (_15602_, _15594_, _14521_);
  and _66813_ (_15603_, _15602_, _15601_);
  and _66814_ (_15604_, _15598_, _14527_);
  or _66815_ (_41053_, _15604_, _15603_);
  or _66816_ (_15605_, _15589_, \oc8051_golden_model_1.IRAM[3] [2]);
  and _66817_ (_15606_, _15605_, _15592_);
  or _66818_ (_15607_, _15594_, _14713_);
  and _66819_ (_15608_, _15607_, _15606_);
  and _66820_ (_15609_, _15598_, _14719_);
  or _66821_ (_41054_, _15609_, _15608_);
  or _66822_ (_15610_, _15589_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _66823_ (_15611_, _15610_, _15592_);
  or _66824_ (_15612_, _15594_, _14900_);
  and _66825_ (_15613_, _15612_, _15611_);
  and _66826_ (_15614_, _15598_, _14906_);
  or _66827_ (_41055_, _15614_, _15613_);
  or _66828_ (_15615_, _15589_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _66829_ (_15616_, _15615_, _15592_);
  or _66830_ (_15617_, _15594_, _15090_);
  and _66831_ (_15618_, _15617_, _15616_);
  and _66832_ (_15619_, _15598_, _15097_);
  or _66833_ (_41056_, _15619_, _15618_);
  or _66834_ (_15620_, _15589_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _66835_ (_15621_, _15620_, _15592_);
  or _66836_ (_15622_, _15594_, _15278_);
  and _66837_ (_15623_, _15622_, _15621_);
  and _66838_ (_15624_, _15598_, _15285_);
  or _66839_ (_41058_, _15624_, _15623_);
  or _66840_ (_15625_, _15589_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _66841_ (_15626_, _15625_, _15592_);
  or _66842_ (_15627_, _15594_, _15481_);
  and _66843_ (_15628_, _15627_, _15626_);
  and _66844_ (_15629_, _15598_, _15487_);
  or _66845_ (_41059_, _15629_, _15628_);
  or _66846_ (_15630_, _15589_, \oc8051_golden_model_1.IRAM[3] [7]);
  and _66847_ (_15631_, _15630_, _15592_);
  or _66848_ (_15632_, _15594_, _09226_);
  and _66849_ (_15633_, _15632_, _15631_);
  and _66850_ (_15634_, _15598_, _09259_);
  or _66851_ (_41060_, _15634_, _15633_);
  and _66852_ (_15635_, _07747_, _07593_);
  and _66853_ (_15636_, _15635_, _14154_);
  not _66854_ (_15637_, _15636_);
  or _66855_ (_15638_, _15637_, _14324_);
  not _66856_ (_15639_, _07759_);
  and _66857_ (_15640_, _14158_, _15639_);
  and _66858_ (_15641_, _15640_, _07178_);
  not _66859_ (_15642_, _15641_);
  or _66860_ (_15643_, _15636_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _66861_ (_15644_, _15643_, _15642_);
  and _66862_ (_15645_, _15644_, _15638_);
  and _66863_ (_15646_, _15641_, _14332_);
  or _66864_ (_41063_, _15646_, _15645_);
  or _66865_ (_15647_, _15637_, _14521_);
  or _66866_ (_15648_, _15636_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _66867_ (_15649_, _15648_, _15642_);
  and _66868_ (_15650_, _15649_, _15647_);
  and _66869_ (_15651_, _15641_, _14527_);
  or _66870_ (_41066_, _15651_, _15650_);
  or _66871_ (_15652_, _15637_, _14713_);
  or _66872_ (_15653_, _15636_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _66873_ (_15654_, _15653_, _15642_);
  and _66874_ (_15655_, _15654_, _15652_);
  and _66875_ (_15656_, _15641_, _14719_);
  or _66876_ (_41067_, _15656_, _15655_);
  or _66877_ (_15657_, _15637_, _14900_);
  or _66878_ (_15658_, _15636_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _66879_ (_15659_, _15658_, _15642_);
  and _66880_ (_15660_, _15659_, _15657_);
  and _66881_ (_15661_, _15641_, _14906_);
  or _66882_ (_41068_, _15661_, _15660_);
  or _66883_ (_15662_, _15637_, _15090_);
  or _66884_ (_15663_, _15636_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _66885_ (_15664_, _15663_, _15642_);
  and _66886_ (_15665_, _15664_, _15662_);
  and _66887_ (_15666_, _15641_, _15097_);
  or _66888_ (_41069_, _15666_, _15665_);
  or _66889_ (_15667_, _15637_, _15278_);
  or _66890_ (_15668_, _15636_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _66891_ (_15669_, _15668_, _15642_);
  and _66892_ (_15670_, _15669_, _15667_);
  and _66893_ (_15671_, _15641_, _15285_);
  or _66894_ (_41070_, _15671_, _15670_);
  or _66895_ (_15672_, _15637_, _15481_);
  or _66896_ (_15673_, _15636_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _66897_ (_15674_, _15673_, _15642_);
  and _66898_ (_15675_, _15674_, _15672_);
  and _66899_ (_15676_, _15641_, _15487_);
  or _66900_ (_41071_, _15676_, _15675_);
  or _66901_ (_15677_, _15637_, _09226_);
  or _66902_ (_15678_, _15636_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _66903_ (_15679_, _15678_, _15642_);
  and _66904_ (_15680_, _15679_, _15677_);
  and _66905_ (_15681_, _15641_, _09259_);
  or _66906_ (_41072_, _15681_, _15680_);
  and _66907_ (_15682_, _15635_, _15494_);
  not _66908_ (_15683_, _15682_);
  or _66909_ (_15684_, _15683_, _14324_);
  and _66910_ (_15685_, _15640_, _07476_);
  not _66911_ (_15686_, _15685_);
  or _66912_ (_15687_, _15682_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _66913_ (_15688_, _15687_, _15686_);
  and _66914_ (_15689_, _15688_, _15684_);
  and _66915_ (_15690_, _15685_, _14332_);
  or _66916_ (_41075_, _15690_, _15689_);
  or _66917_ (_15691_, _15683_, _14521_);
  or _66918_ (_15692_, _15682_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _66919_ (_15693_, _15692_, _15686_);
  and _66920_ (_15694_, _15693_, _15691_);
  and _66921_ (_15695_, _15685_, _14527_);
  or _66922_ (_41077_, _15695_, _15694_);
  or _66923_ (_15696_, _15683_, _14713_);
  or _66924_ (_15697_, _15682_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _66925_ (_15698_, _15697_, _15686_);
  and _66926_ (_15699_, _15698_, _15696_);
  and _66927_ (_15700_, _15685_, _14719_);
  or _66928_ (_41078_, _15700_, _15699_);
  or _66929_ (_15701_, _15683_, _14900_);
  or _66930_ (_15702_, _15682_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _66931_ (_15703_, _15702_, _15686_);
  and _66932_ (_15704_, _15703_, _15701_);
  and _66933_ (_15705_, _15685_, _14906_);
  or _66934_ (_41079_, _15705_, _15704_);
  or _66935_ (_15706_, _15683_, _15090_);
  or _66936_ (_15707_, _15682_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _66937_ (_15708_, _15707_, _15686_);
  and _66938_ (_15709_, _15708_, _15706_);
  and _66939_ (_15710_, _15685_, _15097_);
  or _66940_ (_41080_, _15710_, _15709_);
  or _66941_ (_15711_, _15683_, _15278_);
  or _66942_ (_15712_, _15682_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _66943_ (_15713_, _15712_, _15686_);
  and _66944_ (_15714_, _15713_, _15711_);
  and _66945_ (_15715_, _15685_, _15285_);
  or _66946_ (_41081_, _15715_, _15714_);
  or _66947_ (_15716_, _15683_, _15481_);
  or _66948_ (_15717_, _15682_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _66949_ (_15718_, _15717_, _15686_);
  and _66950_ (_15719_, _15718_, _15716_);
  and _66951_ (_15720_, _15685_, _15487_);
  or _66952_ (_41083_, _15720_, _15719_);
  or _66953_ (_15721_, _15683_, _09226_);
  or _66954_ (_15722_, _15682_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _66955_ (_15723_, _15722_, _15686_);
  and _66956_ (_15724_, _15723_, _15721_);
  and _66957_ (_15725_, _15685_, _09259_);
  or _66958_ (_41084_, _15725_, _15724_);
  and _66959_ (_15726_, _15635_, _15542_);
  not _66960_ (_15727_, _15726_);
  or _66961_ (_15728_, _15727_, _14324_);
  and _66962_ (_15729_, _15640_, _08449_);
  not _66963_ (_15730_, _15729_);
  or _66964_ (_15731_, _15726_, \oc8051_golden_model_1.IRAM[6] [0]);
  and _66965_ (_15732_, _15731_, _15730_);
  and _66966_ (_15733_, _15732_, _15728_);
  and _66967_ (_15734_, _15729_, _14332_);
  or _66968_ (_41088_, _15734_, _15733_);
  or _66969_ (_15735_, _15727_, _14521_);
  or _66970_ (_15736_, _15726_, \oc8051_golden_model_1.IRAM[6] [1]);
  and _66971_ (_15737_, _15736_, _15730_);
  and _66972_ (_15738_, _15737_, _15735_);
  and _66973_ (_15739_, _15729_, _14527_);
  or _66974_ (_41089_, _15739_, _15738_);
  or _66975_ (_15740_, _15727_, _14713_);
  or _66976_ (_15741_, _15726_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _66977_ (_15742_, _15741_, _15730_);
  and _66978_ (_15743_, _15742_, _15740_);
  and _66979_ (_15744_, _15729_, _14719_);
  or _66980_ (_41090_, _15744_, _15743_);
  or _66981_ (_15745_, _15727_, _14900_);
  or _66982_ (_15746_, _15726_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _66983_ (_15747_, _15746_, _15730_);
  and _66984_ (_15748_, _15747_, _15745_);
  and _66985_ (_15749_, _15729_, _14906_);
  or _66986_ (_41091_, _15749_, _15748_);
  or _66987_ (_15750_, _15727_, _15090_);
  or _66988_ (_15751_, _15726_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _66989_ (_15752_, _15751_, _15730_);
  and _66990_ (_15753_, _15752_, _15750_);
  and _66991_ (_15754_, _15729_, _15097_);
  or _66992_ (_41092_, _15754_, _15753_);
  or _66993_ (_15755_, _15727_, _15278_);
  or _66994_ (_15756_, _15726_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _66995_ (_15757_, _15756_, _15730_);
  and _66996_ (_15758_, _15757_, _15755_);
  and _66997_ (_15759_, _15729_, _15285_);
  or _66998_ (_41094_, _15759_, _15758_);
  or _66999_ (_15760_, _15727_, _15481_);
  or _67000_ (_15761_, _15726_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _67001_ (_15762_, _15761_, _15730_);
  and _67002_ (_15763_, _15762_, _15760_);
  and _67003_ (_15764_, _15729_, _15487_);
  or _67004_ (_41095_, _15764_, _15763_);
  or _67005_ (_15765_, _15727_, _09226_);
  or _67006_ (_15766_, _15726_, \oc8051_golden_model_1.IRAM[6] [7]);
  and _67007_ (_15767_, _15766_, _15730_);
  and _67008_ (_15768_, _15767_, _15765_);
  and _67009_ (_15769_, _15729_, _09259_);
  or _67010_ (_41096_, _15769_, _15768_);
  and _67011_ (_15770_, _15640_, _07177_);
  not _67012_ (_15771_, _15770_);
  or _67013_ (_15772_, _15771_, _14332_);
  and _67014_ (_15773_, _15635_, _07421_);
  and _67015_ (_15774_, _15773_, _14324_);
  nor _67016_ (_15775_, _15773_, _07007_);
  or _67017_ (_15776_, _15775_, _15770_);
  or _67018_ (_15777_, _15776_, _15774_);
  and _67019_ (_41100_, _15777_, _15772_);
  nor _67020_ (_15778_, _15773_, _07207_);
  and _67021_ (_15779_, _15773_, _14521_);
  or _67022_ (_15780_, _15779_, _15778_);
  and _67023_ (_15781_, _15780_, _15771_);
  and _67024_ (_15782_, _15770_, _14527_);
  or _67025_ (_41101_, _15782_, _15781_);
  or _67026_ (_15783_, _15773_, \oc8051_golden_model_1.IRAM[7] [2]);
  and _67027_ (_15784_, _15783_, _15771_);
  not _67028_ (_15785_, _15773_);
  or _67029_ (_15786_, _15785_, _14713_);
  and _67030_ (_15787_, _15786_, _15784_);
  and _67031_ (_15788_, _15770_, _14719_);
  or _67032_ (_41102_, _15788_, _15787_);
  or _67033_ (_15789_, _15773_, \oc8051_golden_model_1.IRAM[7] [3]);
  and _67034_ (_15790_, _15789_, _15771_);
  or _67035_ (_15791_, _15785_, _14900_);
  and _67036_ (_15792_, _15791_, _15790_);
  and _67037_ (_15793_, _15770_, _14906_);
  or _67038_ (_41103_, _15793_, _15792_);
  or _67039_ (_15794_, _15773_, \oc8051_golden_model_1.IRAM[7] [4]);
  and _67040_ (_15795_, _15794_, _15771_);
  or _67041_ (_15796_, _15785_, _15090_);
  and _67042_ (_15797_, _15796_, _15795_);
  and _67043_ (_15798_, _15770_, _15097_);
  or _67044_ (_41104_, _15798_, _15797_);
  or _67045_ (_15799_, _15773_, \oc8051_golden_model_1.IRAM[7] [5]);
  and _67046_ (_15800_, _15799_, _15771_);
  or _67047_ (_15801_, _15785_, _15278_);
  and _67048_ (_15802_, _15801_, _15800_);
  and _67049_ (_15803_, _15770_, _15285_);
  or _67050_ (_41106_, _15803_, _15802_);
  or _67051_ (_15804_, _15773_, \oc8051_golden_model_1.IRAM[7] [6]);
  and _67052_ (_15805_, _15804_, _15771_);
  or _67053_ (_15806_, _15785_, _15481_);
  and _67054_ (_15807_, _15806_, _15805_);
  and _67055_ (_15808_, _15770_, _15487_);
  or _67056_ (_41107_, _15808_, _15807_);
  or _67057_ (_15809_, _15773_, \oc8051_golden_model_1.IRAM[7] [7]);
  and _67058_ (_15810_, _15809_, _15771_);
  or _67059_ (_15811_, _15785_, _09226_);
  and _67060_ (_15812_, _15811_, _15810_);
  and _67061_ (_15813_, _15770_, _09259_);
  or _67062_ (_41108_, _15813_, _15812_);
  and _67063_ (_15814_, _14151_, _07746_);
  and _67064_ (_15815_, _15814_, _14154_);
  not _67065_ (_15816_, _15815_);
  or _67066_ (_15817_, _15816_, _14324_);
  or _67067_ (_15818_, _15815_, \oc8051_golden_model_1.IRAM[8] [0]);
  not _67068_ (_15819_, _07755_);
  and _67069_ (_15820_, _07765_, _15819_);
  and _67070_ (_15821_, _15820_, _07178_);
  not _67071_ (_15822_, _15821_);
  and _67072_ (_15823_, _15822_, _15818_);
  and _67073_ (_15824_, _15823_, _15817_);
  and _67074_ (_15825_, _15821_, _14332_);
  or _67075_ (_41112_, _15825_, _15824_);
  or _67076_ (_15826_, _15816_, _14521_);
  or _67077_ (_15827_, _15815_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _67078_ (_15828_, _15827_, _15822_);
  and _67079_ (_15829_, _15828_, _15826_);
  and _67080_ (_15830_, _15821_, _14527_);
  or _67081_ (_41114_, _15830_, _15829_);
  or _67082_ (_15831_, _15816_, _14713_);
  nand _67083_ (_15832_, _07765_, _07753_);
  or _67084_ (_15833_, _15815_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _67085_ (_15834_, _15833_, _15832_);
  and _67086_ (_15835_, _15834_, _15831_);
  and _67087_ (_15836_, _15821_, _14719_);
  or _67088_ (_41115_, _15836_, _15835_);
  or _67089_ (_15837_, _15816_, _14900_);
  or _67090_ (_15838_, _15815_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _67091_ (_15839_, _15838_, _15832_);
  and _67092_ (_15840_, _15839_, _15837_);
  and _67093_ (_15841_, _15821_, _14906_);
  or _67094_ (_41116_, _15841_, _15840_);
  or _67095_ (_15842_, _15816_, _15090_);
  or _67096_ (_15843_, _15815_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _67097_ (_15844_, _15843_, _15832_);
  and _67098_ (_15845_, _15844_, _15842_);
  and _67099_ (_15846_, _15821_, _15097_);
  or _67100_ (_41117_, _15846_, _15845_);
  or _67101_ (_15847_, _15816_, _15278_);
  or _67102_ (_15848_, _15815_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _67103_ (_15849_, _15848_, _15832_);
  and _67104_ (_15850_, _15849_, _15847_);
  and _67105_ (_15851_, _15821_, _15285_);
  or _67106_ (_41118_, _15851_, _15850_);
  or _67107_ (_15852_, _15816_, _15481_);
  or _67108_ (_15853_, _15815_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _67109_ (_15854_, _15853_, _15832_);
  and _67110_ (_15855_, _15854_, _15852_);
  and _67111_ (_15856_, _15821_, _15487_);
  or _67112_ (_41120_, _15856_, _15855_);
  and _67113_ (_15857_, _15815_, _09226_);
  or _67114_ (_15858_, _15815_, _07899_);
  nand _67115_ (_15859_, _15858_, _15832_);
  or _67116_ (_15860_, _15859_, _15857_);
  or _67117_ (_15861_, _15822_, _09259_);
  and _67118_ (_41121_, _15861_, _15860_);
  and _67119_ (_15862_, _15814_, _15494_);
  not _67120_ (_15863_, _15862_);
  or _67121_ (_15864_, _15863_, _14324_);
  or _67122_ (_15865_, _15862_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _67123_ (_15866_, _15820_, _07476_);
  not _67124_ (_15867_, _15866_);
  and _67125_ (_15868_, _15867_, _15865_);
  and _67126_ (_15869_, _15868_, _15864_);
  and _67127_ (_15870_, _15866_, _14332_);
  or _67128_ (_41123_, _15870_, _15869_);
  or _67129_ (_15871_, _15863_, _14521_);
  or _67130_ (_15872_, _15862_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _67131_ (_15873_, _15872_, _15867_);
  and _67132_ (_15874_, _15873_, _15871_);
  and _67133_ (_15875_, _15866_, _14527_);
  or _67134_ (_41124_, _15875_, _15874_);
  or _67135_ (_15876_, _15863_, _14713_);
  nand _67136_ (_15877_, _07765_, _07477_);
  or _67137_ (_15878_, _15862_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _67138_ (_15879_, _15878_, _15877_);
  and _67139_ (_15880_, _15879_, _15876_);
  and _67140_ (_15881_, _15866_, _14719_);
  or _67141_ (_41125_, _15881_, _15880_);
  or _67142_ (_15882_, _15863_, _14900_);
  or _67143_ (_15883_, _15862_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _67144_ (_15884_, _15883_, _15877_);
  and _67145_ (_15885_, _15884_, _15882_);
  and _67146_ (_15886_, _15866_, _14906_);
  or _67147_ (_41126_, _15886_, _15885_);
  or _67148_ (_15887_, _15863_, _15090_);
  or _67149_ (_15888_, _15862_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _67150_ (_15889_, _15888_, _15877_);
  and _67151_ (_15890_, _15889_, _15887_);
  and _67152_ (_15891_, _15866_, _15097_);
  or _67153_ (_41127_, _15891_, _15890_);
  or _67154_ (_15892_, _15863_, _15278_);
  or _67155_ (_15893_, _15862_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _67156_ (_15894_, _15893_, _15877_);
  and _67157_ (_15895_, _15894_, _15892_);
  and _67158_ (_15896_, _15866_, _15285_);
  or _67159_ (_41128_, _15896_, _15895_);
  or _67160_ (_15897_, _15863_, _15481_);
  or _67161_ (_15898_, _15862_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _67162_ (_15899_, _15898_, _15877_);
  and _67163_ (_15900_, _15899_, _15897_);
  and _67164_ (_15901_, _15866_, _15487_);
  or _67165_ (_41131_, _15901_, _15900_);
  and _67166_ (_15902_, _15862_, _09226_);
  or _67167_ (_15903_, _15862_, _07901_);
  nand _67168_ (_15904_, _15903_, _15877_);
  or _67169_ (_15905_, _15904_, _15902_);
  or _67170_ (_15906_, _15867_, _09259_);
  and _67171_ (_41132_, _15906_, _15905_);
  and _67172_ (_15907_, _15814_, _15542_);
  not _67173_ (_15908_, _15907_);
  or _67174_ (_15909_, _15908_, _14324_);
  and _67175_ (_15910_, _15820_, _08449_);
  not _67176_ (_15911_, _15910_);
  or _67177_ (_15912_, _15907_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _67178_ (_15913_, _15912_, _15911_);
  and _67179_ (_15914_, _15913_, _15909_);
  and _67180_ (_15915_, _15910_, _14332_);
  or _67181_ (_41136_, _15915_, _15914_);
  or _67182_ (_15916_, _15908_, _14521_);
  or _67183_ (_15917_, _15907_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _67184_ (_15918_, _15917_, _15911_);
  and _67185_ (_15919_, _15918_, _15916_);
  and _67186_ (_15920_, _15910_, _14527_);
  or _67187_ (_41137_, _15920_, _15919_);
  or _67188_ (_15921_, _15908_, _14713_);
  or _67189_ (_15922_, _15907_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _67190_ (_15923_, _15922_, _15911_);
  and _67191_ (_15924_, _15923_, _15921_);
  and _67192_ (_15925_, _15910_, _14719_);
  or _67193_ (_41138_, _15925_, _15924_);
  or _67194_ (_15926_, _15908_, _14900_);
  or _67195_ (_15927_, _15907_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _67196_ (_15928_, _15927_, _15911_);
  and _67197_ (_15929_, _15928_, _15926_);
  and _67198_ (_15930_, _15910_, _14906_);
  or _67199_ (_41139_, _15930_, _15929_);
  or _67200_ (_15931_, _15908_, _15090_);
  or _67201_ (_15932_, _15907_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _67202_ (_15933_, _15932_, _15911_);
  and _67203_ (_15934_, _15933_, _15931_);
  and _67204_ (_15935_, _15910_, _15097_);
  or _67205_ (_41140_, _15935_, _15934_);
  or _67206_ (_15936_, _15908_, _15278_);
  or _67207_ (_15937_, _15907_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _67208_ (_15938_, _15937_, _15911_);
  and _67209_ (_15939_, _15938_, _15936_);
  and _67210_ (_15940_, _15910_, _15285_);
  or _67211_ (_41142_, _15940_, _15939_);
  or _67212_ (_15941_, _15908_, _15481_);
  or _67213_ (_15942_, _15907_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _67214_ (_15943_, _15942_, _15911_);
  and _67215_ (_15944_, _15943_, _15941_);
  and _67216_ (_15945_, _15910_, _15487_);
  or _67217_ (_41143_, _15945_, _15944_);
  or _67218_ (_15946_, _15908_, _09226_);
  or _67219_ (_15947_, _15907_, \oc8051_golden_model_1.IRAM[10] [7]);
  and _67220_ (_15948_, _15947_, _15911_);
  and _67221_ (_15949_, _15948_, _15946_);
  and _67222_ (_15950_, _15910_, _09259_);
  or _67223_ (_41144_, _15950_, _15949_);
  not _67224_ (_15951_, _07345_);
  and _67225_ (_15952_, _14153_, _15951_);
  and _67226_ (_15953_, _15814_, _15952_);
  not _67227_ (_15954_, _15953_);
  or _67228_ (_15955_, _15954_, _14324_);
  and _67229_ (_15956_, _15820_, _07177_);
  not _67230_ (_15957_, _15956_);
  or _67231_ (_15958_, _15953_, \oc8051_golden_model_1.IRAM[11] [0]);
  and _67232_ (_15959_, _15958_, _15957_);
  and _67233_ (_15960_, _15959_, _15955_);
  and _67234_ (_15961_, _15956_, _14332_);
  or _67235_ (_41148_, _15961_, _15960_);
  or _67236_ (_15962_, _15954_, _14521_);
  or _67237_ (_15963_, _15953_, \oc8051_golden_model_1.IRAM[11] [1]);
  and _67238_ (_15964_, _15963_, _15957_);
  and _67239_ (_15965_, _15964_, _15962_);
  and _67240_ (_15966_, _15956_, _14527_);
  or _67241_ (_41149_, _15966_, _15965_);
  or _67242_ (_15967_, _15954_, _14713_);
  or _67243_ (_15968_, _15953_, \oc8051_golden_model_1.IRAM[11] [2]);
  and _67244_ (_15969_, _15968_, _15957_);
  and _67245_ (_15970_, _15969_, _15967_);
  and _67246_ (_15971_, _15956_, _14719_);
  or _67247_ (_41150_, _15971_, _15970_);
  and _67248_ (_15972_, _15814_, _07421_);
  or _67249_ (_15973_, _15972_, \oc8051_golden_model_1.IRAM[11] [3]);
  and _67250_ (_15974_, _15973_, _15957_);
  not _67251_ (_15975_, _15972_);
  or _67252_ (_15976_, _15975_, _14900_);
  and _67253_ (_15977_, _15976_, _15974_);
  and _67254_ (_15978_, _15956_, _14906_);
  or _67255_ (_41151_, _15978_, _15977_);
  or _67256_ (_15979_, _15972_, \oc8051_golden_model_1.IRAM[11] [4]);
  and _67257_ (_15980_, _15979_, _15957_);
  or _67258_ (_15981_, _15975_, _15090_);
  and _67259_ (_15982_, _15981_, _15980_);
  and _67260_ (_15983_, _15956_, _15097_);
  or _67261_ (_41152_, _15983_, _15982_);
  or _67262_ (_15984_, _15972_, \oc8051_golden_model_1.IRAM[11] [5]);
  and _67263_ (_15985_, _15984_, _15957_);
  or _67264_ (_15986_, _15975_, _15278_);
  and _67265_ (_15987_, _15986_, _15985_);
  and _67266_ (_15988_, _15956_, _15285_);
  or _67267_ (_41153_, _15988_, _15987_);
  or _67268_ (_15989_, _15972_, \oc8051_golden_model_1.IRAM[11] [6]);
  and _67269_ (_15990_, _15989_, _15957_);
  or _67270_ (_15991_, _15975_, _15481_);
  and _67271_ (_15992_, _15991_, _15990_);
  and _67272_ (_15993_, _15956_, _15487_);
  or _67273_ (_41154_, _15993_, _15992_);
  or _67274_ (_15994_, _15972_, \oc8051_golden_model_1.IRAM[11] [7]);
  and _67275_ (_15995_, _15994_, _15957_);
  or _67276_ (_15996_, _15975_, _09226_);
  and _67277_ (_15997_, _15996_, _15995_);
  and _67278_ (_15998_, _15956_, _09259_);
  or _67279_ (_41155_, _15998_, _15997_);
  not _67280_ (_15999_, _07178_);
  nand _67281_ (_16000_, _14158_, _07759_);
  or _67282_ (_16001_, _16000_, _15999_);
  or _67283_ (_16002_, _16001_, _14332_);
  and _67284_ (_16003_, _14154_, _07749_);
  and _67285_ (_16004_, _16003_, _14324_);
  or _67286_ (_16005_, _16003_, _07039_);
  nand _67287_ (_16006_, _16005_, _16001_);
  or _67288_ (_16007_, _16006_, _16004_);
  and _67289_ (_41158_, _16007_, _16002_);
  not _67290_ (_16008_, _07746_);
  and _67291_ (_16009_, _14151_, _16008_);
  and _67292_ (_16010_, _14154_, _16009_);
  not _67293_ (_16011_, _16010_);
  or _67294_ (_16012_, _16011_, _14521_);
  and _67295_ (_16013_, _07766_, _07178_);
  not _67296_ (_16014_, _16013_);
  or _67297_ (_16015_, _16010_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _67298_ (_16016_, _16015_, _16014_);
  and _67299_ (_16017_, _16016_, _16012_);
  and _67300_ (_16018_, _16013_, _14527_);
  or _67301_ (_41159_, _16018_, _16017_);
  or _67302_ (_16019_, _16003_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _67303_ (_16020_, _16019_, _16014_);
  or _67304_ (_16021_, _16011_, _14713_);
  and _67305_ (_16022_, _16021_, _16020_);
  and _67306_ (_16023_, _16013_, _14719_);
  or _67307_ (_41160_, _16023_, _16022_);
  or _67308_ (_16024_, _16003_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _67309_ (_16025_, _16024_, _16014_);
  or _67310_ (_16026_, _16011_, _14900_);
  and _67311_ (_16027_, _16026_, _16025_);
  and _67312_ (_16028_, _16013_, _14906_);
  or _67313_ (_41162_, _16028_, _16027_);
  or _67314_ (_16029_, _16003_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _67315_ (_16030_, _16029_, _16014_);
  or _67316_ (_16031_, _16011_, _15090_);
  and _67317_ (_16032_, _16031_, _16030_);
  and _67318_ (_16033_, _16013_, _15097_);
  or _67319_ (_41163_, _16033_, _16032_);
  or _67320_ (_16034_, _16011_, _15278_);
  or _67321_ (_16035_, _16003_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _67322_ (_16036_, _16035_, _16014_);
  and _67323_ (_16037_, _16036_, _16034_);
  and _67324_ (_16038_, _16013_, _15285_);
  or _67325_ (_41164_, _16038_, _16037_);
  or _67326_ (_16039_, _16003_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _67327_ (_16040_, _16039_, _16014_);
  or _67328_ (_16041_, _16011_, _15481_);
  and _67329_ (_16042_, _16041_, _16040_);
  and _67330_ (_16043_, _16013_, _15487_);
  or _67331_ (_41165_, _16043_, _16042_);
  and _67332_ (_16044_, _16003_, _09226_);
  or _67333_ (_16045_, _16003_, _07913_);
  nand _67334_ (_16046_, _16045_, _16001_);
  or _67335_ (_16047_, _16046_, _16044_);
  or _67336_ (_16048_, _16014_, _09259_);
  and _67337_ (_41166_, _16048_, _16047_);
  and _67338_ (_16049_, _07766_, _07476_);
  not _67339_ (_16050_, _16049_);
  or _67340_ (_16051_, _16050_, _14332_);
  and _67341_ (_16052_, _15494_, _07749_);
  and _67342_ (_16053_, _16052_, _14324_);
  nor _67343_ (_16054_, _16052_, _07041_);
  or _67344_ (_16055_, _16054_, _16049_);
  or _67345_ (_16056_, _16055_, _16053_);
  and _67346_ (_41169_, _16056_, _16051_);
  and _67347_ (_16057_, _15494_, _16009_);
  not _67348_ (_16058_, _16057_);
  or _67349_ (_16059_, _16058_, _14521_);
  or _67350_ (_16060_, _16057_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _67351_ (_16061_, _16060_, _16050_);
  and _67352_ (_16062_, _16061_, _16059_);
  and _67353_ (_16063_, _16049_, _14527_);
  or _67354_ (_41170_, _16063_, _16062_);
  or _67355_ (_16064_, _16052_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _67356_ (_16065_, _16064_, _16050_);
  or _67357_ (_16066_, _16058_, _14713_);
  and _67358_ (_16067_, _16066_, _16065_);
  and _67359_ (_16068_, _16049_, _14719_);
  or _67360_ (_41171_, _16068_, _16067_);
  or _67361_ (_16069_, _16052_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _67362_ (_16070_, _16069_, _16050_);
  or _67363_ (_16071_, _16058_, _14900_);
  and _67364_ (_16072_, _16071_, _16070_);
  and _67365_ (_16073_, _16049_, _14906_);
  or _67366_ (_41173_, _16073_, _16072_);
  or _67367_ (_16074_, _16052_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _67368_ (_16075_, _16074_, _16050_);
  or _67369_ (_16076_, _16058_, _15090_);
  and _67370_ (_16077_, _16076_, _16075_);
  and _67371_ (_16078_, _16049_, _15097_);
  or _67372_ (_41174_, _16078_, _16077_);
  and _67373_ (_16079_, _16049_, _15285_);
  or _67374_ (_16080_, _16052_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _67375_ (_16081_, _16080_, _16050_);
  or _67376_ (_16082_, _16058_, _15278_);
  and _67377_ (_16083_, _16082_, _16081_);
  or _67378_ (_41175_, _16083_, _16079_);
  or _67379_ (_16084_, _16058_, _15481_);
  or _67380_ (_16085_, _16052_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _67381_ (_16086_, _16085_, _16050_);
  and _67382_ (_16087_, _16086_, _16084_);
  and _67383_ (_16088_, _16049_, _15487_);
  or _67384_ (_41176_, _16088_, _16087_);
  and _67385_ (_16089_, _16049_, _09259_);
  or _67386_ (_16090_, _16052_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _67387_ (_16091_, _16090_, _16050_);
  or _67388_ (_16092_, _16058_, _09226_);
  and _67389_ (_16093_, _16092_, _16091_);
  or _67390_ (_41177_, _16093_, _16089_);
  and _67391_ (_16094_, _15542_, _16009_);
  not _67392_ (_16095_, _16094_);
  or _67393_ (_16096_, _16095_, _14324_);
  and _67394_ (_16097_, _15542_, _07749_);
  or _67395_ (_16098_, _16097_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _67396_ (_16099_, _08449_, _07766_);
  not _67397_ (_16100_, _16099_);
  and _67398_ (_16101_, _16100_, _16098_);
  and _67399_ (_16102_, _16101_, _16096_);
  and _67400_ (_16103_, _16099_, _14332_);
  or _67401_ (_41181_, _16103_, _16102_);
  or _67402_ (_16104_, _16095_, _14521_);
  or _67403_ (_16105_, _16094_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _67404_ (_16106_, _16105_, _16100_);
  and _67405_ (_16107_, _16106_, _16104_);
  and _67406_ (_16108_, _16099_, _14527_);
  or _67407_ (_41182_, _16108_, _16107_);
  or _67408_ (_16109_, _16097_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _67409_ (_16110_, _16109_, _16100_);
  or _67410_ (_16111_, _16095_, _14713_);
  and _67411_ (_16112_, _16111_, _16110_);
  and _67412_ (_16113_, _16099_, _14719_);
  or _67413_ (_41184_, _16113_, _16112_);
  or _67414_ (_16114_, _16097_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _67415_ (_16115_, _16114_, _16100_);
  or _67416_ (_16116_, _16095_, _14900_);
  and _67417_ (_16117_, _16116_, _16115_);
  and _67418_ (_16118_, _16099_, _14906_);
  or _67419_ (_41185_, _16118_, _16117_);
  or _67420_ (_16119_, _16095_, _15090_);
  or _67421_ (_16120_, _16097_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _67422_ (_16121_, _16120_, _16100_);
  and _67423_ (_16122_, _16121_, _16119_);
  and _67424_ (_16123_, _16099_, _15097_);
  or _67425_ (_41186_, _16123_, _16122_);
  or _67426_ (_16124_, _16097_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _67427_ (_16125_, _16124_, _16100_);
  or _67428_ (_16126_, _16095_, _15278_);
  and _67429_ (_16127_, _16126_, _16125_);
  and _67430_ (_16128_, _16099_, _15285_);
  or _67431_ (_41187_, _16128_, _16127_);
  or _67432_ (_16129_, _16097_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _67433_ (_16130_, _16129_, _16100_);
  or _67434_ (_16131_, _16095_, _15481_);
  and _67435_ (_16132_, _16131_, _16130_);
  and _67436_ (_16133_, _16099_, _15487_);
  or _67437_ (_41188_, _16133_, _16132_);
  nor _67438_ (_16134_, _16094_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor _67439_ (_16135_, _16095_, _09226_);
  or _67440_ (_16136_, _16135_, _16134_);
  nand _67441_ (_16137_, _16136_, _16100_);
  or _67442_ (_16138_, _16100_, _09259_);
  and _67443_ (_41190_, _16138_, _16137_);
  not _67444_ (_16139_, _07177_);
  or _67445_ (_16140_, _16000_, _16139_);
  or _67446_ (_16141_, _14332_, _16140_);
  and _67447_ (_16142_, _14324_, _07750_);
  or _67448_ (_16143_, _07750_, _07034_);
  nand _67449_ (_16144_, _16143_, _16140_);
  or _67450_ (_16145_, _16144_, _16142_);
  and _67451_ (_41193_, _16145_, _16141_);
  nor _67452_ (_16146_, _07750_, _07237_);
  and _67453_ (_16147_, _14521_, _07750_);
  or _67454_ (_16148_, _16147_, _16146_);
  and _67455_ (_16149_, _16148_, _16140_);
  and _67456_ (_16150_, _14527_, _07767_);
  or _67457_ (_41194_, _16150_, _16149_);
  or _67458_ (_16151_, _07750_, \oc8051_golden_model_1.IRAM[15] [2]);
  and _67459_ (_16152_, _16151_, _07768_);
  or _67460_ (_16153_, _14713_, _07770_);
  and _67461_ (_16154_, _16153_, _16152_);
  and _67462_ (_16155_, _14719_, _07767_);
  or _67463_ (_41196_, _16155_, _16154_);
  or _67464_ (_16156_, _07750_, \oc8051_golden_model_1.IRAM[15] [3]);
  and _67465_ (_16157_, _16156_, _07768_);
  or _67466_ (_16158_, _14900_, _07770_);
  and _67467_ (_16159_, _16158_, _16157_);
  and _67468_ (_16160_, _14906_, _07767_);
  or _67469_ (_41197_, _16160_, _16159_);
  or _67470_ (_16161_, _07750_, \oc8051_golden_model_1.IRAM[15] [4]);
  and _67471_ (_16162_, _16161_, _07768_);
  or _67472_ (_16163_, _15090_, _07770_);
  and _67473_ (_16164_, _16163_, _16162_);
  and _67474_ (_16165_, _15097_, _07767_);
  or _67475_ (_41198_, _16165_, _16164_);
  or _67476_ (_16166_, _07750_, \oc8051_golden_model_1.IRAM[15] [5]);
  and _67477_ (_16167_, _16166_, _07768_);
  or _67478_ (_16168_, _15278_, _07770_);
  and _67479_ (_16169_, _16168_, _16167_);
  and _67480_ (_16170_, _15285_, _07767_);
  or _67481_ (_41199_, _16170_, _16169_);
  or _67482_ (_16171_, _07750_, \oc8051_golden_model_1.IRAM[15] [6]);
  and _67483_ (_16172_, _16171_, _07768_);
  or _67484_ (_16173_, _15481_, _07770_);
  and _67485_ (_16174_, _16173_, _16172_);
  and _67486_ (_16175_, _15487_, _07767_);
  or _67487_ (_41200_, _16175_, _16174_);
  nor _67488_ (_16176_, _01317_, _09899_);
  nor _67489_ (_16177_, _07841_, _09899_);
  and _67490_ (_16178_, _07841_, _07049_);
  or _67491_ (_16179_, _16178_, _16177_);
  or _67492_ (_16180_, _16179_, _07075_);
  nor _67493_ (_16181_, _08211_, _10243_);
  or _67494_ (_16182_, _16181_, _16177_);
  or _67495_ (_16183_, _16182_, _06161_);
  and _67496_ (_16184_, _07841_, \oc8051_golden_model_1.ACC [0]);
  or _67497_ (_16185_, _16184_, _16177_);
  and _67498_ (_16186_, _16185_, _07056_);
  nor _67499_ (_16187_, _07056_, _09899_);
  or _67500_ (_16188_, _16187_, _06160_);
  or _67501_ (_16189_, _16188_, _16186_);
  and _67502_ (_16190_, _16189_, _06157_);
  and _67503_ (_16191_, _16190_, _16183_);
  nor _67504_ (_16192_, _08420_, _09899_);
  and _67505_ (_16193_, _14169_, _08420_);
  or _67506_ (_16194_, _16193_, _16192_);
  and _67507_ (_16195_, _16194_, _06156_);
  or _67508_ (_16196_, _16195_, _16191_);
  or _67509_ (_16197_, _16196_, _06217_);
  and _67510_ (_16198_, _16197_, _16180_);
  or _67511_ (_16199_, _16198_, _06220_);
  or _67512_ (_16200_, _16185_, _06229_);
  and _67513_ (_16201_, _16200_, _06153_);
  and _67514_ (_16202_, _16201_, _16199_);
  and _67515_ (_16203_, _16177_, _06152_);
  or _67516_ (_16204_, _16203_, _06145_);
  or _67517_ (_16205_, _16204_, _16202_);
  or _67518_ (_16206_, _16182_, _06146_);
  and _67519_ (_16207_, _16206_, _16205_);
  or _67520_ (_16208_, _16207_, _09295_);
  nor _67521_ (_16209_, _09793_, _09790_);
  nor _67522_ (_16210_, _16209_, _09795_);
  or _67523_ (_16211_, _16210_, _09301_);
  and _67524_ (_16212_, _16211_, _06140_);
  and _67525_ (_16213_, _16212_, _16208_);
  or _67526_ (_16214_, _16192_, _14170_);
  and _67527_ (_16215_, _16214_, _06139_);
  and _67528_ (_16216_, _16215_, _16194_);
  or _67529_ (_16217_, _16216_, _09842_);
  or _67530_ (_16218_, _16217_, _16213_);
  or _67531_ (_16219_, _16179_, _06132_);
  and _67532_ (_16220_, _16219_, _06117_);
  and _67533_ (_16221_, _16220_, _16218_);
  and _67534_ (_16222_, _09160_, _07841_);
  or _67535_ (_16223_, _16222_, _16177_);
  and _67536_ (_16224_, _16223_, _06116_);
  or _67537_ (_16225_, _16224_, _05787_);
  or _67538_ (_16226_, _16225_, _16221_);
  and _67539_ (_16227_, _14260_, _07841_);
  or _67540_ (_16228_, _16177_, _06114_);
  or _67541_ (_16229_, _16228_, _16227_);
  and _67542_ (_16230_, _16229_, _09861_);
  and _67543_ (_16231_, _16230_, _16226_);
  nand _67544_ (_16232_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  or _67545_ (_16233_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and _67546_ (_16234_, _16233_, _16232_);
  or _67547_ (_16235_, _10209_, _16234_);
  nand _67548_ (_16236_, _10209_, _05855_);
  and _67549_ (_16237_, _16236_, _09855_);
  and _67550_ (_16238_, _16237_, _16235_);
  or _67551_ (_16239_, _16238_, _11136_);
  or _67552_ (_16240_, _16239_, _16231_);
  and _67553_ (_16241_, _14275_, _07841_);
  or _67554_ (_16242_, _16177_, _07127_);
  or _67555_ (_16243_, _16242_, _16241_);
  and _67556_ (_16244_, _07841_, _08708_);
  or _67557_ (_16245_, _16244_, _16177_);
  or _67558_ (_16246_, _16245_, _06111_);
  and _67559_ (_16247_, _16246_, _07125_);
  and _67560_ (_16248_, _16247_, _16243_);
  and _67561_ (_16249_, _16248_, _16240_);
  nor _67562_ (_16250_, _12321_, _10243_);
  or _67563_ (_16251_, _16250_, _16177_);
  nand _67564_ (_16252_, _10276_, _07841_);
  and _67565_ (_16253_, _16252_, _06402_);
  and _67566_ (_16254_, _16253_, _16251_);
  or _67567_ (_16255_, _16254_, _16249_);
  and _67568_ (_16256_, _16255_, _07132_);
  nand _67569_ (_16257_, _16245_, _06306_);
  nor _67570_ (_16258_, _16257_, _16181_);
  or _67571_ (_16259_, _16258_, _06411_);
  or _67572_ (_16260_, _16259_, _16256_);
  nor _67573_ (_16261_, _16177_, _07130_);
  nand _67574_ (_16262_, _16261_, _16252_);
  and _67575_ (_16263_, _16262_, _16260_);
  or _67576_ (_16264_, _16263_, _06303_);
  and _67577_ (_16265_, _14167_, _07841_);
  or _67578_ (_16266_, _16177_, _08819_);
  or _67579_ (_16267_, _16266_, _16265_);
  and _67580_ (_16268_, _16267_, _08824_);
  and _67581_ (_16269_, _16268_, _16264_);
  and _67582_ (_16270_, _16251_, _06396_);
  or _67583_ (_16271_, _16270_, _06433_);
  or _67584_ (_16272_, _16271_, _16269_);
  or _67585_ (_16273_, _16182_, _06829_);
  and _67586_ (_16274_, _16273_, _16272_);
  or _67587_ (_16275_, _16274_, _05748_);
  or _67588_ (_16276_, _16177_, _05749_);
  and _67589_ (_16277_, _16276_, _16275_);
  or _67590_ (_16278_, _16277_, _06440_);
  or _67591_ (_16279_, _16182_, _06444_);
  and _67592_ (_16280_, _16279_, _01317_);
  and _67593_ (_16281_, _16280_, _16278_);
  or _67594_ (_16282_, _16281_, _16176_);
  and _67595_ (_43594_, _16282_, _43100_);
  nor _67596_ (_16283_, _01317_, _09864_);
  nor _67597_ (_16284_, _07841_, _09864_);
  nor _67598_ (_16285_, _10277_, _10243_);
  or _67599_ (_16286_, _16285_, _16284_);
  or _67600_ (_16287_, _16286_, _08824_);
  nor _67601_ (_16288_, _08420_, _09864_);
  and _67602_ (_16289_, _14349_, _08420_);
  or _67603_ (_16290_, _16289_, _16288_);
  and _67604_ (_16291_, _16290_, _06152_);
  and _67605_ (_16292_, _07841_, _07306_);
  or _67606_ (_16293_, _16292_, _16284_);
  or _67607_ (_16294_, _16293_, _07075_);
  or _67608_ (_16295_, _07841_, \oc8051_golden_model_1.B [1]);
  and _67609_ (_16296_, _14363_, _07841_);
  not _67610_ (_16297_, _16296_);
  and _67611_ (_16298_, _16297_, _16295_);
  or _67612_ (_16299_, _16298_, _06161_);
  and _67613_ (_16300_, _07841_, \oc8051_golden_model_1.ACC [1]);
  or _67614_ (_16301_, _16300_, _16284_);
  and _67615_ (_16302_, _16301_, _07056_);
  nor _67616_ (_16303_, _07056_, _09864_);
  or _67617_ (_16304_, _16303_, _06160_);
  or _67618_ (_16305_, _16304_, _16302_);
  and _67619_ (_16306_, _16305_, _06157_);
  and _67620_ (_16307_, _16306_, _16299_);
  and _67621_ (_16308_, _14367_, _08420_);
  or _67622_ (_16309_, _16308_, _16288_);
  and _67623_ (_16310_, _16309_, _06156_);
  or _67624_ (_16311_, _16310_, _06217_);
  or _67625_ (_16312_, _16311_, _16307_);
  and _67626_ (_16313_, _16312_, _16294_);
  or _67627_ (_16314_, _16313_, _06220_);
  or _67628_ (_16315_, _16301_, _06229_);
  and _67629_ (_16316_, _16315_, _06153_);
  and _67630_ (_16317_, _16316_, _16314_);
  or _67631_ (_16318_, _16317_, _16291_);
  and _67632_ (_16319_, _16318_, _06146_);
  and _67633_ (_16320_, _16308_, _14382_);
  or _67634_ (_16321_, _16320_, _16288_);
  and _67635_ (_16322_, _16321_, _06145_);
  or _67636_ (_16323_, _16322_, _09295_);
  or _67637_ (_16324_, _16323_, _16319_);
  nor _67638_ (_16325_, _09798_, _09737_);
  nor _67639_ (_16326_, _16325_, _09799_);
  or _67640_ (_16327_, _16326_, _09301_);
  and _67641_ (_16328_, _16327_, _06140_);
  and _67642_ (_16329_, _16328_, _16324_);
  and _67643_ (_16330_, _14351_, _08420_);
  or _67644_ (_16331_, _16330_, _16288_);
  and _67645_ (_16332_, _16331_, _06139_);
  or _67646_ (_16333_, _16332_, _09842_);
  or _67647_ (_16334_, _16333_, _16329_);
  or _67648_ (_16335_, _16293_, _06132_);
  and _67649_ (_16336_, _16335_, _16334_);
  or _67650_ (_16337_, _16336_, _06116_);
  and _67651_ (_16338_, _09115_, _07841_);
  or _67652_ (_16339_, _16284_, _06117_);
  or _67653_ (_16340_, _16339_, _16338_);
  and _67654_ (_16341_, _16340_, _06114_);
  and _67655_ (_16342_, _16341_, _16337_);
  or _67656_ (_16343_, _14442_, _10243_);
  and _67657_ (_16344_, _16295_, _05787_);
  and _67658_ (_16345_, _16344_, _16343_);
  or _67659_ (_16346_, _16345_, _09855_);
  or _67660_ (_16347_, _16346_, _16342_);
  and _67661_ (_16348_, _10209_, _10155_);
  nor _67662_ (_16349_, _10204_, _10203_);
  or _67663_ (_16350_, _16349_, _10205_);
  nor _67664_ (_16351_, _16350_, _10209_);
  or _67665_ (_16352_, _16351_, _16348_);
  or _67666_ (_16353_, _16352_, _09861_);
  and _67667_ (_16354_, _16353_, _06111_);
  and _67668_ (_16355_, _16354_, _16347_);
  nand _67669_ (_16356_, _07841_, _06945_);
  and _67670_ (_16357_, _16356_, _06110_);
  and _67671_ (_16358_, _16357_, _16295_);
  or _67672_ (_16359_, _16358_, _16355_);
  and _67673_ (_16360_, _16359_, _07127_);
  or _67674_ (_16361_, _14346_, _10243_);
  and _67675_ (_16362_, _16295_, _06297_);
  and _67676_ (_16363_, _16362_, _16361_);
  or _67677_ (_16364_, _16363_, _06402_);
  or _67678_ (_16365_, _16364_, _16360_);
  and _67679_ (_16366_, _10278_, _07841_);
  or _67680_ (_16367_, _16366_, _16284_);
  or _67681_ (_16368_, _16367_, _07125_);
  and _67682_ (_16369_, _16368_, _07132_);
  and _67683_ (_16370_, _16369_, _16365_);
  or _67684_ (_16371_, _14344_, _10243_);
  and _67685_ (_16372_, _16295_, _06306_);
  and _67686_ (_16373_, _16372_, _16371_);
  or _67687_ (_16374_, _16373_, _06411_);
  or _67688_ (_16375_, _16374_, _16370_);
  and _67689_ (_16376_, _16300_, _08176_);
  or _67690_ (_16377_, _16284_, _07130_);
  or _67691_ (_16378_, _16377_, _16376_);
  and _67692_ (_16379_, _16378_, _08819_);
  and _67693_ (_16380_, _16379_, _16375_);
  or _67694_ (_16381_, _16356_, _08176_);
  and _67695_ (_16382_, _16295_, _06303_);
  and _67696_ (_16383_, _16382_, _16381_);
  or _67697_ (_16384_, _16383_, _06396_);
  or _67698_ (_16385_, _16384_, _16380_);
  and _67699_ (_16386_, _16385_, _16287_);
  or _67700_ (_16387_, _16386_, _06433_);
  or _67701_ (_16388_, _16298_, _06829_);
  and _67702_ (_16389_, _16388_, _05749_);
  and _67703_ (_16390_, _16389_, _16387_);
  and _67704_ (_16391_, _16290_, _05748_);
  or _67705_ (_16392_, _16391_, _06440_);
  or _67706_ (_16393_, _16392_, _16390_);
  or _67707_ (_16394_, _16284_, _06444_);
  or _67708_ (_16395_, _16394_, _16296_);
  and _67709_ (_16396_, _16395_, _01317_);
  and _67710_ (_16397_, _16396_, _16393_);
  or _67711_ (_16398_, _16397_, _16283_);
  and _67712_ (_43595_, _16398_, _43100_);
  nor _67713_ (_16399_, _01317_, _09919_);
  nor _67714_ (_16400_, _07841_, _09919_);
  and _67715_ (_16401_, _07841_, _07708_);
  or _67716_ (_16402_, _16401_, _16400_);
  or _67717_ (_16403_, _16402_, _06132_);
  and _67718_ (_16404_, _14538_, _08420_);
  and _67719_ (_16405_, _16404_, _14569_);
  nor _67720_ (_16406_, _08420_, _09919_);
  or _67721_ (_16407_, _16406_, _06146_);
  or _67722_ (_16408_, _16407_, _16405_);
  or _67723_ (_16409_, _16402_, _07075_);
  and _67724_ (_16410_, _14542_, _07841_);
  or _67725_ (_16411_, _16410_, _16400_);
  or _67726_ (_16412_, _16411_, _06161_);
  and _67727_ (_16413_, _07841_, \oc8051_golden_model_1.ACC [2]);
  or _67728_ (_16414_, _16413_, _16400_);
  and _67729_ (_16415_, _16414_, _07056_);
  nor _67730_ (_16416_, _07056_, _09919_);
  or _67731_ (_16417_, _16416_, _06160_);
  or _67732_ (_16418_, _16417_, _16415_);
  and _67733_ (_16419_, _16418_, _06157_);
  and _67734_ (_16420_, _16419_, _16412_);
  or _67735_ (_16421_, _16406_, _16404_);
  and _67736_ (_16422_, _16421_, _06156_);
  or _67737_ (_16423_, _16422_, _06217_);
  or _67738_ (_16424_, _16423_, _16420_);
  and _67739_ (_16425_, _16424_, _16409_);
  or _67740_ (_16426_, _16425_, _06220_);
  or _67741_ (_16427_, _16414_, _06229_);
  and _67742_ (_16428_, _16427_, _06153_);
  and _67743_ (_16429_, _16428_, _16426_);
  and _67744_ (_16430_, _14536_, _08420_);
  or _67745_ (_16431_, _16430_, _16406_);
  and _67746_ (_16432_, _16431_, _06152_);
  or _67747_ (_16433_, _16432_, _06145_);
  or _67748_ (_16434_, _16433_, _16429_);
  and _67749_ (_16435_, _16434_, _16408_);
  or _67750_ (_16436_, _16435_, _09295_);
  or _67751_ (_16437_, _09801_, _09679_);
  and _67752_ (_16438_, _16437_, _09802_);
  or _67753_ (_16439_, _16438_, _09301_);
  and _67754_ (_16440_, _16439_, _06140_);
  and _67755_ (_16441_, _16440_, _16436_);
  and _67756_ (_16442_, _14583_, _08420_);
  or _67757_ (_16443_, _16442_, _16406_);
  and _67758_ (_16444_, _16443_, _06139_);
  or _67759_ (_16445_, _16444_, _09842_);
  or _67760_ (_16446_, _16445_, _16441_);
  and _67761_ (_16447_, _16446_, _16403_);
  or _67762_ (_16448_, _16447_, _06116_);
  and _67763_ (_16449_, _09211_, _07841_);
  or _67764_ (_16450_, _16400_, _06117_);
  or _67765_ (_16451_, _16450_, _16449_);
  and _67766_ (_16452_, _16451_, _16448_);
  or _67767_ (_16453_, _16452_, _05787_);
  and _67768_ (_16454_, _14630_, _07841_);
  or _67769_ (_16455_, _16400_, _06114_);
  or _67770_ (_16456_, _16455_, _16454_);
  and _67771_ (_16457_, _16456_, _09861_);
  and _67772_ (_16458_, _16457_, _16453_);
  nor _67773_ (_16459_, _10205_, _10156_);
  not _67774_ (_16460_, _16459_);
  and _67775_ (_16461_, _16460_, _10149_);
  nor _67776_ (_16462_, _16460_, _10149_);
  nor _67777_ (_16463_, _16462_, _16461_);
  or _67778_ (_16464_, _16463_, _10209_);
  nand _67779_ (_16465_, _10209_, _10146_);
  and _67780_ (_16466_, _16465_, _09855_);
  and _67781_ (_16467_, _16466_, _16464_);
  or _67782_ (_16468_, _16467_, _11136_);
  or _67783_ (_16469_, _16468_, _16458_);
  and _67784_ (_16470_, _14646_, _07841_);
  or _67785_ (_16471_, _16400_, _07127_);
  or _67786_ (_16472_, _16471_, _16470_);
  and _67787_ (_16473_, _07841_, _08768_);
  or _67788_ (_16474_, _16473_, _16400_);
  or _67789_ (_16475_, _16474_, _06111_);
  and _67790_ (_16476_, _16475_, _07125_);
  and _67791_ (_16477_, _16476_, _16472_);
  and _67792_ (_16478_, _16477_, _16469_);
  and _67793_ (_16479_, _10282_, _07841_);
  or _67794_ (_16480_, _16479_, _16400_);
  and _67795_ (_16481_, _16480_, _06402_);
  or _67796_ (_16482_, _16481_, _16478_);
  and _67797_ (_16483_, _16482_, _07132_);
  or _67798_ (_16484_, _16400_, _08248_);
  and _67799_ (_16485_, _16474_, _06306_);
  and _67800_ (_16486_, _16485_, _16484_);
  or _67801_ (_16487_, _16486_, _16483_);
  and _67802_ (_16488_, _16487_, _07130_);
  and _67803_ (_16489_, _16414_, _06411_);
  and _67804_ (_16490_, _16489_, _16484_);
  or _67805_ (_16491_, _16490_, _06303_);
  or _67806_ (_16492_, _16491_, _16488_);
  and _67807_ (_16493_, _14643_, _07841_);
  or _67808_ (_16494_, _16400_, _08819_);
  or _67809_ (_16495_, _16494_, _16493_);
  and _67810_ (_16496_, _16495_, _08824_);
  and _67811_ (_16497_, _16496_, _16492_);
  nor _67812_ (_16498_, _10281_, _10243_);
  or _67813_ (_16499_, _16498_, _16400_);
  and _67814_ (_16500_, _16499_, _06396_);
  or _67815_ (_16501_, _16500_, _06433_);
  or _67816_ (_16502_, _16501_, _16497_);
  or _67817_ (_16503_, _16411_, _06829_);
  and _67818_ (_16504_, _16503_, _05749_);
  and _67819_ (_16505_, _16504_, _16502_);
  and _67820_ (_16506_, _16431_, _05748_);
  or _67821_ (_16507_, _16506_, _06440_);
  or _67822_ (_16508_, _16507_, _16505_);
  and _67823_ (_16509_, _14710_, _07841_);
  or _67824_ (_16510_, _16400_, _06444_);
  or _67825_ (_16511_, _16510_, _16509_);
  and _67826_ (_16512_, _16511_, _01317_);
  and _67827_ (_16513_, _16512_, _16508_);
  or _67828_ (_16514_, _16513_, _16399_);
  and _67829_ (_43596_, _16514_, _43100_);
  nor _67830_ (_16515_, _01317_, _09951_);
  nor _67831_ (_16516_, _07841_, _09951_);
  and _67832_ (_16517_, _14825_, _07841_);
  or _67833_ (_16518_, _16517_, _16516_);
  and _67834_ (_16519_, _16518_, _05787_);
  nor _67835_ (_16520_, _08420_, _09951_);
  and _67836_ (_16521_, _14735_, _08420_);
  or _67837_ (_16522_, _16521_, _16520_);
  or _67838_ (_16523_, _16520_, _14764_);
  and _67839_ (_16524_, _16523_, _16522_);
  or _67840_ (_16525_, _16524_, _06146_);
  and _67841_ (_16526_, _14738_, _07841_);
  or _67842_ (_16527_, _16526_, _16516_);
  or _67843_ (_16528_, _16527_, _06161_);
  and _67844_ (_16529_, _07841_, \oc8051_golden_model_1.ACC [3]);
  or _67845_ (_16530_, _16529_, _16516_);
  and _67846_ (_16531_, _16530_, _07056_);
  nor _67847_ (_16532_, _07056_, _09951_);
  or _67848_ (_16533_, _16532_, _06160_);
  or _67849_ (_16534_, _16533_, _16531_);
  and _67850_ (_16535_, _16534_, _06157_);
  and _67851_ (_16536_, _16535_, _16528_);
  and _67852_ (_16537_, _16522_, _06156_);
  or _67853_ (_16538_, _16537_, _06217_);
  or _67854_ (_16539_, _16538_, _16536_);
  and _67855_ (_16540_, _07841_, _07544_);
  or _67856_ (_16541_, _16540_, _16516_);
  or _67857_ (_16542_, _16541_, _07075_);
  and _67858_ (_16543_, _16542_, _16539_);
  or _67859_ (_16544_, _16543_, _06220_);
  or _67860_ (_16545_, _16530_, _06229_);
  and _67861_ (_16546_, _16545_, _06153_);
  and _67862_ (_16547_, _16546_, _16544_);
  and _67863_ (_16548_, _14731_, _08420_);
  or _67864_ (_16549_, _16548_, _16520_);
  and _67865_ (_16550_, _16549_, _06152_);
  or _67866_ (_16551_, _16550_, _06145_);
  or _67867_ (_16552_, _16551_, _16547_);
  and _67868_ (_16553_, _16552_, _16525_);
  or _67869_ (_16554_, _16553_, _09295_);
  nor _67870_ (_16555_, _09805_, _09621_);
  nor _67871_ (_16556_, _16555_, _09807_);
  or _67872_ (_16557_, _16556_, _09301_);
  and _67873_ (_16558_, _16557_, _06140_);
  and _67874_ (_16559_, _16558_, _16554_);
  and _67875_ (_16560_, _14732_, _08420_);
  or _67876_ (_16561_, _16560_, _16520_);
  and _67877_ (_16562_, _16561_, _06139_);
  or _67878_ (_16563_, _16562_, _09842_);
  or _67879_ (_16564_, _16563_, _16559_);
  or _67880_ (_16565_, _16541_, _06132_);
  and _67881_ (_16566_, _16565_, _16564_);
  or _67882_ (_16567_, _16566_, _06116_);
  and _67883_ (_16568_, _09210_, _07841_);
  or _67884_ (_16569_, _16516_, _06117_);
  or _67885_ (_16570_, _16569_, _16568_);
  and _67886_ (_16571_, _16570_, _06114_);
  and _67887_ (_16572_, _16571_, _16567_);
  or _67888_ (_16573_, _16572_, _16519_);
  and _67889_ (_16574_, _16573_, _09861_);
  nor _67890_ (_16575_, _16461_, _10148_);
  nor _67891_ (_16576_, _16575_, _10140_);
  and _67892_ (_16577_, _16575_, _10140_);
  or _67893_ (_16578_, _16577_, _16576_);
  or _67894_ (_16579_, _16578_, _10209_);
  not _67895_ (_16580_, _10209_);
  or _67896_ (_16581_, _16580_, _10137_);
  and _67897_ (_16582_, _16581_, _09855_);
  and _67898_ (_16583_, _16582_, _16579_);
  or _67899_ (_16584_, _16583_, _11136_);
  or _67900_ (_16585_, _16584_, _16574_);
  and _67901_ (_16586_, _14727_, _07841_);
  or _67902_ (_16587_, _16516_, _07127_);
  or _67903_ (_16588_, _16587_, _16586_);
  and _67904_ (_16589_, _07841_, _08712_);
  or _67905_ (_16590_, _16589_, _16516_);
  or _67906_ (_16591_, _16590_, _06111_);
  and _67907_ (_16592_, _16591_, _07125_);
  and _67908_ (_16593_, _16592_, _16588_);
  and _67909_ (_16594_, _16593_, _16585_);
  and _67910_ (_16595_, _12318_, _07841_);
  or _67911_ (_16596_, _16595_, _16516_);
  and _67912_ (_16597_, _16596_, _06402_);
  or _67913_ (_16598_, _16597_, _16594_);
  and _67914_ (_16599_, _16598_, _07132_);
  or _67915_ (_16600_, _16516_, _08140_);
  and _67916_ (_16601_, _16590_, _06306_);
  and _67917_ (_16602_, _16601_, _16600_);
  or _67918_ (_16603_, _16602_, _16599_);
  and _67919_ (_16604_, _16603_, _07130_);
  and _67920_ (_16605_, _16530_, _06411_);
  and _67921_ (_16606_, _16605_, _16600_);
  or _67922_ (_16607_, _16606_, _06303_);
  or _67923_ (_16608_, _16607_, _16604_);
  and _67924_ (_16609_, _14724_, _07841_);
  or _67925_ (_16610_, _16516_, _08819_);
  or _67926_ (_16611_, _16610_, _16609_);
  and _67927_ (_16612_, _16611_, _08824_);
  and _67928_ (_16613_, _16612_, _16608_);
  nor _67929_ (_16614_, _10273_, _10243_);
  or _67930_ (_16615_, _16614_, _16516_);
  and _67931_ (_16616_, _16615_, _06396_);
  or _67932_ (_16617_, _16616_, _06433_);
  or _67933_ (_16618_, _16617_, _16613_);
  or _67934_ (_16619_, _16527_, _06829_);
  and _67935_ (_16620_, _16619_, _05749_);
  and _67936_ (_16621_, _16620_, _16618_);
  and _67937_ (_16622_, _16549_, _05748_);
  or _67938_ (_16623_, _16622_, _06440_);
  or _67939_ (_16624_, _16623_, _16621_);
  and _67940_ (_16625_, _14897_, _07841_);
  or _67941_ (_16626_, _16516_, _06444_);
  or _67942_ (_16627_, _16626_, _16625_);
  and _67943_ (_16628_, _16627_, _01317_);
  and _67944_ (_16629_, _16628_, _16624_);
  or _67945_ (_16630_, _16629_, _16515_);
  and _67946_ (_43598_, _16630_, _43100_);
  nor _67947_ (_16631_, _01317_, _09876_);
  nor _67948_ (_16632_, _07841_, _09876_);
  and _67949_ (_16633_, _15013_, _07841_);
  or _67950_ (_16634_, _16633_, _16632_);
  and _67951_ (_16635_, _16634_, _05787_);
  and _67952_ (_16636_, _08336_, _07841_);
  or _67953_ (_16637_, _16636_, _16632_);
  or _67954_ (_16638_, _16637_, _06132_);
  nor _67955_ (_16639_, _08420_, _09876_);
  and _67956_ (_16640_, _14942_, _08420_);
  or _67957_ (_16641_, _16640_, _16639_);
  and _67958_ (_16642_, _16641_, _06152_);
  and _67959_ (_16643_, _14928_, _07841_);
  or _67960_ (_16644_, _16643_, _16632_);
  or _67961_ (_16645_, _16644_, _06161_);
  and _67962_ (_16646_, _07841_, \oc8051_golden_model_1.ACC [4]);
  or _67963_ (_16647_, _16646_, _16632_);
  and _67964_ (_16648_, _16647_, _07056_);
  nor _67965_ (_16649_, _07056_, _09876_);
  or _67966_ (_16650_, _16649_, _06160_);
  or _67967_ (_16651_, _16650_, _16648_);
  and _67968_ (_16652_, _16651_, _06157_);
  and _67969_ (_16653_, _16652_, _16645_);
  and _67970_ (_16654_, _14932_, _08420_);
  or _67971_ (_16655_, _16654_, _16639_);
  and _67972_ (_16656_, _16655_, _06156_);
  or _67973_ (_16657_, _16656_, _06217_);
  or _67974_ (_16658_, _16657_, _16653_);
  or _67975_ (_16659_, _16637_, _07075_);
  and _67976_ (_16660_, _16659_, _16658_);
  or _67977_ (_16661_, _16660_, _06220_);
  or _67978_ (_16662_, _16647_, _06229_);
  and _67979_ (_16663_, _16662_, _06153_);
  and _67980_ (_16664_, _16663_, _16661_);
  or _67981_ (_16665_, _16664_, _16642_);
  and _67982_ (_16666_, _16665_, _06146_);
  or _67983_ (_16667_, _16639_, _14949_);
  and _67984_ (_16668_, _16655_, _06145_);
  and _67985_ (_16669_, _16668_, _16667_);
  or _67986_ (_16670_, _16669_, _09295_);
  or _67987_ (_16671_, _16670_, _16666_);
  or _67988_ (_16672_, _09811_, _09808_);
  and _67989_ (_16673_, _16672_, _09813_);
  or _67990_ (_16674_, _16673_, _09301_);
  and _67991_ (_16675_, _16674_, _06140_);
  and _67992_ (_16676_, _16675_, _16671_);
  and _67993_ (_16677_, _14966_, _08420_);
  or _67994_ (_16678_, _16677_, _16639_);
  and _67995_ (_16679_, _16678_, _06139_);
  or _67996_ (_16680_, _16679_, _09842_);
  or _67997_ (_16681_, _16680_, _16676_);
  and _67998_ (_16682_, _16681_, _16638_);
  or _67999_ (_16683_, _16682_, _06116_);
  and _68000_ (_16684_, _09209_, _07841_);
  or _68001_ (_16685_, _16632_, _06117_);
  or _68002_ (_16686_, _16685_, _16684_);
  and _68003_ (_16687_, _16686_, _06114_);
  and _68004_ (_16688_, _16687_, _16683_);
  or _68005_ (_16689_, _16688_, _16635_);
  and _68006_ (_16690_, _16689_, _09861_);
  or _68007_ (_16691_, _16580_, _10175_);
  nor _68008_ (_16692_, _16575_, _10139_);
  or _68009_ (_16693_, _16692_, _10138_);
  nand _68010_ (_16694_, _16693_, _10178_);
  or _68011_ (_16695_, _16693_, _10178_);
  and _68012_ (_16696_, _16695_, _16694_);
  or _68013_ (_16697_, _16696_, _10209_);
  and _68014_ (_16698_, _16697_, _09855_);
  and _68015_ (_16699_, _16698_, _16691_);
  or _68016_ (_16700_, _16699_, _11136_);
  or _68017_ (_16701_, _16700_, _16690_);
  and _68018_ (_16702_, _15029_, _07841_);
  or _68019_ (_16703_, _16632_, _07127_);
  or _68020_ (_16704_, _16703_, _16702_);
  and _68021_ (_16705_, _08715_, _07841_);
  or _68022_ (_16706_, _16705_, _16632_);
  or _68023_ (_16707_, _16706_, _06111_);
  and _68024_ (_16708_, _16707_, _07125_);
  and _68025_ (_16709_, _16708_, _16704_);
  and _68026_ (_16710_, _16709_, _16701_);
  and _68027_ (_16711_, _10289_, _07841_);
  or _68028_ (_16712_, _16711_, _16632_);
  and _68029_ (_16713_, _16712_, _06402_);
  or _68030_ (_16714_, _16713_, _16710_);
  and _68031_ (_16715_, _16714_, _07132_);
  or _68032_ (_16716_, _16632_, _08339_);
  and _68033_ (_16717_, _16706_, _06306_);
  and _68034_ (_16718_, _16717_, _16716_);
  or _68035_ (_16719_, _16718_, _16715_);
  and _68036_ (_16720_, _16719_, _07130_);
  and _68037_ (_16721_, _16647_, _06411_);
  and _68038_ (_16722_, _16721_, _16716_);
  or _68039_ (_16723_, _16722_, _06303_);
  or _68040_ (_16724_, _16723_, _16720_);
  and _68041_ (_16725_, _15026_, _07841_);
  or _68042_ (_16726_, _16632_, _08819_);
  or _68043_ (_16727_, _16726_, _16725_);
  and _68044_ (_16728_, _16727_, _08824_);
  and _68045_ (_16729_, _16728_, _16724_);
  nor _68046_ (_16730_, _10288_, _10243_);
  or _68047_ (_16731_, _16730_, _16632_);
  and _68048_ (_16732_, _16731_, _06396_);
  or _68049_ (_16733_, _16732_, _06433_);
  or _68050_ (_16734_, _16733_, _16729_);
  or _68051_ (_16735_, _16644_, _06829_);
  and _68052_ (_16736_, _16735_, _05749_);
  and _68053_ (_16737_, _16736_, _16734_);
  and _68054_ (_16738_, _16641_, _05748_);
  or _68055_ (_16739_, _16738_, _06440_);
  or _68056_ (_16740_, _16739_, _16737_);
  and _68057_ (_16741_, _15087_, _07841_);
  or _68058_ (_16742_, _16632_, _06444_);
  or _68059_ (_16743_, _16742_, _16741_);
  and _68060_ (_16744_, _16743_, _01317_);
  and _68061_ (_16745_, _16744_, _16740_);
  or _68062_ (_16746_, _16745_, _16631_);
  and _68063_ (_43599_, _16746_, _43100_);
  nor _68064_ (_16747_, _01317_, _09877_);
  nor _68065_ (_16748_, _07841_, _09877_);
  and _68066_ (_16749_, _15203_, _07841_);
  or _68067_ (_16750_, _16749_, _16748_);
  and _68068_ (_16751_, _16750_, _05787_);
  and _68069_ (_16752_, _08101_, _07841_);
  or _68070_ (_16753_, _16752_, _16748_);
  or _68071_ (_16754_, _16753_, _06132_);
  nor _68072_ (_16755_, _08420_, _09877_);
  and _68073_ (_16756_, _15104_, _08420_);
  or _68074_ (_16757_, _16756_, _16755_);
  and _68075_ (_16758_, _16757_, _06152_);
  and _68076_ (_16759_, _15119_, _07841_);
  or _68077_ (_16760_, _16759_, _16748_);
  or _68078_ (_16761_, _16760_, _06161_);
  and _68079_ (_16762_, _07841_, \oc8051_golden_model_1.ACC [5]);
  or _68080_ (_16763_, _16762_, _16748_);
  and _68081_ (_16764_, _16763_, _07056_);
  nor _68082_ (_16765_, _07056_, _09877_);
  or _68083_ (_16766_, _16765_, _06160_);
  or _68084_ (_16767_, _16766_, _16764_);
  and _68085_ (_16768_, _16767_, _06157_);
  and _68086_ (_16769_, _16768_, _16761_);
  and _68087_ (_16770_, _15123_, _08420_);
  or _68088_ (_16771_, _16770_, _16755_);
  and _68089_ (_16772_, _16771_, _06156_);
  or _68090_ (_16773_, _16772_, _06217_);
  or _68091_ (_16774_, _16773_, _16769_);
  or _68092_ (_16775_, _16753_, _07075_);
  and _68093_ (_16776_, _16775_, _16774_);
  or _68094_ (_16777_, _16776_, _06220_);
  or _68095_ (_16778_, _16763_, _06229_);
  and _68096_ (_16779_, _16778_, _06153_);
  and _68097_ (_16780_, _16779_, _16777_);
  or _68098_ (_16781_, _16780_, _16758_);
  and _68099_ (_16782_, _16781_, _06146_);
  or _68100_ (_16783_, _16755_, _15138_);
  and _68101_ (_16784_, _16771_, _06145_);
  and _68102_ (_16785_, _16784_, _16783_);
  or _68103_ (_16786_, _16785_, _09295_);
  or _68104_ (_16787_, _16786_, _16782_);
  or _68105_ (_16788_, _09492_, _09493_);
  and _68106_ (_16789_, _16788_, _09814_);
  nor _68107_ (_16790_, _16789_, _09816_);
  or _68108_ (_16791_, _16790_, _09301_);
  and _68109_ (_16792_, _16791_, _06140_);
  and _68110_ (_16793_, _16792_, _16787_);
  and _68111_ (_16794_, _15155_, _08420_);
  or _68112_ (_16795_, _16794_, _16755_);
  and _68113_ (_16796_, _16795_, _06139_);
  or _68114_ (_16797_, _16796_, _09842_);
  or _68115_ (_16798_, _16797_, _16793_);
  and _68116_ (_16799_, _16798_, _16754_);
  or _68117_ (_16800_, _16799_, _06116_);
  and _68118_ (_16801_, _09208_, _07841_);
  or _68119_ (_16802_, _16748_, _06117_);
  or _68120_ (_16803_, _16802_, _16801_);
  and _68121_ (_16804_, _16803_, _06114_);
  and _68122_ (_16805_, _16804_, _16800_);
  or _68123_ (_16806_, _16805_, _16751_);
  and _68124_ (_16807_, _16806_, _09861_);
  not _68125_ (_16808_, _10177_);
  and _68126_ (_16809_, _16694_, _16808_);
  nor _68127_ (_16810_, _16809_, _10189_);
  and _68128_ (_16811_, _16809_, _10189_);
  or _68129_ (_16812_, _16811_, _16810_);
  nor _68130_ (_16813_, _10209_, _09861_);
  and _68131_ (_16814_, _16813_, _16812_);
  and _68132_ (_16815_, _10186_, _09855_);
  and _68133_ (_16816_, _16815_, _10209_);
  or _68134_ (_16817_, _16816_, _11136_);
  or _68135_ (_16818_, _16817_, _16814_);
  or _68136_ (_16819_, _16818_, _16807_);
  and _68137_ (_16820_, _15219_, _07841_);
  or _68138_ (_16821_, _16748_, _07127_);
  or _68139_ (_16822_, _16821_, _16820_);
  and _68140_ (_16823_, _08736_, _07841_);
  or _68141_ (_16824_, _16823_, _16748_);
  or _68142_ (_16825_, _16824_, _06111_);
  and _68143_ (_16826_, _16825_, _07125_);
  and _68144_ (_16827_, _16826_, _16822_);
  and _68145_ (_16828_, _16827_, _16819_);
  and _68146_ (_16829_, _12325_, _07841_);
  or _68147_ (_16830_, _16829_, _16748_);
  and _68148_ (_16831_, _16830_, _06402_);
  or _68149_ (_16832_, _16831_, _16828_);
  and _68150_ (_16833_, _16832_, _07132_);
  or _68151_ (_16834_, _16748_, _08104_);
  and _68152_ (_16835_, _16824_, _06306_);
  and _68153_ (_16836_, _16835_, _16834_);
  or _68154_ (_16837_, _16836_, _16833_);
  and _68155_ (_16838_, _16837_, _07130_);
  and _68156_ (_16839_, _16763_, _06411_);
  and _68157_ (_16840_, _16839_, _16834_);
  or _68158_ (_16841_, _16840_, _06303_);
  or _68159_ (_16842_, _16841_, _16838_);
  and _68160_ (_16843_, _15216_, _07841_);
  or _68161_ (_16844_, _16748_, _08819_);
  or _68162_ (_16845_, _16844_, _16843_);
  and _68163_ (_16846_, _16845_, _08824_);
  and _68164_ (_16847_, _16846_, _16842_);
  nor _68165_ (_16848_, _10269_, _10243_);
  or _68166_ (_16849_, _16848_, _16748_);
  and _68167_ (_16850_, _16849_, _06396_);
  or _68168_ (_16851_, _16850_, _06433_);
  or _68169_ (_16852_, _16851_, _16847_);
  or _68170_ (_16853_, _16760_, _06829_);
  and _68171_ (_16854_, _16853_, _05749_);
  and _68172_ (_16855_, _16854_, _16852_);
  and _68173_ (_16856_, _16757_, _05748_);
  or _68174_ (_16857_, _16856_, _06440_);
  or _68175_ (_16858_, _16857_, _16855_);
  and _68176_ (_16859_, _15275_, _07841_);
  or _68177_ (_16860_, _16748_, _06444_);
  or _68178_ (_16861_, _16860_, _16859_);
  and _68179_ (_16862_, _16861_, _01317_);
  and _68180_ (_16863_, _16862_, _16858_);
  or _68181_ (_16864_, _16863_, _16747_);
  and _68182_ (_43600_, _16864_, _43100_);
  nor _68183_ (_16865_, _01317_, _10120_);
  nor _68184_ (_16866_, _07841_, _10120_);
  and _68185_ (_16867_, _15395_, _07841_);
  or _68186_ (_16868_, _16867_, _16866_);
  and _68187_ (_16869_, _16868_, _05787_);
  and _68188_ (_16870_, _08012_, _07841_);
  or _68189_ (_16871_, _16870_, _16866_);
  or _68190_ (_16872_, _16871_, _06132_);
  nor _68191_ (_16873_, _08420_, _10120_);
  and _68192_ (_16874_, _15297_, _08420_);
  or _68193_ (_16875_, _16874_, _16873_);
  and _68194_ (_16876_, _16875_, _06152_);
  and _68195_ (_16877_, _15300_, _07841_);
  or _68196_ (_16878_, _16877_, _16866_);
  or _68197_ (_16879_, _16878_, _06161_);
  and _68198_ (_16880_, _07841_, \oc8051_golden_model_1.ACC [6]);
  or _68199_ (_16881_, _16880_, _16866_);
  and _68200_ (_16882_, _16881_, _07056_);
  nor _68201_ (_16883_, _07056_, _10120_);
  or _68202_ (_16884_, _16883_, _06160_);
  or _68203_ (_16885_, _16884_, _16882_);
  and _68204_ (_16886_, _16885_, _06157_);
  and _68205_ (_16887_, _16886_, _16879_);
  and _68206_ (_16888_, _15316_, _08420_);
  or _68207_ (_16889_, _16888_, _16873_);
  and _68208_ (_16890_, _16889_, _06156_);
  or _68209_ (_16891_, _16890_, _06217_);
  or _68210_ (_16892_, _16891_, _16887_);
  or _68211_ (_16893_, _16871_, _07075_);
  and _68212_ (_16894_, _16893_, _16892_);
  or _68213_ (_16895_, _16894_, _06220_);
  or _68214_ (_16896_, _16881_, _06229_);
  and _68215_ (_16897_, _16896_, _06153_);
  and _68216_ (_16898_, _16897_, _16895_);
  or _68217_ (_16899_, _16898_, _16876_);
  and _68218_ (_16900_, _16899_, _06146_);
  or _68219_ (_16901_, _16873_, _15331_);
  and _68220_ (_16902_, _16889_, _06145_);
  and _68221_ (_16903_, _16902_, _16901_);
  or _68222_ (_16904_, _16903_, _09295_);
  or _68223_ (_16905_, _16904_, _16900_);
  nor _68224_ (_16906_, _09834_, _09817_);
  nor _68225_ (_16907_, _16906_, _09835_);
  or _68226_ (_16908_, _16907_, _09301_);
  and _68227_ (_16909_, _16908_, _06140_);
  and _68228_ (_16910_, _16909_, _16905_);
  and _68229_ (_16911_, _15348_, _08420_);
  or _68230_ (_16912_, _16911_, _16873_);
  and _68231_ (_16913_, _16912_, _06139_);
  or _68232_ (_16914_, _16913_, _09842_);
  or _68233_ (_16915_, _16914_, _16910_);
  and _68234_ (_16916_, _16915_, _16872_);
  or _68235_ (_16917_, _16916_, _06116_);
  and _68236_ (_16918_, _09207_, _07841_);
  or _68237_ (_16919_, _16866_, _06117_);
  or _68238_ (_16920_, _16919_, _16918_);
  and _68239_ (_16921_, _16920_, _06114_);
  and _68240_ (_16922_, _16921_, _16917_);
  or _68241_ (_16923_, _16922_, _16869_);
  and _68242_ (_16924_, _16923_, _09861_);
  nor _68243_ (_16925_, _16809_, _10187_);
  or _68244_ (_16926_, _16925_, _10188_);
  and _68245_ (_16927_, _16926_, _10169_);
  nor _68246_ (_16928_, _16926_, _10169_);
  or _68247_ (_16929_, _16928_, _16927_);
  or _68248_ (_16930_, _16929_, _10209_);
  or _68249_ (_16931_, _16580_, _10126_);
  and _68250_ (_16932_, _16931_, _09855_);
  and _68251_ (_16933_, _16932_, _16930_);
  or _68252_ (_16934_, _16933_, _11136_);
  or _68253_ (_16935_, _16934_, _16924_);
  and _68254_ (_16936_, _15413_, _07841_);
  or _68255_ (_16937_, _16866_, _07127_);
  or _68256_ (_16938_, _16937_, _16936_);
  and _68257_ (_16939_, _15402_, _07841_);
  or _68258_ (_16940_, _16939_, _16866_);
  or _68259_ (_16941_, _16940_, _06111_);
  and _68260_ (_16942_, _16941_, _07125_);
  and _68261_ (_16943_, _16942_, _16938_);
  and _68262_ (_16944_, _16943_, _16935_);
  and _68263_ (_16945_, _10295_, _07841_);
  or _68264_ (_16946_, _16945_, _16866_);
  and _68265_ (_16947_, _16946_, _06402_);
  or _68266_ (_16948_, _16947_, _16944_);
  and _68267_ (_16949_, _16948_, _07132_);
  or _68268_ (_16950_, _16866_, _08015_);
  and _68269_ (_16951_, _16940_, _06306_);
  and _68270_ (_16952_, _16951_, _16950_);
  or _68271_ (_16953_, _16952_, _16949_);
  and _68272_ (_16954_, _16953_, _07130_);
  and _68273_ (_16955_, _16881_, _06411_);
  and _68274_ (_16956_, _16955_, _16950_);
  or _68275_ (_16957_, _16956_, _06303_);
  or _68276_ (_16958_, _16957_, _16954_);
  and _68277_ (_16959_, _15410_, _07841_);
  or _68278_ (_16960_, _16866_, _08819_);
  or _68279_ (_16961_, _16960_, _16959_);
  and _68280_ (_16962_, _16961_, _08824_);
  and _68281_ (_16963_, _16962_, _16958_);
  nor _68282_ (_16964_, _10294_, _10243_);
  or _68283_ (_16965_, _16964_, _16866_);
  and _68284_ (_16966_, _16965_, _06396_);
  or _68285_ (_16967_, _16966_, _06433_);
  or _68286_ (_16968_, _16967_, _16963_);
  or _68287_ (_16969_, _16878_, _06829_);
  and _68288_ (_16970_, _16969_, _05749_);
  and _68289_ (_16971_, _16970_, _16968_);
  and _68290_ (_16972_, _16875_, _05748_);
  or _68291_ (_16973_, _16972_, _06440_);
  or _68292_ (_16974_, _16973_, _16971_);
  and _68293_ (_16975_, _15478_, _07841_);
  or _68294_ (_16976_, _16866_, _06444_);
  or _68295_ (_16977_, _16976_, _16975_);
  and _68296_ (_16978_, _16977_, _01317_);
  and _68297_ (_16979_, _16978_, _16974_);
  or _68298_ (_16980_, _16979_, _16865_);
  and _68299_ (_43601_, _16980_, _43100_);
  nor _68300_ (_16981_, _01317_, _05855_);
  nand _68301_ (_16982_, _10262_, _08430_);
  nand _68302_ (_16983_, _12322_, _06169_);
  and _68303_ (_16984_, _16983_, _10265_);
  nor _68304_ (_16985_, _07049_, \oc8051_golden_model_1.ACC [0]);
  nor _68305_ (_16986_, _10985_, _16985_);
  not _68306_ (_16987_, _10962_);
  and _68307_ (_16988_, _16987_, _16986_);
  and _68308_ (_16989_, _14167_, _07809_);
  nor _68309_ (_16990_, _07809_, _05855_);
  or _68310_ (_16991_, _16990_, _08819_);
  or _68311_ (_16992_, _16991_, _16989_);
  nor _68312_ (_16993_, _09160_, \oc8051_golden_model_1.ACC [0]);
  nand _68313_ (_16994_, _10841_, _16993_);
  and _68314_ (_16995_, _14275_, _07809_);
  or _68315_ (_16996_, _16990_, _07127_);
  or _68316_ (_16997_, _16996_, _16995_);
  nand _68317_ (_16998_, _06107_, _05801_);
  and _68318_ (_16999_, _14260_, _07809_);
  or _68319_ (_17000_, _16999_, _16990_);
  and _68320_ (_17001_, _17000_, _05787_);
  and _68321_ (_17002_, _07809_, _07049_);
  or _68322_ (_17003_, _17002_, _16990_);
  or _68323_ (_17004_, _17003_, _06132_);
  nor _68324_ (_17005_, _10627_, _05855_);
  or _68325_ (_17006_, _17005_, _10628_);
  or _68326_ (_17007_, _17006_, _12380_);
  or _68327_ (_17008_, _10458_, _07049_);
  nor _68328_ (_17009_, _10473_, _07064_);
  or _68329_ (_17010_, _17009_, _09160_);
  not _68330_ (_17011_, _10471_);
  and _68331_ (_17012_, _17011_, _07049_);
  or _68332_ (_17013_, _06653_, \oc8051_golden_model_1.ACC [0]);
  nand _68333_ (_17014_, _06653_, \oc8051_golden_model_1.ACC [0]);
  and _68334_ (_17015_, _17014_, _17013_);
  and _68335_ (_17016_, _17015_, _10471_);
  or _68336_ (_17017_, _17016_, _10473_);
  or _68337_ (_17018_, _17017_, _17012_);
  and _68338_ (_17019_, _17018_, _05772_);
  or _68339_ (_17020_, _17019_, _07064_);
  and _68340_ (_17021_, _17020_, _06161_);
  and _68341_ (_17022_, _17021_, _17010_);
  not _68342_ (_17023_, _07809_);
  nor _68343_ (_17024_, _08211_, _17023_);
  nor _68344_ (_17025_, _17024_, _16990_);
  nor _68345_ (_17026_, _17025_, _06161_);
  or _68346_ (_17027_, _17026_, _06156_);
  or _68347_ (_17028_, _17027_, _17022_);
  and _68348_ (_17029_, _14169_, _08409_);
  nor _68349_ (_17030_, _08409_, _05855_);
  or _68350_ (_17031_, _17030_, _06157_);
  or _68351_ (_17032_, _17031_, _17029_);
  and _68352_ (_17033_, _17032_, _07075_);
  and _68353_ (_17034_, _17033_, _17028_);
  and _68354_ (_17035_, _17003_, _06217_);
  or _68355_ (_17036_, _17035_, _10516_);
  or _68356_ (_17037_, _17036_, _17034_);
  and _68357_ (_17038_, _17037_, _17008_);
  or _68358_ (_17039_, _17038_, _07081_);
  or _68359_ (_17040_, _09160_, _07082_);
  and _68360_ (_17041_, _17040_, _06229_);
  and _68361_ (_17042_, _17041_, _17039_);
  and _68362_ (_17043_, _08211_, _06220_);
  or _68363_ (_17044_, _17043_, _10525_);
  or _68364_ (_17045_, _17044_, _17042_);
  nand _68365_ (_17046_, _10525_, _09902_);
  and _68366_ (_17047_, _17046_, _17045_);
  or _68367_ (_17048_, _17047_, _06152_);
  or _68368_ (_17049_, _16990_, _06153_);
  and _68369_ (_17050_, _17049_, _06146_);
  nand _68370_ (_17051_, _17050_, _17048_);
  or _68371_ (_17052_, _17025_, _06146_);
  and _68372_ (_17053_, _17052_, _09301_);
  and _68373_ (_17054_, _17053_, _17051_);
  nand _68374_ (_17055_, _16232_, _09295_);
  nand _68375_ (_17056_, _17055_, _10554_);
  nor _68376_ (_17057_, _17056_, _17054_);
  nor _68377_ (_17058_, _10354_, _05855_);
  nor _68378_ (_17059_, _17058_, _10562_);
  or _68379_ (_17060_, _17059_, _10554_);
  nand _68380_ (_17061_, _17060_, _12380_);
  or _68381_ (_17062_, _17061_, _17057_);
  and _68382_ (_17063_, _17062_, _17007_);
  or _68383_ (_17064_, _17063_, _06260_);
  nor _68384_ (_17065_, _10434_, _05855_);
  or _68385_ (_17066_, _17065_, _10435_);
  or _68386_ (_17067_, _17066_, _06265_);
  and _68387_ (_17068_, _17067_, _10388_);
  and _68388_ (_17069_, _17068_, _17064_);
  nor _68389_ (_17070_, _10701_, _05855_);
  or _68390_ (_17071_, _17070_, _10702_);
  and _68391_ (_17072_, _17071_, _10387_);
  or _68392_ (_17073_, _17072_, _05870_);
  or _68393_ (_17074_, _17073_, _17069_);
  nand _68394_ (_17075_, _06107_, _05870_);
  and _68395_ (_17076_, _17075_, _06140_);
  and _68396_ (_17077_, _17076_, _17074_);
  and _68397_ (_17078_, _14171_, _08409_);
  or _68398_ (_17079_, _17078_, _17030_);
  and _68399_ (_17080_, _17079_, _06139_);
  or _68400_ (_17081_, _17080_, _09842_);
  or _68401_ (_17082_, _17081_, _17077_);
  and _68402_ (_17083_, _17082_, _17004_);
  or _68403_ (_17084_, _17083_, _06116_);
  and _68404_ (_17085_, _09160_, _07809_);
  or _68405_ (_17086_, _16990_, _06117_);
  or _68406_ (_17087_, _17086_, _17085_);
  and _68407_ (_17088_, _17087_, _06114_);
  and _68408_ (_17089_, _17088_, _17084_);
  or _68409_ (_17090_, _17089_, _17001_);
  and _68410_ (_17091_, _17090_, _09861_);
  or _68411_ (_17092_, _16813_, _05801_);
  or _68412_ (_17093_, _17092_, _17091_);
  and _68413_ (_17094_, _17093_, _16998_);
  or _68414_ (_17095_, _17094_, _06110_);
  and _68415_ (_17096_, _07809_, _08708_);
  or _68416_ (_17097_, _17096_, _16990_);
  or _68417_ (_17098_, _17097_, _06111_);
  and _68418_ (_17099_, _17098_, _10752_);
  and _68419_ (_17100_, _17099_, _17095_);
  nor _68420_ (_17101_, _10752_, _06107_);
  or _68421_ (_17102_, _17101_, _06558_);
  or _68422_ (_17103_, _17102_, _17100_);
  or _68423_ (_17104_, _16986_, _10762_);
  and _68424_ (_17105_, _06288_, _06399_);
  nor _68425_ (_17106_, _17105_, _10768_);
  and _68426_ (_17107_, _17106_, _17104_);
  and _68427_ (_17108_, _17107_, _17103_);
  not _68428_ (_17109_, _17106_);
  and _68429_ (_17110_, _17109_, _16986_);
  or _68430_ (_17111_, _17110_, _06771_);
  or _68431_ (_17112_, _17111_, _17108_);
  not _68432_ (_17113_, _06771_);
  or _68433_ (_17114_, _16986_, _17113_);
  and _68434_ (_17115_, _17114_, _17112_);
  or _68435_ (_17116_, _17115_, _10775_);
  nor _68436_ (_17117_, _11027_, _16993_);
  or _68437_ (_17118_, _10776_, _17117_);
  and _68438_ (_17119_, _17118_, _17116_);
  or _68439_ (_17120_, _17119_, _06400_);
  nand _68440_ (_17121_, _12322_, _06400_);
  and _68441_ (_17122_, _17121_, _10788_);
  and _68442_ (_17123_, _17122_, _17120_);
  and _68443_ (_17124_, _10787_, _12339_);
  or _68444_ (_17125_, _17124_, _06297_);
  or _68445_ (_17126_, _17125_, _17123_);
  and _68446_ (_17127_, _17126_, _16997_);
  or _68447_ (_17128_, _17127_, _06402_);
  or _68448_ (_17129_, _16990_, _07125_);
  and _68449_ (_17130_, _17129_, _10808_);
  and _68450_ (_17131_, _17130_, _17128_);
  and _68451_ (_17132_, _10812_, _10985_);
  or _68452_ (_17133_, _17132_, _10811_);
  or _68453_ (_17134_, _17133_, _17131_);
  or _68454_ (_17135_, _10816_, _11027_);
  and _68455_ (_17136_, _17135_, _06410_);
  and _68456_ (_17137_, _17136_, _17134_);
  or _68457_ (_17138_, _10820_, _10276_);
  and _68458_ (_17139_, _17138_, _10822_);
  or _68459_ (_17140_, _17139_, _17137_);
  or _68460_ (_17141_, _10826_, _11067_);
  and _68461_ (_17142_, _17141_, _07132_);
  and _68462_ (_17143_, _17142_, _17140_);
  nand _68463_ (_17144_, _17097_, _06306_);
  nor _68464_ (_17145_, _17144_, _17024_);
  or _68465_ (_17146_, _17145_, _06524_);
  or _68466_ (_17147_, _17146_, _17143_);
  and _68467_ (_17148_, _06957_, _05840_);
  or _68468_ (_17149_, _17148_, _06555_);
  not _68469_ (_17150_, _17149_);
  nand _68470_ (_17151_, _16985_, _06524_);
  and _68471_ (_17152_, _17151_, _17150_);
  and _68472_ (_17153_, _17152_, _17147_);
  and _68473_ (_17154_, _06684_, _05840_);
  and _68474_ (_17155_, _06288_, _05840_);
  or _68475_ (_17156_, _17155_, _17154_);
  nor _68476_ (_17157_, _17150_, _16985_);
  or _68477_ (_17158_, _17157_, _17156_);
  or _68478_ (_17159_, _17158_, _17153_);
  and _68479_ (_17160_, _06273_, _05840_);
  not _68480_ (_17161_, _17160_);
  nand _68481_ (_17162_, _17156_, _16985_);
  and _68482_ (_17163_, _17162_, _17161_);
  and _68483_ (_17164_, _17163_, _17159_);
  nor _68484_ (_17165_, _16985_, _17161_);
  or _68485_ (_17166_, _17165_, _10841_);
  or _68486_ (_17167_, _17166_, _17164_);
  and _68487_ (_17168_, _17167_, _16994_);
  or _68488_ (_17169_, _17168_, _06394_);
  nand _68489_ (_17170_, _12321_, _06394_);
  and _68490_ (_17171_, _17170_, _10851_);
  and _68491_ (_17172_, _17171_, _17169_);
  nor _68492_ (_17173_, _10851_, _12338_);
  or _68493_ (_17174_, _17173_, _06303_);
  or _68494_ (_17175_, _17174_, _17172_);
  and _68495_ (_17176_, _17175_, _16992_);
  or _68496_ (_17177_, _17176_, _10858_);
  nand _68497_ (_17178_, _17059_, _10858_);
  and _68498_ (_17179_, _17178_, _10867_);
  and _68499_ (_17180_, _17179_, _17177_);
  and _68500_ (_17181_, _10865_, _17006_);
  or _68501_ (_17182_, _17181_, _06406_);
  or _68502_ (_17183_, _17182_, _17180_);
  or _68503_ (_17184_, _17066_, _06407_);
  and _68504_ (_17185_, _17184_, _10927_);
  and _68505_ (_17186_, _17185_, _17183_);
  and _68506_ (_17187_, _10895_, _17071_);
  or _68507_ (_17188_, _17187_, _10925_);
  or _68508_ (_17189_, _17188_, _17186_);
  nand _68509_ (_17190_, _10925_, _10693_);
  and _68510_ (_17191_, _17190_, _10962_);
  and _68511_ (_17192_, _17191_, _17189_);
  or _68512_ (_17193_, _17192_, _16988_);
  and _68513_ (_17194_, _17193_, _10957_);
  and _68514_ (_17195_, _06284_, _05825_);
  and _68515_ (_17196_, _16986_, _10956_);
  or _68516_ (_17197_, _17196_, _17195_);
  or _68517_ (_17198_, _17197_, _17194_);
  and _68518_ (_17199_, _06281_, _05825_);
  not _68519_ (_17200_, _17199_);
  not _68520_ (_17201_, _17195_);
  or _68521_ (_17202_, _17201_, _17117_);
  and _68522_ (_17203_, _17202_, _17200_);
  and _68523_ (_17204_, _17203_, _17198_);
  and _68524_ (_17205_, _17117_, _17199_);
  or _68525_ (_17206_, _17205_, _06169_);
  or _68526_ (_17207_, _17206_, _17204_);
  and _68527_ (_17208_, _17207_, _16984_);
  and _68528_ (_17209_, _12339_, _10264_);
  or _68529_ (_17210_, _17209_, _10262_);
  or _68530_ (_17211_, _17210_, _17208_);
  and _68531_ (_17212_, _17211_, _16982_);
  or _68532_ (_17213_, _17212_, _06433_);
  nand _68533_ (_17214_, _17025_, _06433_);
  and _68534_ (_17215_, _17214_, _11090_);
  and _68535_ (_17216_, _17215_, _17213_);
  nor _68536_ (_17217_, _11094_, _05855_);
  nor _68537_ (_17218_, _17217_, _12719_);
  or _68538_ (_17219_, _17218_, _17216_);
  nand _68539_ (_17220_, _11094_, _05887_);
  and _68540_ (_17221_, _17220_, _05749_);
  and _68541_ (_17222_, _17221_, _17219_);
  and _68542_ (_17223_, _16990_, _05748_);
  or _68543_ (_17224_, _17223_, _06440_);
  or _68544_ (_17225_, _17224_, _17222_);
  nand _68545_ (_17226_, _17025_, _06440_);
  and _68546_ (_17227_, _17226_, _11113_);
  and _68547_ (_17228_, _17227_, _17225_);
  nor _68548_ (_17229_, _11119_, _05855_);
  nor _68549_ (_17230_, _17229_, _12744_);
  or _68550_ (_17231_, _17230_, _17228_);
  nand _68551_ (_17232_, _11119_, _05887_);
  and _68552_ (_17233_, _17232_, _01317_);
  and _68553_ (_17234_, _17233_, _17231_);
  or _68554_ (_17235_, _17234_, _16981_);
  and _68555_ (_43603_, _17235_, _43100_);
  nor _68556_ (_17236_, _01317_, _05887_);
  or _68557_ (_17237_, _10906_, _10905_);
  nor _68558_ (_17238_, _10907_, _06407_);
  and _68559_ (_17239_, _17238_, _17237_);
  and _68560_ (_17240_, _06284_, _06300_);
  not _68561_ (_17241_, _17240_);
  not _68562_ (_17242_, _10841_);
  or _68563_ (_17243_, _17242_, _11024_);
  nor _68564_ (_17244_, _10835_, _17154_);
  nor _68565_ (_17245_, _10983_, _17160_);
  or _68566_ (_17246_, _17245_, _17244_);
  or _68567_ (_17247_, _10816_, _11023_);
  not _68568_ (_17248_, _10984_);
  and _68569_ (_17249_, _17106_, _10762_);
  nor _68570_ (_17250_, _17249_, _17248_);
  nor _68571_ (_17251_, _07809_, _05887_);
  and _68572_ (_17252_, _07809_, _07306_);
  or _68573_ (_17253_, _17252_, _17251_);
  or _68574_ (_17254_, _17253_, _06132_);
  or _68575_ (_17255_, _10458_, _07306_);
  or _68576_ (_17256_, _17009_, _09115_);
  and _68577_ (_17257_, _17011_, _07306_);
  or _68578_ (_17258_, _06653_, \oc8051_golden_model_1.ACC [1]);
  nand _68579_ (_17259_, _06653_, \oc8051_golden_model_1.ACC [1]);
  and _68580_ (_17260_, _17259_, _17258_);
  and _68581_ (_17261_, _17260_, _10471_);
  or _68582_ (_17262_, _17261_, _10473_);
  or _68583_ (_17263_, _17262_, _17257_);
  and _68584_ (_17264_, _17263_, _05772_);
  or _68585_ (_17265_, _17264_, _07064_);
  and _68586_ (_17266_, _17265_, _17256_);
  or _68587_ (_17267_, _17266_, _06160_);
  or _68588_ (_17268_, _07809_, \oc8051_golden_model_1.ACC [1]);
  and _68589_ (_17269_, _14363_, _07809_);
  not _68590_ (_17270_, _17269_);
  and _68591_ (_17271_, _17270_, _17268_);
  or _68592_ (_17272_, _17271_, _06161_);
  and _68593_ (_17273_, _17272_, _17267_);
  or _68594_ (_17274_, _17273_, _10490_);
  nor _68595_ (_17275_, _10494_, \oc8051_golden_model_1.PSW [6]);
  nor _68596_ (_17276_, _17275_, \oc8051_golden_model_1.ACC [1]);
  and _68597_ (_17277_, _17275_, \oc8051_golden_model_1.ACC [1]);
  nor _68598_ (_17278_, _17277_, _17276_);
  nand _68599_ (_17279_, _17278_, _10490_);
  and _68600_ (_17280_, _17279_, _06221_);
  and _68601_ (_17281_, _17280_, _17274_);
  nor _68602_ (_17282_, _08409_, _05887_);
  and _68603_ (_17283_, _14367_, _08409_);
  or _68604_ (_17284_, _17283_, _17282_);
  and _68605_ (_17285_, _17284_, _06156_);
  and _68606_ (_17286_, _17253_, _06217_);
  or _68607_ (_17287_, _17286_, _10516_);
  or _68608_ (_17288_, _17287_, _17285_);
  or _68609_ (_17289_, _17288_, _17281_);
  and _68610_ (_17290_, _17289_, _17255_);
  or _68611_ (_17291_, _17290_, _07081_);
  or _68612_ (_17292_, _09115_, _07082_);
  and _68613_ (_17293_, _17292_, _06229_);
  and _68614_ (_17294_, _17293_, _17291_);
  nor _68615_ (_17295_, _08175_, _06229_);
  or _68616_ (_17296_, _17295_, _10525_);
  or _68617_ (_17297_, _17296_, _17294_);
  nand _68618_ (_17298_, _10525_, _09930_);
  and _68619_ (_17299_, _17298_, _17297_);
  or _68620_ (_17300_, _17299_, _06152_);
  and _68621_ (_17301_, _14349_, _08409_);
  or _68622_ (_17302_, _17301_, _17282_);
  or _68623_ (_17303_, _17302_, _06153_);
  and _68624_ (_17304_, _17303_, _06146_);
  and _68625_ (_17305_, _17304_, _17300_);
  or _68626_ (_17306_, _17282_, _14382_);
  and _68627_ (_17307_, _17284_, _06145_);
  and _68628_ (_17308_, _17307_, _17306_);
  or _68629_ (_17309_, _17308_, _09295_);
  or _68630_ (_17310_, _17309_, _17305_);
  nor _68631_ (_17311_, _09771_, _09770_);
  or _68632_ (_17312_, _17311_, _09772_);
  nand _68633_ (_17313_, _17312_, _09295_);
  and _68634_ (_17314_, _17313_, _10554_);
  and _68635_ (_17315_, _17314_, _17310_);
  nor _68636_ (_17316_, _10345_, _05855_);
  or _68637_ (_17317_, _17316_, _10353_);
  or _68638_ (_17318_, _17317_, _17248_);
  nand _68639_ (_17319_, _17317_, _17248_);
  and _68640_ (_17320_, _17319_, _17318_);
  and _68641_ (_17321_, _17320_, _10557_);
  or _68642_ (_17322_, _17321_, _17315_);
  and _68643_ (_17323_, _17322_, _12380_);
  nor _68644_ (_17324_, _10621_, _05855_);
  or _68645_ (_17325_, _17324_, _10626_);
  nor _68646_ (_17326_, _17325_, _11026_);
  and _68647_ (_17327_, _17325_, _11026_);
  or _68648_ (_17328_, _17327_, _17326_);
  and _68649_ (_17329_, _17328_, _12379_);
  or _68650_ (_17330_, _17329_, _17323_);
  and _68651_ (_17331_, _17330_, _06265_);
  nor _68652_ (_17332_, _10389_, _05855_);
  or _68653_ (_17333_, _17332_, _10433_);
  nor _68654_ (_17334_, _17333_, _10278_);
  and _68655_ (_17335_, _17333_, _10278_);
  or _68656_ (_17336_, _17335_, _10387_);
  or _68657_ (_17337_, _17336_, _17334_);
  and _68658_ (_17338_, _17337_, _12386_);
  or _68659_ (_17339_, _17338_, _17331_);
  nor _68660_ (_17340_, _06107_, \oc8051_golden_model_1.ACC [0]);
  nor _68661_ (_17341_, _17340_, _11066_);
  and _68662_ (_17342_, _17340_, _11066_);
  nor _68663_ (_17343_, _17342_, _17341_);
  or _68664_ (_17344_, _12339_, _10693_);
  and _68665_ (_17345_, _17344_, _17343_);
  and _68666_ (_17346_, _12340_, \oc8051_golden_model_1.PSW [7]);
  or _68667_ (_17347_, _17346_, _17345_);
  or _68668_ (_17348_, _17347_, _10388_);
  and _68669_ (_17349_, _17348_, _17339_);
  or _68670_ (_17350_, _17349_, _05870_);
  nand _68671_ (_17351_, _06912_, _05870_);
  and _68672_ (_17352_, _17351_, _06140_);
  and _68673_ (_17353_, _17352_, _17350_);
  and _68674_ (_17354_, _14351_, _08409_);
  or _68675_ (_17355_, _17354_, _17282_);
  and _68676_ (_17356_, _17355_, _06139_);
  or _68677_ (_17357_, _17356_, _09842_);
  or _68678_ (_17358_, _17357_, _17353_);
  and _68679_ (_17359_, _17358_, _17254_);
  or _68680_ (_17360_, _17359_, _06116_);
  and _68681_ (_17361_, _09115_, _07809_);
  or _68682_ (_17362_, _17251_, _06117_);
  or _68683_ (_17363_, _17362_, _17361_);
  and _68684_ (_17364_, _17363_, _06114_);
  and _68685_ (_17365_, _17364_, _17360_);
  or _68686_ (_17366_, _14442_, _17023_);
  and _68687_ (_17367_, _17268_, _05787_);
  and _68688_ (_17368_, _17367_, _17366_);
  or _68689_ (_17369_, _17368_, _09855_);
  or _68690_ (_17370_, _17369_, _17365_);
  or _68691_ (_17371_, _10115_, _09861_);
  and _68692_ (_17372_, _17371_, _17370_);
  or _68693_ (_17373_, _17372_, _05801_);
  nand _68694_ (_17374_, _06912_, _05801_);
  and _68695_ (_17375_, _17374_, _06111_);
  and _68696_ (_17377_, _17375_, _17373_);
  nand _68697_ (_17378_, _07809_, _06945_);
  and _68698_ (_17379_, _17378_, _06110_);
  and _68699_ (_17380_, _17379_, _17268_);
  or _68700_ (_17381_, _17380_, _10751_);
  or _68701_ (_17382_, _17381_, _17377_);
  nand _68702_ (_17383_, _10751_, _06912_);
  and _68703_ (_17384_, _17383_, _17249_);
  and _68704_ (_17385_, _17384_, _17382_);
  or _68705_ (_17386_, _17385_, _17250_);
  and _68706_ (_17388_, _17386_, _17113_);
  and _68707_ (_17389_, _10984_, _06771_);
  or _68708_ (_17390_, _17389_, _10775_);
  or _68709_ (_17391_, _17390_, _17388_);
  or _68710_ (_17392_, _10776_, _11026_);
  and _68711_ (_17393_, _17392_, _17391_);
  or _68712_ (_17394_, _17393_, _06400_);
  or _68713_ (_17395_, _10278_, _06401_);
  and _68714_ (_17396_, _17395_, _10788_);
  and _68715_ (_17397_, _17396_, _17394_);
  and _68716_ (_17399_, _10787_, _11066_);
  or _68717_ (_17400_, _17399_, _17397_);
  and _68718_ (_17401_, _17400_, _07127_);
  or _68719_ (_17402_, _14346_, _17023_);
  and _68720_ (_17403_, _17268_, _06297_);
  and _68721_ (_17404_, _17403_, _17402_);
  or _68722_ (_17405_, _17404_, _06402_);
  or _68723_ (_17406_, _17405_, _17401_);
  and _68724_ (_17407_, _06122_, _06408_);
  not _68725_ (_17408_, _17407_);
  or _68726_ (_17410_, _17251_, _07125_);
  and _68727_ (_17411_, _17410_, _17408_);
  and _68728_ (_17412_, _17411_, _17406_);
  and _68729_ (_17413_, _17407_, _10982_);
  or _68730_ (_17414_, _17413_, _06965_);
  or _68731_ (_17415_, _17414_, _17412_);
  not _68732_ (_17416_, _10807_);
  not _68733_ (_17417_, _06965_);
  or _68734_ (_17418_, _10982_, _17417_);
  and _68735_ (_17419_, _17418_, _17416_);
  and _68736_ (_17421_, _17419_, _17415_);
  and _68737_ (_17422_, _10807_, _10982_);
  or _68738_ (_17423_, _17422_, _10811_);
  or _68739_ (_17424_, _17423_, _17421_);
  and _68740_ (_17425_, _17424_, _17247_);
  or _68741_ (_17426_, _17425_, _06409_);
  or _68742_ (_17427_, _10275_, _06410_);
  and _68743_ (_17428_, _17427_, _10826_);
  and _68744_ (_17429_, _17428_, _17426_);
  and _68745_ (_17430_, _10820_, _11064_);
  or _68746_ (_17432_, _17430_, _17429_);
  and _68747_ (_17433_, _17432_, _07132_);
  or _68748_ (_17434_, _14344_, _17023_);
  and _68749_ (_17435_, _17268_, _06306_);
  and _68750_ (_17436_, _17435_, _17434_);
  or _68751_ (_17437_, _17436_, _06524_);
  or _68752_ (_17438_, _17437_, _17433_);
  nand _68753_ (_17439_, _10983_, _06524_);
  and _68754_ (_17440_, _17439_, _17150_);
  and _68755_ (_17441_, _17440_, _17438_);
  nor _68756_ (_17442_, _17150_, _10983_);
  or _68757_ (_17443_, _17442_, _17156_);
  or _68758_ (_17444_, _17443_, _17441_);
  and _68759_ (_17445_, _17444_, _17246_);
  nor _68760_ (_17446_, _10983_, _17161_);
  or _68761_ (_17447_, _17446_, _10841_);
  or _68762_ (_17448_, _17447_, _17445_);
  and _68763_ (_17449_, _17448_, _17243_);
  or _68764_ (_17450_, _17449_, _06394_);
  nand _68765_ (_17451_, _10277_, _06394_);
  and _68766_ (_17452_, _17451_, _10851_);
  and _68767_ (_17453_, _17452_, _17450_);
  nor _68768_ (_17454_, _10851_, _11065_);
  or _68769_ (_17455_, _17454_, _17453_);
  and _68770_ (_17456_, _17455_, _08819_);
  or _68771_ (_17457_, _17378_, _08176_);
  and _68772_ (_17458_, _17268_, _06303_);
  and _68773_ (_17459_, _17458_, _17457_);
  or _68774_ (_17460_, _17459_, _10858_);
  or _68775_ (_17461_, _17460_, _17456_);
  nor _68776_ (_17462_, _10355_, _10352_);
  nor _68777_ (_17463_, _17462_, _10356_);
  or _68778_ (_17464_, _17463_, _10380_);
  and _68779_ (_17465_, _17464_, _17461_);
  and _68780_ (_17466_, _17465_, _17241_);
  nor _68781_ (_17467_, _10876_, _10875_);
  nor _68782_ (_17468_, _17467_, _10877_);
  and _68783_ (_17469_, _17468_, _17240_);
  or _68784_ (_17470_, _17469_, _17466_);
  or _68785_ (_17471_, _17470_, _06792_);
  or _68786_ (_17472_, _17468_, _06793_);
  and _68787_ (_17473_, _17472_, _06407_);
  and _68788_ (_17474_, _17473_, _17471_);
  or _68789_ (_17475_, _17474_, _17239_);
  and _68790_ (_17476_, _17475_, _10927_);
  nor _68791_ (_17477_, _10936_, _10935_);
  nor _68792_ (_17478_, _17477_, _10937_);
  and _68793_ (_17479_, _17478_, _10895_);
  or _68794_ (_17480_, _17479_, _10925_);
  or _68795_ (_17481_, _17480_, _17476_);
  nand _68796_ (_17482_, _10925_, _05855_);
  and _68797_ (_17483_, _17482_, _10963_);
  and _68798_ (_17484_, _17483_, _17481_);
  or _68799_ (_17485_, _10985_, _10984_);
  nor _68800_ (_17486_, _10986_, _10963_);
  and _68801_ (_17487_, _17486_, _17485_);
  or _68802_ (_17488_, _17487_, _11003_);
  or _68803_ (_17489_, _17488_, _17484_);
  nor _68804_ (_17490_, _11027_, _11026_);
  nor _68805_ (_17491_, _17490_, _11028_);
  or _68806_ (_17492_, _17491_, _11041_);
  and _68807_ (_17493_, _17492_, _06171_);
  and _68808_ (_17494_, _17493_, _17489_);
  nor _68809_ (_17495_, _10278_, _10276_);
  nor _68810_ (_17496_, _17495_, _10279_);
  or _68811_ (_17497_, _17496_, _10264_);
  and _68812_ (_17498_, _17497_, _12691_);
  or _68813_ (_17499_, _17498_, _17494_);
  nor _68814_ (_17500_, _11067_, _11066_);
  nor _68815_ (_17501_, _17500_, _11068_);
  or _68816_ (_17502_, _17501_, _10265_);
  and _68817_ (_17503_, _17502_, _12693_);
  and _68818_ (_17504_, _17503_, _17499_);
  and _68819_ (_17505_, _10262_, \oc8051_golden_model_1.ACC [0]);
  or _68820_ (_17506_, _17505_, _06433_);
  or _68821_ (_17507_, _17506_, _17504_);
  or _68822_ (_17508_, _17271_, _06829_);
  and _68823_ (_17509_, _17508_, _11090_);
  and _68824_ (_17510_, _17509_, _17507_);
  nor _68825_ (_17511_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor _68826_ (_17512_, _11120_, _17511_);
  nor _68827_ (_17513_, _17512_, _11090_);
  or _68828_ (_17514_, _17513_, _11094_);
  or _68829_ (_17515_, _17514_, _17510_);
  nand _68830_ (_17516_, _11094_, _09981_);
  and _68831_ (_17517_, _17516_, _05749_);
  and _68832_ (_17518_, _17517_, _17515_);
  and _68833_ (_17519_, _17302_, _05748_);
  or _68834_ (_17520_, _17519_, _06440_);
  or _68835_ (_17521_, _17520_, _17518_);
  or _68836_ (_17522_, _17269_, _17251_);
  or _68837_ (_17523_, _17522_, _06444_);
  and _68838_ (_17524_, _17523_, _11113_);
  and _68839_ (_17525_, _17524_, _17521_);
  and _68840_ (_17526_, _17512_, _11112_);
  or _68841_ (_17527_, _17526_, _11119_);
  or _68842_ (_17528_, _17527_, _17525_);
  nand _68843_ (_17529_, _11119_, _09981_);
  and _68844_ (_17530_, _17529_, _01317_);
  and _68845_ (_17531_, _17530_, _17528_);
  or _68846_ (_17532_, _17531_, _17236_);
  and _68847_ (_43604_, _17532_, _43100_);
  nor _68848_ (_17533_, _01317_, _09981_);
  nand _68849_ (_17534_, _10262_, _05887_);
  and _68850_ (_17535_, _10283_, _10280_);
  nor _68851_ (_17536_, _17535_, _10284_);
  or _68852_ (_17537_, _17536_, _06171_);
  and _68853_ (_17538_, _17537_, _10265_);
  nand _68854_ (_17539_, _10908_, _10427_);
  nor _68855_ (_17540_, _10909_, _06407_);
  and _68856_ (_17541_, _17540_, _17539_);
  nand _68857_ (_17542_, _10357_, _10344_);
  nor _68858_ (_17543_, _10380_, _10358_);
  and _68859_ (_17544_, _17543_, _17542_);
  nand _68860_ (_17545_, _10848_, _11062_);
  and _68861_ (_17546_, _06122_, _05840_);
  nand _68862_ (_17547_, _17546_, _10979_);
  and _68863_ (_17548_, _14646_, _07809_);
  nor _68864_ (_17549_, _07809_, _09981_);
  or _68865_ (_17550_, _17549_, _07127_);
  or _68866_ (_17551_, _17550_, _17548_);
  or _68867_ (_17552_, _10776_, _11021_);
  nor _68868_ (_17553_, _10752_, _06625_);
  and _68869_ (_17554_, _07809_, _07708_);
  or _68870_ (_17555_, _17554_, _17549_);
  or _68871_ (_17556_, _17555_, _06132_);
  and _68872_ (_17557_, _08175_, \oc8051_golden_model_1.ACC [1]);
  and _68873_ (_17558_, _08211_, _05855_);
  nor _68874_ (_17559_, _17558_, _13920_);
  nor _68875_ (_17560_, _17559_, _17557_);
  nor _68876_ (_17561_, _17560_, _10282_);
  and _68877_ (_17562_, _17560_, _10282_);
  nor _68878_ (_17563_, _17562_, _17561_);
  and _68879_ (_17564_, _12323_, \oc8051_golden_model_1.PSW [7]);
  or _68880_ (_17565_, _17564_, _17563_);
  nand _68881_ (_17566_, _17564_, _17563_);
  and _68882_ (_17567_, _17566_, _17565_);
  or _68883_ (_17568_, _17567_, _06265_);
  and _68884_ (_17569_, _17568_, _10388_);
  or _68885_ (_17570_, _10458_, _07708_);
  nor _68886_ (_17571_, _08409_, _09981_);
  and _68887_ (_17572_, _14538_, _08409_);
  or _68888_ (_17573_, _17572_, _17571_);
  or _68889_ (_17574_, _17573_, _06157_);
  and _68890_ (_17575_, _17574_, _07075_);
  and _68891_ (_17576_, _14542_, _07809_);
  or _68892_ (_17577_, _17576_, _17549_);
  and _68893_ (_17578_, _17577_, _06160_);
  or _68894_ (_17579_, _17009_, _09211_);
  and _68895_ (_17580_, _17011_, _07708_);
  or _68896_ (_17581_, _06653_, \oc8051_golden_model_1.ACC [2]);
  nand _68897_ (_17582_, _06653_, \oc8051_golden_model_1.ACC [2]);
  and _68898_ (_17583_, _17582_, _17581_);
  and _68899_ (_17584_, _17583_, _10471_);
  or _68900_ (_17585_, _17584_, _10473_);
  or _68901_ (_17586_, _17585_, _17580_);
  and _68902_ (_17587_, _17586_, _05772_);
  or _68903_ (_17588_, _17587_, _07064_);
  and _68904_ (_17589_, _17588_, _06161_);
  and _68905_ (_17590_, _17589_, _17579_);
  or _68906_ (_17591_, _17590_, _17578_);
  and _68907_ (_17592_, _17591_, _10491_);
  or _68908_ (_17593_, _17276_, \oc8051_golden_model_1.ACC [2]);
  nand _68909_ (_17594_, _17276_, \oc8051_golden_model_1.ACC [2]);
  and _68910_ (_17595_, _17594_, _17593_);
  and _68911_ (_17596_, _17595_, _10490_);
  or _68912_ (_17597_, _17596_, _06156_);
  or _68913_ (_17598_, _17597_, _17592_);
  and _68914_ (_17599_, _17598_, _17575_);
  and _68915_ (_17600_, _17555_, _06217_);
  or _68916_ (_17601_, _17600_, _10516_);
  or _68917_ (_17602_, _17601_, _17599_);
  and _68918_ (_17603_, _17602_, _17570_);
  or _68919_ (_17604_, _17603_, _07081_);
  or _68920_ (_17605_, _09211_, _07082_);
  and _68921_ (_17606_, _17605_, _06229_);
  and _68922_ (_17607_, _17606_, _17604_);
  nor _68923_ (_17608_, _08247_, _06229_);
  or _68924_ (_17609_, _17608_, _10525_);
  or _68925_ (_17610_, _17609_, _17607_);
  nand _68926_ (_17611_, _10525_, _09883_);
  and _68927_ (_17612_, _17611_, _17610_);
  or _68928_ (_17613_, _17612_, _06152_);
  and _68929_ (_17614_, _14536_, _08409_);
  or _68930_ (_17615_, _17614_, _17571_);
  or _68931_ (_17616_, _17615_, _06153_);
  and _68932_ (_17617_, _17616_, _06146_);
  and _68933_ (_17618_, _17617_, _17613_);
  or _68934_ (_17619_, _17571_, _14569_);
  and _68935_ (_17620_, _17573_, _06145_);
  and _68936_ (_17621_, _17620_, _17619_);
  or _68937_ (_17622_, _17621_, _09295_);
  or _68938_ (_17623_, _17622_, _17618_);
  nor _68939_ (_17624_, _09774_, _09772_);
  or _68940_ (_17625_, _17624_, _09775_);
  nand _68941_ (_17626_, _17625_, _09295_);
  and _68942_ (_17627_, _17626_, _10554_);
  and _68943_ (_17628_, _17627_, _17623_);
  and _68944_ (_17629_, _07252_, \oc8051_golden_model_1.ACC [1]);
  and _68945_ (_17630_, _07049_, _05855_);
  nor _68946_ (_17631_, _17630_, _10984_);
  nor _68947_ (_17632_, _17631_, _17629_);
  nor _68948_ (_17633_, _10980_, _17632_);
  and _68949_ (_17634_, _10980_, _17632_);
  nor _68950_ (_17635_, _17634_, _17633_);
  nor _68951_ (_17636_, _16986_, _10984_);
  and _68952_ (_17637_, _17636_, \oc8051_golden_model_1.PSW [7]);
  nand _68953_ (_17638_, _17637_, _17635_);
  or _68954_ (_17639_, _17637_, _17635_);
  and _68955_ (_17640_, _17639_, _10557_);
  and _68956_ (_17641_, _17640_, _17638_);
  or _68957_ (_17642_, _17641_, _10580_);
  or _68958_ (_17643_, _17642_, _17628_);
  or _68959_ (_17644_, _09115_, _05887_);
  and _68960_ (_17645_, _09160_, _05855_);
  or _68961_ (_17646_, _17645_, _11026_);
  and _68962_ (_17647_, _17646_, _17644_);
  nor _68963_ (_17648_, _11021_, _17647_);
  and _68964_ (_17649_, _11021_, _17647_);
  nor _68965_ (_17650_, _17649_, _17648_);
  nor _68966_ (_17651_, _17117_, _11026_);
  not _68967_ (_17652_, _17651_);
  or _68968_ (_17653_, _17652_, _17650_);
  and _68969_ (_17654_, _17653_, \oc8051_golden_model_1.PSW [7]);
  nor _68970_ (_17655_, _17650_, \oc8051_golden_model_1.PSW [7]);
  nor _68971_ (_17656_, _17655_, _17654_);
  and _68972_ (_17657_, _17652_, _17650_);
  or _68973_ (_17658_, _17657_, _17656_);
  and _68974_ (_17659_, _17658_, _06276_);
  or _68975_ (_17660_, _17659_, _12380_);
  and _68976_ (_17661_, _17660_, _17643_);
  and _68977_ (_17662_, _17658_, _06709_);
  or _68978_ (_17663_, _17662_, _06260_);
  or _68979_ (_17664_, _17663_, _17661_);
  and _68980_ (_17665_, _17664_, _17569_);
  nor _68981_ (_17666_, _17341_, _13944_);
  nor _68982_ (_17667_, _11063_, _17666_);
  and _68983_ (_17668_, _11063_, _17666_);
  nor _68984_ (_17669_, _17668_, _17667_);
  nand _68985_ (_17670_, _17346_, _17669_);
  or _68986_ (_17671_, _17346_, _17669_);
  and _68987_ (_17672_, _17671_, _17670_);
  and _68988_ (_17673_, _17672_, _10387_);
  or _68989_ (_17674_, _17673_, _05870_);
  or _68990_ (_17675_, _17674_, _17665_);
  nand _68991_ (_17676_, _06625_, _05870_);
  and _68992_ (_17677_, _17676_, _06140_);
  and _68993_ (_17678_, _17677_, _17675_);
  and _68994_ (_17679_, _14583_, _08409_);
  or _68995_ (_17680_, _17679_, _17571_);
  and _68996_ (_17681_, _17680_, _06139_);
  or _68997_ (_17682_, _17681_, _09842_);
  or _68998_ (_17683_, _17682_, _17678_);
  and _68999_ (_17684_, _17683_, _17556_);
  or _69000_ (_17685_, _17684_, _06116_);
  and _69001_ (_17686_, _09211_, _07809_);
  or _69002_ (_17687_, _17549_, _06117_);
  or _69003_ (_17688_, _17687_, _17686_);
  and _69004_ (_17689_, _17688_, _06114_);
  and _69005_ (_17690_, _17689_, _17685_);
  and _69006_ (_17691_, _14630_, _07809_);
  or _69007_ (_17692_, _17691_, _17549_);
  and _69008_ (_17693_, _17692_, _05787_);
  or _69009_ (_17694_, _17693_, _09855_);
  or _69010_ (_17695_, _17694_, _17690_);
  or _69011_ (_17696_, _10052_, _09861_);
  and _69012_ (_17697_, _17696_, _05802_);
  and _69013_ (_17698_, _17697_, _17695_);
  nor _69014_ (_17699_, _06625_, _05802_);
  or _69015_ (_17700_, _17699_, _06110_);
  or _69016_ (_17701_, _17700_, _17698_);
  and _69017_ (_17702_, _07809_, _08768_);
  or _69018_ (_17703_, _17702_, _17549_);
  or _69019_ (_17704_, _17703_, _06111_);
  and _69020_ (_17705_, _17704_, _10752_);
  and _69021_ (_17706_, _17705_, _17701_);
  or _69022_ (_17707_, _17706_, _17553_);
  and _69023_ (_17708_, _17707_, _10762_);
  and _69024_ (_17709_, _06957_, _06399_);
  or _69025_ (_17710_, _17709_, _06574_);
  and _69026_ (_17711_, _10980_, _06558_);
  or _69027_ (_17712_, _17711_, _17710_);
  or _69028_ (_17713_, _17712_, _17708_);
  and _69029_ (_17714_, _06684_, _06399_);
  nor _69030_ (_17715_, _10772_, _17714_);
  nand _69031_ (_17716_, _17710_, _10981_);
  and _69032_ (_17717_, _17716_, _17715_);
  and _69033_ (_17718_, _17717_, _17713_);
  nor _69034_ (_17719_, _17715_, _10981_);
  or _69035_ (_17720_, _17719_, _10775_);
  or _69036_ (_17721_, _17720_, _17718_);
  and _69037_ (_17722_, _17721_, _17552_);
  or _69038_ (_17723_, _17722_, _06400_);
  or _69039_ (_17724_, _10282_, _06401_);
  and _69040_ (_17725_, _17724_, _10788_);
  and _69041_ (_17726_, _17725_, _17723_);
  and _69042_ (_17727_, _10787_, _11063_);
  or _69043_ (_17728_, _17727_, _06297_);
  or _69044_ (_17729_, _17728_, _17726_);
  and _69045_ (_17730_, _17729_, _17551_);
  or _69046_ (_17731_, _17730_, _06402_);
  or _69047_ (_17732_, _17549_, _07125_);
  and _69048_ (_17733_, _17732_, _10808_);
  and _69049_ (_17734_, _17733_, _17731_);
  and _69050_ (_17735_, _10812_, _10978_);
  or _69051_ (_17736_, _17735_, _10811_);
  or _69052_ (_17737_, _17736_, _17734_);
  or _69053_ (_17738_, _10816_, _11018_);
  and _69054_ (_17739_, _17738_, _06410_);
  and _69055_ (_17740_, _17739_, _17737_);
  or _69056_ (_17741_, _10820_, _10274_);
  and _69057_ (_17742_, _17741_, _10822_);
  or _69058_ (_17743_, _17742_, _17740_);
  or _69059_ (_17744_, _10826_, _11061_);
  and _69060_ (_17745_, _17744_, _07132_);
  and _69061_ (_17746_, _17745_, _17743_);
  nand _69062_ (_17747_, _17703_, _06306_);
  nor _69063_ (_17748_, _17747_, _10281_);
  or _69064_ (_17749_, _17748_, _17546_);
  or _69065_ (_17750_, _17749_, _17746_);
  nand _69066_ (_17751_, _17750_, _17547_);
  nor _69067_ (_17752_, _17156_, _17148_);
  nand _69068_ (_17753_, _17752_, _17751_);
  not _69069_ (_17754_, _17752_);
  nand _69070_ (_17755_, _17754_, _10979_);
  and _69071_ (_17756_, _17755_, _17161_);
  and _69072_ (_17757_, _17756_, _17753_);
  nor _69073_ (_17758_, _10979_, _17161_);
  or _69074_ (_17759_, _17758_, _10841_);
  or _69075_ (_17760_, _17759_, _17757_);
  or _69076_ (_17761_, _17242_, _11019_);
  and _69077_ (_17762_, _17761_, _06395_);
  and _69078_ (_17763_, _17762_, _17760_);
  nand _69079_ (_17764_, _10851_, _10281_);
  and _69080_ (_17765_, _17764_, _10850_);
  or _69081_ (_17766_, _17765_, _17763_);
  and _69082_ (_17767_, _17766_, _17545_);
  or _69083_ (_17768_, _17767_, _06303_);
  and _69084_ (_17769_, _14643_, _07809_);
  or _69085_ (_17770_, _17549_, _08819_);
  or _69086_ (_17771_, _17770_, _17769_);
  and _69087_ (_17772_, _17771_, _10380_);
  and _69088_ (_17773_, _17772_, _17768_);
  or _69089_ (_17774_, _17773_, _17544_);
  and _69090_ (_17775_, _17774_, _17241_);
  and _69091_ (_17776_, _10878_, _10619_);
  nor _69092_ (_17777_, _17776_, _10879_);
  and _69093_ (_17778_, _17777_, _17240_);
  or _69094_ (_17779_, _17778_, _17775_);
  or _69095_ (_17780_, _17779_, _06792_);
  or _69096_ (_17781_, _17777_, _06793_);
  and _69097_ (_17782_, _17781_, _06407_);
  and _69098_ (_17783_, _17782_, _17780_);
  or _69099_ (_17784_, _17783_, _17541_);
  nand _69100_ (_17785_, _17784_, _10927_);
  and _69101_ (_17786_, _10938_, _10691_);
  or _69102_ (_17787_, _10939_, _10927_);
  or _69103_ (_17788_, _17787_, _17786_);
  and _69104_ (_17789_, _17788_, _10926_);
  and _69105_ (_17790_, _17789_, _17785_);
  nand _69106_ (_17791_, _10925_, _05887_);
  nand _69107_ (_17792_, _17791_, _10963_);
  or _69108_ (_17793_, _17792_, _17790_);
  and _69109_ (_17794_, _10987_, _10981_);
  or _69110_ (_17795_, _17794_, _10988_);
  or _69111_ (_17796_, _17795_, _10963_);
  and _69112_ (_17797_, _17796_, _17201_);
  and _69113_ (_17798_, _17797_, _17793_);
  and _69114_ (_17799_, _11029_, _11022_);
  or _69115_ (_17800_, _17799_, _11030_);
  or _69116_ (_17801_, _17800_, _05707_);
  and _69117_ (_17802_, _17801_, _11003_);
  nor _69118_ (_17803_, _17802_, _17798_);
  or _69119_ (_17804_, _17800_, _17200_);
  nand _69120_ (_17805_, _17804_, _06171_);
  or _69121_ (_17806_, _17805_, _17803_);
  and _69122_ (_17807_, _17806_, _17538_);
  or _69123_ (_17808_, _11070_, _11063_);
  nor _69124_ (_17809_, _11071_, _10265_);
  and _69125_ (_17810_, _17809_, _17808_);
  or _69126_ (_17811_, _17810_, _10262_);
  or _69127_ (_17812_, _17811_, _17807_);
  and _69128_ (_17813_, _17812_, _17534_);
  or _69129_ (_17814_, _17813_, _06433_);
  or _69130_ (_17815_, _17577_, _06829_);
  and _69131_ (_17816_, _17815_, _11090_);
  and _69132_ (_17817_, _17816_, _17814_);
  nor _69133_ (_17818_, _17511_, _09981_);
  or _69134_ (_17819_, _17818_, _11095_);
  nor _69135_ (_17820_, _17819_, _11094_);
  nor _69136_ (_17821_, _17820_, _12719_);
  or _69137_ (_17822_, _17821_, _17817_);
  nand _69138_ (_17823_, _11094_, _10028_);
  and _69139_ (_17824_, _17823_, _05749_);
  and _69140_ (_17825_, _17824_, _17822_);
  and _69141_ (_17826_, _17615_, _05748_);
  or _69142_ (_17827_, _17826_, _06440_);
  or _69143_ (_17828_, _17827_, _17825_);
  and _69144_ (_17829_, _14710_, _07809_);
  or _69145_ (_17830_, _17829_, _17549_);
  or _69146_ (_17831_, _17830_, _06444_);
  and _69147_ (_17832_, _17831_, _11113_);
  and _69148_ (_17833_, _17832_, _17828_);
  nor _69149_ (_17834_, _11120_, \oc8051_golden_model_1.ACC [2]);
  nor _69150_ (_17835_, _17834_, _11121_);
  and _69151_ (_17836_, _17835_, _11112_);
  or _69152_ (_17837_, _17836_, _11119_);
  or _69153_ (_17838_, _17837_, _17833_);
  nand _69154_ (_17839_, _11119_, _10028_);
  and _69155_ (_17840_, _17839_, _01317_);
  and _69156_ (_17841_, _17840_, _17838_);
  or _69157_ (_17842_, _17841_, _17533_);
  and _69158_ (_43605_, _17842_, _43100_);
  nor _69159_ (_17843_, _01317_, _10028_);
  and _69160_ (_17844_, _10359_, _10337_);
  nor _69161_ (_17845_, _17844_, _10360_);
  or _69162_ (_17846_, _17845_, _10380_);
  not _69163_ (_17847_, _10835_);
  nor _69164_ (_17848_, _17847_, _10977_);
  or _69165_ (_17849_, _17848_, _10841_);
  nand _69166_ (_17850_, _10977_, _06524_);
  and _69167_ (_17851_, _10976_, _06965_);
  and _69168_ (_17852_, _17407_, _10976_);
  and _69169_ (_17853_, _14727_, _07809_);
  nor _69170_ (_17854_, _07809_, _10028_);
  or _69171_ (_17855_, _17854_, _07127_);
  or _69172_ (_17856_, _17855_, _17853_);
  nor _69173_ (_17857_, _10752_, _06070_);
  and _69174_ (_17858_, _07809_, _07544_);
  or _69175_ (_17859_, _17858_, _17854_);
  or _69176_ (_17860_, _17859_, _06132_);
  or _69177_ (_17861_, _10458_, _07544_);
  nor _69178_ (_17862_, _08409_, _10028_);
  and _69179_ (_17863_, _14735_, _08409_);
  or _69180_ (_17864_, _17863_, _17862_);
  or _69181_ (_17865_, _17864_, _06157_);
  and _69182_ (_17866_, _17865_, _07075_);
  and _69183_ (_17867_, _14738_, _07809_);
  or _69184_ (_17868_, _17867_, _17854_);
  and _69185_ (_17869_, _17868_, _06160_);
  or _69186_ (_17870_, _17009_, _09210_);
  and _69187_ (_17871_, _17011_, _07544_);
  or _69188_ (_17872_, _06653_, \oc8051_golden_model_1.ACC [3]);
  nand _69189_ (_17873_, _06653_, \oc8051_golden_model_1.ACC [3]);
  and _69190_ (_17874_, _17873_, _17872_);
  and _69191_ (_17875_, _17874_, _10471_);
  or _69192_ (_17876_, _17875_, _10473_);
  or _69193_ (_17877_, _17876_, _17871_);
  and _69194_ (_17878_, _17877_, _05772_);
  or _69195_ (_17879_, _17878_, _07064_);
  and _69196_ (_17880_, _17879_, _06161_);
  and _69197_ (_17881_, _17880_, _17870_);
  or _69198_ (_17882_, _17881_, _17869_);
  and _69199_ (_17883_, _17882_, _10491_);
  not _69200_ (_17884_, \oc8051_golden_model_1.PSW [6]);
  nor _69201_ (_17885_, _10493_, _17884_);
  nor _69202_ (_17886_, _17885_, \oc8051_golden_model_1.ACC [3]);
  nor _69203_ (_17887_, _17886_, _10494_);
  and _69204_ (_17888_, _17887_, _10490_);
  or _69205_ (_17889_, _17888_, _06156_);
  or _69206_ (_17890_, _17889_, _17883_);
  and _69207_ (_17891_, _17890_, _17866_);
  and _69208_ (_17892_, _17859_, _06217_);
  or _69209_ (_17893_, _17892_, _10516_);
  or _69210_ (_17894_, _17893_, _17891_);
  and _69211_ (_17895_, _17894_, _17861_);
  or _69212_ (_17896_, _17895_, _07081_);
  or _69213_ (_17897_, _09210_, _07082_);
  and _69214_ (_17898_, _17897_, _06229_);
  and _69215_ (_17899_, _17898_, _17896_);
  nor _69216_ (_17900_, _08139_, _06229_);
  or _69217_ (_17901_, _17900_, _10525_);
  or _69218_ (_17902_, _17901_, _17899_);
  nand _69219_ (_17903_, _10525_, _08430_);
  and _69220_ (_17904_, _17903_, _17902_);
  or _69221_ (_17905_, _17904_, _06152_);
  and _69222_ (_17906_, _14731_, _08409_);
  or _69223_ (_17907_, _17906_, _17862_);
  or _69224_ (_17908_, _17907_, _06153_);
  and _69225_ (_17909_, _17908_, _06146_);
  and _69226_ (_17910_, _17909_, _17905_);
  or _69227_ (_17911_, _17862_, _14764_);
  and _69228_ (_17912_, _17864_, _06145_);
  and _69229_ (_17913_, _17912_, _17911_);
  or _69230_ (_17914_, _17913_, _09295_);
  or _69231_ (_17915_, _17914_, _17910_);
  nor _69232_ (_17916_, _09777_, _09775_);
  or _69233_ (_17917_, _17916_, _09778_);
  nand _69234_ (_17918_, _17917_, _09295_);
  and _69235_ (_17919_, _17918_, _10554_);
  and _69236_ (_17920_, _17919_, _17915_);
  and _69237_ (_17921_, _07657_, \oc8051_golden_model_1.ACC [2]);
  nor _69238_ (_17922_, _17633_, _17921_);
  nor _69239_ (_17923_, _10976_, _10977_);
  nor _69240_ (_17924_, _17923_, _17922_);
  and _69241_ (_17925_, _17923_, _17922_);
  nor _69242_ (_17926_, _17925_, _17924_);
  not _69243_ (_17927_, _17636_);
  nor _69244_ (_17928_, _17927_, _17635_);
  nand _69245_ (_17929_, _17928_, \oc8051_golden_model_1.PSW [7]);
  and _69246_ (_17930_, _17929_, _17926_);
  not _69247_ (_17931_, _17928_);
  nor _69248_ (_17932_, _17931_, _17926_);
  and _69249_ (_17933_, _17932_, \oc8051_golden_model_1.PSW [7]);
  or _69250_ (_17934_, _17933_, _17930_);
  and _69251_ (_17935_, _17934_, _10557_);
  or _69252_ (_17936_, _17935_, _12379_);
  or _69253_ (_17937_, _17936_, _17920_);
  and _69254_ (_17938_, _09070_, \oc8051_golden_model_1.ACC [2]);
  nor _69255_ (_17939_, _17648_, _17938_);
  nor _69256_ (_17940_, _11016_, _11017_);
  not _69257_ (_17941_, _17940_);
  nand _69258_ (_17942_, _17941_, _17939_);
  or _69259_ (_17943_, _17941_, _17939_);
  and _69260_ (_17944_, _17943_, _17942_);
  or _69261_ (_17945_, _17944_, _10693_);
  nand _69262_ (_17946_, _17944_, _10693_);
  and _69263_ (_17947_, _17946_, _17945_);
  nand _69264_ (_17948_, _17947_, _17654_);
  or _69265_ (_17949_, _17947_, _17654_);
  and _69266_ (_17950_, _17949_, _17948_);
  or _69267_ (_17951_, _17950_, _12380_);
  and _69268_ (_17952_, _17951_, _06265_);
  and _69269_ (_17953_, _17952_, _17937_);
  and _69270_ (_17954_, _12324_, \oc8051_golden_model_1.PSW [7]);
  and _69271_ (_17955_, _08247_, \oc8051_golden_model_1.ACC [2]);
  nor _69272_ (_17956_, _17561_, _17955_);
  nor _69273_ (_17957_, _17956_, _12318_);
  and _69274_ (_17958_, _17956_, _12318_);
  nor _69275_ (_17959_, _17958_, _17957_);
  not _69276_ (_17960_, _12323_);
  or _69277_ (_17961_, _17960_, _17563_);
  or _69278_ (_17962_, _17961_, _10693_);
  and _69279_ (_17963_, _17962_, _17959_);
  or _69280_ (_17964_, _17963_, _10387_);
  or _69281_ (_17965_, _17964_, _17954_);
  and _69282_ (_17966_, _17965_, _12386_);
  or _69283_ (_17967_, _17966_, _17953_);
  and _69284_ (_17968_, _12341_, \oc8051_golden_model_1.PSW [7]);
  and _69285_ (_17969_, _06625_, \oc8051_golden_model_1.ACC [2]);
  nor _69286_ (_17970_, _17667_, _17969_);
  nor _69287_ (_17971_, _12336_, _17970_);
  and _69288_ (_17972_, _12336_, _17970_);
  nor _69289_ (_17973_, _17972_, _17971_);
  not _69290_ (_17974_, _12340_);
  or _69291_ (_17975_, _17974_, _17669_);
  or _69292_ (_17976_, _17975_, _10693_);
  and _69293_ (_17977_, _17976_, _17973_);
  or _69294_ (_17978_, _17977_, _10388_);
  or _69295_ (_17979_, _17978_, _17968_);
  and _69296_ (_17980_, _17979_, _17967_);
  or _69297_ (_17981_, _17980_, _05870_);
  nand _69298_ (_17982_, _06070_, _05870_);
  and _69299_ (_17983_, _17982_, _06140_);
  and _69300_ (_17984_, _17983_, _17981_);
  and _69301_ (_17985_, _14732_, _08409_);
  or _69302_ (_17986_, _17985_, _17862_);
  and _69303_ (_17987_, _17986_, _06139_);
  or _69304_ (_17988_, _17987_, _09842_);
  or _69305_ (_17989_, _17988_, _17984_);
  and _69306_ (_17990_, _17989_, _17860_);
  or _69307_ (_17991_, _17990_, _06116_);
  and _69308_ (_17992_, _09210_, _07809_);
  or _69309_ (_17993_, _17854_, _06117_);
  or _69310_ (_17994_, _17993_, _17992_);
  and _69311_ (_17995_, _17994_, _06114_);
  and _69312_ (_17996_, _17995_, _17991_);
  and _69313_ (_17997_, _14825_, _07809_);
  or _69314_ (_17998_, _17997_, _17854_);
  and _69315_ (_17999_, _17998_, _05787_);
  or _69316_ (_18001_, _17999_, _09855_);
  or _69317_ (_18002_, _18001_, _17996_);
  or _69318_ (_18003_, _09998_, _09861_);
  and _69319_ (_18004_, _18003_, _05802_);
  and _69320_ (_18005_, _18004_, _18002_);
  nor _69321_ (_18006_, _06070_, _05802_);
  or _69322_ (_18007_, _18006_, _06110_);
  or _69323_ (_18008_, _18007_, _18005_);
  and _69324_ (_18009_, _07809_, _08712_);
  or _69325_ (_18010_, _18009_, _17854_);
  or _69326_ (_18011_, _18010_, _06111_);
  and _69327_ (_18012_, _18011_, _10752_);
  and _69328_ (_18013_, _18012_, _18008_);
  or _69329_ (_18014_, _18013_, _17857_);
  and _69330_ (_18015_, _18014_, _10762_);
  and _69331_ (_18016_, _17923_, _06558_);
  or _69332_ (_18017_, _18016_, _17109_);
  or _69333_ (_18018_, _18017_, _18015_);
  or _69334_ (_18019_, _17106_, _17923_);
  and _69335_ (_18020_, _18019_, _17113_);
  and _69336_ (_18021_, _18020_, _18018_);
  and _69337_ (_18022_, _17923_, _06771_);
  or _69338_ (_18023_, _18022_, _18021_);
  and _69339_ (_18024_, _18023_, _10776_);
  and _69340_ (_18025_, _10775_, _17940_);
  or _69341_ (_18026_, _18025_, _06400_);
  or _69342_ (_18027_, _18026_, _18024_);
  or _69343_ (_18028_, _12318_, _06401_);
  and _69344_ (_18029_, _18028_, _10788_);
  and _69345_ (_18030_, _18029_, _18027_);
  and _69346_ (_18031_, _10787_, _12336_);
  or _69347_ (_18032_, _18031_, _06297_);
  or _69348_ (_18033_, _18032_, _18030_);
  and _69349_ (_18034_, _18033_, _17856_);
  or _69350_ (_18035_, _18034_, _06402_);
  or _69351_ (_18036_, _17854_, _07125_);
  and _69352_ (_18037_, _18036_, _17408_);
  and _69353_ (_18038_, _18037_, _18035_);
  or _69354_ (_18039_, _18038_, _17852_);
  and _69355_ (_18040_, _18039_, _17417_);
  or _69356_ (_18041_, _18040_, _17851_);
  and _69357_ (_18042_, _18041_, _17416_);
  and _69358_ (_18043_, _10807_, _10976_);
  or _69359_ (_18044_, _18043_, _10811_);
  or _69360_ (_18045_, _18044_, _18042_);
  or _69361_ (_18046_, _10816_, _11016_);
  and _69362_ (_18047_, _18046_, _06410_);
  and _69363_ (_18048_, _18047_, _18045_);
  and _69364_ (_18049_, _10272_, _06409_);
  or _69365_ (_18050_, _18049_, _10820_);
  or _69366_ (_18051_, _18050_, _18048_);
  or _69367_ (_18052_, _10826_, _11059_);
  and _69368_ (_18053_, _18052_, _07132_);
  and _69369_ (_18054_, _18053_, _18051_);
  nand _69370_ (_18055_, _18010_, _06306_);
  nor _69371_ (_18056_, _18055_, _10273_);
  or _69372_ (_18057_, _18056_, _06524_);
  or _69373_ (_18058_, _18057_, _18054_);
  and _69374_ (_18059_, _18058_, _17850_);
  or _69375_ (_18060_, _18059_, _06555_);
  nand _69376_ (_18061_, _10977_, _06555_);
  and _69377_ (_18062_, _18061_, _18060_);
  or _69378_ (_18063_, _18062_, _06975_);
  nand _69379_ (_18064_, _10977_, _06975_);
  and _69380_ (_18065_, _18064_, _17847_);
  and _69381_ (_18066_, _18065_, _18063_);
  or _69382_ (_18067_, _18066_, _17849_);
  nand _69383_ (_18068_, _10841_, _11017_);
  and _69384_ (_18069_, _18068_, _06395_);
  and _69385_ (_18070_, _18069_, _18067_);
  nand _69386_ (_18071_, _10851_, _10273_);
  and _69387_ (_18072_, _18071_, _10850_);
  or _69388_ (_18073_, _18072_, _18070_);
  nand _69389_ (_18074_, _10848_, _11060_);
  and _69390_ (_18075_, _18074_, _08819_);
  and _69391_ (_18076_, _18075_, _18073_);
  and _69392_ (_18077_, _14724_, _07809_);
  or _69393_ (_18078_, _18077_, _17854_);
  and _69394_ (_18079_, _18078_, _06303_);
  or _69395_ (_18080_, _18079_, _10858_);
  or _69396_ (_18081_, _18080_, _18076_);
  and _69397_ (_18082_, _18081_, _17846_);
  or _69398_ (_18083_, _18082_, _10865_);
  and _69399_ (_18084_, _10880_, _10613_);
  nor _69400_ (_18085_, _18084_, _10881_);
  or _69401_ (_18086_, _18085_, _10867_);
  and _69402_ (_18087_, _18086_, _06407_);
  and _69403_ (_18088_, _18087_, _18083_);
  nand _69404_ (_18089_, _10910_, _10422_);
  nor _69405_ (_18090_, _10911_, _06407_);
  and _69406_ (_18091_, _18090_, _18089_);
  or _69407_ (_18092_, _18091_, _10895_);
  or _69408_ (_18093_, _18092_, _18088_);
  and _69409_ (_18094_, _10940_, _10685_);
  nor _69410_ (_18095_, _18094_, _10941_);
  or _69411_ (_18096_, _18095_, _10927_);
  and _69412_ (_18097_, _18096_, _10926_);
  and _69413_ (_18098_, _18097_, _18093_);
  nand _69414_ (_18099_, _10925_, \oc8051_golden_model_1.ACC [2]);
  nand _69415_ (_18100_, _18099_, _10963_);
  or _69416_ (_18101_, _18100_, _18098_);
  and _69417_ (_18102_, _10989_, _17923_);
  nor _69418_ (_18103_, _10989_, _17923_);
  or _69419_ (_18104_, _18103_, _18102_);
  or _69420_ (_18105_, _18104_, _10963_);
  and _69421_ (_18106_, _18105_, _18101_);
  or _69422_ (_18107_, _18106_, _11003_);
  and _69423_ (_18108_, _11031_, _17940_);
  nor _69424_ (_18109_, _11031_, _17940_);
  or _69425_ (_18110_, _18109_, _11041_);
  or _69426_ (_18111_, _18110_, _18108_);
  and _69427_ (_18112_, _18111_, _06171_);
  and _69428_ (_18113_, _18112_, _18107_);
  and _69429_ (_18114_, _12318_, _10285_);
  nor _69430_ (_18115_, _12318_, _10285_);
  or _69431_ (_18116_, _18115_, _10264_);
  or _69432_ (_18117_, _18116_, _18114_);
  and _69433_ (_18118_, _18117_, _12691_);
  or _69434_ (_18119_, _18118_, _18113_);
  and _69435_ (_18120_, _11072_, _12336_);
  nor _69436_ (_18121_, _11072_, _12336_);
  or _69437_ (_18122_, _18121_, _18120_);
  or _69438_ (_18123_, _18122_, _10265_);
  and _69439_ (_18124_, _18123_, _12693_);
  and _69440_ (_18125_, _18124_, _18119_);
  and _69441_ (_18126_, _10262_, \oc8051_golden_model_1.ACC [2]);
  or _69442_ (_18127_, _18126_, _06433_);
  or _69443_ (_18128_, _18127_, _18125_);
  or _69444_ (_18129_, _17868_, _06829_);
  and _69445_ (_18130_, _18129_, _11090_);
  and _69446_ (_18131_, _18130_, _18128_);
  nor _69447_ (_18132_, _11095_, _10028_);
  or _69448_ (_18133_, _18132_, _11096_);
  and _69449_ (_18134_, _18133_, _11089_);
  or _69450_ (_18135_, _18134_, _11094_);
  or _69451_ (_18136_, _18135_, _18131_);
  nand _69452_ (_18137_, _11094_, _09902_);
  and _69453_ (_18138_, _18137_, _05749_);
  and _69454_ (_18139_, _18138_, _18136_);
  and _69455_ (_18140_, _17907_, _05748_);
  or _69456_ (_18141_, _18140_, _06440_);
  or _69457_ (_18142_, _18141_, _18139_);
  and _69458_ (_18143_, _14897_, _07809_);
  or _69459_ (_18144_, _17854_, _06444_);
  or _69460_ (_18145_, _18144_, _18143_);
  and _69461_ (_18146_, _18145_, _11113_);
  and _69462_ (_18147_, _18146_, _18142_);
  nor _69463_ (_18148_, _11121_, \oc8051_golden_model_1.ACC [3]);
  nor _69464_ (_18149_, _18148_, _11122_);
  and _69465_ (_18150_, _18149_, _11112_);
  or _69466_ (_18151_, _18150_, _11119_);
  or _69467_ (_18152_, _18151_, _18147_);
  nand _69468_ (_18153_, _11119_, _09902_);
  and _69469_ (_18154_, _18153_, _01317_);
  and _69470_ (_18155_, _18154_, _18152_);
  or _69471_ (_18156_, _18155_, _17843_);
  and _69472_ (_43606_, _18156_, _43100_);
  nor _69473_ (_18157_, _01317_, _09902_);
  nand _69474_ (_18158_, _10262_, _10028_);
  or _69475_ (_18159_, _10289_, _10287_);
  and _69476_ (_18160_, _10290_, _06169_);
  and _69477_ (_18161_, _18160_, _18159_);
  or _69478_ (_18162_, _11033_, _11015_);
  and _69479_ (_18163_, _18162_, _11034_);
  or _69480_ (_18164_, _18163_, _17201_);
  or _69481_ (_18165_, _10912_, _10416_);
  and _69482_ (_18166_, _18165_, _10913_);
  or _69483_ (_18167_, _18166_, _06407_);
  and _69484_ (_18168_, _18167_, _10927_);
  nand _69485_ (_18169_, _10848_, _11057_);
  or _69486_ (_18170_, _06965_, _06554_);
  and _69487_ (_18171_, _18170_, _10972_);
  not _69488_ (_18172_, _17105_);
  and _69489_ (_18173_, _18172_, _06772_);
  nor _69490_ (_18174_, _06722_, _05833_);
  and _69491_ (_18175_, _06123_, _06399_);
  nor _69492_ (_18176_, _18175_, _18174_);
  not _69493_ (_18177_, _18176_);
  and _69494_ (_18178_, _06128_, _06399_);
  nor _69495_ (_18179_, _18178_, _18177_);
  and _69496_ (_18180_, _18179_, _18173_);
  and _69497_ (_18181_, _06277_, _06399_);
  not _69498_ (_18182_, _18181_);
  nor _69499_ (_18183_, _10752_, _06876_);
  nor _69500_ (_18184_, _07809_, _09902_);
  and _69501_ (_18185_, _08336_, _07809_);
  or _69502_ (_18186_, _18185_, _18184_);
  or _69503_ (_18187_, _18186_, _06132_);
  nand _69504_ (_18188_, _17948_, _17945_);
  and _69505_ (_18189_, _09210_, _10028_);
  or _69506_ (_18191_, _09210_, _10028_);
  and _69507_ (_18192_, _18191_, _17939_);
  or _69508_ (_18193_, _18192_, _18189_);
  nor _69509_ (_18194_, _11015_, _18193_);
  not _69510_ (_18195_, _18194_);
  nand _69511_ (_18196_, _11015_, _18193_);
  and _69512_ (_18197_, _18196_, _18195_);
  nand _69513_ (_18198_, _18197_, \oc8051_golden_model_1.PSW [7]);
  or _69514_ (_18199_, _18197_, \oc8051_golden_model_1.PSW [7]);
  and _69515_ (_18200_, _18199_, _18198_);
  or _69516_ (_18202_, _18200_, _18188_);
  nand _69517_ (_18203_, _18200_, _18188_);
  and _69518_ (_18204_, _12379_, _18203_);
  and _69519_ (_18205_, _18204_, _18202_);
  nor _69520_ (_18206_, _17932_, _10693_);
  and _69521_ (_18207_, _07544_, _10028_);
  or _69522_ (_18208_, _07544_, _10028_);
  and _69523_ (_18209_, _18208_, _17922_);
  or _69524_ (_18210_, _18209_, _18207_);
  nor _69525_ (_18211_, _10975_, _18210_);
  and _69526_ (_18213_, _10975_, _18210_);
  nor _69527_ (_18214_, _18213_, _18211_);
  and _69528_ (_18215_, _18214_, \oc8051_golden_model_1.PSW [7]);
  nor _69529_ (_18216_, _18214_, \oc8051_golden_model_1.PSW [7]);
  nor _69530_ (_18217_, _18216_, _18215_);
  and _69531_ (_18218_, _18217_, _18206_);
  nor _69532_ (_18219_, _18217_, _18206_);
  nor _69533_ (_18220_, _18219_, _18218_);
  and _69534_ (_18221_, _18220_, _10557_);
  or _69535_ (_18222_, _10458_, _08336_);
  nor _69536_ (_18224_, _08409_, _09902_);
  and _69537_ (_18225_, _14932_, _08409_);
  or _69538_ (_18226_, _18225_, _18224_);
  or _69539_ (_18227_, _18226_, _06157_);
  and _69540_ (_18228_, _18227_, _07075_);
  and _69541_ (_18229_, _14928_, _07809_);
  or _69542_ (_18230_, _18229_, _18184_);
  and _69543_ (_18231_, _18230_, _06160_);
  or _69544_ (_18232_, _10474_, _09209_);
  and _69545_ (_18233_, _17011_, _08336_);
  or _69546_ (_18235_, _06653_, \oc8051_golden_model_1.ACC [4]);
  nand _69547_ (_18236_, _06653_, \oc8051_golden_model_1.ACC [4]);
  and _69548_ (_18237_, _18236_, _18235_);
  and _69549_ (_18238_, _18237_, _10471_);
  or _69550_ (_18239_, _18238_, _10473_);
  or _69551_ (_18240_, _18239_, _18233_);
  and _69552_ (_18241_, _18240_, _10484_);
  and _69553_ (_18242_, _18241_, _18232_);
  or _69554_ (_18243_, _18242_, _18231_);
  and _69555_ (_18244_, _18243_, _10491_);
  nor _69556_ (_18246_, _10494_, \oc8051_golden_model_1.ACC [4]);
  nor _69557_ (_18247_, _18246_, _10495_);
  and _69558_ (_18248_, _18247_, _10490_);
  or _69559_ (_18249_, _18248_, _06156_);
  or _69560_ (_18250_, _18249_, _18244_);
  and _69561_ (_18251_, _18250_, _18228_);
  and _69562_ (_18252_, _18186_, _06217_);
  or _69563_ (_18253_, _18252_, _10516_);
  or _69564_ (_18254_, _18253_, _18251_);
  and _69565_ (_18255_, _18254_, _18222_);
  or _69566_ (_18257_, _18255_, _07081_);
  or _69567_ (_18258_, _09209_, _07082_);
  and _69568_ (_18259_, _18258_, _06229_);
  and _69569_ (_18260_, _18259_, _18257_);
  nor _69570_ (_18261_, _08338_, _06229_);
  or _69571_ (_18262_, _18261_, _10525_);
  or _69572_ (_18263_, _18262_, _18260_);
  nand _69573_ (_18264_, _10525_, _05855_);
  and _69574_ (_18265_, _18264_, _18263_);
  or _69575_ (_18266_, _18265_, _06152_);
  and _69576_ (_18268_, _14942_, _08409_);
  or _69577_ (_18269_, _18268_, _18224_);
  or _69578_ (_18270_, _18269_, _06153_);
  and _69579_ (_18271_, _18270_, _06146_);
  and _69580_ (_18272_, _18271_, _18266_);
  or _69581_ (_18273_, _18224_, _14949_);
  and _69582_ (_18274_, _18226_, _06145_);
  and _69583_ (_18275_, _18274_, _18273_);
  or _69584_ (_18276_, _18275_, _09295_);
  or _69585_ (_18277_, _18276_, _18272_);
  nor _69586_ (_18279_, _09780_, _09778_);
  nor _69587_ (_18280_, _18279_, _09781_);
  or _69588_ (_18281_, _18280_, _09301_);
  and _69589_ (_18282_, _18281_, _10554_);
  and _69590_ (_18283_, _18282_, _18277_);
  or _69591_ (_18284_, _18283_, _18221_);
  and _69592_ (_18285_, _18284_, _12380_);
  or _69593_ (_18286_, _18285_, _18205_);
  and _69594_ (_18287_, _18286_, _06265_);
  nor _69595_ (_18288_, _12324_, _10693_);
  or _69596_ (_18290_, _17956_, _13917_);
  and _69597_ (_18291_, _18290_, _13915_);
  nor _69598_ (_18292_, _18291_, _10289_);
  and _69599_ (_18293_, _18291_, _10289_);
  nor _69600_ (_18294_, _18293_, _18292_);
  and _69601_ (_18295_, _18294_, \oc8051_golden_model_1.PSW [7]);
  nor _69602_ (_18296_, _18294_, \oc8051_golden_model_1.PSW [7]);
  nor _69603_ (_18297_, _18296_, _18295_);
  or _69604_ (_18298_, _18297_, _18288_);
  and _69605_ (_18299_, _18297_, _18288_);
  nor _69606_ (_18301_, _18299_, _06265_);
  and _69607_ (_18302_, _18301_, _18298_);
  or _69608_ (_18303_, _18302_, _18287_);
  and _69609_ (_18304_, _18303_, _10388_);
  nor _69610_ (_18305_, _12341_, _10693_);
  or _69611_ (_18306_, _17970_, _13950_);
  and _69612_ (_18307_, _18306_, _13949_);
  nor _69613_ (_18308_, _11058_, _18307_);
  and _69614_ (_18309_, _11058_, _18307_);
  nor _69615_ (_18310_, _18309_, _18308_);
  and _69616_ (_18312_, _18310_, \oc8051_golden_model_1.PSW [7]);
  nor _69617_ (_18313_, _18310_, \oc8051_golden_model_1.PSW [7]);
  nor _69618_ (_18314_, _18313_, _18312_);
  or _69619_ (_18315_, _18314_, _18305_);
  and _69620_ (_18316_, _18314_, _18305_);
  nor _69621_ (_18317_, _18316_, _10388_);
  and _69622_ (_18318_, _18317_, _18315_);
  or _69623_ (_18319_, _18318_, _05870_);
  or _69624_ (_18320_, _18319_, _18304_);
  nand _69625_ (_18321_, _06876_, _05870_);
  and _69626_ (_18323_, _18321_, _06140_);
  and _69627_ (_18324_, _18323_, _18320_);
  and _69628_ (_18325_, _14966_, _08409_);
  or _69629_ (_18326_, _18325_, _18224_);
  and _69630_ (_18327_, _18326_, _06139_);
  or _69631_ (_18328_, _18327_, _09842_);
  or _69632_ (_18329_, _18328_, _18324_);
  and _69633_ (_18330_, _18329_, _18187_);
  or _69634_ (_18331_, _18330_, _06116_);
  and _69635_ (_18332_, _09209_, _07809_);
  or _69636_ (_18334_, _18184_, _06117_);
  or _69637_ (_18335_, _18334_, _18332_);
  and _69638_ (_18336_, _18335_, _06114_);
  and _69639_ (_18337_, _18336_, _18331_);
  and _69640_ (_18338_, _15013_, _07809_);
  or _69641_ (_18339_, _18338_, _18184_);
  and _69642_ (_18340_, _18339_, _05787_);
  or _69643_ (_18341_, _18340_, _09855_);
  or _69644_ (_18342_, _18341_, _18337_);
  or _69645_ (_18343_, _09947_, _09861_);
  and _69646_ (_18345_, _18343_, _05802_);
  and _69647_ (_18346_, _18345_, _18342_);
  nor _69648_ (_18347_, _06876_, _05802_);
  or _69649_ (_18348_, _18347_, _06110_);
  or _69650_ (_18349_, _18348_, _18346_);
  and _69651_ (_18350_, _08715_, _07809_);
  or _69652_ (_18351_, _18350_, _18184_);
  or _69653_ (_18352_, _18351_, _06111_);
  and _69654_ (_18353_, _18352_, _10752_);
  and _69655_ (_18354_, _18353_, _18349_);
  or _69656_ (_18356_, _18354_, _18183_);
  and _69657_ (_18357_, _18356_, _18182_);
  and _69658_ (_18358_, _10975_, _18181_);
  nor _69659_ (_18359_, _18358_, _18357_);
  nand _69660_ (_18360_, _18359_, _18180_);
  or _69661_ (_18361_, _18180_, _10975_);
  and _69662_ (_18362_, _18361_, _10776_);
  and _69663_ (_18363_, _18362_, _18360_);
  and _69664_ (_18364_, _10775_, _11015_);
  or _69665_ (_18365_, _18364_, _06400_);
  or _69666_ (_18366_, _18365_, _18363_);
  or _69667_ (_18367_, _10289_, _06401_);
  and _69668_ (_18368_, _18367_, _18366_);
  and _69669_ (_18369_, _18368_, _10788_);
  and _69670_ (_18370_, _10787_, _11058_);
  or _69671_ (_18371_, _18370_, _06297_);
  or _69672_ (_18372_, _18371_, _18369_);
  and _69673_ (_18373_, _15029_, _07809_);
  or _69674_ (_18374_, _18184_, _07127_);
  or _69675_ (_18375_, _18374_, _18373_);
  and _69676_ (_18377_, _18375_, _07125_);
  and _69677_ (_18378_, _18377_, _18372_);
  and _69678_ (_18379_, _18184_, _06402_);
  or _69679_ (_18380_, _18379_, _06557_);
  or _69680_ (_18381_, _18380_, _18378_);
  and _69681_ (_18382_, _10972_, _05742_);
  or _69682_ (_18383_, _18382_, _17408_);
  and _69683_ (_18384_, _18383_, _17417_);
  and _69684_ (_18385_, _18384_, _18381_);
  or _69685_ (_18386_, _18385_, _18171_);
  and _69686_ (_18388_, _18386_, _17416_);
  and _69687_ (_18389_, _10807_, _10972_);
  or _69688_ (_18390_, _18389_, _10811_);
  or _69689_ (_18391_, _18390_, _18388_);
  or _69690_ (_18392_, _10816_, _11012_);
  and _69691_ (_18393_, _18392_, _06410_);
  and _69692_ (_18394_, _18393_, _18391_);
  or _69693_ (_18395_, _10820_, _10270_);
  and _69694_ (_18396_, _18395_, _10822_);
  or _69695_ (_18397_, _18396_, _18394_);
  or _69696_ (_18399_, _10826_, _11055_);
  and _69697_ (_18400_, _18399_, _07132_);
  and _69698_ (_18401_, _18400_, _18397_);
  nand _69699_ (_18402_, _18351_, _06306_);
  nor _69700_ (_18403_, _18402_, _10288_);
  or _69701_ (_18404_, _18403_, _06524_);
  or _69702_ (_18405_, _18404_, _18401_);
  not _69703_ (_18406_, _06524_);
  or _69704_ (_18407_, _10973_, _18406_);
  and _69705_ (_18408_, _18407_, _10837_);
  and _69706_ (_18410_, _18408_, _18405_);
  not _69707_ (_18411_, _10837_);
  and _69708_ (_18412_, _18411_, _10973_);
  or _69709_ (_18413_, _18412_, _10841_);
  or _69710_ (_18414_, _18413_, _18410_);
  or _69711_ (_18415_, _17242_, _11014_);
  and _69712_ (_18416_, _18415_, _06395_);
  and _69713_ (_18417_, _18416_, _18414_);
  nand _69714_ (_18418_, _10851_, _10288_);
  and _69715_ (_18419_, _18418_, _10850_);
  or _69716_ (_18421_, _18419_, _18417_);
  and _69717_ (_18422_, _18421_, _18169_);
  or _69718_ (_18423_, _18422_, _06303_);
  and _69719_ (_18424_, _15026_, _07809_);
  or _69720_ (_18425_, _18184_, _08819_);
  or _69721_ (_18426_, _18425_, _18424_);
  and _69722_ (_18427_, _18426_, _10380_);
  and _69723_ (_18428_, _18427_, _18423_);
  or _69724_ (_18429_, _10361_, _10330_);
  and _69725_ (_18430_, _18429_, _10362_);
  and _69726_ (_18432_, _18430_, _10858_);
  or _69727_ (_18433_, _18432_, _17240_);
  or _69728_ (_18434_, _18433_, _18428_);
  or _69729_ (_18435_, _10882_, _10606_);
  and _69730_ (_18436_, _18435_, _10883_);
  and _69731_ (_18437_, _18436_, _06276_);
  or _69732_ (_18438_, _18437_, _10867_);
  and _69733_ (_18439_, _18438_, _18434_);
  and _69734_ (_18440_, _18436_, _06792_);
  or _69735_ (_18441_, _18440_, _06406_);
  or _69736_ (_18443_, _18441_, _18439_);
  and _69737_ (_18444_, _18443_, _18168_);
  or _69738_ (_18445_, _10942_, _10679_);
  and _69739_ (_18446_, _10943_, _10895_);
  and _69740_ (_18447_, _18446_, _18445_);
  or _69741_ (_18448_, _18447_, _10925_);
  or _69742_ (_18449_, _18448_, _18444_);
  nand _69743_ (_18450_, _10925_, _10028_);
  and _69744_ (_18451_, _18450_, _10963_);
  and _69745_ (_18452_, _18451_, _18449_);
  not _69746_ (_18454_, _10963_);
  nor _69747_ (_18455_, _10991_, _10975_);
  nor _69748_ (_18456_, _18455_, _10992_);
  and _69749_ (_18457_, _18456_, _18454_);
  or _69750_ (_18458_, _18457_, _17195_);
  or _69751_ (_18459_, _18458_, _18452_);
  and _69752_ (_18460_, _18459_, _18164_);
  or _69753_ (_18461_, _18460_, _17199_);
  or _69754_ (_18462_, _18163_, _17200_);
  and _69755_ (_18463_, _18462_, _06171_);
  and _69756_ (_18465_, _18463_, _18461_);
  or _69757_ (_18466_, _18465_, _18161_);
  and _69758_ (_18467_, _18466_, _10265_);
  or _69759_ (_18468_, _11074_, _11058_);
  and _69760_ (_18469_, _11075_, _10264_);
  and _69761_ (_18470_, _18469_, _18468_);
  or _69762_ (_18471_, _18470_, _10262_);
  or _69763_ (_18472_, _18471_, _18467_);
  and _69764_ (_18473_, _18472_, _18158_);
  or _69765_ (_18474_, _18473_, _06433_);
  or _69766_ (_18476_, _18230_, _06829_);
  and _69767_ (_18477_, _18476_, _11090_);
  and _69768_ (_18478_, _18477_, _18474_);
  nor _69769_ (_18479_, _11096_, _09902_);
  or _69770_ (_18480_, _18479_, _11097_);
  and _69771_ (_18481_, _18480_, _11089_);
  or _69772_ (_18482_, _18481_, _11094_);
  or _69773_ (_18483_, _18482_, _18478_);
  nand _69774_ (_18484_, _11094_, _09930_);
  and _69775_ (_18485_, _18484_, _05749_);
  and _69776_ (_18487_, _18485_, _18483_);
  and _69777_ (_18488_, _18269_, _05748_);
  or _69778_ (_18489_, _18488_, _06440_);
  or _69779_ (_18490_, _18489_, _18487_);
  and _69780_ (_18491_, _15087_, _07809_);
  or _69781_ (_18492_, _18184_, _06444_);
  or _69782_ (_18493_, _18492_, _18491_);
  and _69783_ (_18494_, _18493_, _11113_);
  and _69784_ (_18495_, _18494_, _18490_);
  nor _69785_ (_18496_, _11122_, \oc8051_golden_model_1.ACC [4]);
  nor _69786_ (_18498_, _18496_, _11123_);
  and _69787_ (_18499_, _18498_, _11112_);
  or _69788_ (_18500_, _18499_, _11119_);
  or _69789_ (_18501_, _18500_, _18495_);
  nand _69790_ (_18502_, _11119_, _09930_);
  and _69791_ (_18503_, _18502_, _01317_);
  and _69792_ (_18504_, _18503_, _18501_);
  or _69793_ (_18505_, _18504_, _18157_);
  and _69794_ (_43607_, _18505_, _43100_);
  nor _69795_ (_18506_, _01317_, _09930_);
  and _69796_ (_18508_, _10363_, _10323_);
  nor _69797_ (_18509_, _18508_, _10364_);
  or _69798_ (_18510_, _18509_, _10380_);
  and _69799_ (_18511_, _15219_, _07809_);
  nor _69800_ (_18512_, _07809_, _09930_);
  or _69801_ (_18513_, _18512_, _07127_);
  or _69802_ (_18514_, _18513_, _18511_);
  nor _69803_ (_18515_, _10971_, _10970_);
  nor _69804_ (_18516_, _18178_, _10772_);
  not _69805_ (_18517_, _18516_);
  and _69806_ (_18519_, _18517_, _18515_);
  nor _69807_ (_18520_, _10752_, _06477_);
  and _69808_ (_18521_, _08101_, _07809_);
  or _69809_ (_18522_, _18521_, _18512_);
  or _69810_ (_18523_, _18522_, _06132_);
  and _69811_ (_18524_, _06876_, \oc8051_golden_model_1.ACC [4]);
  nor _69812_ (_18525_, _18308_, _18524_);
  nor _69813_ (_18526_, _12342_, _18525_);
  and _69814_ (_18527_, _12342_, _18525_);
  nor _69815_ (_18528_, _18527_, _18526_);
  and _69816_ (_18530_, _18528_, \oc8051_golden_model_1.PSW [7]);
  nor _69817_ (_18531_, _18528_, \oc8051_golden_model_1.PSW [7]);
  nor _69818_ (_18532_, _18531_, _18530_);
  nor _69819_ (_18533_, _18316_, _18312_);
  not _69820_ (_18534_, _18533_);
  and _69821_ (_18535_, _18534_, _18532_);
  nor _69822_ (_18536_, _18534_, _18532_);
  nor _69823_ (_18537_, _18536_, _18535_);
  or _69824_ (_18538_, _18537_, _10388_);
  and _69825_ (_18539_, _08980_, \oc8051_golden_model_1.ACC [4]);
  nor _69826_ (_18541_, _18194_, _18539_);
  or _69827_ (_18542_, _11011_, _18541_);
  nand _69828_ (_18543_, _11011_, _18541_);
  and _69829_ (_18544_, _18543_, _18542_);
  or _69830_ (_18545_, _18544_, _10693_);
  nand _69831_ (_18546_, _18544_, _10693_);
  and _69832_ (_18547_, _18546_, _18545_);
  nand _69833_ (_18548_, _18203_, _18198_);
  nand _69834_ (_18549_, _18548_, _18547_);
  or _69835_ (_18550_, _18548_, _18547_);
  and _69836_ (_18552_, _18550_, _18549_);
  or _69837_ (_18553_, _18552_, _12380_);
  or _69838_ (_18554_, _10458_, _08101_);
  or _69839_ (_18555_, _10474_, _09208_);
  and _69840_ (_18556_, _17011_, _08101_);
  or _69841_ (_18557_, _06653_, \oc8051_golden_model_1.ACC [5]);
  nand _69842_ (_18558_, _06653_, \oc8051_golden_model_1.ACC [5]);
  and _69843_ (_18559_, _18558_, _18557_);
  and _69844_ (_18560_, _18559_, _10471_);
  or _69845_ (_18561_, _18560_, _10473_);
  or _69846_ (_18563_, _18561_, _18556_);
  and _69847_ (_18564_, _18563_, _10484_);
  and _69848_ (_18565_, _18564_, _18555_);
  and _69849_ (_18566_, _15119_, _07809_);
  or _69850_ (_18567_, _18566_, _18512_);
  and _69851_ (_18568_, _18567_, _06160_);
  or _69852_ (_18569_, _18568_, _10490_);
  or _69853_ (_18570_, _18569_, _18565_);
  nor _69854_ (_18571_, _13858_, _10502_);
  nand _69855_ (_18572_, _13858_, _10502_);
  nand _69856_ (_18574_, _18572_, _10490_);
  or _69857_ (_18575_, _18574_, _18571_);
  and _69858_ (_18576_, _18575_, _06221_);
  and _69859_ (_18577_, _18576_, _18570_);
  nor _69860_ (_18578_, _08409_, _09930_);
  and _69861_ (_18579_, _15123_, _08409_);
  or _69862_ (_18580_, _18579_, _18578_);
  and _69863_ (_18581_, _18580_, _06156_);
  and _69864_ (_18582_, _18522_, _06217_);
  or _69865_ (_18583_, _18582_, _10516_);
  or _69866_ (_18585_, _18583_, _18581_);
  or _69867_ (_18586_, _18585_, _18577_);
  and _69868_ (_18587_, _18586_, _18554_);
  or _69869_ (_18588_, _18587_, _07081_);
  or _69870_ (_18589_, _09208_, _07082_);
  and _69871_ (_18590_, _18589_, _06229_);
  and _69872_ (_18591_, _18590_, _18588_);
  nor _69873_ (_18592_, _08103_, _06229_);
  or _69874_ (_18593_, _18592_, _10525_);
  or _69875_ (_18594_, _18593_, _18591_);
  nand _69876_ (_18596_, _10525_, _05887_);
  and _69877_ (_18597_, _18596_, _18594_);
  or _69878_ (_18598_, _18597_, _06152_);
  and _69879_ (_18599_, _15104_, _08409_);
  or _69880_ (_18600_, _18599_, _18578_);
  or _69881_ (_18601_, _18600_, _06153_);
  and _69882_ (_18602_, _18601_, _06146_);
  and _69883_ (_18603_, _18602_, _18598_);
  or _69884_ (_18604_, _18578_, _15138_);
  and _69885_ (_18605_, _18580_, _06145_);
  and _69886_ (_18607_, _18605_, _18604_);
  or _69887_ (_18608_, _18607_, _18603_);
  and _69888_ (_18609_, _18608_, _09301_);
  or _69889_ (_18610_, _09783_, _09781_);
  nor _69890_ (_18611_, _09784_, _09301_);
  and _69891_ (_18612_, _18611_, _18610_);
  nor _69892_ (_18613_, _06129_, _05803_);
  or _69893_ (_18614_, _18613_, _10547_);
  or _69894_ (_18615_, _18614_, _18612_);
  or _69895_ (_18616_, _18615_, _18609_);
  and _69896_ (_18618_, _06119_, _05790_);
  not _69897_ (_18619_, _18618_);
  and _69898_ (_18620_, _08349_, \oc8051_golden_model_1.ACC [4]);
  nor _69899_ (_18621_, _18211_, _18620_);
  nor _69900_ (_18622_, _18515_, _18621_);
  and _69901_ (_18623_, _18515_, _18621_);
  nor _69902_ (_18624_, _18623_, _18622_);
  and _69903_ (_18625_, _18624_, \oc8051_golden_model_1.PSW [7]);
  nor _69904_ (_18626_, _18624_, \oc8051_golden_model_1.PSW [7]);
  nor _69905_ (_18627_, _18626_, _18625_);
  nor _69906_ (_18629_, _18218_, _18215_);
  not _69907_ (_18630_, _18629_);
  and _69908_ (_18631_, _18630_, _18627_);
  nor _69909_ (_18632_, _18630_, _18627_);
  nor _69910_ (_18633_, _18632_, _18631_);
  and _69911_ (_18634_, _18633_, _18619_);
  or _69912_ (_18635_, _18634_, _10554_);
  and _69913_ (_18636_, _18635_, _18616_);
  and _69914_ (_18637_, _18633_, _18618_);
  or _69915_ (_18638_, _18637_, _12379_);
  or _69916_ (_18640_, _18638_, _18636_);
  and _69917_ (_18641_, _18640_, _06265_);
  and _69918_ (_18642_, _18641_, _18553_);
  and _69919_ (_18643_, _08338_, \oc8051_golden_model_1.ACC [4]);
  nor _69920_ (_18644_, _18292_, _18643_);
  nor _69921_ (_18645_, _18644_, _12325_);
  and _69922_ (_18646_, _18644_, _12325_);
  nor _69923_ (_18647_, _18646_, _18645_);
  and _69924_ (_18648_, _18647_, \oc8051_golden_model_1.PSW [7]);
  nor _69925_ (_18649_, _18647_, \oc8051_golden_model_1.PSW [7]);
  nor _69926_ (_18651_, _18649_, _18648_);
  nor _69927_ (_18652_, _18299_, _18295_);
  not _69928_ (_18653_, _18652_);
  or _69929_ (_18654_, _18653_, _18651_);
  and _69930_ (_18655_, _18653_, _18651_);
  nor _69931_ (_18656_, _18655_, _06265_);
  and _69932_ (_18657_, _18656_, _18654_);
  or _69933_ (_18658_, _18657_, _10387_);
  or _69934_ (_18659_, _18658_, _18642_);
  and _69935_ (_18660_, _18659_, _18538_);
  or _69936_ (_18661_, _18660_, _05870_);
  nand _69937_ (_18662_, _06477_, _05870_);
  and _69938_ (_18663_, _18662_, _06140_);
  and _69939_ (_18664_, _18663_, _18661_);
  and _69940_ (_18665_, _15155_, _08409_);
  or _69941_ (_18666_, _18665_, _18578_);
  and _69942_ (_18667_, _18666_, _06139_);
  or _69943_ (_18668_, _18667_, _09842_);
  or _69944_ (_18669_, _18668_, _18664_);
  and _69945_ (_18670_, _18669_, _18523_);
  or _69946_ (_18673_, _18670_, _06116_);
  and _69947_ (_18674_, _09208_, _07809_);
  or _69948_ (_18675_, _18512_, _06117_);
  or _69949_ (_18676_, _18675_, _18674_);
  and _69950_ (_18677_, _18676_, _06114_);
  and _69951_ (_18678_, _18677_, _18673_);
  and _69952_ (_18679_, _15203_, _07809_);
  or _69953_ (_18680_, _18679_, _18512_);
  and _69954_ (_18681_, _18680_, _05787_);
  or _69955_ (_18682_, _18681_, _09855_);
  or _69956_ (_18684_, _18682_, _18678_);
  or _69957_ (_18685_, _09916_, _09861_);
  and _69958_ (_18686_, _18685_, _05802_);
  and _69959_ (_18687_, _18686_, _18684_);
  nor _69960_ (_18688_, _06477_, _05802_);
  or _69961_ (_18689_, _18688_, _06110_);
  or _69962_ (_18690_, _18689_, _18687_);
  and _69963_ (_18691_, _08736_, _07809_);
  or _69964_ (_18692_, _18691_, _18512_);
  or _69965_ (_18693_, _18692_, _06111_);
  and _69966_ (_18694_, _18693_, _10752_);
  and _69967_ (_18695_, _18694_, _18690_);
  or _69968_ (_18696_, _18695_, _18520_);
  and _69969_ (_18697_, _18696_, _10762_);
  and _69970_ (_18698_, _18515_, _06558_);
  or _69971_ (_18699_, _18698_, _06574_);
  or _69972_ (_18700_, _18699_, _18697_);
  not _69973_ (_18701_, _06574_);
  or _69974_ (_18702_, _18515_, _18701_);
  and _69975_ (_18703_, _18702_, _18516_);
  and _69976_ (_18706_, _18703_, _18700_);
  or _69977_ (_18707_, _18706_, _18519_);
  and _69978_ (_18708_, _18707_, _10776_);
  nor _69979_ (_18709_, _10776_, _11011_);
  or _69980_ (_18710_, _18709_, _06400_);
  or _69981_ (_18711_, _18710_, _18708_);
  or _69982_ (_18712_, _12325_, _06401_);
  and _69983_ (_18713_, _18712_, _10788_);
  and _69984_ (_18714_, _18713_, _18711_);
  and _69985_ (_18715_, _10787_, _12342_);
  or _69986_ (_18717_, _18715_, _06297_);
  or _69987_ (_18718_, _18717_, _18714_);
  and _69988_ (_18719_, _18718_, _18514_);
  or _69989_ (_18720_, _18719_, _06402_);
  and _69990_ (_18721_, _06957_, _06408_);
  not _69991_ (_18722_, _18721_);
  and _69992_ (_18723_, _06684_, _06408_);
  and _69993_ (_18724_, _06288_, _06408_);
  nor _69994_ (_18725_, _18724_, _18723_);
  and _69995_ (_18726_, _18725_, _18722_);
  and _69996_ (_18727_, _18726_, _17408_);
  or _69997_ (_18728_, _18512_, _07125_);
  and _69998_ (_18729_, _18728_, _18727_);
  and _69999_ (_18730_, _18729_, _18720_);
  and _70000_ (_18731_, _06273_, _06408_);
  or _70001_ (_18732_, _10970_, _18731_);
  and _70002_ (_18733_, _18732_, _10812_);
  or _70003_ (_18734_, _18733_, _18730_);
  not _70004_ (_18735_, _18731_);
  or _70005_ (_18736_, _10970_, _18735_);
  and _70006_ (_18739_, _18736_, _18734_);
  or _70007_ (_18740_, _18739_, _10811_);
  or _70008_ (_18741_, _10816_, _11009_);
  and _70009_ (_18742_, _18741_, _06410_);
  and _70010_ (_18743_, _18742_, _18740_);
  or _70011_ (_18744_, _10820_, _10268_);
  and _70012_ (_18745_, _18744_, _10822_);
  or _70013_ (_18746_, _18745_, _18743_);
  or _70014_ (_18747_, _10826_, _11053_);
  and _70015_ (_18748_, _18747_, _07132_);
  and _70016_ (_18750_, _18748_, _18746_);
  nand _70017_ (_18751_, _18692_, _06306_);
  nor _70018_ (_18752_, _18751_, _10269_);
  or _70019_ (_18753_, _18752_, _06524_);
  or _70020_ (_18754_, _18753_, _18750_);
  nand _70021_ (_18755_, _10971_, _06524_);
  and _70022_ (_18756_, _18755_, _17150_);
  and _70023_ (_18757_, _18756_, _18754_);
  nor _70024_ (_18758_, _17150_, _10971_);
  or _70025_ (_18759_, _18758_, _17156_);
  or _70026_ (_18760_, _18759_, _18757_);
  nand _70027_ (_18761_, _17156_, _10971_);
  and _70028_ (_18762_, _18761_, _17161_);
  and _70029_ (_18763_, _18762_, _18760_);
  nor _70030_ (_18764_, _10971_, _17161_);
  or _70031_ (_18765_, _18764_, _10841_);
  or _70032_ (_18766_, _18765_, _18763_);
  nand _70033_ (_18767_, _10841_, _09930_);
  or _70034_ (_18768_, _18767_, _09208_);
  and _70035_ (_18769_, _18768_, _06395_);
  and _70036_ (_18772_, _18769_, _18766_);
  nand _70037_ (_18773_, _10851_, _10269_);
  and _70038_ (_18774_, _18773_, _10850_);
  or _70039_ (_18775_, _18774_, _18772_);
  nand _70040_ (_18776_, _10848_, _11054_);
  and _70041_ (_18777_, _18776_, _08819_);
  and _70042_ (_18778_, _18777_, _18775_);
  and _70043_ (_18779_, _15216_, _07809_);
  or _70044_ (_18780_, _18779_, _18512_);
  and _70045_ (_18781_, _18780_, _06303_);
  or _70046_ (_18783_, _18781_, _10858_);
  or _70047_ (_18784_, _18783_, _18778_);
  and _70048_ (_18785_, _18784_, _18510_);
  or _70049_ (_18786_, _18785_, _10865_);
  and _70050_ (_18787_, _10884_, _10599_);
  nor _70051_ (_18788_, _18787_, _10885_);
  or _70052_ (_18789_, _18788_, _10867_);
  and _70053_ (_18790_, _18789_, _06407_);
  and _70054_ (_18791_, _18790_, _18786_);
  and _70055_ (_18792_, _10914_, _10410_);
  nor _70056_ (_18793_, _18792_, _10915_);
  or _70057_ (_18794_, _18793_, _10895_);
  and _70058_ (_18795_, _18794_, _10897_);
  or _70059_ (_18796_, _18795_, _18791_);
  and _70060_ (_18797_, _10944_, _10676_);
  nor _70061_ (_18798_, _18797_, _10945_);
  or _70062_ (_18799_, _18798_, _10927_);
  and _70063_ (_18800_, _18799_, _10926_);
  and _70064_ (_18801_, _18800_, _18796_);
  nand _70065_ (_18802_, _10925_, \oc8051_golden_model_1.ACC [4]);
  nand _70066_ (_18805_, _18802_, _10963_);
  or _70067_ (_18806_, _18805_, _18801_);
  and _70068_ (_18807_, _10993_, _18515_);
  nor _70069_ (_18808_, _10993_, _18515_);
  or _70070_ (_18809_, _18808_, _18807_);
  or _70071_ (_18810_, _18809_, _10963_);
  and _70072_ (_18811_, _18810_, _18806_);
  or _70073_ (_18812_, _18811_, _11003_);
  and _70074_ (_18813_, _11035_, _11011_);
  nor _70075_ (_18814_, _18813_, _11036_);
  or _70076_ (_18816_, _18814_, _11041_);
  and _70077_ (_18817_, _18816_, _06171_);
  and _70078_ (_18818_, _18817_, _18812_);
  and _70079_ (_18819_, _12325_, _10291_);
  nor _70080_ (_18820_, _12325_, _10291_);
  or _70081_ (_18821_, _18820_, _10264_);
  or _70082_ (_18822_, _18821_, _18819_);
  and _70083_ (_18823_, _18822_, _12691_);
  or _70084_ (_18824_, _18823_, _18818_);
  and _70085_ (_18825_, _11076_, _12342_);
  nor _70086_ (_18826_, _11076_, _12342_);
  or _70087_ (_18827_, _18826_, _10265_);
  or _70088_ (_18828_, _18827_, _18825_);
  and _70089_ (_18829_, _18828_, _12693_);
  and _70090_ (_18830_, _18829_, _18824_);
  and _70091_ (_18831_, _10262_, \oc8051_golden_model_1.ACC [4]);
  or _70092_ (_18832_, _18831_, _06433_);
  or _70093_ (_18833_, _18832_, _18830_);
  or _70094_ (_18834_, _18567_, _06829_);
  and _70095_ (_18835_, _18834_, _11090_);
  and _70096_ (_18838_, _18835_, _18833_);
  nor _70097_ (_18839_, _11097_, _09930_);
  or _70098_ (_18840_, _18839_, _11098_);
  and _70099_ (_18841_, _18840_, _11089_);
  or _70100_ (_18842_, _18841_, _11094_);
  or _70101_ (_18843_, _18842_, _18838_);
  nand _70102_ (_18844_, _11094_, _09883_);
  and _70103_ (_18845_, _18844_, _05749_);
  and _70104_ (_18846_, _18845_, _18843_);
  and _70105_ (_18847_, _18600_, _05748_);
  or _70106_ (_18849_, _18847_, _06440_);
  or _70107_ (_18850_, _18849_, _18846_);
  and _70108_ (_18851_, _15275_, _07809_);
  or _70109_ (_18852_, _18512_, _06444_);
  or _70110_ (_18853_, _18852_, _18851_);
  and _70111_ (_18854_, _18853_, _11113_);
  and _70112_ (_18855_, _18854_, _18850_);
  nor _70113_ (_18856_, _11123_, \oc8051_golden_model_1.ACC [5]);
  nor _70114_ (_18857_, _18856_, _11124_);
  and _70115_ (_18858_, _18857_, _11112_);
  or _70116_ (_18859_, _18858_, _11119_);
  or _70117_ (_18860_, _18859_, _18855_);
  nand _70118_ (_18861_, _11119_, _09883_);
  and _70119_ (_18862_, _18861_, _01317_);
  and _70120_ (_18863_, _18862_, _18860_);
  or _70121_ (_18864_, _18863_, _18506_);
  and _70122_ (_43608_, _18864_, _43100_);
  nor _70123_ (_18865_, _01317_, _09883_);
  nor _70124_ (_18866_, _11037_, _11008_);
  nor _70125_ (_18867_, _18866_, _11038_);
  or _70126_ (_18870_, _18867_, _17201_);
  nor _70127_ (_18871_, _10916_, _10448_);
  nor _70128_ (_18872_, _18871_, _10917_);
  or _70129_ (_18873_, _18872_, _06407_);
  and _70130_ (_18874_, _18873_, _10927_);
  nand _70131_ (_18875_, _10848_, _11051_);
  or _70132_ (_18876_, _10967_, _18406_);
  and _70133_ (_18877_, _15413_, _07809_);
  nor _70134_ (_18878_, _07809_, _09883_);
  or _70135_ (_18879_, _18878_, _07127_);
  or _70136_ (_18881_, _18879_, _18877_);
  and _70137_ (_18882_, _18178_, _10969_);
  and _70138_ (_18883_, _15395_, _07809_);
  or _70139_ (_18884_, _18883_, _18878_);
  and _70140_ (_18885_, _18884_, _05787_);
  and _70141_ (_18886_, _08012_, _07809_);
  or _70142_ (_18887_, _18886_, _18878_);
  or _70143_ (_18888_, _18887_, _06132_);
  or _70144_ (_18889_, _09208_, _09930_);
  and _70145_ (_18890_, _09208_, _09930_);
  or _70146_ (_18892_, _18541_, _18890_);
  and _70147_ (_18893_, _18892_, _18889_);
  nor _70148_ (_18894_, _18893_, _11008_);
  and _70149_ (_18895_, _18893_, _11008_);
  nor _70150_ (_18896_, _18895_, _18894_);
  and _70151_ (_18897_, _18549_, _18545_);
  nand _70152_ (_18898_, _18897_, \oc8051_golden_model_1.PSW [7]);
  nor _70153_ (_18899_, _18898_, _18896_);
  and _70154_ (_18900_, _18898_, _18896_);
  or _70155_ (_18901_, _18900_, _18899_);
  or _70156_ (_18903_, _18901_, _12380_);
  or _70157_ (_18904_, _10458_, _08012_);
  or _70158_ (_18905_, _10474_, _09207_);
  and _70159_ (_18906_, _17011_, _08012_);
  or _70160_ (_18907_, _06653_, \oc8051_golden_model_1.ACC [6]);
  nand _70161_ (_18908_, _06653_, \oc8051_golden_model_1.ACC [6]);
  and _70162_ (_18909_, _18908_, _18907_);
  and _70163_ (_18910_, _18909_, _10471_);
  or _70164_ (_18911_, _18910_, _10473_);
  or _70165_ (_18912_, _18911_, _18906_);
  and _70166_ (_18914_, _18912_, _10484_);
  and _70167_ (_18915_, _18914_, _18905_);
  and _70168_ (_18916_, _15300_, _07809_);
  or _70169_ (_18917_, _18916_, _18878_);
  and _70170_ (_18918_, _18917_, _06160_);
  or _70171_ (_18919_, _18918_, _10490_);
  or _70172_ (_18920_, _18919_, _18915_);
  not _70173_ (_18921_, _10504_);
  nor _70174_ (_18922_, _18571_, _18921_);
  nand _70175_ (_18923_, _10508_, _10505_);
  nand _70176_ (_18925_, _18923_, _10490_);
  or _70177_ (_18926_, _18925_, _18922_);
  and _70178_ (_18927_, _18926_, _06221_);
  and _70179_ (_18928_, _18927_, _18920_);
  nor _70180_ (_18929_, _08409_, _09883_);
  and _70181_ (_18930_, _15316_, _08409_);
  or _70182_ (_18931_, _18930_, _18929_);
  and _70183_ (_18932_, _18931_, _06156_);
  and _70184_ (_18933_, _18887_, _06217_);
  or _70185_ (_18934_, _18933_, _10516_);
  or _70186_ (_18936_, _18934_, _18932_);
  or _70187_ (_18937_, _18936_, _18928_);
  and _70188_ (_18938_, _18937_, _18904_);
  or _70189_ (_18939_, _18938_, _07081_);
  or _70190_ (_18940_, _09207_, _07082_);
  and _70191_ (_18941_, _18940_, _06229_);
  and _70192_ (_18942_, _18941_, _18939_);
  nor _70193_ (_18943_, _08014_, _06229_);
  or _70194_ (_18944_, _18943_, _10525_);
  or _70195_ (_18945_, _18944_, _18942_);
  nand _70196_ (_18947_, _10525_, _09981_);
  and _70197_ (_18948_, _18947_, _18945_);
  or _70198_ (_18949_, _18948_, _06152_);
  and _70199_ (_18950_, _15297_, _08409_);
  or _70200_ (_18951_, _18950_, _18929_);
  or _70201_ (_18952_, _18951_, _06153_);
  and _70202_ (_18953_, _18952_, _06146_);
  and _70203_ (_18954_, _18953_, _18949_);
  or _70204_ (_18955_, _18929_, _15331_);
  and _70205_ (_18956_, _18931_, _06145_);
  and _70206_ (_18958_, _18956_, _18955_);
  or _70207_ (_18959_, _18958_, _09295_);
  or _70208_ (_18960_, _18959_, _18954_);
  nor _70209_ (_18961_, _09786_, _09784_);
  nor _70210_ (_18962_, _18961_, _09787_);
  or _70211_ (_18963_, _18962_, _09301_);
  and _70212_ (_18964_, _18963_, _10554_);
  and _70213_ (_18965_, _18964_, _18960_);
  or _70214_ (_18966_, _08101_, _09930_);
  and _70215_ (_18967_, _08101_, _09930_);
  or _70216_ (_18969_, _18621_, _18967_);
  and _70217_ (_18970_, _18969_, _18966_);
  nor _70218_ (_18971_, _18970_, _10969_);
  and _70219_ (_18972_, _18970_, _10969_);
  nor _70220_ (_18973_, _18972_, _18971_);
  nor _70221_ (_18974_, _18631_, _18625_);
  and _70222_ (_18975_, _18974_, \oc8051_golden_model_1.PSW [7]);
  or _70223_ (_18976_, _18975_, _18973_);
  nand _70224_ (_18977_, _18975_, _18973_);
  and _70225_ (_18978_, _18977_, _18976_);
  nand _70226_ (_18980_, _18978_, _10557_);
  nand _70227_ (_18981_, _18980_, _12380_);
  or _70228_ (_18982_, _18981_, _18965_);
  and _70229_ (_18983_, _18982_, _06265_);
  and _70230_ (_18984_, _18983_, _18903_);
  nor _70231_ (_18985_, _18655_, _18648_);
  or _70232_ (_18986_, _18644_, _13929_);
  and _70233_ (_18987_, _18986_, _13927_);
  nor _70234_ (_18988_, _18987_, _10295_);
  and _70235_ (_18989_, _18987_, _10295_);
  nor _70236_ (_18991_, _18989_, _18988_);
  nor _70237_ (_18992_, _18991_, _10693_);
  and _70238_ (_18993_, _18991_, _10693_);
  nor _70239_ (_18994_, _18993_, _18992_);
  nand _70240_ (_18995_, _18994_, _18985_);
  or _70241_ (_18996_, _18994_, _18985_);
  and _70242_ (_18997_, _18996_, _06260_);
  and _70243_ (_18998_, _18997_, _18995_);
  or _70244_ (_18999_, _18998_, _18984_);
  and _70245_ (_19000_, _18999_, _10388_);
  or _70246_ (_19002_, _18525_, _13957_);
  and _70247_ (_19003_, _19002_, _13956_);
  nor _70248_ (_19004_, _19003_, _11052_);
  and _70249_ (_19005_, _19003_, _11052_);
  nor _70250_ (_19006_, _19005_, _19004_);
  nor _70251_ (_19007_, _18535_, _18530_);
  and _70252_ (_19008_, _19007_, \oc8051_golden_model_1.PSW [7]);
  or _70253_ (_19009_, _19008_, _19006_);
  nand _70254_ (_19010_, _19008_, _19006_);
  and _70255_ (_19011_, _19010_, _10387_);
  and _70256_ (_19013_, _19011_, _19009_);
  or _70257_ (_19014_, _19013_, _05870_);
  or _70258_ (_19015_, _19014_, _19000_);
  nand _70259_ (_19016_, _06203_, _05870_);
  and _70260_ (_19017_, _19016_, _06140_);
  and _70261_ (_19018_, _19017_, _19015_);
  and _70262_ (_19019_, _15348_, _08409_);
  or _70263_ (_19020_, _19019_, _18929_);
  and _70264_ (_19021_, _19020_, _06139_);
  or _70265_ (_19022_, _19021_, _09842_);
  or _70266_ (_19024_, _19022_, _19018_);
  and _70267_ (_19025_, _19024_, _18888_);
  or _70268_ (_19026_, _19025_, _06116_);
  and _70269_ (_19027_, _09207_, _07809_);
  or _70270_ (_19028_, _18878_, _06117_);
  or _70271_ (_19029_, _19028_, _19027_);
  and _70272_ (_19030_, _19029_, _06114_);
  and _70273_ (_19031_, _19030_, _19026_);
  or _70274_ (_19032_, _19031_, _18885_);
  and _70275_ (_19033_, _19032_, _11922_);
  nor _70276_ (_19035_, _06203_, _05802_);
  not _70277_ (_19036_, _09888_);
  nor _70278_ (_19037_, _19036_, _09884_);
  and _70279_ (_19038_, _19037_, _05799_);
  and _70280_ (_19039_, _19038_, _09855_);
  or _70281_ (_19040_, _19039_, _19035_);
  or _70282_ (_19041_, _19040_, _19033_);
  and _70283_ (_19042_, _19041_, _06111_);
  and _70284_ (_19043_, _15402_, _07809_);
  or _70285_ (_19044_, _19043_, _18878_);
  and _70286_ (_19046_, _19044_, _06110_);
  or _70287_ (_19047_, _19046_, _10751_);
  or _70288_ (_19048_, _19047_, _19042_);
  nand _70289_ (_19049_, _10751_, _06203_);
  and _70290_ (_19050_, _19049_, _18182_);
  and _70291_ (_19051_, _19050_, _19048_);
  and _70292_ (_19052_, _10969_, _18181_);
  nor _70293_ (_19053_, _19052_, _19051_);
  or _70294_ (_19054_, _19053_, _18174_);
  nand _70295_ (_19055_, _10969_, _18174_);
  and _70296_ (_19057_, _19055_, _19054_);
  nor _70297_ (_19058_, _19057_, _18175_);
  and _70298_ (_19059_, _10969_, _18175_);
  or _70299_ (_19060_, _19059_, _06574_);
  or _70300_ (_19061_, _19060_, _19058_);
  nor _70301_ (_19062_, _10969_, _18701_);
  or _70302_ (_19063_, _19062_, _17709_);
  nor _70303_ (_19064_, _19063_, _17714_);
  and _70304_ (_19065_, _19064_, _19061_);
  or _70305_ (_19066_, _19065_, _18882_);
  and _70306_ (_19068_, _19066_, _18172_);
  and _70307_ (_19069_, _17105_, _10969_);
  or _70308_ (_19070_, _19069_, _06771_);
  or _70309_ (_19071_, _19070_, _19068_);
  or _70310_ (_19072_, _10969_, _17113_);
  and _70311_ (_19073_, _19072_, _10776_);
  and _70312_ (_19074_, _19073_, _19071_);
  and _70313_ (_19075_, _10775_, _11008_);
  or _70314_ (_19076_, _19075_, _06400_);
  or _70315_ (_19077_, _19076_, _19074_);
  or _70316_ (_19079_, _10295_, _06401_);
  and _70317_ (_19080_, _19079_, _10788_);
  and _70318_ (_19081_, _19080_, _19077_);
  and _70319_ (_19082_, _10787_, _11052_);
  or _70320_ (_19083_, _19082_, _06297_);
  or _70321_ (_19084_, _19083_, _19081_);
  and _70322_ (_19085_, _19084_, _18881_);
  or _70323_ (_19086_, _19085_, _06402_);
  or _70324_ (_19087_, _18878_, _07125_);
  and _70325_ (_19088_, _19087_, _10808_);
  and _70326_ (_19090_, _19088_, _19086_);
  and _70327_ (_19091_, _10812_, _10966_);
  or _70328_ (_19092_, _19091_, _10811_);
  or _70329_ (_19093_, _19092_, _19090_);
  or _70330_ (_19094_, _10816_, _11005_);
  and _70331_ (_19095_, _19094_, _06410_);
  and _70332_ (_19096_, _19095_, _19093_);
  and _70333_ (_19097_, _10266_, _06409_);
  or _70334_ (_19098_, _19097_, _10820_);
  or _70335_ (_19099_, _19098_, _19096_);
  or _70336_ (_19101_, _10826_, _11049_);
  and _70337_ (_19102_, _19101_, _07132_);
  and _70338_ (_19103_, _19102_, _19099_);
  nand _70339_ (_19104_, _19044_, _06306_);
  nor _70340_ (_19105_, _19104_, _10294_);
  or _70341_ (_19106_, _19105_, _06524_);
  or _70342_ (_19107_, _19106_, _19103_);
  and _70343_ (_19108_, _19107_, _18876_);
  or _70344_ (_19109_, _19108_, _06555_);
  nor _70345_ (_19110_, _10967_, _10834_);
  nor _70346_ (_19112_, _19110_, _06975_);
  and _70347_ (_19113_, _19112_, _19109_);
  and _70348_ (_19114_, _10967_, _06975_);
  or _70349_ (_19115_, _19114_, _19113_);
  and _70350_ (_19116_, _19115_, _17847_);
  and _70351_ (_19117_, _10835_, _10967_);
  or _70352_ (_19118_, _19117_, _10841_);
  or _70353_ (_19119_, _19118_, _19116_);
  or _70354_ (_19120_, _17242_, _11006_);
  and _70355_ (_19121_, _19120_, _06395_);
  and _70356_ (_19123_, _19121_, _19119_);
  nand _70357_ (_19124_, _10851_, _10294_);
  and _70358_ (_19125_, _19124_, _10850_);
  or _70359_ (_19126_, _19125_, _19123_);
  and _70360_ (_19127_, _19126_, _18875_);
  or _70361_ (_19128_, _19127_, _06303_);
  and _70362_ (_19129_, _15410_, _07809_);
  or _70363_ (_19130_, _18878_, _08819_);
  or _70364_ (_19131_, _19130_, _19129_);
  and _70365_ (_19132_, _19131_, _10380_);
  and _70366_ (_19134_, _19132_, _19128_);
  or _70367_ (_19135_, _10365_, _10316_);
  and _70368_ (_19136_, _10858_, _10366_);
  and _70369_ (_19137_, _19136_, _19135_);
  or _70370_ (_19138_, _19137_, _19134_);
  or _70371_ (_19139_, _19138_, _17240_);
  or _70372_ (_19140_, _10886_, _10641_);
  and _70373_ (_19141_, _19140_, _10887_);
  and _70374_ (_19142_, _19141_, _06276_);
  or _70375_ (_19143_, _19142_, _10867_);
  and _70376_ (_19145_, _19143_, _19139_);
  and _70377_ (_19146_, _19141_, _06792_);
  or _70378_ (_19147_, _19146_, _06406_);
  or _70379_ (_19148_, _19147_, _19145_);
  and _70380_ (_19149_, _19148_, _18874_);
  or _70381_ (_19150_, _10946_, _10714_);
  nor _70382_ (_19151_, _10947_, _10927_);
  and _70383_ (_19152_, _19151_, _19150_);
  or _70384_ (_19153_, _19152_, _10925_);
  or _70385_ (_19154_, _19153_, _19149_);
  nand _70386_ (_19156_, _10925_, _09930_);
  and _70387_ (_19157_, _19156_, _10963_);
  and _70388_ (_19158_, _19157_, _19154_);
  nor _70389_ (_19159_, _10995_, _10969_);
  nor _70390_ (_19160_, _19159_, _10996_);
  and _70391_ (_19161_, _19160_, _18454_);
  or _70392_ (_19162_, _19161_, _17195_);
  or _70393_ (_19163_, _19162_, _19158_);
  and _70394_ (_19164_, _19163_, _18870_);
  or _70395_ (_19165_, _19164_, _17199_);
  or _70396_ (_19167_, _18867_, _17200_);
  and _70397_ (_19168_, _19167_, _06171_);
  and _70398_ (_19169_, _19168_, _19165_);
  or _70399_ (_19170_, _10295_, _10293_);
  and _70400_ (_19171_, _19170_, _10296_);
  or _70401_ (_19172_, _19171_, _10264_);
  and _70402_ (_19173_, _19172_, _12691_);
  or _70403_ (_19174_, _19173_, _19169_);
  or _70404_ (_19175_, _11078_, _11052_);
  and _70405_ (_19176_, _19175_, _11079_);
  or _70406_ (_19178_, _19176_, _10265_);
  and _70407_ (_19179_, _19178_, _12693_);
  and _70408_ (_19180_, _19179_, _19174_);
  and _70409_ (_19181_, _10262_, \oc8051_golden_model_1.ACC [5]);
  or _70410_ (_19182_, _19181_, _06433_);
  or _70411_ (_19183_, _19182_, _19180_);
  or _70412_ (_19184_, _18917_, _06829_);
  and _70413_ (_19185_, _19184_, _11090_);
  and _70414_ (_19186_, _19185_, _19183_);
  nor _70415_ (_19187_, _11098_, _09883_);
  or _70416_ (_19189_, _19187_, _11099_);
  and _70417_ (_19190_, _19189_, _11089_);
  or _70418_ (_19191_, _19190_, _11094_);
  or _70419_ (_19192_, _19191_, _19186_);
  nand _70420_ (_19193_, _11094_, _08430_);
  and _70421_ (_19194_, _19193_, _05749_);
  and _70422_ (_19195_, _19194_, _19192_);
  and _70423_ (_19196_, _18951_, _05748_);
  or _70424_ (_19197_, _19196_, _06440_);
  or _70425_ (_19198_, _19197_, _19195_);
  and _70426_ (_19200_, _15478_, _07809_);
  or _70427_ (_19201_, _18878_, _06444_);
  or _70428_ (_19202_, _19201_, _19200_);
  and _70429_ (_19203_, _19202_, _11113_);
  and _70430_ (_19204_, _19203_, _19198_);
  nor _70431_ (_19205_, _11124_, \oc8051_golden_model_1.ACC [6]);
  nor _70432_ (_19206_, _19205_, _11125_);
  and _70433_ (_19207_, _19206_, _11112_);
  or _70434_ (_19208_, _19207_, _11119_);
  or _70435_ (_19209_, _19208_, _19204_);
  nand _70436_ (_19211_, _11119_, _08430_);
  and _70437_ (_19212_, _19211_, _01317_);
  and _70438_ (_19213_, _19212_, _19209_);
  or _70439_ (_19214_, _19213_, _18865_);
  and _70440_ (_43609_, _19214_, _43100_);
  not _70441_ (_19215_, \oc8051_golden_model_1.PCON [0]);
  nor _70442_ (_19216_, _01317_, _19215_);
  and _70443_ (_19217_, _07856_, \oc8051_golden_model_1.ACC [0]);
  and _70444_ (_19218_, _19217_, _08211_);
  nor _70445_ (_19219_, _07856_, _19215_);
  or _70446_ (_19221_, _19219_, _07130_);
  or _70447_ (_19222_, _19221_, _19218_);
  nor _70448_ (_19223_, _08211_, _11137_);
  or _70449_ (_19224_, _19223_, _19219_);
  or _70450_ (_19225_, _19224_, _06161_);
  or _70451_ (_19226_, _19219_, _19217_);
  and _70452_ (_19227_, _19226_, _07056_);
  nor _70453_ (_19228_, _07056_, _19215_);
  or _70454_ (_19229_, _19228_, _06160_);
  or _70455_ (_19230_, _19229_, _19227_);
  and _70456_ (_19232_, _19230_, _07075_);
  and _70457_ (_19233_, _19232_, _19225_);
  and _70458_ (_19234_, _07856_, _07049_);
  or _70459_ (_19235_, _19234_, _19219_);
  and _70460_ (_19236_, _19235_, _06217_);
  or _70461_ (_19237_, _19236_, _19233_);
  and _70462_ (_19238_, _19237_, _06229_);
  and _70463_ (_19239_, _19226_, _06220_);
  or _70464_ (_19240_, _19239_, _09842_);
  or _70465_ (_19241_, _19240_, _19238_);
  or _70466_ (_19243_, _19235_, _06132_);
  and _70467_ (_19244_, _19243_, _19241_);
  or _70468_ (_19245_, _19244_, _06116_);
  and _70469_ (_19246_, _09160_, _07856_);
  or _70470_ (_19247_, _19219_, _06117_);
  or _70471_ (_19248_, _19247_, _19246_);
  and _70472_ (_19249_, _19248_, _19245_);
  or _70473_ (_19250_, _19249_, _05787_);
  and _70474_ (_19251_, _14260_, _07856_);
  or _70475_ (_19252_, _19219_, _06114_);
  or _70476_ (_19254_, _19252_, _19251_);
  and _70477_ (_19255_, _19254_, _06111_);
  and _70478_ (_19256_, _19255_, _19250_);
  and _70479_ (_19257_, _07856_, _08708_);
  or _70480_ (_19258_, _19257_, _19219_);
  and _70481_ (_19259_, _19258_, _06110_);
  or _70482_ (_19260_, _19259_, _06297_);
  or _70483_ (_19261_, _19260_, _19256_);
  and _70484_ (_19262_, _14275_, _07856_);
  or _70485_ (_19263_, _19262_, _19219_);
  or _70486_ (_19265_, _19263_, _07127_);
  and _70487_ (_19266_, _19265_, _07125_);
  and _70488_ (_19267_, _19266_, _19261_);
  nor _70489_ (_19268_, _12321_, _11137_);
  or _70490_ (_19269_, _19268_, _19219_);
  nor _70491_ (_19270_, _19218_, _07125_);
  and _70492_ (_19271_, _19270_, _19269_);
  or _70493_ (_19272_, _19271_, _19267_);
  and _70494_ (_19273_, _19272_, _07132_);
  nand _70495_ (_19274_, _19258_, _06306_);
  nor _70496_ (_19276_, _19274_, _19223_);
  or _70497_ (_19277_, _19276_, _06411_);
  or _70498_ (_19278_, _19277_, _19273_);
  and _70499_ (_19279_, _19278_, _19222_);
  or _70500_ (_19280_, _19279_, _06303_);
  and _70501_ (_19281_, _14167_, _07856_);
  or _70502_ (_19282_, _19219_, _08819_);
  or _70503_ (_19283_, _19282_, _19281_);
  and _70504_ (_19284_, _19283_, _08824_);
  and _70505_ (_19285_, _19284_, _19280_);
  not _70506_ (_19287_, _06630_);
  and _70507_ (_19288_, _19269_, _06396_);
  or _70508_ (_19289_, _19288_, _19287_);
  or _70509_ (_19290_, _19289_, _19285_);
  or _70510_ (_19291_, _19224_, _06630_);
  and _70511_ (_19292_, _19291_, _01317_);
  and _70512_ (_19293_, _19292_, _19290_);
  or _70513_ (_19294_, _19293_, _19216_);
  and _70514_ (_43611_, _19294_, _43100_);
  not _70515_ (_19295_, \oc8051_golden_model_1.PCON [1]);
  nor _70516_ (_19297_, _01317_, _19295_);
  or _70517_ (_19298_, _14442_, _11137_);
  or _70518_ (_19299_, _07856_, \oc8051_golden_model_1.PCON [1]);
  and _70519_ (_19300_, _19299_, _05787_);
  and _70520_ (_19301_, _19300_, _19298_);
  and _70521_ (_19302_, _09115_, _07856_);
  nor _70522_ (_19303_, _07856_, _19295_);
  or _70523_ (_19304_, _19303_, _06117_);
  or _70524_ (_19305_, _19304_, _19302_);
  and _70525_ (_19306_, _07856_, _07306_);
  or _70526_ (_19308_, _19306_, _19303_);
  or _70527_ (_19309_, _19308_, _06132_);
  and _70528_ (_19310_, _14363_, _07856_);
  not _70529_ (_19311_, _19310_);
  and _70530_ (_19312_, _19311_, _19299_);
  or _70531_ (_19313_, _19312_, _06161_);
  and _70532_ (_19314_, _07856_, \oc8051_golden_model_1.ACC [1]);
  or _70533_ (_19315_, _19314_, _19303_);
  and _70534_ (_19316_, _19315_, _07056_);
  nor _70535_ (_19317_, _07056_, _19295_);
  or _70536_ (_19319_, _19317_, _06160_);
  or _70537_ (_19320_, _19319_, _19316_);
  and _70538_ (_19321_, _19320_, _07075_);
  and _70539_ (_19322_, _19321_, _19313_);
  and _70540_ (_19323_, _19308_, _06217_);
  or _70541_ (_19324_, _19323_, _19322_);
  and _70542_ (_19325_, _19324_, _06229_);
  and _70543_ (_19326_, _19315_, _06220_);
  or _70544_ (_19327_, _19326_, _09842_);
  or _70545_ (_19328_, _19327_, _19325_);
  and _70546_ (_19330_, _19328_, _19309_);
  or _70547_ (_19331_, _19330_, _06116_);
  and _70548_ (_19332_, _19331_, _06114_);
  and _70549_ (_19333_, _19332_, _19305_);
  or _70550_ (_19334_, _19333_, _19301_);
  and _70551_ (_19335_, _19334_, _06298_);
  or _70552_ (_19336_, _14346_, _11137_);
  and _70553_ (_19337_, _19299_, _06297_);
  and _70554_ (_19338_, _19337_, _19336_);
  nand _70555_ (_19339_, _07856_, _06945_);
  and _70556_ (_19341_, _19299_, _06110_);
  and _70557_ (_19342_, _19341_, _19339_);
  or _70558_ (_19343_, _19342_, _06402_);
  or _70559_ (_19344_, _19343_, _19338_);
  or _70560_ (_19345_, _19344_, _19335_);
  and _70561_ (_19346_, _10278_, _07856_);
  or _70562_ (_19347_, _19346_, _19303_);
  or _70563_ (_19348_, _19347_, _07125_);
  and _70564_ (_19349_, _19348_, _07132_);
  and _70565_ (_19350_, _19349_, _19345_);
  or _70566_ (_19352_, _14344_, _11137_);
  and _70567_ (_19353_, _19299_, _06306_);
  and _70568_ (_19354_, _19353_, _19352_);
  or _70569_ (_19355_, _19354_, _06411_);
  or _70570_ (_19356_, _19355_, _19350_);
  and _70571_ (_19357_, _19314_, _08176_);
  or _70572_ (_19358_, _19303_, _07130_);
  or _70573_ (_19359_, _19358_, _19357_);
  and _70574_ (_19360_, _19359_, _08819_);
  and _70575_ (_19361_, _19360_, _19356_);
  or _70576_ (_19363_, _19339_, _08176_);
  and _70577_ (_19364_, _19299_, _06303_);
  and _70578_ (_19365_, _19364_, _19363_);
  or _70579_ (_19366_, _19365_, _06396_);
  or _70580_ (_19367_, _19366_, _19361_);
  nor _70581_ (_19368_, _10277_, _11137_);
  or _70582_ (_19369_, _19368_, _19303_);
  or _70583_ (_19370_, _19369_, _08824_);
  and _70584_ (_19371_, _19370_, _19367_);
  and _70585_ (_19372_, _19371_, _06829_);
  and _70586_ (_19374_, _19312_, _06433_);
  or _70587_ (_19375_, _19374_, _06440_);
  or _70588_ (_19376_, _19375_, _19372_);
  or _70589_ (_19377_, _19303_, _06444_);
  or _70590_ (_19378_, _19377_, _19310_);
  and _70591_ (_19379_, _19378_, _01317_);
  and _70592_ (_19380_, _19379_, _19376_);
  or _70593_ (_19381_, _19380_, _19297_);
  and _70594_ (_43612_, _19381_, _43100_);
  not _70595_ (_19382_, \oc8051_golden_model_1.PCON [2]);
  nor _70596_ (_19384_, _01317_, _19382_);
  nor _70597_ (_19385_, _07856_, _19382_);
  and _70598_ (_19386_, _07856_, _07708_);
  or _70599_ (_19387_, _19386_, _19385_);
  or _70600_ (_19388_, _19387_, _06132_);
  and _70601_ (_19389_, _14542_, _07856_);
  or _70602_ (_19390_, _19389_, _19385_);
  and _70603_ (_19391_, _19390_, _06160_);
  nor _70604_ (_19392_, _07056_, _19382_);
  and _70605_ (_19393_, _07856_, \oc8051_golden_model_1.ACC [2]);
  or _70606_ (_19395_, _19393_, _19385_);
  and _70607_ (_19396_, _19395_, _07056_);
  or _70608_ (_19397_, _19396_, _19392_);
  and _70609_ (_19398_, _19397_, _06161_);
  or _70610_ (_19399_, _19398_, _06217_);
  or _70611_ (_19400_, _19399_, _19391_);
  or _70612_ (_19401_, _19387_, _07075_);
  and _70613_ (_19402_, _19401_, _06229_);
  and _70614_ (_19403_, _19402_, _19400_);
  and _70615_ (_19404_, _19395_, _06220_);
  or _70616_ (_19406_, _19404_, _09842_);
  or _70617_ (_19407_, _19406_, _19403_);
  and _70618_ (_19408_, _19407_, _19388_);
  or _70619_ (_19409_, _19408_, _06116_);
  and _70620_ (_19410_, _09211_, _07856_);
  or _70621_ (_19411_, _19385_, _06117_);
  or _70622_ (_19412_, _19411_, _19410_);
  and _70623_ (_19413_, _19412_, _19409_);
  or _70624_ (_19414_, _19413_, _05787_);
  and _70625_ (_19415_, _14630_, _07856_);
  or _70626_ (_19417_, _19415_, _19385_);
  or _70627_ (_19418_, _19417_, _06114_);
  and _70628_ (_19419_, _19418_, _06111_);
  and _70629_ (_19420_, _19419_, _19414_);
  and _70630_ (_19421_, _07856_, _08768_);
  or _70631_ (_19422_, _19421_, _19385_);
  and _70632_ (_19423_, _19422_, _06110_);
  or _70633_ (_19424_, _19423_, _06297_);
  or _70634_ (_19425_, _19424_, _19420_);
  and _70635_ (_19426_, _14646_, _07856_);
  or _70636_ (_19428_, _19385_, _07127_);
  or _70637_ (_19429_, _19428_, _19426_);
  and _70638_ (_19430_, _19429_, _07125_);
  and _70639_ (_19431_, _19430_, _19425_);
  and _70640_ (_19432_, _10282_, _07856_);
  or _70641_ (_19433_, _19432_, _19385_);
  and _70642_ (_19434_, _19433_, _06402_);
  or _70643_ (_19435_, _19434_, _19431_);
  and _70644_ (_19436_, _19435_, _07132_);
  or _70645_ (_19437_, _19385_, _08248_);
  and _70646_ (_19439_, _19422_, _06306_);
  and _70647_ (_19440_, _19439_, _19437_);
  or _70648_ (_19441_, _19440_, _19436_);
  and _70649_ (_19442_, _19441_, _07130_);
  and _70650_ (_19443_, _19395_, _06411_);
  and _70651_ (_19444_, _19443_, _19437_);
  or _70652_ (_19445_, _19444_, _06303_);
  or _70653_ (_19446_, _19445_, _19442_);
  and _70654_ (_19447_, _14643_, _07856_);
  or _70655_ (_19448_, _19385_, _08819_);
  or _70656_ (_19450_, _19448_, _19447_);
  and _70657_ (_19451_, _19450_, _08824_);
  and _70658_ (_19452_, _19451_, _19446_);
  nor _70659_ (_19453_, _10281_, _11137_);
  or _70660_ (_19454_, _19453_, _19385_);
  and _70661_ (_19455_, _19454_, _06396_);
  or _70662_ (_19456_, _19455_, _19452_);
  and _70663_ (_19457_, _19456_, _06829_);
  and _70664_ (_19458_, _19390_, _06433_);
  or _70665_ (_19459_, _19458_, _06440_);
  or _70666_ (_19461_, _19459_, _19457_);
  and _70667_ (_19462_, _14710_, _07856_);
  or _70668_ (_19463_, _19385_, _06444_);
  or _70669_ (_19464_, _19463_, _19462_);
  and _70670_ (_19465_, _19464_, _01317_);
  and _70671_ (_19466_, _19465_, _19461_);
  or _70672_ (_19467_, _19466_, _19384_);
  and _70673_ (_43613_, _19467_, _43100_);
  and _70674_ (_19468_, _11137_, \oc8051_golden_model_1.PCON [3]);
  and _70675_ (_19469_, _14738_, _07856_);
  or _70676_ (_19471_, _19469_, _19468_);
  or _70677_ (_19472_, _19471_, _06161_);
  and _70678_ (_19473_, _07856_, \oc8051_golden_model_1.ACC [3]);
  or _70679_ (_19474_, _19473_, _19468_);
  and _70680_ (_19475_, _19474_, _07056_);
  and _70681_ (_19476_, _07057_, \oc8051_golden_model_1.PCON [3]);
  or _70682_ (_19477_, _19476_, _06160_);
  or _70683_ (_19478_, _19477_, _19475_);
  and _70684_ (_19479_, _19478_, _07075_);
  and _70685_ (_19480_, _19479_, _19472_);
  and _70686_ (_19482_, _07856_, _07544_);
  or _70687_ (_19483_, _19482_, _19468_);
  and _70688_ (_19484_, _19483_, _06217_);
  or _70689_ (_19485_, _19484_, _19480_);
  and _70690_ (_19486_, _19485_, _06229_);
  and _70691_ (_19487_, _19474_, _06220_);
  or _70692_ (_19488_, _19487_, _09842_);
  or _70693_ (_19489_, _19488_, _19486_);
  or _70694_ (_19490_, _19483_, _06132_);
  and _70695_ (_19491_, _19490_, _06117_);
  and _70696_ (_19493_, _19491_, _19489_);
  and _70697_ (_19494_, _09210_, _07856_);
  or _70698_ (_19495_, _19494_, _19468_);
  and _70699_ (_19496_, _19495_, _06116_);
  or _70700_ (_19497_, _19496_, _05787_);
  or _70701_ (_19498_, _19497_, _19493_);
  and _70702_ (_19499_, _14825_, _07856_);
  or _70703_ (_19500_, _19499_, _19468_);
  or _70704_ (_19501_, _19500_, _06114_);
  and _70705_ (_19502_, _19501_, _06111_);
  and _70706_ (_19504_, _19502_, _19498_);
  and _70707_ (_19505_, _07856_, _08712_);
  or _70708_ (_19506_, _19505_, _19468_);
  and _70709_ (_19507_, _19506_, _06110_);
  or _70710_ (_19508_, _19507_, _06297_);
  or _70711_ (_19509_, _19508_, _19504_);
  and _70712_ (_19510_, _14727_, _07856_);
  or _70713_ (_19511_, _19510_, _19468_);
  or _70714_ (_19512_, _19511_, _07127_);
  and _70715_ (_19513_, _19512_, _07125_);
  and _70716_ (_19515_, _19513_, _19509_);
  and _70717_ (_19516_, _12318_, _07856_);
  or _70718_ (_19517_, _19516_, _19468_);
  and _70719_ (_19518_, _19517_, _06402_);
  or _70720_ (_19519_, _19518_, _19515_);
  and _70721_ (_19520_, _19519_, _07132_);
  or _70722_ (_19521_, _19468_, _08140_);
  and _70723_ (_19522_, _19506_, _06306_);
  and _70724_ (_19523_, _19522_, _19521_);
  or _70725_ (_19524_, _19523_, _19520_);
  and _70726_ (_19526_, _19524_, _07130_);
  and _70727_ (_19527_, _19474_, _06411_);
  and _70728_ (_19528_, _19527_, _19521_);
  or _70729_ (_19529_, _19528_, _06303_);
  or _70730_ (_19530_, _19529_, _19526_);
  and _70731_ (_19531_, _14724_, _07856_);
  or _70732_ (_19532_, _19468_, _08819_);
  or _70733_ (_19533_, _19532_, _19531_);
  and _70734_ (_19534_, _19533_, _08824_);
  and _70735_ (_19535_, _19534_, _19530_);
  nor _70736_ (_19537_, _10273_, _11137_);
  or _70737_ (_19538_, _19537_, _19468_);
  and _70738_ (_19539_, _19538_, _06396_);
  or _70739_ (_19540_, _19539_, _06433_);
  or _70740_ (_19541_, _19540_, _19535_);
  or _70741_ (_19542_, _19471_, _06829_);
  and _70742_ (_19543_, _19542_, _06444_);
  and _70743_ (_19544_, _19543_, _19541_);
  and _70744_ (_19545_, _14897_, _07856_);
  or _70745_ (_19546_, _19545_, _19468_);
  and _70746_ (_19548_, _19546_, _06440_);
  or _70747_ (_19549_, _19548_, _01321_);
  or _70748_ (_19550_, _19549_, _19544_);
  or _70749_ (_19551_, _01317_, \oc8051_golden_model_1.PCON [3]);
  and _70750_ (_19552_, _19551_, _43100_);
  and _70751_ (_43614_, _19552_, _19550_);
  and _70752_ (_19553_, _11137_, \oc8051_golden_model_1.PCON [4]);
  and _70753_ (_19554_, _08336_, _07856_);
  or _70754_ (_19555_, _19554_, _19553_);
  or _70755_ (_19556_, _19555_, _06132_);
  and _70756_ (_19558_, _14928_, _07856_);
  or _70757_ (_19559_, _19558_, _19553_);
  or _70758_ (_19560_, _19559_, _06161_);
  and _70759_ (_19561_, _07856_, \oc8051_golden_model_1.ACC [4]);
  or _70760_ (_19562_, _19561_, _19553_);
  and _70761_ (_19563_, _19562_, _07056_);
  and _70762_ (_19564_, _07057_, \oc8051_golden_model_1.PCON [4]);
  or _70763_ (_19565_, _19564_, _06160_);
  or _70764_ (_19566_, _19565_, _19563_);
  and _70765_ (_19567_, _19566_, _07075_);
  and _70766_ (_19569_, _19567_, _19560_);
  and _70767_ (_19570_, _19555_, _06217_);
  or _70768_ (_19571_, _19570_, _19569_);
  and _70769_ (_19572_, _19571_, _06229_);
  and _70770_ (_19573_, _19562_, _06220_);
  or _70771_ (_19574_, _19573_, _09842_);
  or _70772_ (_19575_, _19574_, _19572_);
  and _70773_ (_19576_, _19575_, _19556_);
  or _70774_ (_19577_, _19576_, _06116_);
  and _70775_ (_19578_, _09209_, _07856_);
  or _70776_ (_19580_, _19553_, _06117_);
  or _70777_ (_19581_, _19580_, _19578_);
  and _70778_ (_19582_, _19581_, _06114_);
  and _70779_ (_19583_, _19582_, _19577_);
  and _70780_ (_19584_, _15013_, _07856_);
  or _70781_ (_19585_, _19584_, _19553_);
  and _70782_ (_19586_, _19585_, _05787_);
  or _70783_ (_19587_, _19586_, _19583_);
  or _70784_ (_19588_, _19587_, _11136_);
  and _70785_ (_19589_, _15029_, _07856_);
  or _70786_ (_19591_, _19553_, _07127_);
  or _70787_ (_19592_, _19591_, _19589_);
  and _70788_ (_19593_, _08715_, _07856_);
  or _70789_ (_19594_, _19593_, _19553_);
  or _70790_ (_19595_, _19594_, _06111_);
  and _70791_ (_19596_, _19595_, _07125_);
  and _70792_ (_19597_, _19596_, _19592_);
  and _70793_ (_19598_, _19597_, _19588_);
  and _70794_ (_19599_, _10289_, _07856_);
  or _70795_ (_19600_, _19599_, _19553_);
  and _70796_ (_19602_, _19600_, _06402_);
  or _70797_ (_19603_, _19602_, _19598_);
  and _70798_ (_19604_, _19603_, _07132_);
  or _70799_ (_19605_, _19553_, _08339_);
  and _70800_ (_19606_, _19594_, _06306_);
  and _70801_ (_19607_, _19606_, _19605_);
  or _70802_ (_19608_, _19607_, _19604_);
  and _70803_ (_19609_, _19608_, _07130_);
  and _70804_ (_19610_, _19562_, _06411_);
  and _70805_ (_19611_, _19610_, _19605_);
  or _70806_ (_19613_, _19611_, _06303_);
  or _70807_ (_19614_, _19613_, _19609_);
  and _70808_ (_19615_, _15026_, _07856_);
  or _70809_ (_19616_, _19553_, _08819_);
  or _70810_ (_19617_, _19616_, _19615_);
  and _70811_ (_19618_, _19617_, _08824_);
  and _70812_ (_19619_, _19618_, _19614_);
  nor _70813_ (_19620_, _10288_, _11137_);
  or _70814_ (_19621_, _19620_, _19553_);
  and _70815_ (_19622_, _19621_, _06396_);
  or _70816_ (_19624_, _19622_, _06433_);
  or _70817_ (_19625_, _19624_, _19619_);
  or _70818_ (_19626_, _19559_, _06829_);
  and _70819_ (_19627_, _19626_, _06444_);
  and _70820_ (_19628_, _19627_, _19625_);
  and _70821_ (_19629_, _15087_, _07856_);
  or _70822_ (_19630_, _19629_, _19553_);
  and _70823_ (_19631_, _19630_, _06440_);
  or _70824_ (_19632_, _19631_, _01321_);
  or _70825_ (_19633_, _19632_, _19628_);
  or _70826_ (_19635_, _01317_, \oc8051_golden_model_1.PCON [4]);
  and _70827_ (_19636_, _19635_, _43100_);
  and _70828_ (_43615_, _19636_, _19633_);
  and _70829_ (_19637_, _11137_, \oc8051_golden_model_1.PCON [5]);
  or _70830_ (_19638_, _19637_, _08104_);
  and _70831_ (_19639_, _08736_, _07856_);
  or _70832_ (_19640_, _19639_, _19637_);
  and _70833_ (_19641_, _19640_, _06306_);
  and _70834_ (_19642_, _19641_, _19638_);
  and _70835_ (_19643_, _15119_, _07856_);
  or _70836_ (_19645_, _19643_, _19637_);
  or _70837_ (_19646_, _19645_, _06161_);
  and _70838_ (_19647_, _07856_, \oc8051_golden_model_1.ACC [5]);
  or _70839_ (_19648_, _19647_, _19637_);
  and _70840_ (_19649_, _19648_, _07056_);
  and _70841_ (_19650_, _07057_, \oc8051_golden_model_1.PCON [5]);
  or _70842_ (_19651_, _19650_, _06160_);
  or _70843_ (_19652_, _19651_, _19649_);
  and _70844_ (_19653_, _19652_, _07075_);
  and _70845_ (_19654_, _19653_, _19646_);
  and _70846_ (_19656_, _08101_, _07856_);
  or _70847_ (_19657_, _19656_, _19637_);
  and _70848_ (_19658_, _19657_, _06217_);
  or _70849_ (_19659_, _19658_, _19654_);
  and _70850_ (_19660_, _19659_, _06229_);
  and _70851_ (_19661_, _19648_, _06220_);
  or _70852_ (_19662_, _19661_, _09842_);
  or _70853_ (_19663_, _19662_, _19660_);
  or _70854_ (_19664_, _19657_, _06132_);
  and _70855_ (_19665_, _19664_, _19663_);
  or _70856_ (_19667_, _19665_, _06116_);
  and _70857_ (_19668_, _09208_, _07856_);
  or _70858_ (_19669_, _19637_, _06117_);
  or _70859_ (_19670_, _19669_, _19668_);
  and _70860_ (_19671_, _19670_, _06114_);
  and _70861_ (_19672_, _19671_, _19667_);
  and _70862_ (_19673_, _15203_, _07856_);
  or _70863_ (_19674_, _19673_, _19637_);
  and _70864_ (_19675_, _19674_, _05787_);
  or _70865_ (_19676_, _19675_, _11136_);
  or _70866_ (_19678_, _19676_, _19672_);
  and _70867_ (_19679_, _15219_, _07856_);
  or _70868_ (_19680_, _19637_, _07127_);
  or _70869_ (_19681_, _19680_, _19679_);
  or _70870_ (_19682_, _19640_, _06111_);
  and _70871_ (_19683_, _19682_, _07125_);
  and _70872_ (_19684_, _19683_, _19681_);
  and _70873_ (_19685_, _19684_, _19678_);
  and _70874_ (_19686_, _12325_, _07856_);
  or _70875_ (_19687_, _19686_, _19637_);
  and _70876_ (_19689_, _19687_, _06402_);
  or _70877_ (_19690_, _19689_, _19685_);
  and _70878_ (_19691_, _19690_, _07132_);
  or _70879_ (_19692_, _19691_, _19642_);
  and _70880_ (_19693_, _19692_, _07130_);
  and _70881_ (_19694_, _19648_, _06411_);
  and _70882_ (_19695_, _19694_, _19638_);
  or _70883_ (_19696_, _19695_, _06303_);
  or _70884_ (_19697_, _19696_, _19693_);
  and _70885_ (_19698_, _15216_, _07856_);
  or _70886_ (_19700_, _19637_, _08819_);
  or _70887_ (_19701_, _19700_, _19698_);
  and _70888_ (_19702_, _19701_, _08824_);
  and _70889_ (_19703_, _19702_, _19697_);
  nor _70890_ (_19704_, _10269_, _11137_);
  or _70891_ (_19705_, _19704_, _19637_);
  and _70892_ (_19706_, _19705_, _06396_);
  or _70893_ (_19707_, _19706_, _06433_);
  or _70894_ (_19708_, _19707_, _19703_);
  or _70895_ (_19709_, _19645_, _06829_);
  and _70896_ (_19711_, _19709_, _06444_);
  and _70897_ (_19712_, _19711_, _19708_);
  and _70898_ (_19713_, _15275_, _07856_);
  or _70899_ (_19714_, _19713_, _19637_);
  and _70900_ (_19715_, _19714_, _06440_);
  or _70901_ (_19716_, _19715_, _01321_);
  or _70902_ (_19717_, _19716_, _19712_);
  or _70903_ (_19718_, _01317_, \oc8051_golden_model_1.PCON [5]);
  and _70904_ (_19719_, _19718_, _43100_);
  and _70905_ (_43617_, _19719_, _19717_);
  and _70906_ (_19721_, _11137_, \oc8051_golden_model_1.PCON [6]);
  or _70907_ (_19722_, _19721_, _08015_);
  and _70908_ (_19723_, _15402_, _07856_);
  or _70909_ (_19724_, _19723_, _19721_);
  and _70910_ (_19725_, _19724_, _06306_);
  and _70911_ (_19726_, _19725_, _19722_);
  and _70912_ (_19727_, _15300_, _07856_);
  or _70913_ (_19728_, _19727_, _19721_);
  or _70914_ (_19729_, _19728_, _06161_);
  and _70915_ (_19730_, _07856_, \oc8051_golden_model_1.ACC [6]);
  or _70916_ (_19732_, _19730_, _19721_);
  and _70917_ (_19733_, _19732_, _07056_);
  and _70918_ (_19734_, _07057_, \oc8051_golden_model_1.PCON [6]);
  or _70919_ (_19735_, _19734_, _06160_);
  or _70920_ (_19736_, _19735_, _19733_);
  and _70921_ (_19737_, _19736_, _07075_);
  and _70922_ (_19738_, _19737_, _19729_);
  and _70923_ (_19739_, _08012_, _07856_);
  or _70924_ (_19740_, _19739_, _19721_);
  and _70925_ (_19741_, _19740_, _06217_);
  or _70926_ (_19743_, _19741_, _19738_);
  and _70927_ (_19744_, _19743_, _06229_);
  and _70928_ (_19745_, _19732_, _06220_);
  or _70929_ (_19746_, _19745_, _09842_);
  or _70930_ (_19747_, _19746_, _19744_);
  or _70931_ (_19748_, _19740_, _06132_);
  and _70932_ (_19749_, _19748_, _19747_);
  or _70933_ (_19750_, _19749_, _06116_);
  and _70934_ (_19751_, _09207_, _07856_);
  or _70935_ (_19752_, _19721_, _06117_);
  or _70936_ (_19754_, _19752_, _19751_);
  and _70937_ (_19755_, _19754_, _06114_);
  and _70938_ (_19756_, _19755_, _19750_);
  and _70939_ (_19757_, _15395_, _07856_);
  or _70940_ (_19758_, _19757_, _19721_);
  and _70941_ (_19759_, _19758_, _05787_);
  or _70942_ (_19760_, _19759_, _11136_);
  or _70943_ (_19761_, _19760_, _19756_);
  and _70944_ (_19762_, _15413_, _07856_);
  or _70945_ (_19763_, _19721_, _07127_);
  or _70946_ (_19765_, _19763_, _19762_);
  or _70947_ (_19766_, _19724_, _06111_);
  and _70948_ (_19767_, _19766_, _07125_);
  and _70949_ (_19768_, _19767_, _19765_);
  and _70950_ (_19769_, _19768_, _19761_);
  and _70951_ (_19770_, _10295_, _07856_);
  or _70952_ (_19771_, _19770_, _19721_);
  and _70953_ (_19772_, _19771_, _06402_);
  or _70954_ (_19773_, _19772_, _19769_);
  and _70955_ (_19774_, _19773_, _07132_);
  or _70956_ (_19776_, _19774_, _19726_);
  and _70957_ (_19777_, _19776_, _07130_);
  and _70958_ (_19778_, _19732_, _06411_);
  and _70959_ (_19779_, _19778_, _19722_);
  or _70960_ (_19780_, _19779_, _06303_);
  or _70961_ (_19781_, _19780_, _19777_);
  and _70962_ (_19782_, _15410_, _07856_);
  or _70963_ (_19783_, _19721_, _08819_);
  or _70964_ (_19784_, _19783_, _19782_);
  and _70965_ (_19785_, _19784_, _08824_);
  and _70966_ (_19787_, _19785_, _19781_);
  nor _70967_ (_19788_, _10294_, _11137_);
  or _70968_ (_19789_, _19788_, _19721_);
  and _70969_ (_19790_, _19789_, _06396_);
  or _70970_ (_19791_, _19790_, _06433_);
  or _70971_ (_19792_, _19791_, _19787_);
  or _70972_ (_19793_, _19728_, _06829_);
  and _70973_ (_19794_, _19793_, _06444_);
  and _70974_ (_19795_, _19794_, _19792_);
  and _70975_ (_19796_, _15478_, _07856_);
  or _70976_ (_19798_, _19796_, _19721_);
  and _70977_ (_19799_, _19798_, _06440_);
  or _70978_ (_19800_, _19799_, _01321_);
  or _70979_ (_19801_, _19800_, _19795_);
  or _70980_ (_19802_, _01317_, \oc8051_golden_model_1.PCON [6]);
  and _70981_ (_19803_, _19802_, _43100_);
  and _70982_ (_43618_, _19803_, _19801_);
  not _70983_ (_19804_, \oc8051_golden_model_1.TMOD [0]);
  nor _70984_ (_19805_, _01317_, _19804_);
  nand _70985_ (_19806_, _10276_, _07812_);
  nor _70986_ (_19808_, _07812_, _19804_);
  nor _70987_ (_19809_, _19808_, _07130_);
  nand _70988_ (_19810_, _19809_, _19806_);
  and _70989_ (_19811_, _07812_, _07049_);
  or _70990_ (_19812_, _19811_, _19808_);
  or _70991_ (_19813_, _19812_, _06132_);
  nor _70992_ (_19814_, _08211_, _11214_);
  or _70993_ (_19815_, _19814_, _19808_);
  or _70994_ (_19816_, _19815_, _06161_);
  and _70995_ (_19817_, _07812_, \oc8051_golden_model_1.ACC [0]);
  or _70996_ (_19819_, _19817_, _19808_);
  and _70997_ (_19820_, _19819_, _07056_);
  nor _70998_ (_19821_, _07056_, _19804_);
  or _70999_ (_19822_, _19821_, _06160_);
  or _71000_ (_19823_, _19822_, _19820_);
  and _71001_ (_19824_, _19823_, _07075_);
  and _71002_ (_19825_, _19824_, _19816_);
  and _71003_ (_19826_, _19812_, _06217_);
  or _71004_ (_19827_, _19826_, _19825_);
  and _71005_ (_19828_, _19827_, _06229_);
  and _71006_ (_19830_, _19819_, _06220_);
  or _71007_ (_19831_, _19830_, _09842_);
  or _71008_ (_19832_, _19831_, _19828_);
  and _71009_ (_19833_, _19832_, _19813_);
  or _71010_ (_19834_, _19833_, _06116_);
  and _71011_ (_19835_, _09160_, _07812_);
  or _71012_ (_19836_, _19808_, _06117_);
  or _71013_ (_19837_, _19836_, _19835_);
  and _71014_ (_19838_, _19837_, _19834_);
  or _71015_ (_19839_, _19838_, _05787_);
  and _71016_ (_19841_, _14260_, _07812_);
  or _71017_ (_19842_, _19808_, _06114_);
  or _71018_ (_19843_, _19842_, _19841_);
  and _71019_ (_19844_, _19843_, _06111_);
  and _71020_ (_19845_, _19844_, _19839_);
  and _71021_ (_19846_, _07812_, _08708_);
  or _71022_ (_19847_, _19846_, _19808_);
  and _71023_ (_19848_, _19847_, _06110_);
  or _71024_ (_19849_, _19848_, _06297_);
  or _71025_ (_19850_, _19849_, _19845_);
  and _71026_ (_19852_, _14275_, _07812_);
  or _71027_ (_19853_, _19808_, _07127_);
  or _71028_ (_19854_, _19853_, _19852_);
  and _71029_ (_19855_, _19854_, _07125_);
  and _71030_ (_19856_, _19855_, _19850_);
  nor _71031_ (_19857_, _12321_, _11214_);
  or _71032_ (_19858_, _19857_, _19808_);
  and _71033_ (_19859_, _19806_, _06402_);
  and _71034_ (_19860_, _19859_, _19858_);
  or _71035_ (_19861_, _19860_, _19856_);
  and _71036_ (_19864_, _19861_, _07132_);
  nand _71037_ (_19865_, _19847_, _06306_);
  nor _71038_ (_19866_, _19865_, _19814_);
  or _71039_ (_19867_, _19866_, _06411_);
  or _71040_ (_19868_, _19867_, _19864_);
  and _71041_ (_19869_, _19868_, _19810_);
  or _71042_ (_19870_, _19869_, _06303_);
  and _71043_ (_19871_, _14167_, _07812_);
  or _71044_ (_19872_, _19808_, _08819_);
  or _71045_ (_19873_, _19872_, _19871_);
  and _71046_ (_19876_, _19873_, _08824_);
  and _71047_ (_19877_, _19876_, _19870_);
  and _71048_ (_19878_, _19858_, _06396_);
  or _71049_ (_19879_, _19878_, _19287_);
  or _71050_ (_19880_, _19879_, _19877_);
  or _71051_ (_19881_, _19815_, _06630_);
  and _71052_ (_19882_, _19881_, _01317_);
  and _71053_ (_19883_, _19882_, _19880_);
  or _71054_ (_19884_, _19883_, _19805_);
  and _71055_ (_43619_, _19884_, _43100_);
  and _71056_ (_19887_, _11214_, \oc8051_golden_model_1.TMOD [1]);
  nor _71057_ (_19888_, _10277_, _11214_);
  or _71058_ (_19889_, _19888_, _19887_);
  or _71059_ (_19890_, _19889_, _08824_);
  or _71060_ (_19891_, _14442_, _11214_);
  or _71061_ (_19892_, _07812_, \oc8051_golden_model_1.TMOD [1]);
  and _71062_ (_19893_, _19892_, _05787_);
  and _71063_ (_19894_, _19893_, _19891_);
  and _71064_ (_19895_, _09115_, _07812_);
  or _71065_ (_19896_, _19887_, _06117_);
  or _71066_ (_19899_, _19896_, _19895_);
  and _71067_ (_19900_, _14363_, _07812_);
  not _71068_ (_19901_, _19900_);
  and _71069_ (_19902_, _19901_, _19892_);
  or _71070_ (_19903_, _19902_, _06161_);
  and _71071_ (_19904_, _07812_, \oc8051_golden_model_1.ACC [1]);
  or _71072_ (_19905_, _19904_, _19887_);
  and _71073_ (_19906_, _19905_, _07056_);
  and _71074_ (_19907_, _07057_, \oc8051_golden_model_1.TMOD [1]);
  or _71075_ (_19908_, _19907_, _06160_);
  or _71076_ (_19911_, _19908_, _19906_);
  and _71077_ (_19912_, _19911_, _07075_);
  and _71078_ (_19913_, _19912_, _19903_);
  and _71079_ (_19914_, _07812_, _07306_);
  or _71080_ (_19915_, _19914_, _19887_);
  and _71081_ (_19916_, _19915_, _06217_);
  or _71082_ (_19917_, _19916_, _19913_);
  and _71083_ (_19918_, _19917_, _06229_);
  and _71084_ (_19919_, _19905_, _06220_);
  or _71085_ (_19920_, _19919_, _09842_);
  or _71086_ (_19923_, _19920_, _19918_);
  or _71087_ (_19924_, _19915_, _06132_);
  and _71088_ (_19925_, _19924_, _19923_);
  or _71089_ (_19926_, _19925_, _06116_);
  and _71090_ (_19927_, _19926_, _06114_);
  and _71091_ (_19928_, _19927_, _19899_);
  or _71092_ (_19929_, _19928_, _19894_);
  and _71093_ (_19930_, _19929_, _06298_);
  or _71094_ (_19931_, _14346_, _11214_);
  and _71095_ (_19932_, _19931_, _06297_);
  nand _71096_ (_19935_, _07812_, _06945_);
  and _71097_ (_19936_, _19935_, _06110_);
  or _71098_ (_19937_, _19936_, _19932_);
  and _71099_ (_19938_, _19937_, _19892_);
  or _71100_ (_19939_, _19938_, _06402_);
  or _71101_ (_19940_, _19939_, _19930_);
  nand _71102_ (_19941_, _10275_, _07812_);
  and _71103_ (_19942_, _19941_, _19889_);
  or _71104_ (_19943_, _19942_, _07125_);
  and _71105_ (_19944_, _19943_, _07132_);
  and _71106_ (_19946_, _19944_, _19940_);
  or _71107_ (_19947_, _14344_, _11214_);
  and _71108_ (_19948_, _19892_, _06306_);
  and _71109_ (_19949_, _19948_, _19947_);
  or _71110_ (_19950_, _19949_, _06411_);
  or _71111_ (_19951_, _19950_, _19946_);
  nor _71112_ (_19952_, _19887_, _07130_);
  nand _71113_ (_19953_, _19952_, _19941_);
  and _71114_ (_19954_, _19953_, _08819_);
  and _71115_ (_19955_, _19954_, _19951_);
  or _71116_ (_19957_, _19935_, _08176_);
  and _71117_ (_19958_, _19892_, _06303_);
  and _71118_ (_19959_, _19958_, _19957_);
  or _71119_ (_19960_, _19959_, _06396_);
  or _71120_ (_19961_, _19960_, _19955_);
  and _71121_ (_19962_, _19961_, _19890_);
  or _71122_ (_19963_, _19962_, _06433_);
  or _71123_ (_19964_, _19902_, _06829_);
  and _71124_ (_19965_, _19964_, _06444_);
  and _71125_ (_19966_, _19965_, _19963_);
  or _71126_ (_19968_, _19900_, _19887_);
  and _71127_ (_19969_, _19968_, _06440_);
  or _71128_ (_19970_, _19969_, _01321_);
  or _71129_ (_19971_, _19970_, _19966_);
  or _71130_ (_19972_, _01317_, \oc8051_golden_model_1.TMOD [1]);
  and _71131_ (_19973_, _19972_, _43100_);
  and _71132_ (_43621_, _19973_, _19971_);
  and _71133_ (_19974_, _01321_, \oc8051_golden_model_1.TMOD [2]);
  and _71134_ (_19975_, _11214_, \oc8051_golden_model_1.TMOD [2]);
  and _71135_ (_19976_, _09211_, _07812_);
  or _71136_ (_19978_, _19976_, _19975_);
  and _71137_ (_19979_, _19978_, _06116_);
  and _71138_ (_19980_, _14542_, _07812_);
  or _71139_ (_19981_, _19980_, _19975_);
  or _71140_ (_19982_, _19981_, _06161_);
  and _71141_ (_19983_, _07812_, \oc8051_golden_model_1.ACC [2]);
  or _71142_ (_19984_, _19983_, _19975_);
  and _71143_ (_19985_, _19984_, _07056_);
  and _71144_ (_19986_, _07057_, \oc8051_golden_model_1.TMOD [2]);
  or _71145_ (_19987_, _19986_, _06160_);
  or _71146_ (_19989_, _19987_, _19985_);
  and _71147_ (_19990_, _19989_, _07075_);
  and _71148_ (_19991_, _19990_, _19982_);
  and _71149_ (_19992_, _07812_, _07708_);
  or _71150_ (_19993_, _19992_, _19975_);
  and _71151_ (_19994_, _19993_, _06217_);
  or _71152_ (_19995_, _19994_, _19991_);
  and _71153_ (_19996_, _19995_, _06229_);
  and _71154_ (_19997_, _19984_, _06220_);
  or _71155_ (_19998_, _19997_, _09842_);
  or _71156_ (_20000_, _19998_, _19996_);
  or _71157_ (_20001_, _19993_, _06132_);
  and _71158_ (_20002_, _20001_, _06117_);
  and _71159_ (_20003_, _20002_, _20000_);
  or _71160_ (_20004_, _20003_, _05787_);
  or _71161_ (_20005_, _20004_, _19979_);
  and _71162_ (_20006_, _14630_, _07812_);
  or _71163_ (_20007_, _20006_, _19975_);
  or _71164_ (_20008_, _20007_, _06114_);
  and _71165_ (_20009_, _20008_, _06111_);
  and _71166_ (_20011_, _20009_, _20005_);
  and _71167_ (_20012_, _07812_, _08768_);
  or _71168_ (_20013_, _20012_, _19975_);
  and _71169_ (_20014_, _20013_, _06110_);
  or _71170_ (_20015_, _20014_, _06297_);
  or _71171_ (_20016_, _20015_, _20011_);
  and _71172_ (_20017_, _14646_, _07812_);
  or _71173_ (_20018_, _19975_, _07127_);
  or _71174_ (_20019_, _20018_, _20017_);
  and _71175_ (_20020_, _20019_, _07125_);
  and _71176_ (_20022_, _20020_, _20016_);
  and _71177_ (_20023_, _10282_, _07812_);
  or _71178_ (_20024_, _20023_, _19975_);
  and _71179_ (_20025_, _20024_, _06402_);
  or _71180_ (_20026_, _20025_, _20022_);
  and _71181_ (_20027_, _20026_, _07132_);
  or _71182_ (_20028_, _19975_, _08248_);
  and _71183_ (_20029_, _20013_, _06306_);
  and _71184_ (_20030_, _20029_, _20028_);
  or _71185_ (_20031_, _20030_, _20027_);
  and _71186_ (_20033_, _20031_, _07130_);
  and _71187_ (_20034_, _19984_, _06411_);
  and _71188_ (_20035_, _20034_, _20028_);
  or _71189_ (_20036_, _20035_, _06303_);
  or _71190_ (_20037_, _20036_, _20033_);
  and _71191_ (_20038_, _14643_, _07812_);
  or _71192_ (_20039_, _19975_, _08819_);
  or _71193_ (_20040_, _20039_, _20038_);
  and _71194_ (_20041_, _20040_, _08824_);
  and _71195_ (_20042_, _20041_, _20037_);
  nor _71196_ (_20044_, _10281_, _11214_);
  or _71197_ (_20045_, _20044_, _19975_);
  and _71198_ (_20046_, _20045_, _06396_);
  or _71199_ (_20047_, _20046_, _20042_);
  and _71200_ (_20048_, _20047_, _06829_);
  and _71201_ (_20049_, _19981_, _06433_);
  or _71202_ (_20050_, _20049_, _06440_);
  or _71203_ (_20051_, _20050_, _20048_);
  and _71204_ (_20052_, _14710_, _07812_);
  or _71205_ (_20053_, _19975_, _06444_);
  or _71206_ (_20055_, _20053_, _20052_);
  and _71207_ (_20056_, _20055_, _01317_);
  and _71208_ (_20057_, _20056_, _20051_);
  or _71209_ (_20058_, _20057_, _19974_);
  and _71210_ (_43622_, _20058_, _43100_);
  and _71211_ (_20059_, _11214_, \oc8051_golden_model_1.TMOD [3]);
  and _71212_ (_20060_, _14738_, _07812_);
  or _71213_ (_20061_, _20060_, _20059_);
  or _71214_ (_20062_, _20061_, _06161_);
  and _71215_ (_20063_, _07812_, \oc8051_golden_model_1.ACC [3]);
  or _71216_ (_20065_, _20063_, _20059_);
  and _71217_ (_20066_, _20065_, _07056_);
  and _71218_ (_20067_, _07057_, \oc8051_golden_model_1.TMOD [3]);
  or _71219_ (_20068_, _20067_, _06160_);
  or _71220_ (_20069_, _20068_, _20066_);
  and _71221_ (_20070_, _20069_, _07075_);
  and _71222_ (_20071_, _20070_, _20062_);
  and _71223_ (_20072_, _07812_, _07544_);
  or _71224_ (_20073_, _20072_, _20059_);
  and _71225_ (_20074_, _20073_, _06217_);
  or _71226_ (_20076_, _20074_, _20071_);
  and _71227_ (_20077_, _20076_, _06229_);
  and _71228_ (_20078_, _20065_, _06220_);
  or _71229_ (_20079_, _20078_, _09842_);
  or _71230_ (_20080_, _20079_, _20077_);
  or _71231_ (_20081_, _20073_, _06132_);
  and _71232_ (_20082_, _20081_, _20080_);
  or _71233_ (_20083_, _20082_, _06116_);
  and _71234_ (_20084_, _09210_, _07812_);
  or _71235_ (_20085_, _20059_, _06117_);
  or _71236_ (_20087_, _20085_, _20084_);
  and _71237_ (_20088_, _20087_, _06114_);
  and _71238_ (_20089_, _20088_, _20083_);
  and _71239_ (_20090_, _14825_, _07812_);
  or _71240_ (_20091_, _20090_, _20059_);
  and _71241_ (_20092_, _20091_, _05787_);
  or _71242_ (_20093_, _20092_, _11136_);
  or _71243_ (_20094_, _20093_, _20089_);
  and _71244_ (_20095_, _14727_, _07812_);
  or _71245_ (_20096_, _20059_, _07127_);
  or _71246_ (_20098_, _20096_, _20095_);
  and _71247_ (_20099_, _07812_, _08712_);
  or _71248_ (_20100_, _20099_, _20059_);
  or _71249_ (_20101_, _20100_, _06111_);
  and _71250_ (_20102_, _20101_, _07125_);
  and _71251_ (_20103_, _20102_, _20098_);
  and _71252_ (_20104_, _20103_, _20094_);
  and _71253_ (_20105_, _12318_, _07812_);
  or _71254_ (_20106_, _20105_, _20059_);
  and _71255_ (_20107_, _20106_, _06402_);
  or _71256_ (_20109_, _20107_, _20104_);
  and _71257_ (_20110_, _20109_, _07132_);
  or _71258_ (_20111_, _20059_, _08140_);
  and _71259_ (_20112_, _20100_, _06306_);
  and _71260_ (_20113_, _20112_, _20111_);
  or _71261_ (_20114_, _20113_, _20110_);
  and _71262_ (_20115_, _20114_, _07130_);
  and _71263_ (_20116_, _20065_, _06411_);
  and _71264_ (_20117_, _20116_, _20111_);
  or _71265_ (_20118_, _20117_, _06303_);
  or _71266_ (_20120_, _20118_, _20115_);
  and _71267_ (_20121_, _14724_, _07812_);
  or _71268_ (_20122_, _20059_, _08819_);
  or _71269_ (_20123_, _20122_, _20121_);
  and _71270_ (_20124_, _20123_, _08824_);
  and _71271_ (_20125_, _20124_, _20120_);
  nor _71272_ (_20126_, _10273_, _11214_);
  or _71273_ (_20127_, _20126_, _20059_);
  and _71274_ (_20128_, _20127_, _06396_);
  or _71275_ (_20129_, _20128_, _06433_);
  or _71276_ (_20131_, _20129_, _20125_);
  or _71277_ (_20132_, _20061_, _06829_);
  and _71278_ (_20133_, _20132_, _06444_);
  and _71279_ (_20134_, _20133_, _20131_);
  and _71280_ (_20135_, _14897_, _07812_);
  or _71281_ (_20136_, _20135_, _20059_);
  and _71282_ (_20137_, _20136_, _06440_);
  or _71283_ (_20138_, _20137_, _01321_);
  or _71284_ (_20139_, _20138_, _20134_);
  or _71285_ (_20140_, _01317_, \oc8051_golden_model_1.TMOD [3]);
  and _71286_ (_20142_, _20140_, _43100_);
  and _71287_ (_43623_, _20142_, _20139_);
  and _71288_ (_20143_, _11214_, \oc8051_golden_model_1.TMOD [4]);
  and _71289_ (_20144_, _08336_, _07812_);
  or _71290_ (_20145_, _20144_, _20143_);
  or _71291_ (_20146_, _20145_, _06132_);
  and _71292_ (_20147_, _14928_, _07812_);
  or _71293_ (_20148_, _20147_, _20143_);
  or _71294_ (_20149_, _20148_, _06161_);
  and _71295_ (_20150_, _07812_, \oc8051_golden_model_1.ACC [4]);
  or _71296_ (_20152_, _20150_, _20143_);
  and _71297_ (_20153_, _20152_, _07056_);
  and _71298_ (_20154_, _07057_, \oc8051_golden_model_1.TMOD [4]);
  or _71299_ (_20155_, _20154_, _06160_);
  or _71300_ (_20156_, _20155_, _20153_);
  and _71301_ (_20157_, _20156_, _07075_);
  and _71302_ (_20158_, _20157_, _20149_);
  and _71303_ (_20159_, _20145_, _06217_);
  or _71304_ (_20160_, _20159_, _20158_);
  and _71305_ (_20161_, _20160_, _06229_);
  and _71306_ (_20163_, _20152_, _06220_);
  or _71307_ (_20164_, _20163_, _09842_);
  or _71308_ (_20165_, _20164_, _20161_);
  and _71309_ (_20166_, _20165_, _20146_);
  or _71310_ (_20167_, _20166_, _06116_);
  and _71311_ (_20168_, _09209_, _07812_);
  or _71312_ (_20169_, _20143_, _06117_);
  or _71313_ (_20170_, _20169_, _20168_);
  and _71314_ (_20171_, _20170_, _06114_);
  and _71315_ (_20172_, _20171_, _20167_);
  and _71316_ (_20174_, _15013_, _07812_);
  or _71317_ (_20175_, _20174_, _20143_);
  and _71318_ (_20176_, _20175_, _05787_);
  or _71319_ (_20177_, _20176_, _20172_);
  or _71320_ (_20178_, _20177_, _11136_);
  and _71321_ (_20179_, _15029_, _07812_);
  or _71322_ (_20180_, _20143_, _07127_);
  or _71323_ (_20181_, _20180_, _20179_);
  and _71324_ (_20182_, _08715_, _07812_);
  or _71325_ (_20183_, _20182_, _20143_);
  or _71326_ (_20185_, _20183_, _06111_);
  and _71327_ (_20186_, _20185_, _07125_);
  and _71328_ (_20187_, _20186_, _20181_);
  and _71329_ (_20188_, _20187_, _20178_);
  and _71330_ (_20189_, _10289_, _07812_);
  or _71331_ (_20190_, _20189_, _20143_);
  and _71332_ (_20191_, _20190_, _06402_);
  or _71333_ (_20192_, _20191_, _20188_);
  and _71334_ (_20193_, _20192_, _07132_);
  or _71335_ (_20194_, _20143_, _08339_);
  and _71336_ (_20196_, _20183_, _06306_);
  and _71337_ (_20197_, _20196_, _20194_);
  or _71338_ (_20198_, _20197_, _20193_);
  and _71339_ (_20199_, _20198_, _07130_);
  and _71340_ (_20200_, _20152_, _06411_);
  and _71341_ (_20201_, _20200_, _20194_);
  or _71342_ (_20202_, _20201_, _06303_);
  or _71343_ (_20203_, _20202_, _20199_);
  and _71344_ (_20204_, _15026_, _07812_);
  or _71345_ (_20205_, _20143_, _08819_);
  or _71346_ (_20207_, _20205_, _20204_);
  and _71347_ (_20208_, _20207_, _08824_);
  and _71348_ (_20209_, _20208_, _20203_);
  nor _71349_ (_20210_, _10288_, _11214_);
  or _71350_ (_20211_, _20210_, _20143_);
  and _71351_ (_20212_, _20211_, _06396_);
  or _71352_ (_20213_, _20212_, _06433_);
  or _71353_ (_20214_, _20213_, _20209_);
  or _71354_ (_20215_, _20148_, _06829_);
  and _71355_ (_20216_, _20215_, _06444_);
  and _71356_ (_20218_, _20216_, _20214_);
  and _71357_ (_20219_, _15087_, _07812_);
  or _71358_ (_20220_, _20219_, _20143_);
  and _71359_ (_20221_, _20220_, _06440_);
  or _71360_ (_20222_, _20221_, _01321_);
  or _71361_ (_20223_, _20222_, _20218_);
  or _71362_ (_20224_, _01317_, \oc8051_golden_model_1.TMOD [4]);
  and _71363_ (_20225_, _20224_, _43100_);
  and _71364_ (_43624_, _20225_, _20223_);
  and _71365_ (_20226_, _11214_, \oc8051_golden_model_1.TMOD [5]);
  and _71366_ (_20228_, _15119_, _07812_);
  or _71367_ (_20229_, _20228_, _20226_);
  or _71368_ (_20230_, _20229_, _06161_);
  and _71369_ (_20231_, _07812_, \oc8051_golden_model_1.ACC [5]);
  or _71370_ (_20232_, _20231_, _20226_);
  and _71371_ (_20233_, _20232_, _07056_);
  and _71372_ (_20234_, _07057_, \oc8051_golden_model_1.TMOD [5]);
  or _71373_ (_20235_, _20234_, _06160_);
  or _71374_ (_20236_, _20235_, _20233_);
  and _71375_ (_20237_, _20236_, _07075_);
  and _71376_ (_20239_, _20237_, _20230_);
  and _71377_ (_20240_, _08101_, _07812_);
  or _71378_ (_20241_, _20240_, _20226_);
  and _71379_ (_20242_, _20241_, _06217_);
  or _71380_ (_20243_, _20242_, _20239_);
  and _71381_ (_20244_, _20243_, _06229_);
  and _71382_ (_20245_, _20232_, _06220_);
  or _71383_ (_20246_, _20245_, _09842_);
  or _71384_ (_20247_, _20246_, _20244_);
  or _71385_ (_20248_, _20241_, _06132_);
  and _71386_ (_20250_, _20248_, _20247_);
  or _71387_ (_20251_, _20250_, _06116_);
  and _71388_ (_20252_, _09208_, _07812_);
  or _71389_ (_20253_, _20226_, _06117_);
  or _71390_ (_20254_, _20253_, _20252_);
  and _71391_ (_20255_, _20254_, _06114_);
  and _71392_ (_20256_, _20255_, _20251_);
  and _71393_ (_20257_, _15203_, _07812_);
  or _71394_ (_20258_, _20257_, _20226_);
  and _71395_ (_20259_, _20258_, _05787_);
  or _71396_ (_20261_, _20259_, _11136_);
  or _71397_ (_20262_, _20261_, _20256_);
  and _71398_ (_20263_, _15219_, _07812_);
  or _71399_ (_20264_, _20226_, _07127_);
  or _71400_ (_20265_, _20264_, _20263_);
  and _71401_ (_20266_, _08736_, _07812_);
  or _71402_ (_20267_, _20266_, _20226_);
  or _71403_ (_20268_, _20267_, _06111_);
  and _71404_ (_20269_, _20268_, _07125_);
  and _71405_ (_20270_, _20269_, _20265_);
  and _71406_ (_20272_, _20270_, _20262_);
  and _71407_ (_20273_, _12325_, _07812_);
  or _71408_ (_20274_, _20273_, _20226_);
  and _71409_ (_20275_, _20274_, _06402_);
  or _71410_ (_20276_, _20275_, _20272_);
  and _71411_ (_20277_, _20276_, _07132_);
  or _71412_ (_20278_, _20226_, _08104_);
  and _71413_ (_20279_, _20267_, _06306_);
  and _71414_ (_20280_, _20279_, _20278_);
  or _71415_ (_20281_, _20280_, _20277_);
  and _71416_ (_20283_, _20281_, _07130_);
  and _71417_ (_20284_, _20232_, _06411_);
  and _71418_ (_20285_, _20284_, _20278_);
  or _71419_ (_20286_, _20285_, _06303_);
  or _71420_ (_20287_, _20286_, _20283_);
  and _71421_ (_20288_, _15216_, _07812_);
  or _71422_ (_20289_, _20226_, _08819_);
  or _71423_ (_20290_, _20289_, _20288_);
  and _71424_ (_20291_, _20290_, _08824_);
  and _71425_ (_20292_, _20291_, _20287_);
  nor _71426_ (_20294_, _10269_, _11214_);
  or _71427_ (_20295_, _20294_, _20226_);
  and _71428_ (_20296_, _20295_, _06396_);
  or _71429_ (_20297_, _20296_, _06433_);
  or _71430_ (_20298_, _20297_, _20292_);
  or _71431_ (_20299_, _20229_, _06829_);
  and _71432_ (_20300_, _20299_, _06444_);
  and _71433_ (_20301_, _20300_, _20298_);
  and _71434_ (_20302_, _15275_, _07812_);
  or _71435_ (_20303_, _20302_, _20226_);
  and _71436_ (_20305_, _20303_, _06440_);
  or _71437_ (_20306_, _20305_, _01321_);
  or _71438_ (_20307_, _20306_, _20301_);
  or _71439_ (_20308_, _01317_, \oc8051_golden_model_1.TMOD [5]);
  and _71440_ (_20309_, _20308_, _43100_);
  and _71441_ (_43625_, _20309_, _20307_);
  and _71442_ (_20310_, _11214_, \oc8051_golden_model_1.TMOD [6]);
  and _71443_ (_20311_, _15300_, _07812_);
  or _71444_ (_20312_, _20311_, _20310_);
  or _71445_ (_20313_, _20312_, _06161_);
  and _71446_ (_20315_, _07812_, \oc8051_golden_model_1.ACC [6]);
  or _71447_ (_20316_, _20315_, _20310_);
  and _71448_ (_20317_, _20316_, _07056_);
  and _71449_ (_20318_, _07057_, \oc8051_golden_model_1.TMOD [6]);
  or _71450_ (_20319_, _20318_, _06160_);
  or _71451_ (_20320_, _20319_, _20317_);
  and _71452_ (_20321_, _20320_, _07075_);
  and _71453_ (_20322_, _20321_, _20313_);
  and _71454_ (_20323_, _08012_, _07812_);
  or _71455_ (_20324_, _20323_, _20310_);
  and _71456_ (_20326_, _20324_, _06217_);
  or _71457_ (_20327_, _20326_, _20322_);
  and _71458_ (_20328_, _20327_, _06229_);
  and _71459_ (_20329_, _20316_, _06220_);
  or _71460_ (_20330_, _20329_, _09842_);
  or _71461_ (_20331_, _20330_, _20328_);
  or _71462_ (_20332_, _20324_, _06132_);
  and _71463_ (_20333_, _20332_, _20331_);
  or _71464_ (_20334_, _20333_, _06116_);
  and _71465_ (_20335_, _09207_, _07812_);
  or _71466_ (_20337_, _20310_, _06117_);
  or _71467_ (_20338_, _20337_, _20335_);
  and _71468_ (_20339_, _20338_, _06114_);
  and _71469_ (_20340_, _20339_, _20334_);
  and _71470_ (_20341_, _15395_, _07812_);
  or _71471_ (_20342_, _20341_, _20310_);
  and _71472_ (_20343_, _20342_, _05787_);
  or _71473_ (_20344_, _20343_, _11136_);
  or _71474_ (_20345_, _20344_, _20340_);
  and _71475_ (_20346_, _15413_, _07812_);
  or _71476_ (_20348_, _20310_, _07127_);
  or _71477_ (_20349_, _20348_, _20346_);
  and _71478_ (_20350_, _15402_, _07812_);
  or _71479_ (_20351_, _20350_, _20310_);
  or _71480_ (_20352_, _20351_, _06111_);
  and _71481_ (_20353_, _20352_, _07125_);
  and _71482_ (_20354_, _20353_, _20349_);
  and _71483_ (_20355_, _20354_, _20345_);
  and _71484_ (_20356_, _10295_, _07812_);
  or _71485_ (_20357_, _20356_, _20310_);
  and _71486_ (_20359_, _20357_, _06402_);
  or _71487_ (_20360_, _20359_, _20355_);
  and _71488_ (_20361_, _20360_, _07132_);
  or _71489_ (_20362_, _20310_, _08015_);
  and _71490_ (_20363_, _20351_, _06306_);
  and _71491_ (_20364_, _20363_, _20362_);
  or _71492_ (_20365_, _20364_, _20361_);
  and _71493_ (_20366_, _20365_, _07130_);
  and _71494_ (_20367_, _20316_, _06411_);
  and _71495_ (_20368_, _20367_, _20362_);
  or _71496_ (_20370_, _20368_, _06303_);
  or _71497_ (_20371_, _20370_, _20366_);
  and _71498_ (_20372_, _15410_, _07812_);
  or _71499_ (_20373_, _20310_, _08819_);
  or _71500_ (_20374_, _20373_, _20372_);
  and _71501_ (_20375_, _20374_, _08824_);
  and _71502_ (_20376_, _20375_, _20371_);
  nor _71503_ (_20377_, _10294_, _11214_);
  or _71504_ (_20378_, _20377_, _20310_);
  and _71505_ (_20379_, _20378_, _06396_);
  or _71506_ (_20381_, _20379_, _06433_);
  or _71507_ (_20382_, _20381_, _20376_);
  or _71508_ (_20383_, _20312_, _06829_);
  and _71509_ (_20384_, _20383_, _06444_);
  and _71510_ (_20385_, _20384_, _20382_);
  and _71511_ (_20386_, _15478_, _07812_);
  or _71512_ (_20387_, _20386_, _20310_);
  and _71513_ (_20388_, _20387_, _06440_);
  or _71514_ (_20389_, _20388_, _01321_);
  or _71515_ (_20390_, _20389_, _20385_);
  or _71516_ (_20392_, _01317_, \oc8051_golden_model_1.TMOD [6]);
  and _71517_ (_20393_, _20392_, _43100_);
  and _71518_ (_43626_, _20393_, _20390_);
  not _71519_ (_20394_, \oc8051_golden_model_1.DPL [0]);
  nor _71520_ (_20395_, _01317_, _20394_);
  nand _71521_ (_20396_, _10276_, _07849_);
  nor _71522_ (_20397_, _07849_, _20394_);
  nor _71523_ (_20398_, _20397_, _07130_);
  nand _71524_ (_20399_, _20398_, _20396_);
  and _71525_ (_20400_, _07849_, _07049_);
  or _71526_ (_20402_, _20400_, _20397_);
  or _71527_ (_20403_, _20402_, _06132_);
  and _71528_ (_20404_, _07849_, \oc8051_golden_model_1.ACC [0]);
  or _71529_ (_20405_, _20404_, _20397_);
  or _71530_ (_20406_, _20405_, _06229_);
  nor _71531_ (_20407_, _08211_, _11371_);
  or _71532_ (_20408_, _20407_, _20397_);
  or _71533_ (_20409_, _20408_, _06161_);
  and _71534_ (_20410_, _20405_, _07056_);
  nor _71535_ (_20411_, _07056_, _20394_);
  or _71536_ (_20413_, _20411_, _06160_);
  or _71537_ (_20414_, _20413_, _20410_);
  and _71538_ (_20415_, _20414_, _07075_);
  and _71539_ (_20416_, _20415_, _20409_);
  and _71540_ (_20417_, _20402_, _06217_);
  or _71541_ (_20418_, _20417_, _06220_);
  or _71542_ (_20419_, _20418_, _20416_);
  and _71543_ (_20420_, _20419_, _20406_);
  or _71544_ (_20421_, _20420_, _11311_);
  nand _71545_ (_20422_, _11311_, \oc8051_golden_model_1.DPL [0]);
  and _71546_ (_20424_, _20422_, _11296_);
  and _71547_ (_20425_, _20424_, _20421_);
  nor _71548_ (_20426_, _06758_, _11296_);
  or _71549_ (_20427_, _20426_, _09842_);
  or _71550_ (_20428_, _20427_, _20425_);
  and _71551_ (_20429_, _20428_, _20403_);
  or _71552_ (_20430_, _20429_, _06116_);
  and _71553_ (_20431_, _09160_, _07849_);
  or _71554_ (_20432_, _20397_, _06117_);
  or _71555_ (_20433_, _20432_, _20431_);
  and _71556_ (_20435_, _20433_, _20430_);
  or _71557_ (_20436_, _20435_, _05787_);
  and _71558_ (_20437_, _14260_, _07849_);
  or _71559_ (_20438_, _20437_, _20397_);
  or _71560_ (_20439_, _20438_, _06114_);
  and _71561_ (_20440_, _20439_, _06111_);
  and _71562_ (_20441_, _20440_, _20436_);
  and _71563_ (_20442_, _07849_, _08708_);
  or _71564_ (_20443_, _20442_, _20397_);
  and _71565_ (_20444_, _20443_, _06110_);
  or _71566_ (_20446_, _20444_, _06297_);
  or _71567_ (_20447_, _20446_, _20441_);
  and _71568_ (_20448_, _14275_, _07849_);
  or _71569_ (_20449_, _20448_, _20397_);
  or _71570_ (_20450_, _20449_, _07127_);
  and _71571_ (_20451_, _20450_, _07125_);
  and _71572_ (_20452_, _20451_, _20447_);
  nor _71573_ (_20453_, _12321_, _11371_);
  or _71574_ (_20454_, _20453_, _20397_);
  and _71575_ (_20455_, _20396_, _06402_);
  and _71576_ (_20457_, _20455_, _20454_);
  or _71577_ (_20458_, _20457_, _20452_);
  and _71578_ (_20459_, _20458_, _07132_);
  nand _71579_ (_20460_, _20443_, _06306_);
  nor _71580_ (_20461_, _20460_, _20407_);
  or _71581_ (_20462_, _20461_, _06411_);
  or _71582_ (_20463_, _20462_, _20459_);
  and _71583_ (_20464_, _20463_, _20399_);
  or _71584_ (_20465_, _20464_, _06303_);
  and _71585_ (_20466_, _14167_, _07849_);
  or _71586_ (_20468_, _20397_, _08819_);
  or _71587_ (_20469_, _20468_, _20466_);
  and _71588_ (_20470_, _20469_, _08824_);
  and _71589_ (_20471_, _20470_, _20465_);
  and _71590_ (_20472_, _20454_, _06396_);
  or _71591_ (_20473_, _20472_, _19287_);
  or _71592_ (_20474_, _20473_, _20471_);
  or _71593_ (_20475_, _20408_, _06630_);
  and _71594_ (_20476_, _20475_, _01317_);
  and _71595_ (_20477_, _20476_, _20474_);
  or _71596_ (_20479_, _20477_, _20395_);
  and _71597_ (_43628_, _20479_, _43100_);
  not _71598_ (_20480_, \oc8051_golden_model_1.DPL [1]);
  nor _71599_ (_20481_, _01317_, _20480_);
  and _71600_ (_20482_, _09115_, _07849_);
  nor _71601_ (_20483_, _07849_, _20480_);
  or _71602_ (_20484_, _20483_, _20482_);
  and _71603_ (_20485_, _20484_, _06116_);
  or _71604_ (_20486_, _07849_, \oc8051_golden_model_1.DPL [1]);
  and _71605_ (_20487_, _14363_, _07849_);
  not _71606_ (_20489_, _20487_);
  and _71607_ (_20490_, _20489_, _20486_);
  or _71608_ (_20491_, _20490_, _06161_);
  and _71609_ (_20492_, _07849_, \oc8051_golden_model_1.ACC [1]);
  or _71610_ (_20493_, _20492_, _20483_);
  and _71611_ (_20494_, _20493_, _07056_);
  nor _71612_ (_20495_, _07056_, _20480_);
  or _71613_ (_20496_, _20495_, _06160_);
  or _71614_ (_20497_, _20496_, _20494_);
  and _71615_ (_20498_, _20497_, _07075_);
  and _71616_ (_20500_, _20498_, _20491_);
  and _71617_ (_20501_, _07849_, _07306_);
  or _71618_ (_20502_, _20501_, _20483_);
  and _71619_ (_20503_, _20502_, _06217_);
  or _71620_ (_20504_, _20503_, _06220_);
  or _71621_ (_20505_, _20504_, _20500_);
  or _71622_ (_20506_, _20493_, _06229_);
  and _71623_ (_20507_, _20506_, _11312_);
  and _71624_ (_20508_, _20507_, _20505_);
  nor _71625_ (_20509_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor _71626_ (_20511_, _20509_, _11316_);
  and _71627_ (_20512_, _20511_, _11311_);
  or _71628_ (_20513_, _20512_, _20508_);
  and _71629_ (_20514_, _20513_, _11296_);
  nor _71630_ (_20515_, _06945_, _11296_);
  or _71631_ (_20516_, _20515_, _09842_);
  or _71632_ (_20517_, _20516_, _20514_);
  or _71633_ (_20518_, _20502_, _06132_);
  and _71634_ (_20519_, _20518_, _06117_);
  and _71635_ (_20520_, _20519_, _20517_);
  or _71636_ (_20522_, _20520_, _20485_);
  and _71637_ (_20523_, _20522_, _06114_);
  or _71638_ (_20524_, _14442_, _11371_);
  and _71639_ (_20525_, _20486_, _05787_);
  and _71640_ (_20526_, _20525_, _20524_);
  or _71641_ (_20527_, _20526_, _20523_);
  and _71642_ (_20528_, _20527_, _06298_);
  or _71643_ (_20529_, _14346_, _11371_);
  and _71644_ (_20530_, _20529_, _06297_);
  nand _71645_ (_20531_, _07849_, _06945_);
  and _71646_ (_20533_, _20531_, _06110_);
  or _71647_ (_20534_, _20533_, _20530_);
  and _71648_ (_20535_, _20534_, _20486_);
  or _71649_ (_20536_, _20535_, _06402_);
  or _71650_ (_20537_, _20536_, _20528_);
  nor _71651_ (_20538_, _10277_, _11371_);
  or _71652_ (_20539_, _20538_, _20483_);
  nand _71653_ (_20540_, _10275_, _07849_);
  and _71654_ (_20541_, _20540_, _20539_);
  or _71655_ (_20542_, _20541_, _07125_);
  and _71656_ (_20544_, _20542_, _07132_);
  and _71657_ (_20545_, _20544_, _20537_);
  or _71658_ (_20546_, _14344_, _11371_);
  and _71659_ (_20547_, _20486_, _06306_);
  and _71660_ (_20548_, _20547_, _20546_);
  or _71661_ (_20549_, _20548_, _06411_);
  or _71662_ (_20550_, _20549_, _20545_);
  nor _71663_ (_20551_, _20483_, _07130_);
  nand _71664_ (_20552_, _20551_, _20540_);
  and _71665_ (_20553_, _20552_, _08819_);
  and _71666_ (_20555_, _20553_, _20550_);
  or _71667_ (_20556_, _20531_, _08176_);
  and _71668_ (_20557_, _20486_, _06303_);
  and _71669_ (_20558_, _20557_, _20556_);
  or _71670_ (_20559_, _20558_, _06396_);
  or _71671_ (_20560_, _20559_, _20555_);
  or _71672_ (_20561_, _20539_, _08824_);
  and _71673_ (_20562_, _20561_, _06829_);
  and _71674_ (_20563_, _20562_, _20560_);
  and _71675_ (_20564_, _20490_, _06433_);
  or _71676_ (_20566_, _20564_, _06440_);
  or _71677_ (_20567_, _20566_, _20563_);
  or _71678_ (_20568_, _20483_, _06444_);
  or _71679_ (_20569_, _20568_, _20487_);
  and _71680_ (_20570_, _20569_, _01317_);
  and _71681_ (_20571_, _20570_, _20567_);
  or _71682_ (_20572_, _20571_, _20481_);
  and _71683_ (_43629_, _20572_, _43100_);
  not _71684_ (_20573_, \oc8051_golden_model_1.DPL [2]);
  nor _71685_ (_20574_, _01317_, _20573_);
  nor _71686_ (_20576_, _07849_, _20573_);
  or _71687_ (_20577_, _20576_, _08248_);
  and _71688_ (_20578_, _07849_, _08768_);
  or _71689_ (_20579_, _20578_, _20576_);
  and _71690_ (_20580_, _20579_, _06306_);
  and _71691_ (_20581_, _20580_, _20577_);
  and _71692_ (_20582_, _07849_, _07708_);
  or _71693_ (_20583_, _20582_, _20576_);
  or _71694_ (_20584_, _20583_, _07075_);
  and _71695_ (_20585_, _14542_, _07849_);
  or _71696_ (_20587_, _20585_, _20576_);
  and _71697_ (_20588_, _20587_, _06160_);
  nor _71698_ (_20589_, _07056_, _20573_);
  and _71699_ (_20590_, _07849_, \oc8051_golden_model_1.ACC [2]);
  or _71700_ (_20591_, _20590_, _20576_);
  and _71701_ (_20592_, _20591_, _07056_);
  or _71702_ (_20593_, _20592_, _20589_);
  and _71703_ (_20594_, _20593_, _06161_);
  or _71704_ (_20595_, _20594_, _06217_);
  or _71705_ (_20596_, _20595_, _20588_);
  and _71706_ (_20598_, _20596_, _20584_);
  or _71707_ (_20599_, _20598_, _06220_);
  or _71708_ (_20600_, _20591_, _06229_);
  and _71709_ (_20601_, _20600_, _11312_);
  and _71710_ (_20602_, _20601_, _20599_);
  nor _71711_ (_20603_, _11316_, \oc8051_golden_model_1.DPL [2]);
  nor _71712_ (_20604_, _20603_, _11317_);
  and _71713_ (_20605_, _20604_, _11311_);
  or _71714_ (_20606_, _20605_, _20602_);
  and _71715_ (_20607_, _20606_, _11296_);
  nor _71716_ (_20609_, _06521_, _11296_);
  or _71717_ (_20610_, _20609_, _09842_);
  or _71718_ (_20611_, _20610_, _20607_);
  or _71719_ (_20612_, _20583_, _06132_);
  and _71720_ (_20613_, _20612_, _20611_);
  or _71721_ (_20614_, _20613_, _06116_);
  and _71722_ (_20615_, _09211_, _07849_);
  or _71723_ (_20616_, _20576_, _06117_);
  or _71724_ (_20617_, _20616_, _20615_);
  and _71725_ (_20618_, _20617_, _06114_);
  and _71726_ (_20620_, _20618_, _20614_);
  and _71727_ (_20621_, _14630_, _07849_);
  or _71728_ (_20622_, _20621_, _20576_);
  and _71729_ (_20623_, _20622_, _05787_);
  or _71730_ (_20624_, _20623_, _11136_);
  or _71731_ (_20625_, _20624_, _20620_);
  and _71732_ (_20626_, _14646_, _07849_);
  or _71733_ (_20627_, _20576_, _07127_);
  or _71734_ (_20628_, _20627_, _20626_);
  or _71735_ (_20629_, _20579_, _06111_);
  and _71736_ (_20631_, _20629_, _07125_);
  and _71737_ (_20632_, _20631_, _20628_);
  and _71738_ (_20633_, _20632_, _20625_);
  and _71739_ (_20634_, _10282_, _07849_);
  or _71740_ (_20635_, _20634_, _20576_);
  and _71741_ (_20636_, _20635_, _06402_);
  or _71742_ (_20637_, _20636_, _20633_);
  and _71743_ (_20638_, _20637_, _07132_);
  or _71744_ (_20639_, _20638_, _20581_);
  and _71745_ (_20640_, _20639_, _07130_);
  and _71746_ (_20642_, _20591_, _06411_);
  and _71747_ (_20643_, _20642_, _20577_);
  or _71748_ (_20644_, _20643_, _06303_);
  or _71749_ (_20645_, _20644_, _20640_);
  and _71750_ (_20646_, _14643_, _07849_);
  or _71751_ (_20647_, _20576_, _08819_);
  or _71752_ (_20648_, _20647_, _20646_);
  and _71753_ (_20649_, _20648_, _08824_);
  and _71754_ (_20650_, _20649_, _20645_);
  nor _71755_ (_20651_, _10281_, _11371_);
  or _71756_ (_20653_, _20651_, _20576_);
  and _71757_ (_20654_, _20653_, _06396_);
  or _71758_ (_20655_, _20654_, _20650_);
  and _71759_ (_20656_, _20655_, _06829_);
  and _71760_ (_20657_, _20587_, _06433_);
  or _71761_ (_20658_, _20657_, _06440_);
  or _71762_ (_20659_, _20658_, _20656_);
  and _71763_ (_20660_, _14710_, _07849_);
  or _71764_ (_20661_, _20576_, _06444_);
  or _71765_ (_20662_, _20661_, _20660_);
  and _71766_ (_20664_, _20662_, _01317_);
  and _71767_ (_20665_, _20664_, _20659_);
  or _71768_ (_20666_, _20665_, _20574_);
  and _71769_ (_43630_, _20666_, _43100_);
  and _71770_ (_20667_, _11371_, \oc8051_golden_model_1.DPL [3]);
  or _71771_ (_20668_, _20667_, _08140_);
  and _71772_ (_20669_, _07849_, _08712_);
  or _71773_ (_20670_, _20669_, _20667_);
  and _71774_ (_20671_, _20670_, _06306_);
  and _71775_ (_20672_, _20671_, _20668_);
  and _71776_ (_20674_, _14738_, _07849_);
  or _71777_ (_20675_, _20674_, _20667_);
  or _71778_ (_20676_, _20675_, _06161_);
  and _71779_ (_20677_, _07849_, \oc8051_golden_model_1.ACC [3]);
  or _71780_ (_20678_, _20677_, _20667_);
  and _71781_ (_20679_, _20678_, _07056_);
  and _71782_ (_20680_, _07057_, \oc8051_golden_model_1.DPL [3]);
  or _71783_ (_20681_, _20680_, _06160_);
  or _71784_ (_20682_, _20681_, _20679_);
  and _71785_ (_20683_, _20682_, _07075_);
  and _71786_ (_20685_, _20683_, _20676_);
  and _71787_ (_20686_, _07849_, _07544_);
  or _71788_ (_20687_, _20686_, _20667_);
  and _71789_ (_20688_, _20687_, _06217_);
  or _71790_ (_20689_, _20688_, _06220_);
  or _71791_ (_20690_, _20689_, _20685_);
  or _71792_ (_20691_, _20678_, _06229_);
  and _71793_ (_20692_, _20691_, _11312_);
  and _71794_ (_20693_, _20692_, _20690_);
  nor _71795_ (_20694_, _11317_, \oc8051_golden_model_1.DPL [3]);
  nor _71796_ (_20696_, _20694_, _11318_);
  and _71797_ (_20697_, _20696_, _11311_);
  or _71798_ (_20698_, _20697_, _20693_);
  and _71799_ (_20699_, _20698_, _11296_);
  nor _71800_ (_20700_, _06389_, _11296_);
  or _71801_ (_20701_, _20700_, _09842_);
  or _71802_ (_20702_, _20701_, _20699_);
  or _71803_ (_20703_, _20687_, _06132_);
  and _71804_ (_20704_, _20703_, _20702_);
  or _71805_ (_20705_, _20704_, _06116_);
  and _71806_ (_20707_, _09210_, _07849_);
  or _71807_ (_20708_, _20667_, _06117_);
  or _71808_ (_20709_, _20708_, _20707_);
  and _71809_ (_20710_, _20709_, _06114_);
  and _71810_ (_20711_, _20710_, _20705_);
  and _71811_ (_20712_, _14825_, _07849_);
  or _71812_ (_20713_, _20712_, _20667_);
  and _71813_ (_20714_, _20713_, _05787_);
  or _71814_ (_20715_, _20714_, _11136_);
  or _71815_ (_20716_, _20715_, _20711_);
  and _71816_ (_20718_, _14727_, _07849_);
  or _71817_ (_20719_, _20667_, _07127_);
  or _71818_ (_20720_, _20719_, _20718_);
  or _71819_ (_20721_, _20670_, _06111_);
  and _71820_ (_20722_, _20721_, _07125_);
  and _71821_ (_20723_, _20722_, _20720_);
  and _71822_ (_20724_, _20723_, _20716_);
  and _71823_ (_20725_, _12318_, _07849_);
  or _71824_ (_20726_, _20725_, _20667_);
  and _71825_ (_20727_, _20726_, _06402_);
  or _71826_ (_20729_, _20727_, _20724_);
  and _71827_ (_20730_, _20729_, _07132_);
  or _71828_ (_20731_, _20730_, _20672_);
  and _71829_ (_20732_, _20731_, _07130_);
  and _71830_ (_20733_, _20678_, _06411_);
  and _71831_ (_20734_, _20733_, _20668_);
  or _71832_ (_20735_, _20734_, _06303_);
  or _71833_ (_20736_, _20735_, _20732_);
  and _71834_ (_20737_, _14724_, _07849_);
  or _71835_ (_20738_, _20667_, _08819_);
  or _71836_ (_20740_, _20738_, _20737_);
  and _71837_ (_20741_, _20740_, _08824_);
  and _71838_ (_20742_, _20741_, _20736_);
  nor _71839_ (_20743_, _10273_, _11371_);
  or _71840_ (_20744_, _20743_, _20667_);
  and _71841_ (_20745_, _20744_, _06396_);
  or _71842_ (_20746_, _20745_, _06433_);
  or _71843_ (_20747_, _20746_, _20742_);
  or _71844_ (_20748_, _20675_, _06829_);
  and _71845_ (_20749_, _20748_, _06444_);
  and _71846_ (_20751_, _20749_, _20747_);
  and _71847_ (_20752_, _14897_, _07849_);
  or _71848_ (_20753_, _20752_, _20667_);
  and _71849_ (_20754_, _20753_, _06440_);
  or _71850_ (_20755_, _20754_, _01321_);
  or _71851_ (_20756_, _20755_, _20751_);
  or _71852_ (_20757_, _01317_, \oc8051_golden_model_1.DPL [3]);
  and _71853_ (_20758_, _20757_, _43100_);
  and _71854_ (_43631_, _20758_, _20756_);
  and _71855_ (_20759_, _11371_, \oc8051_golden_model_1.DPL [4]);
  and _71856_ (_20760_, _08336_, _07849_);
  or _71857_ (_20761_, _20760_, _20759_);
  or _71858_ (_20762_, _20761_, _06132_);
  and _71859_ (_20763_, _14928_, _07849_);
  or _71860_ (_20764_, _20763_, _20759_);
  or _71861_ (_20765_, _20764_, _06161_);
  and _71862_ (_20766_, _07849_, \oc8051_golden_model_1.ACC [4]);
  or _71863_ (_20767_, _20766_, _20759_);
  and _71864_ (_20768_, _20767_, _07056_);
  and _71865_ (_20769_, _07057_, \oc8051_golden_model_1.DPL [4]);
  or _71866_ (_20771_, _20769_, _06160_);
  or _71867_ (_20772_, _20771_, _20768_);
  and _71868_ (_20773_, _20772_, _07075_);
  and _71869_ (_20774_, _20773_, _20765_);
  and _71870_ (_20775_, _20761_, _06217_);
  or _71871_ (_20776_, _20775_, _06220_);
  or _71872_ (_20777_, _20776_, _20774_);
  or _71873_ (_20778_, _20767_, _06229_);
  and _71874_ (_20779_, _20778_, _11312_);
  and _71875_ (_20780_, _20779_, _20777_);
  nor _71876_ (_20783_, _11318_, \oc8051_golden_model_1.DPL [4]);
  nor _71877_ (_20784_, _20783_, _11319_);
  and _71878_ (_20785_, _20784_, _11311_);
  or _71879_ (_20786_, _20785_, _20780_);
  and _71880_ (_20787_, _20786_, _11296_);
  nor _71881_ (_20788_, _08670_, _11296_);
  or _71882_ (_20789_, _20788_, _09842_);
  or _71883_ (_20790_, _20789_, _20787_);
  and _71884_ (_20791_, _20790_, _20762_);
  or _71885_ (_20792_, _20791_, _06116_);
  and _71886_ (_20794_, _09209_, _07849_);
  or _71887_ (_20795_, _20759_, _06117_);
  or _71888_ (_20796_, _20795_, _20794_);
  and _71889_ (_20797_, _20796_, _06114_);
  and _71890_ (_20798_, _20797_, _20792_);
  and _71891_ (_20799_, _15013_, _07849_);
  or _71892_ (_20800_, _20799_, _20759_);
  and _71893_ (_20801_, _20800_, _05787_);
  or _71894_ (_20802_, _20801_, _20798_);
  or _71895_ (_20803_, _20802_, _11136_);
  and _71896_ (_20804_, _15029_, _07849_);
  or _71897_ (_20805_, _20759_, _07127_);
  or _71898_ (_20806_, _20805_, _20804_);
  and _71899_ (_20807_, _08715_, _07849_);
  or _71900_ (_20808_, _20807_, _20759_);
  or _71901_ (_20809_, _20808_, _06111_);
  and _71902_ (_20810_, _20809_, _07125_);
  and _71903_ (_20811_, _20810_, _20806_);
  and _71904_ (_20812_, _20811_, _20803_);
  and _71905_ (_20813_, _10289_, _07849_);
  or _71906_ (_20815_, _20813_, _20759_);
  and _71907_ (_20816_, _20815_, _06402_);
  or _71908_ (_20817_, _20816_, _20812_);
  and _71909_ (_20818_, _20817_, _07132_);
  or _71910_ (_20819_, _20759_, _08339_);
  and _71911_ (_20820_, _20808_, _06306_);
  and _71912_ (_20821_, _20820_, _20819_);
  or _71913_ (_20822_, _20821_, _20818_);
  and _71914_ (_20823_, _20822_, _07130_);
  and _71915_ (_20824_, _20767_, _06411_);
  and _71916_ (_20827_, _20824_, _20819_);
  or _71917_ (_20828_, _20827_, _06303_);
  or _71918_ (_20829_, _20828_, _20823_);
  and _71919_ (_20830_, _15026_, _07849_);
  or _71920_ (_20831_, _20759_, _08819_);
  or _71921_ (_20832_, _20831_, _20830_);
  and _71922_ (_20833_, _20832_, _08824_);
  and _71923_ (_20834_, _20833_, _20829_);
  nor _71924_ (_20835_, _10288_, _11371_);
  or _71925_ (_20836_, _20835_, _20759_);
  and _71926_ (_20837_, _20836_, _06396_);
  or _71927_ (_20838_, _20837_, _06433_);
  or _71928_ (_20839_, _20838_, _20834_);
  or _71929_ (_20840_, _20764_, _06829_);
  and _71930_ (_20841_, _20840_, _06444_);
  and _71931_ (_20842_, _20841_, _20839_);
  and _71932_ (_20843_, _15087_, _07849_);
  or _71933_ (_20844_, _20843_, _20759_);
  and _71934_ (_20845_, _20844_, _06440_);
  or _71935_ (_20846_, _20845_, _01321_);
  or _71936_ (_20848_, _20846_, _20842_);
  or _71937_ (_20849_, _01317_, \oc8051_golden_model_1.DPL [4]);
  and _71938_ (_20850_, _20849_, _43100_);
  and _71939_ (_43632_, _20850_, _20848_);
  and _71940_ (_20851_, _11371_, \oc8051_golden_model_1.DPL [5]);
  and _71941_ (_20852_, _08101_, _07849_);
  or _71942_ (_20853_, _20852_, _20851_);
  or _71943_ (_20854_, _20853_, _06132_);
  and _71944_ (_20855_, _15119_, _07849_);
  or _71945_ (_20856_, _20855_, _20851_);
  or _71946_ (_20859_, _20856_, _06161_);
  and _71947_ (_20860_, _07849_, \oc8051_golden_model_1.ACC [5]);
  or _71948_ (_20861_, _20860_, _20851_);
  and _71949_ (_20862_, _20861_, _07056_);
  and _71950_ (_20863_, _07057_, \oc8051_golden_model_1.DPL [5]);
  or _71951_ (_20864_, _20863_, _06160_);
  or _71952_ (_20865_, _20864_, _20862_);
  and _71953_ (_20866_, _20865_, _07075_);
  and _71954_ (_20867_, _20866_, _20859_);
  and _71955_ (_20868_, _20853_, _06217_);
  or _71956_ (_20870_, _20868_, _06220_);
  or _71957_ (_20871_, _20870_, _20867_);
  or _71958_ (_20872_, _20861_, _06229_);
  and _71959_ (_20873_, _20872_, _11312_);
  and _71960_ (_20874_, _20873_, _20871_);
  nor _71961_ (_20875_, _11319_, \oc8051_golden_model_1.DPL [5]);
  nor _71962_ (_20876_, _20875_, _11320_);
  and _71963_ (_20877_, _20876_, _11311_);
  or _71964_ (_20878_, _20877_, _20874_);
  and _71965_ (_20879_, _20878_, _11296_);
  nor _71966_ (_20881_, _08701_, _11296_);
  or _71967_ (_20882_, _20881_, _09842_);
  or _71968_ (_20883_, _20882_, _20879_);
  and _71969_ (_20884_, _20883_, _20854_);
  or _71970_ (_20885_, _20884_, _06116_);
  and _71971_ (_20886_, _09208_, _07849_);
  or _71972_ (_20887_, _20851_, _06117_);
  or _71973_ (_20888_, _20887_, _20886_);
  and _71974_ (_20889_, _20888_, _06114_);
  and _71975_ (_20890_, _20889_, _20885_);
  and _71976_ (_20892_, _15203_, _07849_);
  or _71977_ (_20893_, _20892_, _20851_);
  and _71978_ (_20894_, _20893_, _05787_);
  or _71979_ (_20895_, _20894_, _20890_);
  or _71980_ (_20896_, _20895_, _11136_);
  and _71981_ (_20897_, _15219_, _07849_);
  or _71982_ (_20898_, _20851_, _07127_);
  or _71983_ (_20899_, _20898_, _20897_);
  and _71984_ (_20900_, _08736_, _07849_);
  or _71985_ (_20901_, _20900_, _20851_);
  or _71986_ (_20902_, _20901_, _06111_);
  and _71987_ (_20903_, _20902_, _07125_);
  and _71988_ (_20904_, _20903_, _20899_);
  and _71989_ (_20905_, _20904_, _20896_);
  and _71990_ (_20906_, _12325_, _07849_);
  or _71991_ (_20907_, _20906_, _20851_);
  and _71992_ (_20908_, _20907_, _06402_);
  or _71993_ (_20909_, _20908_, _20905_);
  and _71994_ (_20910_, _20909_, _07132_);
  or _71995_ (_20911_, _20851_, _08104_);
  and _71996_ (_20914_, _20901_, _06306_);
  and _71997_ (_20915_, _20914_, _20911_);
  or _71998_ (_20916_, _20915_, _20910_);
  and _71999_ (_20917_, _20916_, _07130_);
  and _72000_ (_20918_, _20861_, _06411_);
  and _72001_ (_20919_, _20918_, _20911_);
  or _72002_ (_20920_, _20919_, _06303_);
  or _72003_ (_20921_, _20920_, _20917_);
  and _72004_ (_20922_, _15216_, _07849_);
  or _72005_ (_20923_, _20851_, _08819_);
  or _72006_ (_20925_, _20923_, _20922_);
  and _72007_ (_20926_, _20925_, _08824_);
  and _72008_ (_20927_, _20926_, _20921_);
  nor _72009_ (_20928_, _10269_, _11371_);
  or _72010_ (_20929_, _20928_, _20851_);
  and _72011_ (_20930_, _20929_, _06396_);
  or _72012_ (_20931_, _20930_, _06433_);
  or _72013_ (_20932_, _20931_, _20927_);
  or _72014_ (_20933_, _20856_, _06829_);
  and _72015_ (_20934_, _20933_, _06444_);
  and _72016_ (_20936_, _20934_, _20932_);
  and _72017_ (_20937_, _15275_, _07849_);
  or _72018_ (_20938_, _20937_, _20851_);
  and _72019_ (_20939_, _20938_, _06440_);
  or _72020_ (_20940_, _20939_, _01321_);
  or _72021_ (_20941_, _20940_, _20936_);
  or _72022_ (_20942_, _01317_, \oc8051_golden_model_1.DPL [5]);
  and _72023_ (_20943_, _20942_, _43100_);
  and _72024_ (_43633_, _20943_, _20941_);
  and _72025_ (_20944_, _11371_, \oc8051_golden_model_1.DPL [6]);
  and _72026_ (_20946_, _08012_, _07849_);
  or _72027_ (_20947_, _20946_, _20944_);
  or _72028_ (_20948_, _20947_, _06132_);
  and _72029_ (_20949_, _15300_, _07849_);
  or _72030_ (_20950_, _20949_, _20944_);
  or _72031_ (_20951_, _20950_, _06161_);
  and _72032_ (_20952_, _07849_, \oc8051_golden_model_1.ACC [6]);
  or _72033_ (_20953_, _20952_, _20944_);
  and _72034_ (_20954_, _20953_, _07056_);
  and _72035_ (_20955_, _07057_, \oc8051_golden_model_1.DPL [6]);
  or _72036_ (_20957_, _20955_, _06160_);
  or _72037_ (_20958_, _20957_, _20954_);
  and _72038_ (_20959_, _20958_, _07075_);
  and _72039_ (_20960_, _20959_, _20951_);
  and _72040_ (_20961_, _20947_, _06217_);
  or _72041_ (_20962_, _20961_, _06220_);
  or _72042_ (_20963_, _20962_, _20960_);
  or _72043_ (_20964_, _20953_, _06229_);
  and _72044_ (_20965_, _20964_, _11312_);
  and _72045_ (_20966_, _20965_, _20963_);
  nor _72046_ (_20968_, _11320_, \oc8051_golden_model_1.DPL [6]);
  nor _72047_ (_20969_, _20968_, _11321_);
  and _72048_ (_20970_, _20969_, _11311_);
  or _72049_ (_20971_, _20970_, _20966_);
  and _72050_ (_20972_, _20971_, _11296_);
  nor _72051_ (_20973_, _08638_, _11296_);
  or _72052_ (_20974_, _20973_, _09842_);
  or _72053_ (_20975_, _20974_, _20972_);
  and _72054_ (_20976_, _20975_, _20948_);
  or _72055_ (_20977_, _20976_, _06116_);
  and _72056_ (_20979_, _09207_, _07849_);
  or _72057_ (_20980_, _20944_, _06117_);
  or _72058_ (_20981_, _20980_, _20979_);
  and _72059_ (_20982_, _20981_, _06114_);
  and _72060_ (_20983_, _20982_, _20977_);
  and _72061_ (_20984_, _15395_, _07849_);
  or _72062_ (_20985_, _20984_, _20944_);
  and _72063_ (_20986_, _20985_, _05787_);
  or _72064_ (_20987_, _20986_, _20983_);
  or _72065_ (_20988_, _20987_, _11136_);
  and _72066_ (_20990_, _15413_, _07849_);
  or _72067_ (_20991_, _20944_, _07127_);
  or _72068_ (_20992_, _20991_, _20990_);
  and _72069_ (_20993_, _15402_, _07849_);
  or _72070_ (_20994_, _20993_, _20944_);
  or _72071_ (_20995_, _20994_, _06111_);
  and _72072_ (_20996_, _20995_, _07125_);
  and _72073_ (_20997_, _20996_, _20992_);
  and _72074_ (_20998_, _20997_, _20988_);
  and _72075_ (_20999_, _10295_, _07849_);
  or _72076_ (_21001_, _20999_, _20944_);
  and _72077_ (_21002_, _21001_, _06402_);
  or _72078_ (_21003_, _21002_, _20998_);
  and _72079_ (_21004_, _21003_, _07132_);
  or _72080_ (_21005_, _20944_, _08015_);
  and _72081_ (_21006_, _20994_, _06306_);
  and _72082_ (_21007_, _21006_, _21005_);
  or _72083_ (_21008_, _21007_, _21004_);
  and _72084_ (_21009_, _21008_, _07130_);
  and _72085_ (_21010_, _20953_, _06411_);
  and _72086_ (_21012_, _21010_, _21005_);
  or _72087_ (_21013_, _21012_, _06303_);
  or _72088_ (_21014_, _21013_, _21009_);
  and _72089_ (_21015_, _15410_, _07849_);
  or _72090_ (_21016_, _20944_, _08819_);
  or _72091_ (_21017_, _21016_, _21015_);
  and _72092_ (_21018_, _21017_, _08824_);
  and _72093_ (_21019_, _21018_, _21014_);
  nor _72094_ (_21020_, _10294_, _11371_);
  or _72095_ (_21021_, _21020_, _20944_);
  and _72096_ (_21023_, _21021_, _06396_);
  or _72097_ (_21024_, _21023_, _06433_);
  or _72098_ (_21025_, _21024_, _21019_);
  or _72099_ (_21026_, _20950_, _06829_);
  and _72100_ (_21027_, _21026_, _06444_);
  and _72101_ (_21028_, _21027_, _21025_);
  and _72102_ (_21029_, _15478_, _07849_);
  or _72103_ (_21030_, _21029_, _20944_);
  and _72104_ (_21031_, _21030_, _06440_);
  or _72105_ (_21032_, _21031_, _01321_);
  or _72106_ (_21033_, _21032_, _21028_);
  or _72107_ (_21034_, _01317_, \oc8051_golden_model_1.DPL [6]);
  and _72108_ (_21035_, _21034_, _43100_);
  and _72109_ (_43634_, _21035_, _21033_);
  nor _72110_ (_21036_, _01317_, _12434_);
  nor _72111_ (_21037_, _11390_, _12434_);
  and _72112_ (_21038_, _11390_, \oc8051_golden_model_1.ACC [0]);
  and _72113_ (_21039_, _21038_, _08211_);
  or _72114_ (_21040_, _21039_, _21037_);
  or _72115_ (_21041_, _21040_, _07130_);
  nor _72116_ (_21044_, _08211_, _11468_);
  or _72117_ (_21045_, _21044_, _21037_);
  or _72118_ (_21046_, _21045_, _06161_);
  or _72119_ (_21047_, _21038_, _21037_);
  and _72120_ (_21048_, _21047_, _07056_);
  nor _72121_ (_21049_, _07056_, _12434_);
  or _72122_ (_21050_, _21049_, _06160_);
  or _72123_ (_21051_, _21050_, _21048_);
  and _72124_ (_21052_, _21051_, _07075_);
  and _72125_ (_21053_, _21052_, _21046_);
  and _72126_ (_21055_, _07852_, _07049_);
  or _72127_ (_21056_, _21055_, _21037_);
  and _72128_ (_21057_, _21056_, _06217_);
  or _72129_ (_21058_, _21057_, _06220_);
  or _72130_ (_21059_, _21058_, _21053_);
  or _72131_ (_21060_, _21047_, _06229_);
  and _72132_ (_21061_, _21060_, _11312_);
  and _72133_ (_21062_, _21061_, _21059_);
  nor _72134_ (_21063_, _11323_, \oc8051_golden_model_1.DPH [0]);
  nor _72135_ (_21064_, _21063_, _11412_);
  and _72136_ (_21066_, _21064_, _11311_);
  or _72137_ (_21067_, _21066_, _21062_);
  and _72138_ (_21068_, _21067_, _11296_);
  nor _72139_ (_21069_, _11296_, _06107_);
  or _72140_ (_21070_, _21069_, _09842_);
  or _72141_ (_21071_, _21070_, _21068_);
  or _72142_ (_21072_, _21056_, _06132_);
  and _72143_ (_21073_, _21072_, _21071_);
  or _72144_ (_21074_, _21073_, _06116_);
  and _72145_ (_21075_, _09160_, _11390_);
  or _72146_ (_21077_, _21037_, _06117_);
  or _72147_ (_21078_, _21077_, _21075_);
  and _72148_ (_21079_, _21078_, _21074_);
  or _72149_ (_21080_, _21079_, _05787_);
  and _72150_ (_21081_, _14260_, _11390_);
  or _72151_ (_21082_, _21081_, _21037_);
  or _72152_ (_21083_, _21082_, _06114_);
  and _72153_ (_21084_, _21083_, _06111_);
  and _72154_ (_21085_, _21084_, _21080_);
  and _72155_ (_21086_, _11390_, _08708_);
  or _72156_ (_21088_, _21086_, _21037_);
  and _72157_ (_21089_, _21088_, _06110_);
  or _72158_ (_21090_, _21089_, _06297_);
  or _72159_ (_21091_, _21090_, _21085_);
  and _72160_ (_21092_, _14275_, _07852_);
  or _72161_ (_21093_, _21037_, _07127_);
  or _72162_ (_21094_, _21093_, _21092_);
  and _72163_ (_21095_, _21094_, _07125_);
  and _72164_ (_21096_, _21095_, _21091_);
  nor _72165_ (_21097_, _12321_, _11468_);
  or _72166_ (_21099_, _21097_, _21037_);
  nor _72167_ (_21100_, _21039_, _07125_);
  and _72168_ (_21101_, _21100_, _21099_);
  or _72169_ (_21102_, _21101_, _21096_);
  and _72170_ (_21103_, _21102_, _07132_);
  nand _72171_ (_21104_, _21088_, _06306_);
  nor _72172_ (_21105_, _21104_, _21044_);
  or _72173_ (_21106_, _21105_, _06411_);
  or _72174_ (_21107_, _21106_, _21103_);
  and _72175_ (_21108_, _21107_, _21041_);
  or _72176_ (_21110_, _21108_, _06303_);
  and _72177_ (_21111_, _14167_, _07852_);
  or _72178_ (_21112_, _21037_, _08819_);
  or _72179_ (_21113_, _21112_, _21111_);
  and _72180_ (_21114_, _21113_, _08824_);
  and _72181_ (_21115_, _21114_, _21110_);
  and _72182_ (_21116_, _21099_, _06396_);
  or _72183_ (_21117_, _21116_, _19287_);
  or _72184_ (_21118_, _21117_, _21115_);
  or _72185_ (_21119_, _21045_, _06630_);
  and _72186_ (_21121_, _21119_, _01317_);
  and _72187_ (_21122_, _21121_, _21118_);
  or _72188_ (_21123_, _21122_, _21036_);
  and _72189_ (_43636_, _21123_, _43100_);
  not _72190_ (_21124_, \oc8051_golden_model_1.DPH [1]);
  nor _72191_ (_21125_, _11390_, _21124_);
  nor _72192_ (_21126_, _10277_, _11468_);
  or _72193_ (_21127_, _21126_, _21125_);
  or _72194_ (_21128_, _21127_, _08824_);
  or _72195_ (_21129_, _14442_, _11468_);
  or _72196_ (_21131_, _11390_, \oc8051_golden_model_1.DPH [1]);
  and _72197_ (_21132_, _21131_, _05787_);
  and _72198_ (_21133_, _21132_, _21129_);
  and _72199_ (_21134_, _09115_, _11390_);
  or _72200_ (_21135_, _21134_, _21125_);
  and _72201_ (_21136_, _21135_, _06116_);
  and _72202_ (_21137_, _14363_, _07852_);
  not _72203_ (_21138_, _21137_);
  and _72204_ (_21139_, _21138_, _21131_);
  or _72205_ (_21140_, _21139_, _06161_);
  and _72206_ (_21142_, _11390_, \oc8051_golden_model_1.ACC [1]);
  or _72207_ (_21143_, _21142_, _21125_);
  and _72208_ (_21144_, _21143_, _07056_);
  nor _72209_ (_21145_, _07056_, _21124_);
  or _72210_ (_21146_, _21145_, _06160_);
  or _72211_ (_21147_, _21146_, _21144_);
  and _72212_ (_21148_, _21147_, _07075_);
  and _72213_ (_21149_, _21148_, _21140_);
  and _72214_ (_21150_, _07852_, _07306_);
  or _72215_ (_21151_, _21150_, _21125_);
  and _72216_ (_21153_, _21151_, _06217_);
  or _72217_ (_21154_, _21153_, _06220_);
  or _72218_ (_21155_, _21154_, _21149_);
  or _72219_ (_21156_, _21143_, _06229_);
  and _72220_ (_21157_, _21156_, _11312_);
  and _72221_ (_21158_, _21157_, _21155_);
  nor _72222_ (_21159_, _11412_, \oc8051_golden_model_1.DPH [1]);
  nor _72223_ (_21160_, _21159_, _11413_);
  and _72224_ (_21161_, _21160_, _11311_);
  or _72225_ (_21162_, _21161_, _21158_);
  and _72226_ (_21164_, _21162_, _11296_);
  nor _72227_ (_21165_, _06912_, _11296_);
  or _72228_ (_21166_, _21165_, _09842_);
  or _72229_ (_21167_, _21166_, _21164_);
  or _72230_ (_21168_, _21151_, _06132_);
  and _72231_ (_21169_, _21168_, _06117_);
  and _72232_ (_21170_, _21169_, _21167_);
  or _72233_ (_21171_, _21170_, _21136_);
  and _72234_ (_21172_, _21171_, _06114_);
  or _72235_ (_21173_, _21172_, _21133_);
  and _72236_ (_21175_, _21173_, _06298_);
  or _72237_ (_21176_, _14346_, _11468_);
  and _72238_ (_21177_, _21176_, _06297_);
  nand _72239_ (_21178_, _07852_, _06945_);
  and _72240_ (_21179_, _21178_, _06110_);
  or _72241_ (_21180_, _21179_, _21177_);
  and _72242_ (_21181_, _21180_, _21131_);
  or _72243_ (_21182_, _21181_, _06402_);
  or _72244_ (_21183_, _21182_, _21175_);
  nand _72245_ (_21184_, _10275_, _07852_);
  and _72246_ (_21186_, _21184_, _21127_);
  or _72247_ (_21187_, _21186_, _07125_);
  and _72248_ (_21188_, _21187_, _07132_);
  and _72249_ (_21189_, _21188_, _21183_);
  or _72250_ (_21190_, _14344_, _11468_);
  and _72251_ (_21191_, _21131_, _06306_);
  and _72252_ (_21192_, _21191_, _21190_);
  or _72253_ (_21193_, _21192_, _06411_);
  or _72254_ (_21194_, _21193_, _21189_);
  nor _72255_ (_21195_, _21125_, _07130_);
  nand _72256_ (_21197_, _21195_, _21184_);
  and _72257_ (_21198_, _21197_, _08819_);
  and _72258_ (_21199_, _21198_, _21194_);
  or _72259_ (_21200_, _21178_, _08176_);
  and _72260_ (_21201_, _21131_, _06303_);
  and _72261_ (_21202_, _21201_, _21200_);
  or _72262_ (_21203_, _21202_, _06396_);
  or _72263_ (_21204_, _21203_, _21199_);
  and _72264_ (_21205_, _21204_, _21128_);
  or _72265_ (_21206_, _21205_, _06433_);
  or _72266_ (_21207_, _21139_, _06829_);
  and _72267_ (_21208_, _21207_, _06444_);
  and _72268_ (_21209_, _21208_, _21206_);
  or _72269_ (_21210_, _21137_, _21125_);
  and _72270_ (_21211_, _21210_, _06440_);
  or _72271_ (_21212_, _21211_, _01321_);
  or _72272_ (_21213_, _21212_, _21209_);
  or _72273_ (_21214_, _01317_, \oc8051_golden_model_1.DPH [1]);
  and _72274_ (_21215_, _21214_, _43100_);
  and _72275_ (_43637_, _21215_, _21213_);
  and _72276_ (_21218_, _01321_, \oc8051_golden_model_1.DPH [2]);
  and _72277_ (_21219_, _11468_, \oc8051_golden_model_1.DPH [2]);
  and _72278_ (_21220_, _07852_, _07708_);
  or _72279_ (_21221_, _21220_, _21219_);
  or _72280_ (_21222_, _21221_, _06132_);
  and _72281_ (_21223_, _14542_, _07852_);
  or _72282_ (_21224_, _21223_, _21219_);
  or _72283_ (_21225_, _21224_, _06161_);
  and _72284_ (_21226_, _11390_, \oc8051_golden_model_1.ACC [2]);
  or _72285_ (_21227_, _21226_, _21219_);
  and _72286_ (_21229_, _21227_, _07056_);
  and _72287_ (_21230_, _07057_, \oc8051_golden_model_1.DPH [2]);
  or _72288_ (_21231_, _21230_, _06160_);
  or _72289_ (_21232_, _21231_, _21229_);
  and _72290_ (_21233_, _21232_, _07075_);
  and _72291_ (_21234_, _21233_, _21225_);
  and _72292_ (_21235_, _21221_, _06217_);
  or _72293_ (_21236_, _21235_, _06220_);
  or _72294_ (_21237_, _21236_, _21234_);
  or _72295_ (_21238_, _21227_, _06229_);
  and _72296_ (_21240_, _21238_, _11312_);
  and _72297_ (_21241_, _21240_, _21237_);
  or _72298_ (_21242_, _11413_, \oc8051_golden_model_1.DPH [2]);
  nor _72299_ (_21243_, _11414_, _11312_);
  and _72300_ (_21244_, _21243_, _21242_);
  or _72301_ (_21245_, _21244_, _21241_);
  and _72302_ (_21246_, _21245_, _11296_);
  nor _72303_ (_21247_, _06625_, _11296_);
  or _72304_ (_21248_, _21247_, _09842_);
  or _72305_ (_21249_, _21248_, _21246_);
  and _72306_ (_21251_, _21249_, _21222_);
  or _72307_ (_21252_, _21251_, _06116_);
  or _72308_ (_21253_, _21219_, _06117_);
  and _72309_ (_21254_, _09211_, _11390_);
  or _72310_ (_21255_, _21254_, _21253_);
  and _72311_ (_21256_, _21255_, _06114_);
  and _72312_ (_21257_, _21256_, _21252_);
  and _72313_ (_21258_, _14630_, _11390_);
  or _72314_ (_21259_, _21258_, _21219_);
  and _72315_ (_21260_, _21259_, _05787_);
  or _72316_ (_21262_, _21260_, _21257_);
  or _72317_ (_21263_, _21262_, _11136_);
  and _72318_ (_21264_, _14646_, _07852_);
  or _72319_ (_21265_, _21219_, _07127_);
  or _72320_ (_21266_, _21265_, _21264_);
  and _72321_ (_21267_, _11390_, _08768_);
  or _72322_ (_21268_, _21267_, _21219_);
  or _72323_ (_21269_, _21268_, _06111_);
  and _72324_ (_21270_, _21269_, _07125_);
  and _72325_ (_21271_, _21270_, _21266_);
  and _72326_ (_21273_, _21271_, _21263_);
  and _72327_ (_21274_, _10282_, _11390_);
  or _72328_ (_21275_, _21274_, _21219_);
  and _72329_ (_21276_, _21275_, _06402_);
  or _72330_ (_21277_, _21276_, _21273_);
  and _72331_ (_21278_, _21277_, _07132_);
  or _72332_ (_21279_, _21219_, _08248_);
  and _72333_ (_21280_, _21268_, _06306_);
  and _72334_ (_21281_, _21280_, _21279_);
  or _72335_ (_21282_, _21281_, _21278_);
  and _72336_ (_21284_, _21282_, _07130_);
  and _72337_ (_21285_, _21227_, _06411_);
  and _72338_ (_21286_, _21285_, _21279_);
  or _72339_ (_21287_, _21286_, _06303_);
  or _72340_ (_21288_, _21287_, _21284_);
  and _72341_ (_21289_, _14643_, _07852_);
  or _72342_ (_21290_, _21219_, _08819_);
  or _72343_ (_21291_, _21290_, _21289_);
  and _72344_ (_21292_, _21291_, _08824_);
  and _72345_ (_21293_, _21292_, _21288_);
  nor _72346_ (_21295_, _10281_, _11468_);
  or _72347_ (_21296_, _21295_, _21219_);
  and _72348_ (_21297_, _21296_, _06396_);
  or _72349_ (_21298_, _21297_, _21293_);
  and _72350_ (_21299_, _21298_, _06829_);
  and _72351_ (_21300_, _21224_, _06433_);
  or _72352_ (_21301_, _21300_, _06440_);
  or _72353_ (_21302_, _21301_, _21299_);
  and _72354_ (_21303_, _14710_, _07852_);
  or _72355_ (_21304_, _21219_, _06444_);
  or _72356_ (_21306_, _21304_, _21303_);
  and _72357_ (_21307_, _21306_, _01317_);
  and _72358_ (_21308_, _21307_, _21302_);
  or _72359_ (_21309_, _21308_, _21218_);
  and _72360_ (_43638_, _21309_, _43100_);
  and _72361_ (_21310_, _11468_, \oc8051_golden_model_1.DPH [3]);
  or _72362_ (_21311_, _21310_, _08140_);
  and _72363_ (_21312_, _11390_, _08712_);
  or _72364_ (_21313_, _21312_, _21310_);
  and _72365_ (_21314_, _21313_, _06306_);
  and _72366_ (_21316_, _21314_, _21311_);
  and _72367_ (_21317_, _14738_, _07852_);
  or _72368_ (_21318_, _21317_, _21310_);
  or _72369_ (_21319_, _21318_, _06161_);
  and _72370_ (_21320_, _11390_, \oc8051_golden_model_1.ACC [3]);
  or _72371_ (_21321_, _21320_, _21310_);
  and _72372_ (_21322_, _21321_, _07056_);
  and _72373_ (_21323_, _07057_, \oc8051_golden_model_1.DPH [3]);
  or _72374_ (_21324_, _21323_, _06160_);
  or _72375_ (_21325_, _21324_, _21322_);
  and _72376_ (_21327_, _21325_, _07075_);
  and _72377_ (_21328_, _21327_, _21319_);
  and _72378_ (_21329_, _07852_, _07544_);
  or _72379_ (_21330_, _21329_, _21310_);
  and _72380_ (_21331_, _21330_, _06217_);
  or _72381_ (_21332_, _21331_, _06220_);
  or _72382_ (_21333_, _21332_, _21328_);
  or _72383_ (_21334_, _21321_, _06229_);
  and _72384_ (_21335_, _21334_, _11312_);
  and _72385_ (_21336_, _21335_, _21333_);
  or _72386_ (_21338_, _11414_, \oc8051_golden_model_1.DPH [3]);
  nor _72387_ (_21339_, _11415_, _11312_);
  and _72388_ (_21340_, _21339_, _21338_);
  or _72389_ (_21341_, _21340_, _21336_);
  and _72390_ (_21342_, _21341_, _11296_);
  nor _72391_ (_21343_, _11296_, _06070_);
  or _72392_ (_21344_, _21343_, _09842_);
  or _72393_ (_21345_, _21344_, _21342_);
  or _72394_ (_21346_, _21330_, _06132_);
  and _72395_ (_21347_, _21346_, _21345_);
  or _72396_ (_21349_, _21347_, _06116_);
  and _72397_ (_21350_, _09210_, _11390_);
  or _72398_ (_21351_, _21310_, _06117_);
  or _72399_ (_21352_, _21351_, _21350_);
  and _72400_ (_21353_, _21352_, _06114_);
  and _72401_ (_21354_, _21353_, _21349_);
  and _72402_ (_21355_, _14825_, _07852_);
  or _72403_ (_21356_, _21355_, _21310_);
  and _72404_ (_21357_, _21356_, _05787_);
  or _72405_ (_21358_, _21357_, _11136_);
  or _72406_ (_21360_, _21358_, _21354_);
  and _72407_ (_21361_, _14727_, _07852_);
  or _72408_ (_21362_, _21310_, _07127_);
  or _72409_ (_21363_, _21362_, _21361_);
  or _72410_ (_21364_, _21313_, _06111_);
  and _72411_ (_21365_, _21364_, _07125_);
  and _72412_ (_21366_, _21365_, _21363_);
  and _72413_ (_21367_, _21366_, _21360_);
  and _72414_ (_21368_, _12318_, _11390_);
  or _72415_ (_21369_, _21368_, _21310_);
  and _72416_ (_21371_, _21369_, _06402_);
  or _72417_ (_21372_, _21371_, _21367_);
  and _72418_ (_21373_, _21372_, _07132_);
  or _72419_ (_21374_, _21373_, _21316_);
  and _72420_ (_21375_, _21374_, _07130_);
  and _72421_ (_21376_, _21321_, _06411_);
  and _72422_ (_21377_, _21376_, _21311_);
  or _72423_ (_21378_, _21377_, _06303_);
  or _72424_ (_21379_, _21378_, _21375_);
  and _72425_ (_21380_, _14724_, _07852_);
  or _72426_ (_21382_, _21310_, _08819_);
  or _72427_ (_21383_, _21382_, _21380_);
  and _72428_ (_21384_, _21383_, _08824_);
  and _72429_ (_21385_, _21384_, _21379_);
  nor _72430_ (_21386_, _10273_, _11468_);
  or _72431_ (_21387_, _21386_, _21310_);
  and _72432_ (_21388_, _21387_, _06396_);
  or _72433_ (_21389_, _21388_, _06433_);
  or _72434_ (_21390_, _21389_, _21385_);
  or _72435_ (_21391_, _21318_, _06829_);
  and _72436_ (_21393_, _21391_, _06444_);
  and _72437_ (_21394_, _21393_, _21390_);
  and _72438_ (_21395_, _14897_, _07852_);
  or _72439_ (_21396_, _21395_, _21310_);
  and _72440_ (_21397_, _21396_, _06440_);
  or _72441_ (_21398_, _21397_, _01321_);
  or _72442_ (_21399_, _21398_, _21394_);
  or _72443_ (_21400_, _01317_, \oc8051_golden_model_1.DPH [3]);
  and _72444_ (_21401_, _21400_, _43100_);
  and _72445_ (_43640_, _21401_, _21399_);
  not _72446_ (_21402_, \oc8051_golden_model_1.DPH [4]);
  nor _72447_ (_21403_, _11390_, _21402_);
  and _72448_ (_21404_, _08336_, _07852_);
  or _72449_ (_21405_, _21404_, _21403_);
  or _72450_ (_21406_, _21405_, _06132_);
  and _72451_ (_21407_, _14928_, _07852_);
  or _72452_ (_21408_, _21407_, _21403_);
  or _72453_ (_21409_, _21408_, _06161_);
  and _72454_ (_21410_, _11390_, \oc8051_golden_model_1.ACC [4]);
  or _72455_ (_21411_, _21410_, _21403_);
  and _72456_ (_21414_, _21411_, _07056_);
  nor _72457_ (_21415_, _07056_, _21402_);
  or _72458_ (_21416_, _21415_, _06160_);
  or _72459_ (_21417_, _21416_, _21414_);
  and _72460_ (_21418_, _21417_, _07075_);
  and _72461_ (_21419_, _21418_, _21409_);
  and _72462_ (_21420_, _21405_, _06217_);
  or _72463_ (_21421_, _21420_, _06220_);
  or _72464_ (_21422_, _21421_, _21419_);
  or _72465_ (_21423_, _21411_, _06229_);
  and _72466_ (_21425_, _21423_, _11312_);
  and _72467_ (_21426_, _21425_, _21422_);
  or _72468_ (_21427_, _11415_, \oc8051_golden_model_1.DPH [4]);
  nor _72469_ (_21428_, _11416_, _11312_);
  and _72470_ (_21429_, _21428_, _21427_);
  or _72471_ (_21430_, _21429_, _21426_);
  and _72472_ (_21431_, _21430_, _11296_);
  nor _72473_ (_21432_, _06876_, _11296_);
  or _72474_ (_21433_, _21432_, _09842_);
  or _72475_ (_21434_, _21433_, _21431_);
  and _72476_ (_21436_, _21434_, _21406_);
  or _72477_ (_21437_, _21436_, _06116_);
  or _72478_ (_21438_, _21403_, _06117_);
  and _72479_ (_21439_, _09209_, _11390_);
  or _72480_ (_21440_, _21439_, _21438_);
  and _72481_ (_21441_, _21440_, _06114_);
  and _72482_ (_21442_, _21441_, _21437_);
  and _72483_ (_21443_, _15013_, _11390_);
  or _72484_ (_21444_, _21443_, _21403_);
  and _72485_ (_21445_, _21444_, _05787_);
  or _72486_ (_21447_, _21445_, _21442_);
  or _72487_ (_21448_, _21447_, _11136_);
  and _72488_ (_21449_, _15029_, _07852_);
  or _72489_ (_21450_, _21403_, _07127_);
  or _72490_ (_21451_, _21450_, _21449_);
  and _72491_ (_21452_, _08715_, _11390_);
  or _72492_ (_21453_, _21452_, _21403_);
  or _72493_ (_21454_, _21453_, _06111_);
  and _72494_ (_21455_, _21454_, _07125_);
  and _72495_ (_21456_, _21455_, _21451_);
  and _72496_ (_21458_, _21456_, _21448_);
  and _72497_ (_21459_, _10289_, _11390_);
  or _72498_ (_21460_, _21459_, _21403_);
  and _72499_ (_21461_, _21460_, _06402_);
  or _72500_ (_21462_, _21461_, _21458_);
  and _72501_ (_21463_, _21462_, _07132_);
  or _72502_ (_21464_, _21403_, _08339_);
  and _72503_ (_21465_, _21453_, _06306_);
  and _72504_ (_21466_, _21465_, _21464_);
  or _72505_ (_21467_, _21466_, _21463_);
  and _72506_ (_21469_, _21467_, _07130_);
  and _72507_ (_21470_, _21411_, _06411_);
  and _72508_ (_21471_, _21470_, _21464_);
  or _72509_ (_21472_, _21471_, _06303_);
  or _72510_ (_21473_, _21472_, _21469_);
  and _72511_ (_21474_, _15026_, _07852_);
  or _72512_ (_21475_, _21403_, _08819_);
  or _72513_ (_21476_, _21475_, _21474_);
  and _72514_ (_21477_, _21476_, _08824_);
  and _72515_ (_21478_, _21477_, _21473_);
  nor _72516_ (_21480_, _10288_, _11468_);
  or _72517_ (_21481_, _21480_, _21403_);
  and _72518_ (_21482_, _21481_, _06396_);
  or _72519_ (_21483_, _21482_, _06433_);
  or _72520_ (_21484_, _21483_, _21478_);
  or _72521_ (_21485_, _21408_, _06829_);
  and _72522_ (_21486_, _21485_, _06444_);
  and _72523_ (_21487_, _21486_, _21484_);
  and _72524_ (_21488_, _15087_, _07852_);
  or _72525_ (_21489_, _21488_, _21403_);
  and _72526_ (_21491_, _21489_, _06440_);
  or _72527_ (_21492_, _21491_, _01321_);
  or _72528_ (_21493_, _21492_, _21487_);
  or _72529_ (_21494_, _01317_, \oc8051_golden_model_1.DPH [4]);
  and _72530_ (_21495_, _21494_, _43100_);
  and _72531_ (_43641_, _21495_, _21493_);
  and _72532_ (_21496_, _11468_, \oc8051_golden_model_1.DPH [5]);
  and _72533_ (_21497_, _08101_, _07852_);
  or _72534_ (_21498_, _21497_, _21496_);
  or _72535_ (_21499_, _21498_, _06132_);
  and _72536_ (_21501_, _15119_, _07852_);
  or _72537_ (_21502_, _21501_, _21496_);
  or _72538_ (_21503_, _21502_, _06161_);
  and _72539_ (_21504_, _11390_, \oc8051_golden_model_1.ACC [5]);
  or _72540_ (_21505_, _21504_, _21496_);
  and _72541_ (_21506_, _21505_, _07056_);
  and _72542_ (_21507_, _07057_, \oc8051_golden_model_1.DPH [5]);
  or _72543_ (_21508_, _21507_, _06160_);
  or _72544_ (_21509_, _21508_, _21506_);
  and _72545_ (_21510_, _21509_, _07075_);
  and _72546_ (_21512_, _21510_, _21503_);
  and _72547_ (_21513_, _21498_, _06217_);
  or _72548_ (_21514_, _21513_, _06220_);
  or _72549_ (_21515_, _21514_, _21512_);
  or _72550_ (_21516_, _21505_, _06229_);
  and _72551_ (_21517_, _21516_, _11312_);
  and _72552_ (_21518_, _21517_, _21515_);
  or _72553_ (_21519_, _11416_, \oc8051_golden_model_1.DPH [5]);
  nor _72554_ (_21520_, _11417_, _11312_);
  and _72555_ (_21521_, _21520_, _21519_);
  or _72556_ (_21523_, _21521_, _21518_);
  and _72557_ (_21524_, _21523_, _11296_);
  nor _72558_ (_21525_, _06477_, _11296_);
  or _72559_ (_21526_, _21525_, _09842_);
  or _72560_ (_21527_, _21526_, _21524_);
  and _72561_ (_21528_, _21527_, _21499_);
  or _72562_ (_21529_, _21528_, _06116_);
  or _72563_ (_21530_, _21496_, _06117_);
  and _72564_ (_21531_, _09208_, _11390_);
  or _72565_ (_21532_, _21531_, _21530_);
  and _72566_ (_21534_, _21532_, _06114_);
  and _72567_ (_21535_, _21534_, _21529_);
  and _72568_ (_21536_, _15203_, _11390_);
  or _72569_ (_21537_, _21536_, _21496_);
  and _72570_ (_21538_, _21537_, _05787_);
  or _72571_ (_21539_, _21538_, _21535_);
  or _72572_ (_21540_, _21539_, _11136_);
  and _72573_ (_21541_, _15219_, _07852_);
  or _72574_ (_21542_, _21496_, _07127_);
  or _72575_ (_21543_, _21542_, _21541_);
  and _72576_ (_21545_, _08736_, _11390_);
  or _72577_ (_21546_, _21545_, _21496_);
  or _72578_ (_21547_, _21546_, _06111_);
  and _72579_ (_21548_, _21547_, _07125_);
  and _72580_ (_21549_, _21548_, _21543_);
  and _72581_ (_21550_, _21549_, _21540_);
  and _72582_ (_21551_, _12325_, _11390_);
  or _72583_ (_21552_, _21551_, _21496_);
  and _72584_ (_21553_, _21552_, _06402_);
  or _72585_ (_21554_, _21553_, _21550_);
  and _72586_ (_21556_, _21554_, _07132_);
  or _72587_ (_21557_, _21496_, _08104_);
  and _72588_ (_21558_, _21546_, _06306_);
  and _72589_ (_21559_, _21558_, _21557_);
  or _72590_ (_21560_, _21559_, _21556_);
  and _72591_ (_21561_, _21560_, _07130_);
  and _72592_ (_21562_, _21505_, _06411_);
  and _72593_ (_21563_, _21562_, _21557_);
  or _72594_ (_21564_, _21563_, _06303_);
  or _72595_ (_21565_, _21564_, _21561_);
  and _72596_ (_21567_, _15216_, _07852_);
  or _72597_ (_21568_, _21496_, _08819_);
  or _72598_ (_21569_, _21568_, _21567_);
  and _72599_ (_21570_, _21569_, _08824_);
  and _72600_ (_21571_, _21570_, _21565_);
  nor _72601_ (_21572_, _10269_, _11468_);
  or _72602_ (_21573_, _21572_, _21496_);
  and _72603_ (_21574_, _21573_, _06396_);
  or _72604_ (_21575_, _21574_, _06433_);
  or _72605_ (_21576_, _21575_, _21571_);
  or _72606_ (_21578_, _21502_, _06829_);
  and _72607_ (_21579_, _21578_, _06444_);
  and _72608_ (_21580_, _21579_, _21576_);
  and _72609_ (_21581_, _15275_, _07852_);
  or _72610_ (_21582_, _21581_, _21496_);
  and _72611_ (_21583_, _21582_, _06440_);
  or _72612_ (_21584_, _21583_, _01321_);
  or _72613_ (_21585_, _21584_, _21580_);
  or _72614_ (_21586_, _01317_, \oc8051_golden_model_1.DPH [5]);
  and _72615_ (_21587_, _21586_, _43100_);
  and _72616_ (_43642_, _21587_, _21585_);
  not _72617_ (_21589_, \oc8051_golden_model_1.DPH [6]);
  nor _72618_ (_21590_, _11390_, _21589_);
  and _72619_ (_21591_, _08012_, _07852_);
  or _72620_ (_21592_, _21591_, _21590_);
  or _72621_ (_21593_, _21592_, _06132_);
  and _72622_ (_21594_, _15300_, _07852_);
  or _72623_ (_21595_, _21594_, _21590_);
  or _72624_ (_21596_, _21595_, _06161_);
  and _72625_ (_21597_, _11390_, \oc8051_golden_model_1.ACC [6]);
  or _72626_ (_21599_, _21597_, _21590_);
  and _72627_ (_21600_, _21599_, _07056_);
  nor _72628_ (_21601_, _07056_, _21589_);
  or _72629_ (_21602_, _21601_, _06160_);
  or _72630_ (_21603_, _21602_, _21600_);
  and _72631_ (_21604_, _21603_, _07075_);
  and _72632_ (_21605_, _21604_, _21596_);
  and _72633_ (_21606_, _21592_, _06217_);
  or _72634_ (_21607_, _21606_, _06220_);
  or _72635_ (_21608_, _21607_, _21605_);
  or _72636_ (_21610_, _21599_, _06229_);
  and _72637_ (_21611_, _21610_, _11312_);
  and _72638_ (_21612_, _21611_, _21608_);
  or _72639_ (_21613_, _11417_, \oc8051_golden_model_1.DPH [6]);
  nor _72640_ (_21614_, _11418_, _11312_);
  and _72641_ (_21615_, _21614_, _21613_);
  or _72642_ (_21616_, _21615_, _21612_);
  and _72643_ (_21617_, _21616_, _11296_);
  nor _72644_ (_21618_, _11296_, _06203_);
  or _72645_ (_21619_, _21618_, _09842_);
  or _72646_ (_21621_, _21619_, _21617_);
  and _72647_ (_21622_, _21621_, _21593_);
  or _72648_ (_21623_, _21622_, _06116_);
  or _72649_ (_21624_, _21590_, _06117_);
  and _72650_ (_21625_, _09207_, _11390_);
  or _72651_ (_21626_, _21625_, _21624_);
  and _72652_ (_21627_, _21626_, _06114_);
  and _72653_ (_21628_, _21627_, _21623_);
  and _72654_ (_21629_, _15395_, _11390_);
  or _72655_ (_21630_, _21629_, _21590_);
  and _72656_ (_21632_, _21630_, _05787_);
  or _72657_ (_21633_, _21632_, _21628_);
  or _72658_ (_21634_, _21633_, _11136_);
  and _72659_ (_21635_, _15413_, _07852_);
  or _72660_ (_21636_, _21590_, _07127_);
  or _72661_ (_21637_, _21636_, _21635_);
  and _72662_ (_21638_, _15402_, _11390_);
  or _72663_ (_21639_, _21638_, _21590_);
  or _72664_ (_21640_, _21639_, _06111_);
  and _72665_ (_21641_, _21640_, _07125_);
  and _72666_ (_21643_, _21641_, _21637_);
  and _72667_ (_21644_, _21643_, _21634_);
  and _72668_ (_21645_, _10295_, _11390_);
  or _72669_ (_21646_, _21645_, _21590_);
  and _72670_ (_21647_, _21646_, _06402_);
  or _72671_ (_21648_, _21647_, _21644_);
  and _72672_ (_21649_, _21648_, _07132_);
  or _72673_ (_21650_, _21590_, _08015_);
  and _72674_ (_21651_, _21639_, _06306_);
  and _72675_ (_21652_, _21651_, _21650_);
  or _72676_ (_21654_, _21652_, _21649_);
  and _72677_ (_21655_, _21654_, _07130_);
  and _72678_ (_21656_, _21599_, _06411_);
  and _72679_ (_21657_, _21656_, _21650_);
  or _72680_ (_21658_, _21657_, _06303_);
  or _72681_ (_21659_, _21658_, _21655_);
  and _72682_ (_21660_, _15410_, _07852_);
  or _72683_ (_21661_, _21590_, _08819_);
  or _72684_ (_21662_, _21661_, _21660_);
  and _72685_ (_21663_, _21662_, _08824_);
  and _72686_ (_21665_, _21663_, _21659_);
  nor _72687_ (_21666_, _10294_, _11468_);
  or _72688_ (_21667_, _21666_, _21590_);
  and _72689_ (_21668_, _21667_, _06396_);
  or _72690_ (_21669_, _21668_, _06433_);
  or _72691_ (_21670_, _21669_, _21665_);
  or _72692_ (_21671_, _21595_, _06829_);
  and _72693_ (_21672_, _21671_, _06444_);
  and _72694_ (_21673_, _21672_, _21670_);
  and _72695_ (_21674_, _15478_, _07852_);
  or _72696_ (_21676_, _21674_, _21590_);
  and _72697_ (_21677_, _21676_, _06440_);
  or _72698_ (_21678_, _21677_, _01321_);
  or _72699_ (_21679_, _21678_, _21673_);
  or _72700_ (_21680_, _01317_, \oc8051_golden_model_1.DPH [6]);
  and _72701_ (_21681_, _21680_, _43100_);
  and _72702_ (_43643_, _21681_, _21679_);
  not _72703_ (_21682_, \oc8051_golden_model_1.TL1 [0]);
  nor _72704_ (_21683_, _01317_, _21682_);
  nand _72705_ (_21684_, _10276_, _07837_);
  nor _72706_ (_21686_, _07837_, _21682_);
  nor _72707_ (_21687_, _21686_, _07130_);
  nand _72708_ (_21688_, _21687_, _21684_);
  nor _72709_ (_21689_, _08211_, _11484_);
  or _72710_ (_21690_, _21689_, _21686_);
  or _72711_ (_21691_, _21690_, _06161_);
  and _72712_ (_21692_, _07837_, \oc8051_golden_model_1.ACC [0]);
  or _72713_ (_21693_, _21692_, _21686_);
  and _72714_ (_21694_, _21693_, _07056_);
  nor _72715_ (_21695_, _07056_, _21682_);
  or _72716_ (_21697_, _21695_, _06160_);
  or _72717_ (_21698_, _21697_, _21694_);
  and _72718_ (_21699_, _21698_, _07075_);
  and _72719_ (_21700_, _21699_, _21691_);
  and _72720_ (_21701_, _07837_, _07049_);
  or _72721_ (_21702_, _21701_, _21686_);
  and _72722_ (_21703_, _21702_, _06217_);
  or _72723_ (_21704_, _21703_, _21700_);
  and _72724_ (_21705_, _21704_, _06229_);
  and _72725_ (_21706_, _21693_, _06220_);
  or _72726_ (_21708_, _21706_, _09842_);
  or _72727_ (_21709_, _21708_, _21705_);
  or _72728_ (_21710_, _21702_, _06132_);
  and _72729_ (_21711_, _21710_, _21709_);
  or _72730_ (_21712_, _21711_, _06116_);
  and _72731_ (_21713_, _09160_, _07837_);
  or _72732_ (_21714_, _21686_, _06117_);
  or _72733_ (_21715_, _21714_, _21713_);
  and _72734_ (_21716_, _21715_, _21712_);
  or _72735_ (_21717_, _21716_, _05787_);
  and _72736_ (_21719_, _14260_, _07837_);
  or _72737_ (_21720_, _21686_, _06114_);
  or _72738_ (_21721_, _21720_, _21719_);
  and _72739_ (_21722_, _21721_, _06111_);
  and _72740_ (_21723_, _21722_, _21717_);
  and _72741_ (_21724_, _07837_, _08708_);
  or _72742_ (_21725_, _21724_, _21686_);
  and _72743_ (_21726_, _21725_, _06110_);
  or _72744_ (_21727_, _21726_, _06297_);
  or _72745_ (_21728_, _21727_, _21723_);
  and _72746_ (_21730_, _14275_, _07837_);
  or _72747_ (_21731_, _21730_, _21686_);
  or _72748_ (_21732_, _21731_, _07127_);
  and _72749_ (_21733_, _21732_, _07125_);
  and _72750_ (_21734_, _21733_, _21728_);
  nor _72751_ (_21735_, _12321_, _11484_);
  or _72752_ (_21736_, _21735_, _21686_);
  and _72753_ (_21737_, _21684_, _06402_);
  and _72754_ (_21738_, _21737_, _21736_);
  or _72755_ (_21739_, _21738_, _21734_);
  and _72756_ (_21741_, _21739_, _07132_);
  nand _72757_ (_21742_, _21725_, _06306_);
  nor _72758_ (_21743_, _21742_, _21689_);
  or _72759_ (_21744_, _21743_, _06411_);
  or _72760_ (_21745_, _21744_, _21741_);
  and _72761_ (_21746_, _21745_, _21688_);
  or _72762_ (_21747_, _21746_, _06303_);
  and _72763_ (_21748_, _14167_, _07837_);
  or _72764_ (_21749_, _21686_, _08819_);
  or _72765_ (_21750_, _21749_, _21748_);
  and _72766_ (_21751_, _21750_, _08824_);
  and _72767_ (_21752_, _21751_, _21747_);
  and _72768_ (_21753_, _21736_, _06396_);
  or _72769_ (_21754_, _21753_, _19287_);
  or _72770_ (_21755_, _21754_, _21752_);
  or _72771_ (_21756_, _21690_, _06630_);
  and _72772_ (_21757_, _21756_, _01317_);
  and _72773_ (_21758_, _21757_, _21755_);
  or _72774_ (_21759_, _21758_, _21683_);
  and _72775_ (_43645_, _21759_, _43100_);
  not _72776_ (_21762_, \oc8051_golden_model_1.TL1 [1]);
  nor _72777_ (_21763_, _01317_, _21762_);
  and _72778_ (_21764_, _09115_, _07837_);
  nor _72779_ (_21765_, _07837_, _21762_);
  or _72780_ (_21766_, _21765_, _06117_);
  or _72781_ (_21767_, _21766_, _21764_);
  and _72782_ (_21768_, _07837_, _07306_);
  or _72783_ (_21769_, _21768_, _21765_);
  or _72784_ (_21770_, _21769_, _06132_);
  or _72785_ (_21771_, _07837_, \oc8051_golden_model_1.TL1 [1]);
  and _72786_ (_21773_, _14363_, _07837_);
  not _72787_ (_21774_, _21773_);
  and _72788_ (_21775_, _21774_, _21771_);
  or _72789_ (_21776_, _21775_, _06161_);
  and _72790_ (_21777_, _07837_, \oc8051_golden_model_1.ACC [1]);
  or _72791_ (_21778_, _21777_, _21765_);
  and _72792_ (_21779_, _21778_, _07056_);
  nor _72793_ (_21780_, _07056_, _21762_);
  or _72794_ (_21781_, _21780_, _06160_);
  or _72795_ (_21782_, _21781_, _21779_);
  and _72796_ (_21784_, _21782_, _07075_);
  and _72797_ (_21785_, _21784_, _21776_);
  and _72798_ (_21786_, _21769_, _06217_);
  or _72799_ (_21787_, _21786_, _21785_);
  and _72800_ (_21788_, _21787_, _06229_);
  and _72801_ (_21789_, _21778_, _06220_);
  or _72802_ (_21790_, _21789_, _09842_);
  or _72803_ (_21791_, _21790_, _21788_);
  and _72804_ (_21792_, _21791_, _21770_);
  or _72805_ (_21793_, _21792_, _06116_);
  and _72806_ (_21795_, _21793_, _06114_);
  and _72807_ (_21796_, _21795_, _21767_);
  or _72808_ (_21797_, _14442_, _11484_);
  and _72809_ (_21798_, _21771_, _05787_);
  and _72810_ (_21799_, _21798_, _21797_);
  or _72811_ (_21800_, _21799_, _21796_);
  and _72812_ (_21801_, _21800_, _06298_);
  or _72813_ (_21802_, _14346_, _11484_);
  and _72814_ (_21803_, _21802_, _06297_);
  nand _72815_ (_21804_, _07837_, _06945_);
  and _72816_ (_21806_, _21804_, _06110_);
  or _72817_ (_21807_, _21806_, _21803_);
  and _72818_ (_21808_, _21807_, _21771_);
  or _72819_ (_21809_, _21808_, _06402_);
  or _72820_ (_21810_, _21809_, _21801_);
  nor _72821_ (_21811_, _10277_, _11484_);
  or _72822_ (_21812_, _21811_, _21765_);
  nand _72823_ (_21813_, _10275_, _07837_);
  and _72824_ (_21814_, _21813_, _21812_);
  or _72825_ (_21815_, _21814_, _07125_);
  and _72826_ (_21817_, _21815_, _07132_);
  and _72827_ (_21818_, _21817_, _21810_);
  or _72828_ (_21819_, _14344_, _11484_);
  and _72829_ (_21820_, _21771_, _06306_);
  and _72830_ (_21821_, _21820_, _21819_);
  or _72831_ (_21822_, _21821_, _06411_);
  or _72832_ (_21823_, _21822_, _21818_);
  nor _72833_ (_21824_, _21765_, _07130_);
  nand _72834_ (_21825_, _21824_, _21813_);
  and _72835_ (_21826_, _21825_, _08819_);
  and _72836_ (_21828_, _21826_, _21823_);
  or _72837_ (_21829_, _21804_, _08176_);
  and _72838_ (_21830_, _21771_, _06303_);
  and _72839_ (_21831_, _21830_, _21829_);
  or _72840_ (_21832_, _21831_, _06396_);
  or _72841_ (_21833_, _21832_, _21828_);
  or _72842_ (_21834_, _21812_, _08824_);
  and _72843_ (_21835_, _21834_, _06829_);
  and _72844_ (_21836_, _21835_, _21833_);
  and _72845_ (_21837_, _21775_, _06433_);
  or _72846_ (_21839_, _21837_, _06440_);
  or _72847_ (_21840_, _21839_, _21836_);
  or _72848_ (_21841_, _21765_, _06444_);
  or _72849_ (_21842_, _21841_, _21773_);
  and _72850_ (_21843_, _21842_, _01317_);
  and _72851_ (_21844_, _21843_, _21840_);
  or _72852_ (_21845_, _21844_, _21763_);
  and _72853_ (_43646_, _21845_, _43100_);
  and _72854_ (_21846_, _01321_, \oc8051_golden_model_1.TL1 [2]);
  and _72855_ (_21847_, _11484_, \oc8051_golden_model_1.TL1 [2]);
  or _72856_ (_21849_, _21847_, _08248_);
  and _72857_ (_21850_, _07837_, _08768_);
  or _72858_ (_21851_, _21850_, _21847_);
  and _72859_ (_21852_, _21851_, _06306_);
  and _72860_ (_21853_, _21852_, _21849_);
  and _72861_ (_21854_, _09211_, _07837_);
  or _72862_ (_21855_, _21854_, _21847_);
  and _72863_ (_21856_, _21855_, _06116_);
  and _72864_ (_21857_, _14542_, _07837_);
  or _72865_ (_21858_, _21857_, _21847_);
  or _72866_ (_21859_, _21858_, _06161_);
  and _72867_ (_21860_, _07837_, \oc8051_golden_model_1.ACC [2]);
  or _72868_ (_21861_, _21860_, _21847_);
  and _72869_ (_21862_, _21861_, _07056_);
  and _72870_ (_21863_, _07057_, \oc8051_golden_model_1.TL1 [2]);
  or _72871_ (_21864_, _21863_, _06160_);
  or _72872_ (_21865_, _21864_, _21862_);
  and _72873_ (_21866_, _21865_, _07075_);
  and _72874_ (_21867_, _21866_, _21859_);
  and _72875_ (_21868_, _07837_, _07708_);
  or _72876_ (_21871_, _21868_, _21847_);
  and _72877_ (_21872_, _21871_, _06217_);
  or _72878_ (_21873_, _21872_, _21867_);
  and _72879_ (_21874_, _21873_, _06229_);
  and _72880_ (_21875_, _21861_, _06220_);
  or _72881_ (_21876_, _21875_, _09842_);
  or _72882_ (_21877_, _21876_, _21874_);
  or _72883_ (_21878_, _21871_, _06132_);
  and _72884_ (_21879_, _21878_, _06117_);
  and _72885_ (_21880_, _21879_, _21877_);
  or _72886_ (_21882_, _21880_, _05787_);
  or _72887_ (_21883_, _21882_, _21856_);
  and _72888_ (_21884_, _14630_, _07837_);
  or _72889_ (_21885_, _21884_, _21847_);
  or _72890_ (_21886_, _21885_, _06114_);
  and _72891_ (_21887_, _21886_, _06111_);
  and _72892_ (_21888_, _21887_, _21883_);
  and _72893_ (_21889_, _21851_, _06110_);
  or _72894_ (_21890_, _21889_, _06297_);
  or _72895_ (_21891_, _21890_, _21888_);
  and _72896_ (_21893_, _14646_, _07837_);
  or _72897_ (_21894_, _21893_, _21847_);
  or _72898_ (_21895_, _21894_, _07127_);
  and _72899_ (_21896_, _21895_, _07125_);
  and _72900_ (_21897_, _21896_, _21891_);
  and _72901_ (_21898_, _10282_, _07837_);
  or _72902_ (_21899_, _21898_, _21847_);
  and _72903_ (_21900_, _21899_, _06402_);
  or _72904_ (_21901_, _21900_, _21897_);
  and _72905_ (_21902_, _21901_, _07132_);
  or _72906_ (_21904_, _21902_, _21853_);
  and _72907_ (_21905_, _21904_, _07130_);
  and _72908_ (_21906_, _21861_, _06411_);
  and _72909_ (_21907_, _21906_, _21849_);
  or _72910_ (_21908_, _21907_, _06303_);
  or _72911_ (_21909_, _21908_, _21905_);
  and _72912_ (_21910_, _14643_, _07837_);
  or _72913_ (_21911_, _21847_, _08819_);
  or _72914_ (_21912_, _21911_, _21910_);
  and _72915_ (_21913_, _21912_, _08824_);
  and _72916_ (_21915_, _21913_, _21909_);
  nor _72917_ (_21916_, _10281_, _11484_);
  or _72918_ (_21917_, _21916_, _21847_);
  and _72919_ (_21918_, _21917_, _06396_);
  or _72920_ (_21919_, _21918_, _21915_);
  and _72921_ (_21920_, _21919_, _06829_);
  and _72922_ (_21921_, _21858_, _06433_);
  or _72923_ (_21922_, _21921_, _06440_);
  or _72924_ (_21923_, _21922_, _21920_);
  and _72925_ (_21924_, _14710_, _07837_);
  or _72926_ (_21926_, _21847_, _06444_);
  or _72927_ (_21927_, _21926_, _21924_);
  and _72928_ (_21928_, _21927_, _01317_);
  and _72929_ (_21929_, _21928_, _21923_);
  or _72930_ (_21930_, _21929_, _21846_);
  and _72931_ (_43647_, _21930_, _43100_);
  and _72932_ (_21931_, _11484_, \oc8051_golden_model_1.TL1 [3]);
  and _72933_ (_21932_, _14738_, _07837_);
  or _72934_ (_21933_, _21932_, _21931_);
  or _72935_ (_21934_, _21933_, _06161_);
  and _72936_ (_21936_, _07837_, \oc8051_golden_model_1.ACC [3]);
  or _72937_ (_21937_, _21936_, _21931_);
  and _72938_ (_21938_, _21937_, _07056_);
  and _72939_ (_21939_, _07057_, \oc8051_golden_model_1.TL1 [3]);
  or _72940_ (_21940_, _21939_, _06160_);
  or _72941_ (_21941_, _21940_, _21938_);
  and _72942_ (_21942_, _21941_, _07075_);
  and _72943_ (_21943_, _21942_, _21934_);
  and _72944_ (_21944_, _07837_, _07544_);
  or _72945_ (_21945_, _21944_, _21931_);
  and _72946_ (_21947_, _21945_, _06217_);
  or _72947_ (_21948_, _21947_, _21943_);
  and _72948_ (_21949_, _21948_, _06229_);
  and _72949_ (_21950_, _21937_, _06220_);
  or _72950_ (_21951_, _21950_, _09842_);
  or _72951_ (_21952_, _21951_, _21949_);
  or _72952_ (_21953_, _21945_, _06132_);
  and _72953_ (_21954_, _21953_, _21952_);
  or _72954_ (_21955_, _21954_, _06116_);
  and _72955_ (_21956_, _09210_, _07837_);
  or _72956_ (_21958_, _21931_, _06117_);
  or _72957_ (_21959_, _21958_, _21956_);
  and _72958_ (_21960_, _21959_, _06114_);
  and _72959_ (_21961_, _21960_, _21955_);
  and _72960_ (_21962_, _14825_, _07837_);
  or _72961_ (_21963_, _21962_, _21931_);
  and _72962_ (_21964_, _21963_, _05787_);
  or _72963_ (_21965_, _21964_, _11136_);
  or _72964_ (_21966_, _21965_, _21961_);
  and _72965_ (_21967_, _14727_, _07837_);
  or _72966_ (_21969_, _21931_, _07127_);
  or _72967_ (_21970_, _21969_, _21967_);
  and _72968_ (_21971_, _07837_, _08712_);
  or _72969_ (_21972_, _21971_, _21931_);
  or _72970_ (_21973_, _21972_, _06111_);
  and _72971_ (_21974_, _21973_, _07125_);
  and _72972_ (_21975_, _21974_, _21970_);
  and _72973_ (_21976_, _21975_, _21966_);
  and _72974_ (_21977_, _12318_, _07837_);
  or _72975_ (_21978_, _21977_, _21931_);
  and _72976_ (_21980_, _21978_, _06402_);
  or _72977_ (_21981_, _21980_, _21976_);
  and _72978_ (_21982_, _21981_, _07132_);
  or _72979_ (_21983_, _21931_, _08140_);
  and _72980_ (_21984_, _21972_, _06306_);
  and _72981_ (_21985_, _21984_, _21983_);
  or _72982_ (_21986_, _21985_, _21982_);
  and _72983_ (_21987_, _21986_, _07130_);
  and _72984_ (_21988_, _21937_, _06411_);
  and _72985_ (_21989_, _21988_, _21983_);
  or _72986_ (_21991_, _21989_, _06303_);
  or _72987_ (_21992_, _21991_, _21987_);
  and _72988_ (_21993_, _14724_, _07837_);
  or _72989_ (_21994_, _21931_, _08819_);
  or _72990_ (_21995_, _21994_, _21993_);
  and _72991_ (_21996_, _21995_, _08824_);
  and _72992_ (_21997_, _21996_, _21992_);
  nor _72993_ (_21998_, _10273_, _11484_);
  or _72994_ (_21999_, _21998_, _21931_);
  and _72995_ (_22000_, _21999_, _06396_);
  or _72996_ (_22002_, _22000_, _06433_);
  or _72997_ (_22003_, _22002_, _21997_);
  or _72998_ (_22004_, _21933_, _06829_);
  and _72999_ (_22005_, _22004_, _06444_);
  and _73000_ (_22006_, _22005_, _22003_);
  and _73001_ (_22007_, _14897_, _07837_);
  or _73002_ (_22008_, _22007_, _21931_);
  and _73003_ (_22009_, _22008_, _06440_);
  or _73004_ (_22010_, _22009_, _01321_);
  or _73005_ (_22011_, _22010_, _22006_);
  or _73006_ (_22013_, _01317_, \oc8051_golden_model_1.TL1 [3]);
  and _73007_ (_22014_, _22013_, _43100_);
  and _73008_ (_43648_, _22014_, _22011_);
  and _73009_ (_22015_, _11484_, \oc8051_golden_model_1.TL1 [4]);
  and _73010_ (_22016_, _14928_, _07837_);
  or _73011_ (_22017_, _22016_, _22015_);
  or _73012_ (_22018_, _22017_, _06161_);
  and _73013_ (_22019_, _07837_, \oc8051_golden_model_1.ACC [4]);
  or _73014_ (_22020_, _22019_, _22015_);
  and _73015_ (_22021_, _22020_, _07056_);
  and _73016_ (_22023_, _07057_, \oc8051_golden_model_1.TL1 [4]);
  or _73017_ (_22024_, _22023_, _06160_);
  or _73018_ (_22025_, _22024_, _22021_);
  and _73019_ (_22026_, _22025_, _07075_);
  and _73020_ (_22027_, _22026_, _22018_);
  and _73021_ (_22028_, _08336_, _07837_);
  or _73022_ (_22029_, _22028_, _22015_);
  and _73023_ (_22030_, _22029_, _06217_);
  or _73024_ (_22031_, _22030_, _22027_);
  and _73025_ (_22032_, _22031_, _06229_);
  and _73026_ (_22034_, _22020_, _06220_);
  or _73027_ (_22035_, _22034_, _09842_);
  or _73028_ (_22036_, _22035_, _22032_);
  or _73029_ (_22037_, _22029_, _06132_);
  and _73030_ (_22038_, _22037_, _22036_);
  or _73031_ (_22039_, _22038_, _06116_);
  and _73032_ (_22040_, _09209_, _07837_);
  or _73033_ (_22041_, _22015_, _06117_);
  or _73034_ (_22042_, _22041_, _22040_);
  and _73035_ (_22043_, _22042_, _06114_);
  and _73036_ (_22045_, _22043_, _22039_);
  and _73037_ (_22046_, _15013_, _07837_);
  or _73038_ (_22047_, _22046_, _22015_);
  and _73039_ (_22048_, _22047_, _05787_);
  or _73040_ (_22049_, _22048_, _22045_);
  or _73041_ (_22050_, _22049_, _11136_);
  and _73042_ (_22051_, _15029_, _07837_);
  or _73043_ (_22052_, _22015_, _07127_);
  or _73044_ (_22053_, _22052_, _22051_);
  and _73045_ (_22054_, _08715_, _07837_);
  or _73046_ (_22056_, _22054_, _22015_);
  or _73047_ (_22057_, _22056_, _06111_);
  and _73048_ (_22058_, _22057_, _07125_);
  and _73049_ (_22059_, _22058_, _22053_);
  and _73050_ (_22060_, _22059_, _22050_);
  and _73051_ (_22061_, _10289_, _07837_);
  or _73052_ (_22062_, _22061_, _22015_);
  and _73053_ (_22063_, _22062_, _06402_);
  or _73054_ (_22064_, _22063_, _22060_);
  and _73055_ (_22065_, _22064_, _07132_);
  or _73056_ (_22067_, _22015_, _08339_);
  and _73057_ (_22068_, _22056_, _06306_);
  and _73058_ (_22069_, _22068_, _22067_);
  or _73059_ (_22070_, _22069_, _22065_);
  and _73060_ (_22071_, _22070_, _07130_);
  and _73061_ (_22072_, _22020_, _06411_);
  and _73062_ (_22073_, _22072_, _22067_);
  or _73063_ (_22074_, _22073_, _06303_);
  or _73064_ (_22075_, _22074_, _22071_);
  and _73065_ (_22076_, _15026_, _07837_);
  or _73066_ (_22078_, _22015_, _08819_);
  or _73067_ (_22079_, _22078_, _22076_);
  and _73068_ (_22080_, _22079_, _08824_);
  and _73069_ (_22081_, _22080_, _22075_);
  nor _73070_ (_22082_, _10288_, _11484_);
  or _73071_ (_22083_, _22082_, _22015_);
  and _73072_ (_22084_, _22083_, _06396_);
  or _73073_ (_22085_, _22084_, _06433_);
  or _73074_ (_22086_, _22085_, _22081_);
  or _73075_ (_22087_, _22017_, _06829_);
  and _73076_ (_22089_, _22087_, _06444_);
  and _73077_ (_22090_, _22089_, _22086_);
  and _73078_ (_22091_, _15087_, _07837_);
  or _73079_ (_22092_, _22091_, _22015_);
  and _73080_ (_22093_, _22092_, _06440_);
  or _73081_ (_22094_, _22093_, _01321_);
  or _73082_ (_22095_, _22094_, _22090_);
  or _73083_ (_22096_, _01317_, \oc8051_golden_model_1.TL1 [4]);
  and _73084_ (_22097_, _22096_, _43100_);
  and _73085_ (_43649_, _22097_, _22095_);
  and _73086_ (_22099_, _11484_, \oc8051_golden_model_1.TL1 [5]);
  or _73087_ (_22100_, _22099_, _08104_);
  and _73088_ (_22101_, _08736_, _07837_);
  or _73089_ (_22102_, _22101_, _22099_);
  and _73090_ (_22103_, _22102_, _06306_);
  and _73091_ (_22104_, _22103_, _22100_);
  and _73092_ (_22105_, _15119_, _07837_);
  or _73093_ (_22106_, _22105_, _22099_);
  or _73094_ (_22107_, _22106_, _06161_);
  and _73095_ (_22108_, _07837_, \oc8051_golden_model_1.ACC [5]);
  or _73096_ (_22110_, _22108_, _22099_);
  and _73097_ (_22111_, _22110_, _07056_);
  and _73098_ (_22112_, _07057_, \oc8051_golden_model_1.TL1 [5]);
  or _73099_ (_22113_, _22112_, _06160_);
  or _73100_ (_22114_, _22113_, _22111_);
  and _73101_ (_22115_, _22114_, _07075_);
  and _73102_ (_22116_, _22115_, _22107_);
  and _73103_ (_22117_, _08101_, _07837_);
  or _73104_ (_22118_, _22117_, _22099_);
  and _73105_ (_22119_, _22118_, _06217_);
  or _73106_ (_22121_, _22119_, _22116_);
  and _73107_ (_22122_, _22121_, _06229_);
  and _73108_ (_22123_, _22110_, _06220_);
  or _73109_ (_22124_, _22123_, _09842_);
  or _73110_ (_22125_, _22124_, _22122_);
  or _73111_ (_22126_, _22118_, _06132_);
  and _73112_ (_22127_, _22126_, _22125_);
  or _73113_ (_22128_, _22127_, _06116_);
  and _73114_ (_22129_, _09208_, _07837_);
  or _73115_ (_22130_, _22099_, _06117_);
  or _73116_ (_22132_, _22130_, _22129_);
  and _73117_ (_22133_, _22132_, _06114_);
  and _73118_ (_22134_, _22133_, _22128_);
  and _73119_ (_22135_, _15203_, _07837_);
  or _73120_ (_22136_, _22135_, _22099_);
  and _73121_ (_22137_, _22136_, _05787_);
  or _73122_ (_22138_, _22137_, _11136_);
  or _73123_ (_22139_, _22138_, _22134_);
  and _73124_ (_22140_, _15219_, _07837_);
  or _73125_ (_22141_, _22099_, _07127_);
  or _73126_ (_22143_, _22141_, _22140_);
  or _73127_ (_22144_, _22102_, _06111_);
  and _73128_ (_22145_, _22144_, _07125_);
  and _73129_ (_22146_, _22145_, _22143_);
  and _73130_ (_22147_, _22146_, _22139_);
  and _73131_ (_22148_, _12325_, _07837_);
  or _73132_ (_22149_, _22148_, _22099_);
  and _73133_ (_22150_, _22149_, _06402_);
  or _73134_ (_22151_, _22150_, _22147_);
  and _73135_ (_22152_, _22151_, _07132_);
  or _73136_ (_22154_, _22152_, _22104_);
  and _73137_ (_22155_, _22154_, _07130_);
  and _73138_ (_22156_, _22110_, _06411_);
  and _73139_ (_22157_, _22156_, _22100_);
  or _73140_ (_22158_, _22157_, _06303_);
  or _73141_ (_22159_, _22158_, _22155_);
  and _73142_ (_22160_, _15216_, _07837_);
  or _73143_ (_22161_, _22099_, _08819_);
  or _73144_ (_22162_, _22161_, _22160_);
  and _73145_ (_22163_, _22162_, _08824_);
  and _73146_ (_22165_, _22163_, _22159_);
  nor _73147_ (_22166_, _10269_, _11484_);
  or _73148_ (_22167_, _22166_, _22099_);
  and _73149_ (_22168_, _22167_, _06396_);
  or _73150_ (_22169_, _22168_, _06433_);
  or _73151_ (_22170_, _22169_, _22165_);
  or _73152_ (_22171_, _22106_, _06829_);
  and _73153_ (_22172_, _22171_, _06444_);
  and _73154_ (_22173_, _22172_, _22170_);
  and _73155_ (_22174_, _15275_, _07837_);
  or _73156_ (_22176_, _22174_, _22099_);
  and _73157_ (_22177_, _22176_, _06440_);
  or _73158_ (_22178_, _22177_, _01321_);
  or _73159_ (_22179_, _22178_, _22173_);
  or _73160_ (_22180_, _01317_, \oc8051_golden_model_1.TL1 [5]);
  and _73161_ (_22181_, _22180_, _43100_);
  and _73162_ (_43650_, _22181_, _22179_);
  and _73163_ (_22182_, _11484_, \oc8051_golden_model_1.TL1 [6]);
  or _73164_ (_22183_, _22182_, _08015_);
  and _73165_ (_22184_, _15402_, _07837_);
  or _73166_ (_22186_, _22184_, _22182_);
  and _73167_ (_22187_, _22186_, _06306_);
  and _73168_ (_22188_, _22187_, _22183_);
  and _73169_ (_22189_, _15300_, _07837_);
  or _73170_ (_22190_, _22189_, _22182_);
  or _73171_ (_22191_, _22190_, _06161_);
  and _73172_ (_22192_, _07837_, \oc8051_golden_model_1.ACC [6]);
  or _73173_ (_22193_, _22192_, _22182_);
  and _73174_ (_22194_, _22193_, _07056_);
  and _73175_ (_22195_, _07057_, \oc8051_golden_model_1.TL1 [6]);
  or _73176_ (_22197_, _22195_, _06160_);
  or _73177_ (_22198_, _22197_, _22194_);
  and _73178_ (_22199_, _22198_, _07075_);
  and _73179_ (_22200_, _22199_, _22191_);
  and _73180_ (_22201_, _08012_, _07837_);
  or _73181_ (_22202_, _22201_, _22182_);
  and _73182_ (_22203_, _22202_, _06217_);
  or _73183_ (_22204_, _22203_, _22200_);
  and _73184_ (_22205_, _22204_, _06229_);
  and _73185_ (_22206_, _22193_, _06220_);
  or _73186_ (_22208_, _22206_, _09842_);
  or _73187_ (_22209_, _22208_, _22205_);
  or _73188_ (_22210_, _22202_, _06132_);
  and _73189_ (_22211_, _22210_, _22209_);
  or _73190_ (_22212_, _22211_, _06116_);
  and _73191_ (_22213_, _09207_, _07837_);
  or _73192_ (_22214_, _22182_, _06117_);
  or _73193_ (_22215_, _22214_, _22213_);
  and _73194_ (_22216_, _22215_, _06114_);
  and _73195_ (_22217_, _22216_, _22212_);
  and _73196_ (_22220_, _15395_, _07837_);
  or _73197_ (_22221_, _22220_, _22182_);
  and _73198_ (_22222_, _22221_, _05787_);
  or _73199_ (_22223_, _22222_, _11136_);
  or _73200_ (_22224_, _22223_, _22217_);
  and _73201_ (_22225_, _15413_, _07837_);
  or _73202_ (_22226_, _22182_, _07127_);
  or _73203_ (_22227_, _22226_, _22225_);
  or _73204_ (_22228_, _22186_, _06111_);
  and _73205_ (_22229_, _22228_, _07125_);
  and _73206_ (_22231_, _22229_, _22227_);
  and _73207_ (_22232_, _22231_, _22224_);
  and _73208_ (_22233_, _10295_, _07837_);
  or _73209_ (_22234_, _22233_, _22182_);
  and _73210_ (_22235_, _22234_, _06402_);
  or _73211_ (_22236_, _22235_, _22232_);
  and _73212_ (_22237_, _22236_, _07132_);
  or _73213_ (_22238_, _22237_, _22188_);
  and _73214_ (_22239_, _22238_, _07130_);
  and _73215_ (_22240_, _22193_, _06411_);
  and _73216_ (_22242_, _22240_, _22183_);
  or _73217_ (_22243_, _22242_, _06303_);
  or _73218_ (_22244_, _22243_, _22239_);
  and _73219_ (_22245_, _15410_, _07837_);
  or _73220_ (_22246_, _22182_, _08819_);
  or _73221_ (_22247_, _22246_, _22245_);
  and _73222_ (_22248_, _22247_, _08824_);
  and _73223_ (_22249_, _22248_, _22244_);
  nor _73224_ (_22250_, _10294_, _11484_);
  or _73225_ (_22251_, _22250_, _22182_);
  and _73226_ (_22253_, _22251_, _06396_);
  or _73227_ (_22254_, _22253_, _06433_);
  or _73228_ (_22255_, _22254_, _22249_);
  or _73229_ (_22256_, _22190_, _06829_);
  and _73230_ (_22257_, _22256_, _06444_);
  and _73231_ (_22258_, _22257_, _22255_);
  and _73232_ (_22259_, _15478_, _07837_);
  or _73233_ (_22260_, _22259_, _22182_);
  and _73234_ (_22261_, _22260_, _06440_);
  or _73235_ (_22262_, _22261_, _01321_);
  or _73236_ (_22264_, _22262_, _22258_);
  or _73237_ (_22265_, _01317_, \oc8051_golden_model_1.TL1 [6]);
  and _73238_ (_22266_, _22265_, _43100_);
  and _73239_ (_43651_, _22266_, _22264_);
  not _73240_ (_22267_, \oc8051_golden_model_1.TL0 [0]);
  nor _73241_ (_22268_, _01317_, _22267_);
  nand _73242_ (_22269_, _10276_, _07803_);
  nor _73243_ (_22270_, _07803_, _22267_);
  nor _73244_ (_22271_, _22270_, _07130_);
  nand _73245_ (_22272_, _22271_, _22269_);
  and _73246_ (_22274_, _07803_, _07049_);
  or _73247_ (_22275_, _22274_, _22270_);
  or _73248_ (_22276_, _22275_, _06132_);
  nor _73249_ (_22277_, _08211_, _11561_);
  or _73250_ (_22278_, _22277_, _22270_);
  or _73251_ (_22279_, _22278_, _06161_);
  and _73252_ (_22280_, _07803_, \oc8051_golden_model_1.ACC [0]);
  or _73253_ (_22281_, _22280_, _22270_);
  and _73254_ (_22282_, _22281_, _07056_);
  nor _73255_ (_22283_, _07056_, _22267_);
  or _73256_ (_22285_, _22283_, _06160_);
  or _73257_ (_22286_, _22285_, _22282_);
  and _73258_ (_22287_, _22286_, _07075_);
  and _73259_ (_22288_, _22287_, _22279_);
  and _73260_ (_22289_, _22275_, _06217_);
  or _73261_ (_22290_, _22289_, _22288_);
  and _73262_ (_22291_, _22290_, _06229_);
  and _73263_ (_22292_, _22281_, _06220_);
  or _73264_ (_22293_, _22292_, _09842_);
  or _73265_ (_22294_, _22293_, _22291_);
  and _73266_ (_22296_, _22294_, _22276_);
  or _73267_ (_22297_, _22296_, _06116_);
  and _73268_ (_22298_, _09160_, _07803_);
  or _73269_ (_22299_, _22270_, _06117_);
  or _73270_ (_22300_, _22299_, _22298_);
  and _73271_ (_22301_, _22300_, _22297_);
  or _73272_ (_22302_, _22301_, _05787_);
  and _73273_ (_22303_, _14260_, _07803_);
  or _73274_ (_22304_, _22303_, _22270_);
  or _73275_ (_22305_, _22304_, _06114_);
  and _73276_ (_22306_, _22305_, _06111_);
  and _73277_ (_22307_, _22306_, _22302_);
  and _73278_ (_22308_, _07803_, _08708_);
  or _73279_ (_22309_, _22308_, _22270_);
  and _73280_ (_22310_, _22309_, _06110_);
  or _73281_ (_22311_, _22310_, _06297_);
  or _73282_ (_22312_, _22311_, _22307_);
  and _73283_ (_22313_, _14275_, _07803_);
  or _73284_ (_22314_, _22270_, _07127_);
  or _73285_ (_22315_, _22314_, _22313_);
  and _73286_ (_22318_, _22315_, _07125_);
  and _73287_ (_22319_, _22318_, _22312_);
  nor _73288_ (_22320_, _12321_, _11561_);
  or _73289_ (_22321_, _22320_, _22270_);
  and _73290_ (_22322_, _22269_, _06402_);
  and _73291_ (_22323_, _22322_, _22321_);
  or _73292_ (_22324_, _22323_, _22319_);
  and _73293_ (_22325_, _22324_, _07132_);
  nand _73294_ (_22326_, _22309_, _06306_);
  nor _73295_ (_22327_, _22326_, _22277_);
  or _73296_ (_22329_, _22327_, _06411_);
  or _73297_ (_22330_, _22329_, _22325_);
  and _73298_ (_22331_, _22330_, _22272_);
  or _73299_ (_22332_, _22331_, _06303_);
  and _73300_ (_22333_, _14167_, _07803_);
  or _73301_ (_22334_, _22333_, _22270_);
  or _73302_ (_22335_, _22334_, _08819_);
  and _73303_ (_22336_, _22335_, _08824_);
  and _73304_ (_22337_, _22336_, _22332_);
  and _73305_ (_22338_, _22321_, _06396_);
  or _73306_ (_22340_, _22338_, _19287_);
  or _73307_ (_22341_, _22340_, _22337_);
  or _73308_ (_22342_, _22278_, _06630_);
  and _73309_ (_22343_, _22342_, _01317_);
  and _73310_ (_22344_, _22343_, _22341_);
  or _73311_ (_22345_, _22344_, _22268_);
  and _73312_ (_43653_, _22345_, _43100_);
  and _73313_ (_22346_, _11561_, \oc8051_golden_model_1.TL0 [1]);
  nor _73314_ (_22347_, _10277_, _11561_);
  or _73315_ (_22348_, _22347_, _22346_);
  or _73316_ (_22350_, _22348_, _08824_);
  or _73317_ (_22351_, _14442_, _11561_);
  or _73318_ (_22352_, _07803_, \oc8051_golden_model_1.TL0 [1]);
  and _73319_ (_22353_, _22352_, _05787_);
  and _73320_ (_22354_, _22353_, _22351_);
  and _73321_ (_22355_, _09115_, _07803_);
  or _73322_ (_22356_, _22346_, _06117_);
  or _73323_ (_22357_, _22356_, _22355_);
  and _73324_ (_22358_, _14363_, _07803_);
  not _73325_ (_22359_, _22358_);
  and _73326_ (_22361_, _22359_, _22352_);
  or _73327_ (_22362_, _22361_, _06161_);
  and _73328_ (_22363_, _07803_, \oc8051_golden_model_1.ACC [1]);
  or _73329_ (_22364_, _22363_, _22346_);
  and _73330_ (_22365_, _22364_, _07056_);
  and _73331_ (_22366_, _07057_, \oc8051_golden_model_1.TL0 [1]);
  or _73332_ (_22367_, _22366_, _06160_);
  or _73333_ (_22368_, _22367_, _22365_);
  and _73334_ (_22369_, _22368_, _07075_);
  and _73335_ (_22370_, _22369_, _22362_);
  and _73336_ (_22372_, _07803_, _07306_);
  or _73337_ (_22373_, _22372_, _22346_);
  and _73338_ (_22374_, _22373_, _06217_);
  or _73339_ (_22375_, _22374_, _22370_);
  and _73340_ (_22376_, _22375_, _06229_);
  and _73341_ (_22377_, _22364_, _06220_);
  or _73342_ (_22378_, _22377_, _09842_);
  or _73343_ (_22379_, _22378_, _22376_);
  or _73344_ (_22380_, _22373_, _06132_);
  and _73345_ (_22381_, _22380_, _22379_);
  or _73346_ (_22383_, _22381_, _06116_);
  and _73347_ (_22384_, _22383_, _06114_);
  and _73348_ (_22385_, _22384_, _22357_);
  or _73349_ (_22386_, _22385_, _22354_);
  and _73350_ (_22387_, _22386_, _06298_);
  or _73351_ (_22388_, _14346_, _11561_);
  and _73352_ (_22389_, _22388_, _06297_);
  nand _73353_ (_22390_, _07803_, _06945_);
  and _73354_ (_22391_, _22390_, _06110_);
  or _73355_ (_22392_, _22391_, _22389_);
  and _73356_ (_22394_, _22392_, _22352_);
  or _73357_ (_22395_, _22394_, _06402_);
  or _73358_ (_22396_, _22395_, _22387_);
  nand _73359_ (_22397_, _10275_, _07803_);
  and _73360_ (_22398_, _22397_, _22348_);
  or _73361_ (_22399_, _22398_, _07125_);
  and _73362_ (_22400_, _22399_, _07132_);
  and _73363_ (_22401_, _22400_, _22396_);
  or _73364_ (_22402_, _14344_, _11561_);
  and _73365_ (_22403_, _22352_, _06306_);
  and _73366_ (_22405_, _22403_, _22402_);
  or _73367_ (_22406_, _22405_, _06411_);
  or _73368_ (_22407_, _22406_, _22401_);
  nor _73369_ (_22408_, _22346_, _07130_);
  nand _73370_ (_22409_, _22408_, _22397_);
  and _73371_ (_22410_, _22409_, _08819_);
  and _73372_ (_22411_, _22410_, _22407_);
  or _73373_ (_22412_, _22390_, _08176_);
  and _73374_ (_22413_, _22352_, _06303_);
  and _73375_ (_22414_, _22413_, _22412_);
  or _73376_ (_22416_, _22414_, _06396_);
  or _73377_ (_22417_, _22416_, _22411_);
  and _73378_ (_22418_, _22417_, _22350_);
  or _73379_ (_22419_, _22418_, _06433_);
  or _73380_ (_22420_, _22361_, _06829_);
  and _73381_ (_22421_, _22420_, _06444_);
  and _73382_ (_22422_, _22421_, _22419_);
  or _73383_ (_22423_, _22358_, _22346_);
  and _73384_ (_22424_, _22423_, _06440_);
  or _73385_ (_22425_, _22424_, _01321_);
  or _73386_ (_22427_, _22425_, _22422_);
  or _73387_ (_22428_, _01317_, \oc8051_golden_model_1.TL0 [1]);
  and _73388_ (_22429_, _22428_, _43100_);
  and _73389_ (_43654_, _22429_, _22427_);
  and _73390_ (_22430_, _01321_, \oc8051_golden_model_1.TL0 [2]);
  and _73391_ (_22431_, _11561_, \oc8051_golden_model_1.TL0 [2]);
  and _73392_ (_22432_, _09211_, _07803_);
  or _73393_ (_22433_, _22432_, _22431_);
  and _73394_ (_22434_, _22433_, _06116_);
  and _73395_ (_22435_, _14542_, _07803_);
  or _73396_ (_22437_, _22435_, _22431_);
  or _73397_ (_22438_, _22437_, _06161_);
  and _73398_ (_22439_, _07803_, \oc8051_golden_model_1.ACC [2]);
  or _73399_ (_22440_, _22439_, _22431_);
  and _73400_ (_22441_, _22440_, _07056_);
  and _73401_ (_22442_, _07057_, \oc8051_golden_model_1.TL0 [2]);
  or _73402_ (_22443_, _22442_, _06160_);
  or _73403_ (_22444_, _22443_, _22441_);
  and _73404_ (_22445_, _22444_, _07075_);
  and _73405_ (_22446_, _22445_, _22438_);
  and _73406_ (_22448_, _07803_, _07708_);
  or _73407_ (_22449_, _22448_, _22431_);
  and _73408_ (_22450_, _22449_, _06217_);
  or _73409_ (_22451_, _22450_, _22446_);
  and _73410_ (_22452_, _22451_, _06229_);
  and _73411_ (_22453_, _22440_, _06220_);
  or _73412_ (_22454_, _22453_, _09842_);
  or _73413_ (_22455_, _22454_, _22452_);
  or _73414_ (_22456_, _22449_, _06132_);
  and _73415_ (_22457_, _22456_, _06117_);
  and _73416_ (_22459_, _22457_, _22455_);
  or _73417_ (_22460_, _22459_, _05787_);
  or _73418_ (_22461_, _22460_, _22434_);
  and _73419_ (_22462_, _14630_, _07803_);
  or _73420_ (_22463_, _22431_, _06114_);
  or _73421_ (_22464_, _22463_, _22462_);
  and _73422_ (_22465_, _22464_, _06111_);
  and _73423_ (_22466_, _22465_, _22461_);
  and _73424_ (_22467_, _07803_, _08768_);
  or _73425_ (_22468_, _22467_, _22431_);
  and _73426_ (_22470_, _22468_, _06110_);
  or _73427_ (_22471_, _22470_, _06297_);
  or _73428_ (_22472_, _22471_, _22466_);
  and _73429_ (_22473_, _14646_, _07803_);
  or _73430_ (_22474_, _22473_, _22431_);
  or _73431_ (_22475_, _22474_, _07127_);
  and _73432_ (_22476_, _22475_, _07125_);
  and _73433_ (_22477_, _22476_, _22472_);
  and _73434_ (_22478_, _10282_, _07803_);
  or _73435_ (_22479_, _22478_, _22431_);
  and _73436_ (_22481_, _22479_, _06402_);
  or _73437_ (_22482_, _22481_, _22477_);
  and _73438_ (_22483_, _22482_, _07132_);
  or _73439_ (_22484_, _22431_, _08248_);
  and _73440_ (_22485_, _22468_, _06306_);
  and _73441_ (_22486_, _22485_, _22484_);
  or _73442_ (_22487_, _22486_, _22483_);
  and _73443_ (_22488_, _22487_, _07130_);
  and _73444_ (_22489_, _22440_, _06411_);
  and _73445_ (_22490_, _22489_, _22484_);
  or _73446_ (_22492_, _22490_, _06303_);
  or _73447_ (_22493_, _22492_, _22488_);
  and _73448_ (_22494_, _14643_, _07803_);
  or _73449_ (_22495_, _22431_, _08819_);
  or _73450_ (_22496_, _22495_, _22494_);
  and _73451_ (_22497_, _22496_, _08824_);
  and _73452_ (_22498_, _22497_, _22493_);
  nor _73453_ (_22499_, _10281_, _11561_);
  or _73454_ (_22500_, _22499_, _22431_);
  and _73455_ (_22501_, _22500_, _06396_);
  or _73456_ (_22503_, _22501_, _22498_);
  and _73457_ (_22504_, _22503_, _06829_);
  and _73458_ (_22505_, _22437_, _06433_);
  or _73459_ (_22506_, _22505_, _06440_);
  or _73460_ (_22507_, _22506_, _22504_);
  and _73461_ (_22508_, _14710_, _07803_);
  or _73462_ (_22509_, _22431_, _06444_);
  or _73463_ (_22510_, _22509_, _22508_);
  and _73464_ (_22511_, _22510_, _01317_);
  and _73465_ (_22512_, _22511_, _22507_);
  or _73466_ (_22514_, _22512_, _22430_);
  and _73467_ (_43655_, _22514_, _43100_);
  and _73468_ (_22515_, _11561_, \oc8051_golden_model_1.TL0 [3]);
  or _73469_ (_22516_, _22515_, _08140_);
  and _73470_ (_22517_, _07803_, _08712_);
  or _73471_ (_22518_, _22517_, _22515_);
  and _73472_ (_22519_, _22518_, _06306_);
  and _73473_ (_22520_, _22519_, _22516_);
  and _73474_ (_22521_, _14738_, _07803_);
  or _73475_ (_22522_, _22521_, _22515_);
  or _73476_ (_22524_, _22522_, _06161_);
  and _73477_ (_22525_, _07803_, \oc8051_golden_model_1.ACC [3]);
  or _73478_ (_22526_, _22525_, _22515_);
  and _73479_ (_22527_, _22526_, _07056_);
  and _73480_ (_22528_, _07057_, \oc8051_golden_model_1.TL0 [3]);
  or _73481_ (_22529_, _22528_, _06160_);
  or _73482_ (_22530_, _22529_, _22527_);
  and _73483_ (_22531_, _22530_, _07075_);
  and _73484_ (_22532_, _22531_, _22524_);
  and _73485_ (_22533_, _07803_, _07544_);
  or _73486_ (_22535_, _22533_, _22515_);
  and _73487_ (_22536_, _22535_, _06217_);
  or _73488_ (_22537_, _22536_, _22532_);
  and _73489_ (_22538_, _22537_, _06229_);
  and _73490_ (_22539_, _22526_, _06220_);
  or _73491_ (_22540_, _22539_, _09842_);
  or _73492_ (_22541_, _22540_, _22538_);
  or _73493_ (_22542_, _22535_, _06132_);
  and _73494_ (_22543_, _22542_, _06117_);
  and _73495_ (_22544_, _22543_, _22541_);
  and _73496_ (_22546_, _09210_, _07803_);
  or _73497_ (_22547_, _22546_, _22515_);
  and _73498_ (_22548_, _22547_, _06116_);
  or _73499_ (_22549_, _22548_, _05787_);
  or _73500_ (_22550_, _22549_, _22544_);
  and _73501_ (_22551_, _14825_, _07803_);
  or _73502_ (_22552_, _22551_, _22515_);
  or _73503_ (_22553_, _22552_, _06114_);
  and _73504_ (_22554_, _22553_, _06111_);
  and _73505_ (_22555_, _22554_, _22550_);
  and _73506_ (_22557_, _22518_, _06110_);
  or _73507_ (_22558_, _22557_, _06297_);
  or _73508_ (_22559_, _22558_, _22555_);
  and _73509_ (_22560_, _14727_, _07803_);
  or _73510_ (_22561_, _22515_, _07127_);
  or _73511_ (_22562_, _22561_, _22560_);
  and _73512_ (_22563_, _22562_, _07125_);
  and _73513_ (_22564_, _22563_, _22559_);
  and _73514_ (_22565_, _12318_, _07803_);
  or _73515_ (_22566_, _22565_, _22515_);
  and _73516_ (_22568_, _22566_, _06402_);
  or _73517_ (_22569_, _22568_, _22564_);
  and _73518_ (_22570_, _22569_, _07132_);
  or _73519_ (_22571_, _22570_, _22520_);
  and _73520_ (_22572_, _22571_, _07130_);
  and _73521_ (_22573_, _22526_, _06411_);
  and _73522_ (_22574_, _22573_, _22516_);
  or _73523_ (_22575_, _22574_, _06303_);
  or _73524_ (_22576_, _22575_, _22572_);
  and _73525_ (_22577_, _14724_, _07803_);
  or _73526_ (_22579_, _22515_, _08819_);
  or _73527_ (_22580_, _22579_, _22577_);
  and _73528_ (_22581_, _22580_, _08824_);
  and _73529_ (_22582_, _22581_, _22576_);
  nor _73530_ (_22583_, _10273_, _11561_);
  or _73531_ (_22584_, _22583_, _22515_);
  and _73532_ (_22585_, _22584_, _06396_);
  or _73533_ (_22586_, _22585_, _06433_);
  or _73534_ (_22587_, _22586_, _22582_);
  or _73535_ (_22588_, _22522_, _06829_);
  and _73536_ (_22590_, _22588_, _06444_);
  and _73537_ (_22591_, _22590_, _22587_);
  and _73538_ (_22592_, _14897_, _07803_);
  or _73539_ (_22593_, _22592_, _22515_);
  and _73540_ (_22594_, _22593_, _06440_);
  or _73541_ (_22595_, _22594_, _01321_);
  or _73542_ (_22596_, _22595_, _22591_);
  or _73543_ (_22597_, _01317_, \oc8051_golden_model_1.TL0 [3]);
  and _73544_ (_22598_, _22597_, _43100_);
  and _73545_ (_43656_, _22598_, _22596_);
  and _73546_ (_22599_, _11561_, \oc8051_golden_model_1.TL0 [4]);
  and _73547_ (_22600_, _08336_, _07803_);
  or _73548_ (_22601_, _22600_, _22599_);
  or _73549_ (_22602_, _22601_, _06132_);
  and _73550_ (_22603_, _14928_, _07803_);
  or _73551_ (_22604_, _22603_, _22599_);
  or _73552_ (_22605_, _22604_, _06161_);
  and _73553_ (_22606_, _07803_, \oc8051_golden_model_1.ACC [4]);
  or _73554_ (_22607_, _22606_, _22599_);
  and _73555_ (_22608_, _22607_, _07056_);
  and _73556_ (_22611_, _07057_, \oc8051_golden_model_1.TL0 [4]);
  or _73557_ (_22612_, _22611_, _06160_);
  or _73558_ (_22613_, _22612_, _22608_);
  and _73559_ (_22614_, _22613_, _07075_);
  and _73560_ (_22615_, _22614_, _22605_);
  and _73561_ (_22616_, _22601_, _06217_);
  or _73562_ (_22617_, _22616_, _22615_);
  and _73563_ (_22618_, _22617_, _06229_);
  and _73564_ (_22619_, _22607_, _06220_);
  or _73565_ (_22620_, _22619_, _09842_);
  or _73566_ (_22622_, _22620_, _22618_);
  and _73567_ (_22623_, _22622_, _22602_);
  or _73568_ (_22624_, _22623_, _06116_);
  and _73569_ (_22625_, _09209_, _07803_);
  or _73570_ (_22626_, _22599_, _06117_);
  or _73571_ (_22627_, _22626_, _22625_);
  and _73572_ (_22628_, _22627_, _06114_);
  and _73573_ (_22629_, _22628_, _22624_);
  and _73574_ (_22630_, _15013_, _07803_);
  or _73575_ (_22631_, _22630_, _22599_);
  and _73576_ (_22633_, _22631_, _05787_);
  or _73577_ (_22634_, _22633_, _22629_);
  or _73578_ (_22635_, _22634_, _11136_);
  and _73579_ (_22636_, _15029_, _07803_);
  or _73580_ (_22637_, _22599_, _07127_);
  or _73581_ (_22638_, _22637_, _22636_);
  and _73582_ (_22639_, _08715_, _07803_);
  or _73583_ (_22640_, _22639_, _22599_);
  or _73584_ (_22641_, _22640_, _06111_);
  and _73585_ (_22642_, _22641_, _07125_);
  and _73586_ (_22644_, _22642_, _22638_);
  and _73587_ (_22645_, _22644_, _22635_);
  and _73588_ (_22646_, _10289_, _07803_);
  or _73589_ (_22647_, _22646_, _22599_);
  and _73590_ (_22648_, _22647_, _06402_);
  or _73591_ (_22649_, _22648_, _22645_);
  and _73592_ (_22650_, _22649_, _07132_);
  or _73593_ (_22651_, _22599_, _08339_);
  and _73594_ (_22652_, _22640_, _06306_);
  and _73595_ (_22653_, _22652_, _22651_);
  or _73596_ (_22655_, _22653_, _22650_);
  and _73597_ (_22656_, _22655_, _07130_);
  and _73598_ (_22657_, _22607_, _06411_);
  and _73599_ (_22658_, _22657_, _22651_);
  or _73600_ (_22659_, _22658_, _06303_);
  or _73601_ (_22660_, _22659_, _22656_);
  and _73602_ (_22661_, _15026_, _07803_);
  or _73603_ (_22662_, _22599_, _08819_);
  or _73604_ (_22663_, _22662_, _22661_);
  and _73605_ (_22664_, _22663_, _08824_);
  and _73606_ (_22666_, _22664_, _22660_);
  nor _73607_ (_22667_, _10288_, _11561_);
  or _73608_ (_22668_, _22667_, _22599_);
  and _73609_ (_22669_, _22668_, _06396_);
  or _73610_ (_22670_, _22669_, _06433_);
  or _73611_ (_22671_, _22670_, _22666_);
  or _73612_ (_22672_, _22604_, _06829_);
  and _73613_ (_22673_, _22672_, _06444_);
  and _73614_ (_22674_, _22673_, _22671_);
  and _73615_ (_22675_, _15087_, _07803_);
  or _73616_ (_22677_, _22675_, _22599_);
  and _73617_ (_22678_, _22677_, _06440_);
  or _73618_ (_22679_, _22678_, _01321_);
  or _73619_ (_22680_, _22679_, _22674_);
  or _73620_ (_22681_, _01317_, \oc8051_golden_model_1.TL0 [4]);
  and _73621_ (_22682_, _22681_, _43100_);
  and _73622_ (_43657_, _22682_, _22680_);
  and _73623_ (_22683_, _11561_, \oc8051_golden_model_1.TL0 [5]);
  or _73624_ (_22684_, _22683_, _08104_);
  and _73625_ (_22685_, _08736_, _07803_);
  or _73626_ (_22687_, _22685_, _22683_);
  and _73627_ (_22688_, _22687_, _06306_);
  and _73628_ (_22689_, _22688_, _22684_);
  and _73629_ (_22690_, _15119_, _07803_);
  or _73630_ (_22691_, _22690_, _22683_);
  or _73631_ (_22692_, _22691_, _06161_);
  and _73632_ (_22693_, _07803_, \oc8051_golden_model_1.ACC [5]);
  or _73633_ (_22694_, _22693_, _22683_);
  and _73634_ (_22695_, _22694_, _07056_);
  and _73635_ (_22696_, _07057_, \oc8051_golden_model_1.TL0 [5]);
  or _73636_ (_22698_, _22696_, _06160_);
  or _73637_ (_22699_, _22698_, _22695_);
  and _73638_ (_22700_, _22699_, _07075_);
  and _73639_ (_22701_, _22700_, _22692_);
  and _73640_ (_22702_, _08101_, _07803_);
  or _73641_ (_22703_, _22702_, _22683_);
  and _73642_ (_22704_, _22703_, _06217_);
  or _73643_ (_22705_, _22704_, _22701_);
  and _73644_ (_22706_, _22705_, _06229_);
  and _73645_ (_22707_, _22694_, _06220_);
  or _73646_ (_22708_, _22707_, _09842_);
  or _73647_ (_22709_, _22708_, _22706_);
  or _73648_ (_22710_, _22703_, _06132_);
  and _73649_ (_22711_, _22710_, _22709_);
  or _73650_ (_22712_, _22711_, _06116_);
  and _73651_ (_22713_, _09208_, _07803_);
  or _73652_ (_22714_, _22683_, _06117_);
  or _73653_ (_22715_, _22714_, _22713_);
  and _73654_ (_22716_, _22715_, _06114_);
  and _73655_ (_22717_, _22716_, _22712_);
  and _73656_ (_22720_, _15203_, _07803_);
  or _73657_ (_22721_, _22720_, _22683_);
  and _73658_ (_22722_, _22721_, _05787_);
  or _73659_ (_22723_, _22722_, _11136_);
  or _73660_ (_22724_, _22723_, _22717_);
  and _73661_ (_22725_, _15219_, _07803_);
  or _73662_ (_22726_, _22683_, _07127_);
  or _73663_ (_22727_, _22726_, _22725_);
  or _73664_ (_22728_, _22687_, _06111_);
  and _73665_ (_22729_, _22728_, _07125_);
  and _73666_ (_22731_, _22729_, _22727_);
  and _73667_ (_22732_, _22731_, _22724_);
  and _73668_ (_22733_, _12325_, _07803_);
  or _73669_ (_22734_, _22733_, _22683_);
  and _73670_ (_22735_, _22734_, _06402_);
  or _73671_ (_22736_, _22735_, _22732_);
  and _73672_ (_22737_, _22736_, _07132_);
  or _73673_ (_22738_, _22737_, _22689_);
  and _73674_ (_22739_, _22738_, _07130_);
  and _73675_ (_22740_, _22694_, _06411_);
  and _73676_ (_22742_, _22740_, _22684_);
  or _73677_ (_22743_, _22742_, _06303_);
  or _73678_ (_22744_, _22743_, _22739_);
  and _73679_ (_22745_, _15216_, _07803_);
  or _73680_ (_22746_, _22683_, _08819_);
  or _73681_ (_22747_, _22746_, _22745_);
  and _73682_ (_22748_, _22747_, _08824_);
  and _73683_ (_22749_, _22748_, _22744_);
  nor _73684_ (_22750_, _10269_, _11561_);
  or _73685_ (_22751_, _22750_, _22683_);
  and _73686_ (_22753_, _22751_, _06396_);
  or _73687_ (_22754_, _22753_, _06433_);
  or _73688_ (_22755_, _22754_, _22749_);
  or _73689_ (_22756_, _22691_, _06829_);
  and _73690_ (_22757_, _22756_, _06444_);
  and _73691_ (_22758_, _22757_, _22755_);
  and _73692_ (_22759_, _15275_, _07803_);
  or _73693_ (_22760_, _22759_, _22683_);
  and _73694_ (_22761_, _22760_, _06440_);
  or _73695_ (_22762_, _22761_, _01321_);
  or _73696_ (_22764_, _22762_, _22758_);
  or _73697_ (_22765_, _01317_, \oc8051_golden_model_1.TL0 [5]);
  and _73698_ (_22766_, _22765_, _43100_);
  and _73699_ (_43659_, _22766_, _22764_);
  and _73700_ (_22767_, _11561_, \oc8051_golden_model_1.TL0 [6]);
  or _73701_ (_22768_, _22767_, _08015_);
  and _73702_ (_22769_, _15402_, _07803_);
  or _73703_ (_22770_, _22769_, _22767_);
  and _73704_ (_22771_, _22770_, _06306_);
  and _73705_ (_22772_, _22771_, _22768_);
  and _73706_ (_22774_, _15300_, _07803_);
  or _73707_ (_22775_, _22774_, _22767_);
  or _73708_ (_22776_, _22775_, _06161_);
  and _73709_ (_22777_, _07803_, \oc8051_golden_model_1.ACC [6]);
  or _73710_ (_22778_, _22777_, _22767_);
  and _73711_ (_22779_, _22778_, _07056_);
  and _73712_ (_22780_, _07057_, \oc8051_golden_model_1.TL0 [6]);
  or _73713_ (_22781_, _22780_, _06160_);
  or _73714_ (_22782_, _22781_, _22779_);
  and _73715_ (_22783_, _22782_, _07075_);
  and _73716_ (_22785_, _22783_, _22776_);
  and _73717_ (_22786_, _08012_, _07803_);
  or _73718_ (_22787_, _22786_, _22767_);
  and _73719_ (_22788_, _22787_, _06217_);
  or _73720_ (_22789_, _22788_, _22785_);
  and _73721_ (_22790_, _22789_, _06229_);
  and _73722_ (_22791_, _22778_, _06220_);
  or _73723_ (_22792_, _22791_, _09842_);
  or _73724_ (_22793_, _22792_, _22790_);
  or _73725_ (_22794_, _22787_, _06132_);
  and _73726_ (_22796_, _22794_, _22793_);
  or _73727_ (_22797_, _22796_, _06116_);
  and _73728_ (_22798_, _09207_, _07803_);
  or _73729_ (_22799_, _22767_, _06117_);
  or _73730_ (_22800_, _22799_, _22798_);
  and _73731_ (_22801_, _22800_, _06114_);
  and _73732_ (_22802_, _22801_, _22797_);
  and _73733_ (_22803_, _15395_, _07803_);
  or _73734_ (_22804_, _22803_, _22767_);
  and _73735_ (_22805_, _22804_, _05787_);
  or _73736_ (_22807_, _22805_, _11136_);
  or _73737_ (_22808_, _22807_, _22802_);
  and _73738_ (_22809_, _15413_, _07803_);
  or _73739_ (_22810_, _22767_, _07127_);
  or _73740_ (_22811_, _22810_, _22809_);
  or _73741_ (_22812_, _22770_, _06111_);
  and _73742_ (_22813_, _22812_, _07125_);
  and _73743_ (_22814_, _22813_, _22811_);
  and _73744_ (_22815_, _22814_, _22808_);
  and _73745_ (_22816_, _10295_, _07803_);
  or _73746_ (_22818_, _22816_, _22767_);
  and _73747_ (_22819_, _22818_, _06402_);
  or _73748_ (_22820_, _22819_, _22815_);
  and _73749_ (_22821_, _22820_, _07132_);
  or _73750_ (_22822_, _22821_, _22772_);
  and _73751_ (_22823_, _22822_, _07130_);
  and _73752_ (_22824_, _22778_, _06411_);
  and _73753_ (_22825_, _22824_, _22768_);
  or _73754_ (_22826_, _22825_, _06303_);
  or _73755_ (_22827_, _22826_, _22823_);
  and _73756_ (_22829_, _15410_, _07803_);
  or _73757_ (_22830_, _22767_, _08819_);
  or _73758_ (_22831_, _22830_, _22829_);
  and _73759_ (_22832_, _22831_, _08824_);
  and _73760_ (_22833_, _22832_, _22827_);
  nor _73761_ (_22834_, _10294_, _11561_);
  or _73762_ (_22835_, _22834_, _22767_);
  and _73763_ (_22836_, _22835_, _06396_);
  or _73764_ (_22837_, _22836_, _06433_);
  or _73765_ (_22838_, _22837_, _22833_);
  or _73766_ (_22840_, _22775_, _06829_);
  and _73767_ (_22841_, _22840_, _06444_);
  and _73768_ (_22842_, _22841_, _22838_);
  and _73769_ (_22843_, _15478_, _07803_);
  or _73770_ (_22844_, _22843_, _22767_);
  and _73771_ (_22845_, _22844_, _06440_);
  or _73772_ (_22846_, _22845_, _01321_);
  or _73773_ (_22847_, _22846_, _22842_);
  or _73774_ (_22848_, _01317_, \oc8051_golden_model_1.TL0 [6]);
  and _73775_ (_22849_, _22848_, _43100_);
  and _73776_ (_43660_, _22849_, _22847_);
  not _73777_ (_22851_, \oc8051_golden_model_1.TCON [0]);
  nor _73778_ (_22852_, _01317_, _22851_);
  nand _73779_ (_22853_, _10276_, _07788_);
  nor _73780_ (_22854_, _07788_, _22851_);
  nor _73781_ (_22855_, _22854_, _07130_);
  nand _73782_ (_22856_, _22855_, _22853_);
  and _73783_ (_22857_, _07788_, _07049_);
  or _73784_ (_22858_, _22857_, _22854_);
  or _73785_ (_22859_, _22858_, _06132_);
  nor _73786_ (_22861_, _08211_, _11639_);
  or _73787_ (_22862_, _22861_, _22854_);
  or _73788_ (_22863_, _22862_, _06161_);
  and _73789_ (_22864_, _07788_, \oc8051_golden_model_1.ACC [0]);
  or _73790_ (_22865_, _22864_, _22854_);
  and _73791_ (_22866_, _22865_, _07056_);
  nor _73792_ (_22867_, _07056_, _22851_);
  or _73793_ (_22868_, _22867_, _06160_);
  or _73794_ (_22869_, _22868_, _22866_);
  and _73795_ (_22870_, _22869_, _06157_);
  and _73796_ (_22872_, _22870_, _22863_);
  nor _73797_ (_22873_, _08407_, _22851_);
  and _73798_ (_22874_, _14169_, _08407_);
  or _73799_ (_22875_, _22874_, _22873_);
  and _73800_ (_22876_, _22875_, _06156_);
  or _73801_ (_22877_, _22876_, _22872_);
  and _73802_ (_22878_, _22877_, _07075_);
  and _73803_ (_22879_, _22858_, _06217_);
  or _73804_ (_22880_, _22879_, _06220_);
  or _73805_ (_22881_, _22880_, _22878_);
  or _73806_ (_22883_, _22865_, _06229_);
  and _73807_ (_22884_, _22883_, _06153_);
  and _73808_ (_22885_, _22884_, _22881_);
  and _73809_ (_22886_, _22854_, _06152_);
  or _73810_ (_22887_, _22886_, _06145_);
  or _73811_ (_22888_, _22887_, _22885_);
  or _73812_ (_22889_, _22862_, _06146_);
  and _73813_ (_22890_, _22889_, _06140_);
  and _73814_ (_22891_, _22890_, _22888_);
  or _73815_ (_22892_, _22873_, _14170_);
  and _73816_ (_22894_, _22892_, _06139_);
  and _73817_ (_22895_, _22894_, _22875_);
  or _73818_ (_22896_, _22895_, _09842_);
  or _73819_ (_22897_, _22896_, _22891_);
  and _73820_ (_22898_, _22897_, _22859_);
  or _73821_ (_22899_, _22898_, _06116_);
  and _73822_ (_22900_, _09160_, _07788_);
  or _73823_ (_22901_, _22854_, _06117_);
  or _73824_ (_22902_, _22901_, _22900_);
  and _73825_ (_22903_, _22902_, _06114_);
  and _73826_ (_22905_, _22903_, _22899_);
  and _73827_ (_22906_, _14260_, _07788_);
  or _73828_ (_22907_, _22906_, _22854_);
  and _73829_ (_22908_, _22907_, _05787_);
  or _73830_ (_22909_, _22908_, _22905_);
  or _73831_ (_22910_, _22909_, _11136_);
  and _73832_ (_22911_, _14275_, _07788_);
  or _73833_ (_22912_, _22854_, _07127_);
  or _73834_ (_22913_, _22912_, _22911_);
  and _73835_ (_22914_, _07788_, _08708_);
  or _73836_ (_22916_, _22914_, _22854_);
  or _73837_ (_22917_, _22916_, _06111_);
  and _73838_ (_22918_, _22917_, _07125_);
  and _73839_ (_22919_, _22918_, _22913_);
  and _73840_ (_22920_, _22919_, _22910_);
  nor _73841_ (_22921_, _12321_, _11639_);
  or _73842_ (_22922_, _22921_, _22854_);
  and _73843_ (_22923_, _22853_, _06402_);
  and _73844_ (_22924_, _22923_, _22922_);
  or _73845_ (_22925_, _22924_, _22920_);
  and _73846_ (_22926_, _22925_, _07132_);
  nand _73847_ (_22927_, _22916_, _06306_);
  nor _73848_ (_22928_, _22927_, _22861_);
  or _73849_ (_22929_, _22928_, _06411_);
  or _73850_ (_22930_, _22929_, _22926_);
  and _73851_ (_22931_, _22930_, _22856_);
  or _73852_ (_22932_, _22931_, _06303_);
  and _73853_ (_22933_, _14167_, _07788_);
  or _73854_ (_22934_, _22854_, _08819_);
  or _73855_ (_22935_, _22934_, _22933_);
  and _73856_ (_22938_, _22935_, _08824_);
  and _73857_ (_22939_, _22938_, _22932_);
  and _73858_ (_22940_, _22922_, _06396_);
  or _73859_ (_22941_, _22940_, _06433_);
  or _73860_ (_22942_, _22941_, _22939_);
  or _73861_ (_22943_, _22862_, _06829_);
  and _73862_ (_22944_, _22943_, _22942_);
  or _73863_ (_22945_, _22944_, _05748_);
  or _73864_ (_22946_, _22854_, _05749_);
  and _73865_ (_22947_, _22946_, _22945_);
  or _73866_ (_22949_, _22947_, _06440_);
  or _73867_ (_22950_, _22862_, _06444_);
  and _73868_ (_22951_, _22950_, _01317_);
  and _73869_ (_22952_, _22951_, _22949_);
  or _73870_ (_22953_, _22952_, _22852_);
  and _73871_ (_43661_, _22953_, _43100_);
  and _73872_ (_22954_, _01321_, \oc8051_golden_model_1.TCON [1]);
  and _73873_ (_22955_, _11639_, \oc8051_golden_model_1.TCON [1]);
  nor _73874_ (_22956_, _10277_, _11639_);
  or _73875_ (_22957_, _22956_, _22955_);
  or _73876_ (_22959_, _22957_, _08824_);
  or _73877_ (_22960_, _14442_, _11639_);
  or _73878_ (_22961_, _07788_, \oc8051_golden_model_1.TCON [1]);
  and _73879_ (_22962_, _22961_, _05787_);
  and _73880_ (_22963_, _22962_, _22960_);
  and _73881_ (_22964_, _07788_, _07306_);
  or _73882_ (_22965_, _22964_, _22955_);
  or _73883_ (_22966_, _22965_, _07075_);
  and _73884_ (_22967_, _14363_, _07788_);
  not _73885_ (_22968_, _22967_);
  and _73886_ (_22970_, _22968_, _22961_);
  or _73887_ (_22971_, _22970_, _06161_);
  and _73888_ (_22972_, _07788_, \oc8051_golden_model_1.ACC [1]);
  or _73889_ (_22973_, _22972_, _22955_);
  and _73890_ (_22974_, _22973_, _07056_);
  and _73891_ (_22975_, _07057_, \oc8051_golden_model_1.TCON [1]);
  or _73892_ (_22976_, _22975_, _06160_);
  or _73893_ (_22977_, _22976_, _22974_);
  and _73894_ (_22978_, _22977_, _06157_);
  and _73895_ (_22979_, _22978_, _22971_);
  and _73896_ (_22981_, _11644_, \oc8051_golden_model_1.TCON [1]);
  and _73897_ (_22982_, _14367_, _08407_);
  or _73898_ (_22983_, _22982_, _22981_);
  and _73899_ (_22984_, _22983_, _06156_);
  or _73900_ (_22985_, _22984_, _06217_);
  or _73901_ (_22986_, _22985_, _22979_);
  and _73902_ (_22987_, _22986_, _22966_);
  or _73903_ (_22988_, _22987_, _06220_);
  or _73904_ (_22989_, _22973_, _06229_);
  and _73905_ (_22990_, _22989_, _06153_);
  and _73906_ (_22992_, _22990_, _22988_);
  and _73907_ (_22993_, _14349_, _08407_);
  or _73908_ (_22994_, _22993_, _22981_);
  and _73909_ (_22995_, _22994_, _06152_);
  or _73910_ (_22996_, _22995_, _06145_);
  or _73911_ (_22997_, _22996_, _22992_);
  and _73912_ (_22998_, _22982_, _14382_);
  or _73913_ (_22999_, _22981_, _06146_);
  or _73914_ (_23000_, _22999_, _22998_);
  and _73915_ (_23001_, _23000_, _22997_);
  and _73916_ (_23003_, _23001_, _06140_);
  and _73917_ (_23004_, _14351_, _08407_);
  or _73918_ (_23005_, _22981_, _23004_);
  and _73919_ (_23006_, _23005_, _06139_);
  or _73920_ (_23007_, _23006_, _09842_);
  or _73921_ (_23008_, _23007_, _23003_);
  or _73922_ (_23009_, _22965_, _06132_);
  and _73923_ (_23010_, _23009_, _23008_);
  or _73924_ (_23011_, _23010_, _06116_);
  and _73925_ (_23012_, _09115_, _07788_);
  or _73926_ (_23014_, _22955_, _06117_);
  or _73927_ (_23015_, _23014_, _23012_);
  and _73928_ (_23016_, _23015_, _06114_);
  and _73929_ (_23017_, _23016_, _23011_);
  or _73930_ (_23018_, _23017_, _22963_);
  and _73931_ (_23019_, _23018_, _06298_);
  or _73932_ (_23020_, _14346_, _11639_);
  and _73933_ (_23021_, _23020_, _06297_);
  nand _73934_ (_23022_, _07788_, _06945_);
  and _73935_ (_23023_, _23022_, _06110_);
  or _73936_ (_23025_, _23023_, _23021_);
  and _73937_ (_23026_, _23025_, _22961_);
  or _73938_ (_23027_, _23026_, _06402_);
  or _73939_ (_23028_, _23027_, _23019_);
  and _73940_ (_23029_, _10278_, _07788_);
  or _73941_ (_23030_, _23029_, _22955_);
  or _73942_ (_23031_, _23030_, _07125_);
  and _73943_ (_23032_, _23031_, _07132_);
  and _73944_ (_23033_, _23032_, _23028_);
  or _73945_ (_23034_, _14344_, _11639_);
  and _73946_ (_23036_, _22961_, _06306_);
  and _73947_ (_23037_, _23036_, _23034_);
  or _73948_ (_23038_, _23037_, _06411_);
  or _73949_ (_23039_, _23038_, _23033_);
  and _73950_ (_23040_, _22972_, _08176_);
  or _73951_ (_23041_, _22955_, _07130_);
  or _73952_ (_23042_, _23041_, _23040_);
  and _73953_ (_23043_, _23042_, _08819_);
  and _73954_ (_23044_, _23043_, _23039_);
  or _73955_ (_23045_, _23022_, _08176_);
  and _73956_ (_23046_, _22961_, _06303_);
  and _73957_ (_23047_, _23046_, _23045_);
  or _73958_ (_23048_, _23047_, _06396_);
  or _73959_ (_23049_, _23048_, _23044_);
  and _73960_ (_23050_, _23049_, _22959_);
  or _73961_ (_23051_, _23050_, _06433_);
  or _73962_ (_23052_, _22970_, _06829_);
  and _73963_ (_23053_, _23052_, _05749_);
  and _73964_ (_23054_, _23053_, _23051_);
  and _73965_ (_23055_, _22994_, _05748_);
  or _73966_ (_23057_, _23055_, _06440_);
  or _73967_ (_23058_, _23057_, _23054_);
  or _73968_ (_23059_, _22955_, _06444_);
  or _73969_ (_23060_, _23059_, _22967_);
  and _73970_ (_23061_, _23060_, _01317_);
  and _73971_ (_23062_, _23061_, _23058_);
  or _73972_ (_23063_, _23062_, _22954_);
  and _73973_ (_43663_, _23063_, _43100_);
  and _73974_ (_23064_, _01321_, \oc8051_golden_model_1.TCON [2]);
  and _73975_ (_23065_, _11639_, \oc8051_golden_model_1.TCON [2]);
  and _73976_ (_23067_, _07788_, _07708_);
  or _73977_ (_23068_, _23067_, _23065_);
  or _73978_ (_23069_, _23068_, _06132_);
  or _73979_ (_23070_, _23068_, _07075_);
  and _73980_ (_23071_, _14542_, _07788_);
  or _73981_ (_23072_, _23071_, _23065_);
  or _73982_ (_23073_, _23072_, _06161_);
  and _73983_ (_23074_, _07788_, \oc8051_golden_model_1.ACC [2]);
  or _73984_ (_23075_, _23074_, _23065_);
  and _73985_ (_23076_, _23075_, _07056_);
  and _73986_ (_23078_, _07057_, \oc8051_golden_model_1.TCON [2]);
  or _73987_ (_23079_, _23078_, _06160_);
  or _73988_ (_23080_, _23079_, _23076_);
  and _73989_ (_23081_, _23080_, _06157_);
  and _73990_ (_23082_, _23081_, _23073_);
  and _73991_ (_23083_, _11644_, \oc8051_golden_model_1.TCON [2]);
  and _73992_ (_23084_, _14538_, _08407_);
  or _73993_ (_23085_, _23084_, _23083_);
  and _73994_ (_23086_, _23085_, _06156_);
  or _73995_ (_23087_, _23086_, _06217_);
  or _73996_ (_23088_, _23087_, _23082_);
  and _73997_ (_23089_, _23088_, _23070_);
  or _73998_ (_23090_, _23089_, _06220_);
  or _73999_ (_23091_, _23075_, _06229_);
  and _74000_ (_23092_, _23091_, _06153_);
  and _74001_ (_23093_, _23092_, _23090_);
  and _74002_ (_23094_, _14536_, _08407_);
  or _74003_ (_23095_, _23094_, _23083_);
  and _74004_ (_23096_, _23095_, _06152_);
  or _74005_ (_23097_, _23096_, _06145_);
  or _74006_ (_23099_, _23097_, _23093_);
  and _74007_ (_23100_, _23084_, _14569_);
  or _74008_ (_23101_, _23083_, _06146_);
  or _74009_ (_23102_, _23101_, _23100_);
  and _74010_ (_23103_, _23102_, _06140_);
  and _74011_ (_23104_, _23103_, _23099_);
  and _74012_ (_23105_, _14583_, _08407_);
  or _74013_ (_23106_, _23105_, _23083_);
  and _74014_ (_23107_, _23106_, _06139_);
  or _74015_ (_23108_, _23107_, _09842_);
  or _74016_ (_23109_, _23108_, _23104_);
  and _74017_ (_23110_, _23109_, _23069_);
  or _74018_ (_23111_, _23110_, _06116_);
  and _74019_ (_23112_, _09211_, _07788_);
  or _74020_ (_23113_, _23065_, _06117_);
  or _74021_ (_23114_, _23113_, _23112_);
  and _74022_ (_23115_, _23114_, _06114_);
  and _74023_ (_23116_, _23115_, _23111_);
  and _74024_ (_23117_, _14630_, _07788_);
  or _74025_ (_23118_, _23065_, _23117_);
  and _74026_ (_23120_, _23118_, _05787_);
  or _74027_ (_23121_, _23120_, _23116_);
  or _74028_ (_23122_, _23121_, _11136_);
  and _74029_ (_23123_, _14646_, _07788_);
  or _74030_ (_23124_, _23065_, _07127_);
  or _74031_ (_23125_, _23124_, _23123_);
  and _74032_ (_23126_, _07788_, _08768_);
  or _74033_ (_23127_, _23126_, _23065_);
  or _74034_ (_23128_, _23127_, _06111_);
  and _74035_ (_23129_, _23128_, _07125_);
  and _74036_ (_23131_, _23129_, _23125_);
  and _74037_ (_23132_, _23131_, _23122_);
  and _74038_ (_23133_, _10282_, _07788_);
  or _74039_ (_23134_, _23133_, _23065_);
  and _74040_ (_23135_, _23134_, _06402_);
  or _74041_ (_23136_, _23135_, _23132_);
  and _74042_ (_23137_, _23136_, _07132_);
  or _74043_ (_23138_, _23065_, _08248_);
  and _74044_ (_23139_, _23127_, _06306_);
  and _74045_ (_23140_, _23139_, _23138_);
  or _74046_ (_23141_, _23140_, _23137_);
  and _74047_ (_23142_, _23141_, _07130_);
  and _74048_ (_23143_, _23075_, _06411_);
  and _74049_ (_23144_, _23143_, _23138_);
  or _74050_ (_23145_, _23144_, _06303_);
  or _74051_ (_23146_, _23145_, _23142_);
  and _74052_ (_23147_, _14643_, _07788_);
  or _74053_ (_23148_, _23065_, _08819_);
  or _74054_ (_23149_, _23148_, _23147_);
  and _74055_ (_23150_, _23149_, _08824_);
  and _74056_ (_23152_, _23150_, _23146_);
  nor _74057_ (_23153_, _10281_, _11639_);
  or _74058_ (_23154_, _23153_, _23065_);
  and _74059_ (_23155_, _23154_, _06396_);
  or _74060_ (_23156_, _23155_, _06433_);
  or _74061_ (_23157_, _23156_, _23152_);
  or _74062_ (_23158_, _23072_, _06829_);
  and _74063_ (_23159_, _23158_, _05749_);
  and _74064_ (_23160_, _23159_, _23157_);
  and _74065_ (_23161_, _23095_, _05748_);
  or _74066_ (_23163_, _23161_, _06440_);
  or _74067_ (_23164_, _23163_, _23160_);
  and _74068_ (_23165_, _14710_, _07788_);
  or _74069_ (_23166_, _23065_, _06444_);
  or _74070_ (_23167_, _23166_, _23165_);
  and _74071_ (_23168_, _23167_, _01317_);
  and _74072_ (_23169_, _23168_, _23164_);
  or _74073_ (_23170_, _23169_, _23064_);
  and _74074_ (_43664_, _23170_, _43100_);
  and _74075_ (_23171_, _01321_, \oc8051_golden_model_1.TCON [3]);
  and _74076_ (_23172_, _11639_, \oc8051_golden_model_1.TCON [3]);
  and _74077_ (_23173_, _07788_, _07544_);
  or _74078_ (_23174_, _23173_, _23172_);
  or _74079_ (_23175_, _23174_, _06132_);
  and _74080_ (_23176_, _14738_, _07788_);
  or _74081_ (_23177_, _23176_, _23172_);
  or _74082_ (_23178_, _23177_, _06161_);
  and _74083_ (_23179_, _07788_, \oc8051_golden_model_1.ACC [3]);
  or _74084_ (_23180_, _23179_, _23172_);
  and _74085_ (_23181_, _23180_, _07056_);
  and _74086_ (_23182_, _07057_, \oc8051_golden_model_1.TCON [3]);
  or _74087_ (_23183_, _23182_, _06160_);
  or _74088_ (_23184_, _23183_, _23181_);
  and _74089_ (_23185_, _23184_, _06157_);
  and _74090_ (_23186_, _23185_, _23178_);
  and _74091_ (_23187_, _11644_, \oc8051_golden_model_1.TCON [3]);
  and _74092_ (_23188_, _14735_, _08407_);
  or _74093_ (_23189_, _23188_, _23187_);
  and _74094_ (_23190_, _23189_, _06156_);
  or _74095_ (_23191_, _23190_, _06217_);
  or _74096_ (_23194_, _23191_, _23186_);
  or _74097_ (_23195_, _23174_, _07075_);
  and _74098_ (_23196_, _23195_, _23194_);
  or _74099_ (_23197_, _23196_, _06220_);
  or _74100_ (_23198_, _23180_, _06229_);
  and _74101_ (_23199_, _23198_, _06153_);
  and _74102_ (_23200_, _23199_, _23197_);
  and _74103_ (_23201_, _14731_, _08407_);
  or _74104_ (_23202_, _23201_, _23187_);
  and _74105_ (_23203_, _23202_, _06152_);
  or _74106_ (_23204_, _23203_, _06145_);
  or _74107_ (_23205_, _23204_, _23200_);
  or _74108_ (_23206_, _23187_, _14764_);
  and _74109_ (_23207_, _23206_, _23189_);
  or _74110_ (_23208_, _23207_, _06146_);
  and _74111_ (_23209_, _23208_, _06140_);
  and _74112_ (_23210_, _23209_, _23205_);
  and _74113_ (_23211_, _14732_, _08407_);
  or _74114_ (_23212_, _23211_, _23187_);
  and _74115_ (_23213_, _23212_, _06139_);
  or _74116_ (_23215_, _23213_, _09842_);
  or _74117_ (_23216_, _23215_, _23210_);
  and _74118_ (_23217_, _23216_, _23175_);
  or _74119_ (_23218_, _23217_, _06116_);
  and _74120_ (_23219_, _09210_, _07788_);
  or _74121_ (_23220_, _23172_, _06117_);
  or _74122_ (_23221_, _23220_, _23219_);
  and _74123_ (_23222_, _23221_, _06114_);
  and _74124_ (_23223_, _23222_, _23218_);
  and _74125_ (_23224_, _14825_, _07788_);
  or _74126_ (_23226_, _23172_, _23224_);
  and _74127_ (_23227_, _23226_, _05787_);
  or _74128_ (_23228_, _23227_, _23223_);
  or _74129_ (_23229_, _23228_, _11136_);
  and _74130_ (_23230_, _14727_, _07788_);
  or _74131_ (_23231_, _23172_, _07127_);
  or _74132_ (_23232_, _23231_, _23230_);
  and _74133_ (_23233_, _07788_, _08712_);
  or _74134_ (_23234_, _23233_, _23172_);
  or _74135_ (_23235_, _23234_, _06111_);
  and _74136_ (_23236_, _23235_, _07125_);
  and _74137_ (_23237_, _23236_, _23232_);
  and _74138_ (_23238_, _23237_, _23229_);
  and _74139_ (_23239_, _12318_, _07788_);
  or _74140_ (_23240_, _23239_, _23172_);
  and _74141_ (_23241_, _23240_, _06402_);
  or _74142_ (_23242_, _23241_, _23238_);
  and _74143_ (_23243_, _23242_, _07132_);
  or _74144_ (_23244_, _23172_, _08140_);
  and _74145_ (_23245_, _23234_, _06306_);
  and _74146_ (_23247_, _23245_, _23244_);
  or _74147_ (_23248_, _23247_, _23243_);
  and _74148_ (_23249_, _23248_, _07130_);
  and _74149_ (_23250_, _23180_, _06411_);
  and _74150_ (_23251_, _23250_, _23244_);
  or _74151_ (_23252_, _23251_, _06303_);
  or _74152_ (_23253_, _23252_, _23249_);
  and _74153_ (_23254_, _14724_, _07788_);
  or _74154_ (_23255_, _23172_, _08819_);
  or _74155_ (_23256_, _23255_, _23254_);
  and _74156_ (_23258_, _23256_, _08824_);
  and _74157_ (_23259_, _23258_, _23253_);
  nor _74158_ (_23260_, _10273_, _11639_);
  or _74159_ (_23261_, _23260_, _23172_);
  and _74160_ (_23262_, _23261_, _06396_);
  or _74161_ (_23263_, _23262_, _06433_);
  or _74162_ (_23264_, _23263_, _23259_);
  or _74163_ (_23265_, _23177_, _06829_);
  and _74164_ (_23266_, _23265_, _05749_);
  and _74165_ (_23267_, _23266_, _23264_);
  and _74166_ (_23268_, _23202_, _05748_);
  or _74167_ (_23269_, _23268_, _06440_);
  or _74168_ (_23270_, _23269_, _23267_);
  and _74169_ (_23271_, _14897_, _07788_);
  or _74170_ (_23272_, _23172_, _06444_);
  or _74171_ (_23273_, _23272_, _23271_);
  and _74172_ (_23274_, _23273_, _01317_);
  and _74173_ (_23275_, _23274_, _23270_);
  or _74174_ (_23276_, _23275_, _23171_);
  and _74175_ (_43665_, _23276_, _43100_);
  and _74176_ (_23278_, _01321_, \oc8051_golden_model_1.TCON [4]);
  and _74177_ (_23279_, _11639_, \oc8051_golden_model_1.TCON [4]);
  and _74178_ (_23280_, _08336_, _07788_);
  or _74179_ (_23281_, _23280_, _23279_);
  or _74180_ (_23282_, _23281_, _06132_);
  and _74181_ (_23283_, _11644_, \oc8051_golden_model_1.TCON [4]);
  and _74182_ (_23284_, _14942_, _08407_);
  or _74183_ (_23285_, _23284_, _23283_);
  and _74184_ (_23286_, _23285_, _06152_);
  and _74185_ (_23287_, _14928_, _07788_);
  or _74186_ (_23289_, _23287_, _23279_);
  or _74187_ (_23290_, _23289_, _06161_);
  and _74188_ (_23291_, _07788_, \oc8051_golden_model_1.ACC [4]);
  or _74189_ (_23292_, _23291_, _23279_);
  and _74190_ (_23293_, _23292_, _07056_);
  and _74191_ (_23294_, _07057_, \oc8051_golden_model_1.TCON [4]);
  or _74192_ (_23295_, _23294_, _06160_);
  or _74193_ (_23296_, _23295_, _23293_);
  and _74194_ (_23297_, _23296_, _06157_);
  and _74195_ (_23298_, _23297_, _23290_);
  and _74196_ (_23299_, _14932_, _08407_);
  or _74197_ (_23300_, _23299_, _23283_);
  and _74198_ (_23301_, _23300_, _06156_);
  or _74199_ (_23302_, _23301_, _06217_);
  or _74200_ (_23303_, _23302_, _23298_);
  or _74201_ (_23304_, _23281_, _07075_);
  and _74202_ (_23305_, _23304_, _23303_);
  or _74203_ (_23306_, _23305_, _06220_);
  or _74204_ (_23307_, _23292_, _06229_);
  and _74205_ (_23308_, _23307_, _06153_);
  and _74206_ (_23310_, _23308_, _23306_);
  or _74207_ (_23311_, _23310_, _23286_);
  and _74208_ (_23312_, _23311_, _06146_);
  and _74209_ (_23313_, _14950_, _08407_);
  or _74210_ (_23314_, _23313_, _23283_);
  and _74211_ (_23315_, _23314_, _06145_);
  or _74212_ (_23316_, _23315_, _23312_);
  and _74213_ (_23317_, _23316_, _06140_);
  and _74214_ (_23318_, _14966_, _08407_);
  or _74215_ (_23319_, _23318_, _23283_);
  and _74216_ (_23321_, _23319_, _06139_);
  or _74217_ (_23322_, _23321_, _09842_);
  or _74218_ (_23323_, _23322_, _23317_);
  and _74219_ (_23324_, _23323_, _23282_);
  or _74220_ (_23325_, _23324_, _06116_);
  and _74221_ (_23326_, _09209_, _07788_);
  or _74222_ (_23327_, _23279_, _06117_);
  or _74223_ (_23328_, _23327_, _23326_);
  and _74224_ (_23329_, _23328_, _06114_);
  and _74225_ (_23330_, _23329_, _23325_);
  and _74226_ (_23331_, _15013_, _07788_);
  or _74227_ (_23332_, _23331_, _23279_);
  and _74228_ (_23333_, _23332_, _05787_);
  or _74229_ (_23334_, _23333_, _11136_);
  or _74230_ (_23335_, _23334_, _23330_);
  and _74231_ (_23336_, _15029_, _07788_);
  or _74232_ (_23337_, _23279_, _07127_);
  or _74233_ (_23338_, _23337_, _23336_);
  and _74234_ (_23339_, _08715_, _07788_);
  or _74235_ (_23340_, _23339_, _23279_);
  or _74236_ (_23342_, _23340_, _06111_);
  and _74237_ (_23343_, _23342_, _07125_);
  and _74238_ (_23344_, _23343_, _23338_);
  and _74239_ (_23345_, _23344_, _23335_);
  and _74240_ (_23346_, _10289_, _07788_);
  or _74241_ (_23347_, _23346_, _23279_);
  and _74242_ (_23348_, _23347_, _06402_);
  or _74243_ (_23349_, _23348_, _23345_);
  and _74244_ (_23350_, _23349_, _07132_);
  or _74245_ (_23351_, _23279_, _08339_);
  and _74246_ (_23353_, _23340_, _06306_);
  and _74247_ (_23354_, _23353_, _23351_);
  or _74248_ (_23355_, _23354_, _23350_);
  and _74249_ (_23356_, _23355_, _07130_);
  and _74250_ (_23357_, _23292_, _06411_);
  and _74251_ (_23358_, _23357_, _23351_);
  or _74252_ (_23359_, _23358_, _06303_);
  or _74253_ (_23360_, _23359_, _23356_);
  and _74254_ (_23361_, _15026_, _07788_);
  or _74255_ (_23362_, _23279_, _08819_);
  or _74256_ (_23363_, _23362_, _23361_);
  and _74257_ (_23364_, _23363_, _08824_);
  and _74258_ (_23365_, _23364_, _23360_);
  nor _74259_ (_23366_, _10288_, _11639_);
  or _74260_ (_23367_, _23366_, _23279_);
  and _74261_ (_23368_, _23367_, _06396_);
  or _74262_ (_23369_, _23368_, _06433_);
  or _74263_ (_23370_, _23369_, _23365_);
  or _74264_ (_23371_, _23289_, _06829_);
  and _74265_ (_23372_, _23371_, _05749_);
  and _74266_ (_23374_, _23372_, _23370_);
  and _74267_ (_23375_, _23285_, _05748_);
  or _74268_ (_23376_, _23375_, _06440_);
  or _74269_ (_23377_, _23376_, _23374_);
  and _74270_ (_23378_, _15087_, _07788_);
  or _74271_ (_23379_, _23279_, _06444_);
  or _74272_ (_23380_, _23379_, _23378_);
  and _74273_ (_23381_, _23380_, _01317_);
  and _74274_ (_23382_, _23381_, _23377_);
  or _74275_ (_23383_, _23382_, _23278_);
  and _74276_ (_43666_, _23383_, _43100_);
  and _74277_ (_23385_, _01321_, \oc8051_golden_model_1.TCON [5]);
  and _74278_ (_23386_, _11639_, \oc8051_golden_model_1.TCON [5]);
  and _74279_ (_23387_, _15119_, _07788_);
  or _74280_ (_23388_, _23387_, _23386_);
  or _74281_ (_23389_, _23388_, _06161_);
  and _74282_ (_23390_, _07788_, \oc8051_golden_model_1.ACC [5]);
  or _74283_ (_23391_, _23390_, _23386_);
  and _74284_ (_23392_, _23391_, _07056_);
  and _74285_ (_23393_, _07057_, \oc8051_golden_model_1.TCON [5]);
  or _74286_ (_23394_, _23393_, _06160_);
  or _74287_ (_23395_, _23394_, _23392_);
  and _74288_ (_23396_, _23395_, _06157_);
  and _74289_ (_23397_, _23396_, _23389_);
  and _74290_ (_23398_, _11644_, \oc8051_golden_model_1.TCON [5]);
  and _74291_ (_23399_, _15123_, _08407_);
  or _74292_ (_23400_, _23399_, _23398_);
  and _74293_ (_23401_, _23400_, _06156_);
  or _74294_ (_23402_, _23401_, _06217_);
  or _74295_ (_23403_, _23402_, _23397_);
  and _74296_ (_23405_, _08101_, _07788_);
  or _74297_ (_23406_, _23405_, _23386_);
  or _74298_ (_23407_, _23406_, _07075_);
  and _74299_ (_23408_, _23407_, _23403_);
  or _74300_ (_23409_, _23408_, _06220_);
  or _74301_ (_23410_, _23391_, _06229_);
  and _74302_ (_23411_, _23410_, _06153_);
  and _74303_ (_23412_, _23411_, _23409_);
  and _74304_ (_23413_, _15104_, _08407_);
  or _74305_ (_23414_, _23413_, _23398_);
  and _74306_ (_23416_, _23414_, _06152_);
  or _74307_ (_23417_, _23416_, _06145_);
  or _74308_ (_23418_, _23417_, _23412_);
  or _74309_ (_23419_, _23398_, _15138_);
  and _74310_ (_23420_, _23419_, _23400_);
  or _74311_ (_23421_, _23420_, _06146_);
  and _74312_ (_23422_, _23421_, _06140_);
  and _74313_ (_23423_, _23422_, _23418_);
  and _74314_ (_23424_, _15155_, _08407_);
  or _74315_ (_23425_, _23424_, _23398_);
  and _74316_ (_23426_, _23425_, _06139_);
  or _74317_ (_23427_, _23426_, _09842_);
  or _74318_ (_23428_, _23427_, _23423_);
  or _74319_ (_23429_, _23406_, _06132_);
  and _74320_ (_23430_, _23429_, _23428_);
  or _74321_ (_23431_, _23430_, _06116_);
  and _74322_ (_23432_, _09208_, _07788_);
  or _74323_ (_23433_, _23386_, _06117_);
  or _74324_ (_23434_, _23433_, _23432_);
  and _74325_ (_23435_, _23434_, _06114_);
  and _74326_ (_23437_, _23435_, _23431_);
  and _74327_ (_23438_, _15203_, _07788_);
  or _74328_ (_23439_, _23438_, _23386_);
  and _74329_ (_23440_, _23439_, _05787_);
  or _74330_ (_23441_, _23440_, _11136_);
  or _74331_ (_23442_, _23441_, _23437_);
  and _74332_ (_23443_, _15219_, _07788_);
  or _74333_ (_23444_, _23386_, _07127_);
  or _74334_ (_23445_, _23444_, _23443_);
  and _74335_ (_23446_, _08736_, _07788_);
  or _74336_ (_23448_, _23446_, _23386_);
  or _74337_ (_23449_, _23448_, _06111_);
  and _74338_ (_23450_, _23449_, _07125_);
  and _74339_ (_23451_, _23450_, _23445_);
  and _74340_ (_23452_, _23451_, _23442_);
  and _74341_ (_23453_, _12325_, _07788_);
  or _74342_ (_23454_, _23453_, _23386_);
  and _74343_ (_23455_, _23454_, _06402_);
  or _74344_ (_23456_, _23455_, _23452_);
  and _74345_ (_23457_, _23456_, _07132_);
  or _74346_ (_23458_, _23386_, _08104_);
  and _74347_ (_23459_, _23448_, _06306_);
  and _74348_ (_23460_, _23459_, _23458_);
  or _74349_ (_23461_, _23460_, _23457_);
  and _74350_ (_23462_, _23461_, _07130_);
  and _74351_ (_23463_, _23391_, _06411_);
  and _74352_ (_23464_, _23463_, _23458_);
  or _74353_ (_23465_, _23464_, _06303_);
  or _74354_ (_23466_, _23465_, _23462_);
  and _74355_ (_23467_, _15216_, _07788_);
  or _74356_ (_23469_, _23386_, _08819_);
  or _74357_ (_23470_, _23469_, _23467_);
  and _74358_ (_23471_, _23470_, _08824_);
  and _74359_ (_23472_, _23471_, _23466_);
  nor _74360_ (_23473_, _10269_, _11639_);
  or _74361_ (_23474_, _23473_, _23386_);
  and _74362_ (_23475_, _23474_, _06396_);
  or _74363_ (_23476_, _23475_, _06433_);
  or _74364_ (_23477_, _23476_, _23472_);
  or _74365_ (_23478_, _23388_, _06829_);
  and _74366_ (_23480_, _23478_, _05749_);
  and _74367_ (_23481_, _23480_, _23477_);
  and _74368_ (_23482_, _23414_, _05748_);
  or _74369_ (_23483_, _23482_, _06440_);
  or _74370_ (_23484_, _23483_, _23481_);
  and _74371_ (_23485_, _15275_, _07788_);
  or _74372_ (_23486_, _23386_, _06444_);
  or _74373_ (_23487_, _23486_, _23485_);
  and _74374_ (_23488_, _23487_, _01317_);
  and _74375_ (_23489_, _23488_, _23484_);
  or _74376_ (_23491_, _23489_, _23385_);
  and _74377_ (_43667_, _23491_, _43100_);
  and _74378_ (_23492_, _01321_, \oc8051_golden_model_1.TCON [6]);
  and _74379_ (_23493_, _11639_, \oc8051_golden_model_1.TCON [6]);
  and _74380_ (_23494_, _15300_, _07788_);
  or _74381_ (_23495_, _23494_, _23493_);
  or _74382_ (_23496_, _23495_, _06161_);
  and _74383_ (_23497_, _07788_, \oc8051_golden_model_1.ACC [6]);
  or _74384_ (_23498_, _23497_, _23493_);
  and _74385_ (_23499_, _23498_, _07056_);
  and _74386_ (_23500_, _07057_, \oc8051_golden_model_1.TCON [6]);
  or _74387_ (_23501_, _23500_, _06160_);
  or _74388_ (_23502_, _23501_, _23499_);
  and _74389_ (_23503_, _23502_, _06157_);
  and _74390_ (_23504_, _23503_, _23496_);
  and _74391_ (_23505_, _11644_, \oc8051_golden_model_1.TCON [6]);
  and _74392_ (_23506_, _15316_, _08407_);
  or _74393_ (_23507_, _23506_, _23505_);
  and _74394_ (_23508_, _23507_, _06156_);
  or _74395_ (_23509_, _23508_, _06217_);
  or _74396_ (_23511_, _23509_, _23504_);
  and _74397_ (_23512_, _08012_, _07788_);
  or _74398_ (_23513_, _23512_, _23493_);
  or _74399_ (_23514_, _23513_, _07075_);
  and _74400_ (_23515_, _23514_, _23511_);
  or _74401_ (_23516_, _23515_, _06220_);
  or _74402_ (_23517_, _23498_, _06229_);
  and _74403_ (_23518_, _23517_, _06153_);
  and _74404_ (_23519_, _23518_, _23516_);
  and _74405_ (_23520_, _15297_, _08407_);
  or _74406_ (_23522_, _23520_, _23505_);
  and _74407_ (_23523_, _23522_, _06152_);
  or _74408_ (_23524_, _23523_, _06145_);
  or _74409_ (_23525_, _23524_, _23519_);
  or _74410_ (_23526_, _23505_, _15331_);
  and _74411_ (_23527_, _23526_, _23507_);
  or _74412_ (_23528_, _23527_, _06146_);
  and _74413_ (_23529_, _23528_, _06140_);
  and _74414_ (_23530_, _23529_, _23525_);
  and _74415_ (_23531_, _15348_, _08407_);
  or _74416_ (_23533_, _23531_, _23505_);
  and _74417_ (_23534_, _23533_, _06139_);
  or _74418_ (_23535_, _23534_, _09842_);
  or _74419_ (_23536_, _23535_, _23530_);
  or _74420_ (_23537_, _23513_, _06132_);
  and _74421_ (_23538_, _23537_, _23536_);
  or _74422_ (_23539_, _23538_, _06116_);
  and _74423_ (_23540_, _09207_, _07788_);
  or _74424_ (_23541_, _23493_, _06117_);
  or _74425_ (_23542_, _23541_, _23540_);
  and _74426_ (_23543_, _23542_, _06114_);
  and _74427_ (_23544_, _23543_, _23539_);
  and _74428_ (_23545_, _15395_, _07788_);
  or _74429_ (_23546_, _23545_, _23493_);
  and _74430_ (_23547_, _23546_, _05787_);
  or _74431_ (_23548_, _23547_, _11136_);
  or _74432_ (_23549_, _23548_, _23544_);
  and _74433_ (_23550_, _15413_, _07788_);
  or _74434_ (_23551_, _23493_, _07127_);
  or _74435_ (_23552_, _23551_, _23550_);
  and _74436_ (_23554_, _15402_, _07788_);
  or _74437_ (_23555_, _23554_, _23493_);
  or _74438_ (_23556_, _23555_, _06111_);
  and _74439_ (_23557_, _23556_, _07125_);
  and _74440_ (_23558_, _23557_, _23552_);
  and _74441_ (_23559_, _23558_, _23549_);
  and _74442_ (_23560_, _10295_, _07788_);
  or _74443_ (_23561_, _23560_, _23493_);
  and _74444_ (_23562_, _23561_, _06402_);
  or _74445_ (_23563_, _23562_, _23559_);
  and _74446_ (_23565_, _23563_, _07132_);
  or _74447_ (_23566_, _23493_, _08015_);
  and _74448_ (_23567_, _23555_, _06306_);
  and _74449_ (_23568_, _23567_, _23566_);
  or _74450_ (_23569_, _23568_, _23565_);
  and _74451_ (_23570_, _23569_, _07130_);
  and _74452_ (_23571_, _23498_, _06411_);
  and _74453_ (_23572_, _23571_, _23566_);
  or _74454_ (_23573_, _23572_, _06303_);
  or _74455_ (_23574_, _23573_, _23570_);
  and _74456_ (_23575_, _15410_, _07788_);
  or _74457_ (_23576_, _23493_, _08819_);
  or _74458_ (_23577_, _23576_, _23575_);
  and _74459_ (_23578_, _23577_, _08824_);
  and _74460_ (_23579_, _23578_, _23574_);
  nor _74461_ (_23580_, _10294_, _11639_);
  or _74462_ (_23581_, _23580_, _23493_);
  and _74463_ (_23582_, _23581_, _06396_);
  or _74464_ (_23583_, _23582_, _06433_);
  or _74465_ (_23584_, _23583_, _23579_);
  or _74466_ (_23586_, _23495_, _06829_);
  and _74467_ (_23587_, _23586_, _05749_);
  and _74468_ (_23588_, _23587_, _23584_);
  and _74469_ (_23589_, _23522_, _05748_);
  or _74470_ (_23590_, _23589_, _06440_);
  or _74471_ (_23591_, _23590_, _23588_);
  and _74472_ (_23592_, _15478_, _07788_);
  or _74473_ (_23593_, _23493_, _06444_);
  or _74474_ (_23594_, _23593_, _23592_);
  and _74475_ (_23595_, _23594_, _01317_);
  and _74476_ (_23597_, _23595_, _23591_);
  or _74477_ (_23598_, _23597_, _23492_);
  and _74478_ (_43668_, _23598_, _43100_);
  not _74479_ (_23599_, \oc8051_golden_model_1.TH1 [0]);
  nor _74480_ (_23600_, _01317_, _23599_);
  nand _74481_ (_23601_, _10276_, _07817_);
  nor _74482_ (_23602_, _07817_, _23599_);
  nor _74483_ (_23603_, _23602_, _07130_);
  nand _74484_ (_23604_, _23603_, _23601_);
  nor _74485_ (_23605_, _08211_, _11740_);
  or _74486_ (_23607_, _23605_, _23602_);
  or _74487_ (_23608_, _23607_, _06161_);
  and _74488_ (_23609_, _07817_, \oc8051_golden_model_1.ACC [0]);
  or _74489_ (_23610_, _23609_, _23602_);
  and _74490_ (_23611_, _23610_, _07056_);
  nor _74491_ (_23612_, _07056_, _23599_);
  or _74492_ (_23613_, _23612_, _06160_);
  or _74493_ (_23614_, _23613_, _23611_);
  and _74494_ (_23615_, _23614_, _07075_);
  and _74495_ (_23616_, _23615_, _23608_);
  and _74496_ (_23618_, _07817_, _07049_);
  or _74497_ (_23619_, _23618_, _23602_);
  and _74498_ (_23620_, _23619_, _06217_);
  or _74499_ (_23621_, _23620_, _23616_);
  and _74500_ (_23622_, _23621_, _06229_);
  and _74501_ (_23623_, _23610_, _06220_);
  or _74502_ (_23624_, _23623_, _09842_);
  or _74503_ (_23625_, _23624_, _23622_);
  or _74504_ (_23626_, _23619_, _06132_);
  and _74505_ (_23627_, _23626_, _23625_);
  or _74506_ (_23629_, _23627_, _06116_);
  and _74507_ (_23630_, _09160_, _07817_);
  or _74508_ (_23631_, _23602_, _06117_);
  or _74509_ (_23632_, _23631_, _23630_);
  and _74510_ (_23633_, _23632_, _23629_);
  or _74511_ (_23634_, _23633_, _05787_);
  and _74512_ (_23635_, _14260_, _07817_);
  or _74513_ (_23636_, _23635_, _23602_);
  or _74514_ (_23637_, _23636_, _06114_);
  and _74515_ (_23638_, _23637_, _06111_);
  and _74516_ (_23640_, _23638_, _23634_);
  and _74517_ (_23641_, _07817_, _08708_);
  or _74518_ (_23642_, _23641_, _23602_);
  and _74519_ (_23643_, _23642_, _06110_);
  or _74520_ (_23644_, _23643_, _06297_);
  or _74521_ (_23645_, _23644_, _23640_);
  and _74522_ (_23646_, _14275_, _07817_);
  or _74523_ (_23647_, _23602_, _07127_);
  or _74524_ (_23648_, _23647_, _23646_);
  and _74525_ (_23649_, _23648_, _07125_);
  and _74526_ (_23651_, _23649_, _23645_);
  nor _74527_ (_23652_, _12321_, _11740_);
  or _74528_ (_23653_, _23652_, _23602_);
  and _74529_ (_23654_, _23601_, _06402_);
  and _74530_ (_23655_, _23654_, _23653_);
  or _74531_ (_23656_, _23655_, _23651_);
  and _74532_ (_23657_, _23656_, _07132_);
  nand _74533_ (_23658_, _23642_, _06306_);
  nor _74534_ (_23659_, _23658_, _23605_);
  or _74535_ (_23660_, _23659_, _06411_);
  or _74536_ (_23662_, _23660_, _23657_);
  and _74537_ (_23663_, _23662_, _23604_);
  or _74538_ (_23664_, _23663_, _06303_);
  and _74539_ (_23665_, _14167_, _07817_);
  or _74540_ (_23666_, _23602_, _08819_);
  or _74541_ (_23667_, _23666_, _23665_);
  and _74542_ (_23668_, _23667_, _08824_);
  and _74543_ (_23669_, _23668_, _23664_);
  and _74544_ (_23670_, _23653_, _06396_);
  or _74545_ (_23671_, _23670_, _19287_);
  or _74546_ (_23673_, _23671_, _23669_);
  or _74547_ (_23674_, _23607_, _06630_);
  and _74548_ (_23675_, _23674_, _01317_);
  and _74549_ (_23676_, _23675_, _23673_);
  or _74550_ (_23677_, _23676_, _23600_);
  and _74551_ (_43670_, _23677_, _43100_);
  not _74552_ (_23678_, \oc8051_golden_model_1.TH1 [1]);
  nor _74553_ (_23679_, _01317_, _23678_);
  or _74554_ (_23680_, _14442_, _11740_);
  or _74555_ (_23681_, _07817_, \oc8051_golden_model_1.TH1 [1]);
  and _74556_ (_23682_, _23681_, _05787_);
  and _74557_ (_23683_, _23682_, _23680_);
  nor _74558_ (_23684_, _07817_, _23678_);
  and _74559_ (_23685_, _07817_, _07306_);
  or _74560_ (_23686_, _23685_, _23684_);
  or _74561_ (_23687_, _23686_, _06132_);
  and _74562_ (_23688_, _07817_, \oc8051_golden_model_1.ACC [1]);
  or _74563_ (_23689_, _23688_, _23684_);
  and _74564_ (_23690_, _23689_, _06220_);
  or _74565_ (_23691_, _23690_, _09842_);
  and _74566_ (_23692_, _14363_, _07817_);
  not _74567_ (_23693_, _23692_);
  and _74568_ (_23694_, _23693_, _23681_);
  and _74569_ (_23695_, _23694_, _06160_);
  nor _74570_ (_23696_, _07056_, _23678_);
  and _74571_ (_23697_, _23689_, _07056_);
  or _74572_ (_23698_, _23697_, _23696_);
  and _74573_ (_23699_, _23698_, _06161_);
  or _74574_ (_23700_, _23699_, _06217_);
  or _74575_ (_23701_, _23700_, _23695_);
  or _74576_ (_23703_, _23686_, _07075_);
  and _74577_ (_23704_, _23703_, _06229_);
  and _74578_ (_23705_, _23704_, _23701_);
  or _74579_ (_23706_, _23705_, _23691_);
  and _74580_ (_23707_, _23706_, _23687_);
  or _74581_ (_23708_, _23707_, _06116_);
  and _74582_ (_23709_, _23708_, _06114_);
  and _74583_ (_23710_, _09115_, _07817_);
  or _74584_ (_23711_, _23684_, _06117_);
  or _74585_ (_23712_, _23711_, _23710_);
  and _74586_ (_23714_, _23712_, _23709_);
  or _74587_ (_23715_, _23714_, _23683_);
  and _74588_ (_23716_, _23715_, _06298_);
  or _74589_ (_23717_, _14346_, _11740_);
  and _74590_ (_23718_, _23717_, _06297_);
  nand _74591_ (_23719_, _07817_, _06945_);
  and _74592_ (_23720_, _23719_, _06110_);
  or _74593_ (_23721_, _23720_, _23718_);
  and _74594_ (_23722_, _23721_, _23681_);
  or _74595_ (_23723_, _23722_, _06402_);
  or _74596_ (_23725_, _23723_, _23716_);
  nor _74597_ (_23726_, _10277_, _11740_);
  or _74598_ (_23727_, _23726_, _23684_);
  nand _74599_ (_23728_, _10275_, _07817_);
  and _74600_ (_23729_, _23728_, _23727_);
  or _74601_ (_23730_, _23729_, _07125_);
  and _74602_ (_23731_, _23730_, _07132_);
  and _74603_ (_23732_, _23731_, _23725_);
  or _74604_ (_23733_, _14344_, _11740_);
  and _74605_ (_23734_, _23681_, _06306_);
  and _74606_ (_23736_, _23734_, _23733_);
  or _74607_ (_23737_, _23736_, _06411_);
  or _74608_ (_23738_, _23737_, _23732_);
  nor _74609_ (_23739_, _23684_, _07130_);
  nand _74610_ (_23740_, _23739_, _23728_);
  and _74611_ (_23741_, _23740_, _08819_);
  and _74612_ (_23742_, _23741_, _23738_);
  or _74613_ (_23743_, _23719_, _08176_);
  and _74614_ (_23744_, _23681_, _06303_);
  and _74615_ (_23745_, _23744_, _23743_);
  or _74616_ (_23747_, _23745_, _06396_);
  or _74617_ (_23748_, _23747_, _23742_);
  or _74618_ (_23749_, _23727_, _08824_);
  and _74619_ (_23750_, _23749_, _06829_);
  and _74620_ (_23751_, _23750_, _23748_);
  and _74621_ (_23752_, _23694_, _06433_);
  or _74622_ (_23753_, _23752_, _06440_);
  or _74623_ (_23754_, _23753_, _23751_);
  or _74624_ (_23755_, _23684_, _06444_);
  or _74625_ (_23756_, _23755_, _23692_);
  and _74626_ (_23758_, _23756_, _01317_);
  and _74627_ (_23759_, _23758_, _23754_);
  or _74628_ (_23760_, _23759_, _23679_);
  and _74629_ (_43671_, _23760_, _43100_);
  and _74630_ (_23761_, _01321_, \oc8051_golden_model_1.TH1 [2]);
  and _74631_ (_23762_, _11740_, \oc8051_golden_model_1.TH1 [2]);
  or _74632_ (_23763_, _23762_, _08248_);
  and _74633_ (_23764_, _07817_, _08768_);
  or _74634_ (_23765_, _23764_, _23762_);
  and _74635_ (_23766_, _23765_, _06306_);
  and _74636_ (_23768_, _23766_, _23763_);
  and _74637_ (_23769_, _09211_, _07817_);
  or _74638_ (_23770_, _23769_, _23762_);
  and _74639_ (_23771_, _23770_, _06116_);
  and _74640_ (_23772_, _14542_, _07817_);
  or _74641_ (_23773_, _23772_, _23762_);
  or _74642_ (_23774_, _23773_, _06161_);
  and _74643_ (_23775_, _07817_, \oc8051_golden_model_1.ACC [2]);
  or _74644_ (_23776_, _23775_, _23762_);
  and _74645_ (_23777_, _23776_, _07056_);
  and _74646_ (_23779_, _07057_, \oc8051_golden_model_1.TH1 [2]);
  or _74647_ (_23780_, _23779_, _06160_);
  or _74648_ (_23781_, _23780_, _23777_);
  and _74649_ (_23782_, _23781_, _07075_);
  and _74650_ (_23783_, _23782_, _23774_);
  and _74651_ (_23784_, _07817_, _07708_);
  or _74652_ (_23785_, _23784_, _23762_);
  and _74653_ (_23786_, _23785_, _06217_);
  or _74654_ (_23787_, _23786_, _23783_);
  and _74655_ (_23788_, _23787_, _06229_);
  and _74656_ (_23790_, _23776_, _06220_);
  or _74657_ (_23791_, _23790_, _09842_);
  or _74658_ (_23792_, _23791_, _23788_);
  or _74659_ (_23793_, _23785_, _06132_);
  and _74660_ (_23794_, _23793_, _06117_);
  and _74661_ (_23795_, _23794_, _23792_);
  or _74662_ (_23796_, _23795_, _05787_);
  or _74663_ (_23797_, _23796_, _23771_);
  and _74664_ (_23798_, _14630_, _07817_);
  or _74665_ (_23799_, _23798_, _23762_);
  or _74666_ (_23801_, _23799_, _06114_);
  and _74667_ (_23802_, _23801_, _06111_);
  and _74668_ (_23803_, _23802_, _23797_);
  and _74669_ (_23804_, _23765_, _06110_);
  or _74670_ (_23805_, _23804_, _06297_);
  or _74671_ (_23806_, _23805_, _23803_);
  and _74672_ (_23807_, _14646_, _07817_);
  or _74673_ (_23808_, _23762_, _07127_);
  or _74674_ (_23809_, _23808_, _23807_);
  and _74675_ (_23810_, _23809_, _07125_);
  and _74676_ (_23812_, _23810_, _23806_);
  and _74677_ (_23813_, _10282_, _07817_);
  or _74678_ (_23814_, _23813_, _23762_);
  and _74679_ (_23815_, _23814_, _06402_);
  or _74680_ (_23816_, _23815_, _23812_);
  and _74681_ (_23817_, _23816_, _07132_);
  or _74682_ (_23818_, _23817_, _23768_);
  and _74683_ (_23819_, _23818_, _07130_);
  and _74684_ (_23820_, _23776_, _06411_);
  and _74685_ (_23821_, _23820_, _23763_);
  or _74686_ (_23823_, _23821_, _06303_);
  or _74687_ (_23824_, _23823_, _23819_);
  and _74688_ (_23825_, _14643_, _07817_);
  or _74689_ (_23826_, _23762_, _08819_);
  or _74690_ (_23827_, _23826_, _23825_);
  and _74691_ (_23828_, _23827_, _08824_);
  and _74692_ (_23829_, _23828_, _23824_);
  nor _74693_ (_23830_, _10281_, _11740_);
  or _74694_ (_23831_, _23830_, _23762_);
  and _74695_ (_23832_, _23831_, _06396_);
  or _74696_ (_23834_, _23832_, _23829_);
  and _74697_ (_23835_, _23834_, _06829_);
  and _74698_ (_23836_, _23773_, _06433_);
  or _74699_ (_23837_, _23836_, _06440_);
  or _74700_ (_23838_, _23837_, _23835_);
  and _74701_ (_23839_, _14710_, _07817_);
  or _74702_ (_23840_, _23762_, _06444_);
  or _74703_ (_23841_, _23840_, _23839_);
  and _74704_ (_23842_, _23841_, _01317_);
  and _74705_ (_23843_, _23842_, _23838_);
  or _74706_ (_23845_, _23843_, _23761_);
  and _74707_ (_43672_, _23845_, _43100_);
  and _74708_ (_23846_, _11740_, \oc8051_golden_model_1.TH1 [3]);
  and _74709_ (_23847_, _14738_, _07817_);
  or _74710_ (_23848_, _23847_, _23846_);
  or _74711_ (_23849_, _23848_, _06161_);
  and _74712_ (_23850_, _07817_, \oc8051_golden_model_1.ACC [3]);
  or _74713_ (_23851_, _23850_, _23846_);
  and _74714_ (_23852_, _23851_, _07056_);
  and _74715_ (_23853_, _07057_, \oc8051_golden_model_1.TH1 [3]);
  or _74716_ (_23855_, _23853_, _06160_);
  or _74717_ (_23856_, _23855_, _23852_);
  and _74718_ (_23857_, _23856_, _07075_);
  and _74719_ (_23858_, _23857_, _23849_);
  and _74720_ (_23859_, _07817_, _07544_);
  or _74721_ (_23860_, _23859_, _23846_);
  and _74722_ (_23861_, _23860_, _06217_);
  or _74723_ (_23862_, _23861_, _23858_);
  and _74724_ (_23863_, _23862_, _06229_);
  and _74725_ (_23864_, _23851_, _06220_);
  or _74726_ (_23866_, _23864_, _09842_);
  or _74727_ (_23867_, _23866_, _23863_);
  or _74728_ (_23868_, _23860_, _06132_);
  and _74729_ (_23869_, _23868_, _06117_);
  and _74730_ (_23870_, _23869_, _23867_);
  and _74731_ (_23871_, _09210_, _07817_);
  or _74732_ (_23872_, _23871_, _23846_);
  and _74733_ (_23873_, _23872_, _06116_);
  or _74734_ (_23874_, _23873_, _05787_);
  or _74735_ (_23875_, _23874_, _23870_);
  and _74736_ (_23877_, _14825_, _07817_);
  or _74737_ (_23878_, _23846_, _06114_);
  or _74738_ (_23879_, _23878_, _23877_);
  and _74739_ (_23880_, _23879_, _06111_);
  and _74740_ (_23881_, _23880_, _23875_);
  and _74741_ (_23882_, _07817_, _08712_);
  or _74742_ (_23883_, _23882_, _23846_);
  and _74743_ (_23884_, _23883_, _06110_);
  or _74744_ (_23885_, _23884_, _06297_);
  or _74745_ (_23886_, _23885_, _23881_);
  and _74746_ (_23887_, _14727_, _07817_);
  or _74747_ (_23888_, _23887_, _23846_);
  or _74748_ (_23889_, _23888_, _07127_);
  and _74749_ (_23890_, _23889_, _07125_);
  and _74750_ (_23891_, _23890_, _23886_);
  and _74751_ (_23892_, _12318_, _07817_);
  or _74752_ (_23893_, _23892_, _23846_);
  and _74753_ (_23894_, _23893_, _06402_);
  or _74754_ (_23895_, _23894_, _23891_);
  and _74755_ (_23896_, _23895_, _07132_);
  or _74756_ (_23899_, _23846_, _08140_);
  and _74757_ (_23900_, _23883_, _06306_);
  and _74758_ (_23901_, _23900_, _23899_);
  or _74759_ (_23902_, _23901_, _23896_);
  and _74760_ (_23903_, _23902_, _07130_);
  and _74761_ (_23904_, _23851_, _06411_);
  and _74762_ (_23905_, _23904_, _23899_);
  or _74763_ (_23906_, _23905_, _06303_);
  or _74764_ (_23907_, _23906_, _23903_);
  and _74765_ (_23908_, _14724_, _07817_);
  or _74766_ (_23910_, _23846_, _08819_);
  or _74767_ (_23911_, _23910_, _23908_);
  and _74768_ (_23912_, _23911_, _08824_);
  and _74769_ (_23913_, _23912_, _23907_);
  nor _74770_ (_23914_, _10273_, _11740_);
  or _74771_ (_23915_, _23914_, _23846_);
  and _74772_ (_23916_, _23915_, _06396_);
  or _74773_ (_23917_, _23916_, _06433_);
  or _74774_ (_23918_, _23917_, _23913_);
  or _74775_ (_23919_, _23848_, _06829_);
  and _74776_ (_23921_, _23919_, _06444_);
  and _74777_ (_23922_, _23921_, _23918_);
  and _74778_ (_23923_, _14897_, _07817_);
  or _74779_ (_23924_, _23923_, _23846_);
  and _74780_ (_23925_, _23924_, _06440_);
  or _74781_ (_23926_, _23925_, _01321_);
  or _74782_ (_23927_, _23926_, _23922_);
  or _74783_ (_23928_, _01317_, \oc8051_golden_model_1.TH1 [3]);
  and _74784_ (_23929_, _23928_, _43100_);
  and _74785_ (_43673_, _23929_, _23927_);
  and _74786_ (_23931_, _11740_, \oc8051_golden_model_1.TH1 [4]);
  and _74787_ (_23932_, _14928_, _07817_);
  or _74788_ (_23933_, _23932_, _23931_);
  or _74789_ (_23934_, _23933_, _06161_);
  and _74790_ (_23935_, _07817_, \oc8051_golden_model_1.ACC [4]);
  or _74791_ (_23936_, _23935_, _23931_);
  and _74792_ (_23937_, _23936_, _07056_);
  and _74793_ (_23938_, _07057_, \oc8051_golden_model_1.TH1 [4]);
  or _74794_ (_23939_, _23938_, _06160_);
  or _74795_ (_23940_, _23939_, _23937_);
  and _74796_ (_23942_, _23940_, _07075_);
  and _74797_ (_23943_, _23942_, _23934_);
  and _74798_ (_23944_, _08336_, _07817_);
  or _74799_ (_23945_, _23944_, _23931_);
  and _74800_ (_23946_, _23945_, _06217_);
  or _74801_ (_23947_, _23946_, _23943_);
  and _74802_ (_23948_, _23947_, _06229_);
  and _74803_ (_23949_, _23936_, _06220_);
  or _74804_ (_23950_, _23949_, _09842_);
  or _74805_ (_23951_, _23950_, _23948_);
  or _74806_ (_23953_, _23945_, _06132_);
  and _74807_ (_23954_, _23953_, _23951_);
  or _74808_ (_23955_, _23954_, _06116_);
  and _74809_ (_23956_, _09209_, _07817_);
  or _74810_ (_23957_, _23931_, _06117_);
  or _74811_ (_23958_, _23957_, _23956_);
  and _74812_ (_23959_, _23958_, _06114_);
  and _74813_ (_23960_, _23959_, _23955_);
  and _74814_ (_23961_, _15013_, _07817_);
  or _74815_ (_23962_, _23961_, _23931_);
  and _74816_ (_23964_, _23962_, _05787_);
  or _74817_ (_23965_, _23964_, _23960_);
  or _74818_ (_23966_, _23965_, _11136_);
  and _74819_ (_23967_, _15029_, _07817_);
  or _74820_ (_23968_, _23931_, _07127_);
  or _74821_ (_23969_, _23968_, _23967_);
  and _74822_ (_23970_, _08715_, _07817_);
  or _74823_ (_23971_, _23970_, _23931_);
  or _74824_ (_23972_, _23971_, _06111_);
  and _74825_ (_23973_, _23972_, _07125_);
  and _74826_ (_23975_, _23973_, _23969_);
  and _74827_ (_23976_, _23975_, _23966_);
  and _74828_ (_23977_, _10289_, _07817_);
  or _74829_ (_23978_, _23977_, _23931_);
  and _74830_ (_23979_, _23978_, _06402_);
  or _74831_ (_23980_, _23979_, _23976_);
  and _74832_ (_23981_, _23980_, _07132_);
  or _74833_ (_23982_, _23931_, _08339_);
  and _74834_ (_23983_, _23971_, _06306_);
  and _74835_ (_23984_, _23983_, _23982_);
  or _74836_ (_23986_, _23984_, _23981_);
  and _74837_ (_23987_, _23986_, _07130_);
  and _74838_ (_23988_, _23936_, _06411_);
  and _74839_ (_23989_, _23988_, _23982_);
  or _74840_ (_23990_, _23989_, _06303_);
  or _74841_ (_23991_, _23990_, _23987_);
  and _74842_ (_23992_, _15026_, _07817_);
  or _74843_ (_23993_, _23931_, _08819_);
  or _74844_ (_23994_, _23993_, _23992_);
  and _74845_ (_23995_, _23994_, _08824_);
  and _74846_ (_23997_, _23995_, _23991_);
  nor _74847_ (_23998_, _10288_, _11740_);
  or _74848_ (_23999_, _23998_, _23931_);
  and _74849_ (_24000_, _23999_, _06396_);
  or _74850_ (_24001_, _24000_, _06433_);
  or _74851_ (_24002_, _24001_, _23997_);
  or _74852_ (_24003_, _23933_, _06829_);
  and _74853_ (_24004_, _24003_, _06444_);
  and _74854_ (_24005_, _24004_, _24002_);
  and _74855_ (_24006_, _15087_, _07817_);
  or _74856_ (_24008_, _24006_, _23931_);
  and _74857_ (_24009_, _24008_, _06440_);
  or _74858_ (_24010_, _24009_, _01321_);
  or _74859_ (_24011_, _24010_, _24005_);
  or _74860_ (_24012_, _01317_, \oc8051_golden_model_1.TH1 [4]);
  and _74861_ (_24013_, _24012_, _43100_);
  and _74862_ (_43674_, _24013_, _24011_);
  and _74863_ (_24014_, _11740_, \oc8051_golden_model_1.TH1 [5]);
  or _74864_ (_24015_, _24014_, _08104_);
  and _74865_ (_24016_, _08736_, _07817_);
  or _74866_ (_24018_, _24016_, _24014_);
  and _74867_ (_24019_, _24018_, _06306_);
  and _74868_ (_24020_, _24019_, _24015_);
  and _74869_ (_24021_, _15119_, _07817_);
  or _74870_ (_24022_, _24021_, _24014_);
  or _74871_ (_24023_, _24022_, _06161_);
  and _74872_ (_24024_, _07817_, \oc8051_golden_model_1.ACC [5]);
  or _74873_ (_24025_, _24024_, _24014_);
  and _74874_ (_24026_, _24025_, _07056_);
  and _74875_ (_24027_, _07057_, \oc8051_golden_model_1.TH1 [5]);
  or _74876_ (_24029_, _24027_, _06160_);
  or _74877_ (_24030_, _24029_, _24026_);
  and _74878_ (_24031_, _24030_, _07075_);
  and _74879_ (_24032_, _24031_, _24023_);
  and _74880_ (_24033_, _08101_, _07817_);
  or _74881_ (_24034_, _24033_, _24014_);
  and _74882_ (_24035_, _24034_, _06217_);
  or _74883_ (_24036_, _24035_, _24032_);
  and _74884_ (_24037_, _24036_, _06229_);
  and _74885_ (_24038_, _24025_, _06220_);
  or _74886_ (_24040_, _24038_, _09842_);
  or _74887_ (_24041_, _24040_, _24037_);
  or _74888_ (_24042_, _24034_, _06132_);
  and _74889_ (_24043_, _24042_, _24041_);
  or _74890_ (_24044_, _24043_, _06116_);
  and _74891_ (_24045_, _09208_, _07817_);
  or _74892_ (_24046_, _24014_, _06117_);
  or _74893_ (_24047_, _24046_, _24045_);
  and _74894_ (_24048_, _24047_, _06114_);
  and _74895_ (_24049_, _24048_, _24044_);
  and _74896_ (_24051_, _15203_, _07817_);
  or _74897_ (_24052_, _24051_, _24014_);
  and _74898_ (_24053_, _24052_, _05787_);
  or _74899_ (_24054_, _24053_, _11136_);
  or _74900_ (_24055_, _24054_, _24049_);
  and _74901_ (_24056_, _15219_, _07817_);
  or _74902_ (_24057_, _24014_, _07127_);
  or _74903_ (_24058_, _24057_, _24056_);
  or _74904_ (_24059_, _24018_, _06111_);
  and _74905_ (_24060_, _24059_, _07125_);
  and _74906_ (_24062_, _24060_, _24058_);
  and _74907_ (_24063_, _24062_, _24055_);
  and _74908_ (_24064_, _12325_, _07817_);
  or _74909_ (_24065_, _24064_, _24014_);
  and _74910_ (_24066_, _24065_, _06402_);
  or _74911_ (_24067_, _24066_, _24063_);
  and _74912_ (_24068_, _24067_, _07132_);
  or _74913_ (_24069_, _24068_, _24020_);
  and _74914_ (_24070_, _24069_, _07130_);
  and _74915_ (_24071_, _24025_, _06411_);
  and _74916_ (_24072_, _24071_, _24015_);
  or _74917_ (_24073_, _24072_, _06303_);
  or _74918_ (_24074_, _24073_, _24070_);
  and _74919_ (_24075_, _15216_, _07817_);
  or _74920_ (_24076_, _24014_, _08819_);
  or _74921_ (_24077_, _24076_, _24075_);
  and _74922_ (_24078_, _24077_, _08824_);
  and _74923_ (_24079_, _24078_, _24074_);
  nor _74924_ (_24080_, _10269_, _11740_);
  or _74925_ (_24081_, _24080_, _24014_);
  and _74926_ (_24084_, _24081_, _06396_);
  or _74927_ (_24085_, _24084_, _06433_);
  or _74928_ (_24086_, _24085_, _24079_);
  or _74929_ (_24087_, _24022_, _06829_);
  and _74930_ (_24088_, _24087_, _06444_);
  and _74931_ (_24089_, _24088_, _24086_);
  and _74932_ (_24090_, _15275_, _07817_);
  or _74933_ (_24091_, _24090_, _24014_);
  and _74934_ (_24092_, _24091_, _06440_);
  or _74935_ (_24093_, _24092_, _01321_);
  or _74936_ (_24095_, _24093_, _24089_);
  or _74937_ (_24096_, _01317_, \oc8051_golden_model_1.TH1 [5]);
  and _74938_ (_24097_, _24096_, _43100_);
  and _74939_ (_43675_, _24097_, _24095_);
  and _74940_ (_24098_, _11740_, \oc8051_golden_model_1.TH1 [6]);
  and _74941_ (_24099_, _15300_, _07817_);
  or _74942_ (_24100_, _24099_, _24098_);
  or _74943_ (_24101_, _24100_, _06161_);
  and _74944_ (_24102_, _07817_, \oc8051_golden_model_1.ACC [6]);
  or _74945_ (_24103_, _24102_, _24098_);
  and _74946_ (_24105_, _24103_, _07056_);
  and _74947_ (_24106_, _07057_, \oc8051_golden_model_1.TH1 [6]);
  or _74948_ (_24107_, _24106_, _06160_);
  or _74949_ (_24108_, _24107_, _24105_);
  and _74950_ (_24109_, _24108_, _07075_);
  and _74951_ (_24110_, _24109_, _24101_);
  and _74952_ (_24111_, _08012_, _07817_);
  or _74953_ (_24112_, _24111_, _24098_);
  and _74954_ (_24113_, _24112_, _06217_);
  or _74955_ (_24114_, _24113_, _24110_);
  and _74956_ (_24116_, _24114_, _06229_);
  and _74957_ (_24117_, _24103_, _06220_);
  or _74958_ (_24118_, _24117_, _09842_);
  or _74959_ (_24119_, _24118_, _24116_);
  or _74960_ (_24120_, _24112_, _06132_);
  and _74961_ (_24121_, _24120_, _24119_);
  or _74962_ (_24122_, _24121_, _06116_);
  and _74963_ (_24123_, _09207_, _07817_);
  or _74964_ (_24124_, _24098_, _06117_);
  or _74965_ (_24125_, _24124_, _24123_);
  and _74966_ (_24127_, _24125_, _06114_);
  and _74967_ (_24128_, _24127_, _24122_);
  and _74968_ (_24129_, _15395_, _07817_);
  or _74969_ (_24130_, _24129_, _24098_);
  and _74970_ (_24131_, _24130_, _05787_);
  or _74971_ (_24132_, _24131_, _11136_);
  or _74972_ (_24133_, _24132_, _24128_);
  and _74973_ (_24134_, _15413_, _07817_);
  or _74974_ (_24135_, _24098_, _07127_);
  or _74975_ (_24136_, _24135_, _24134_);
  and _74976_ (_24138_, _15402_, _07817_);
  or _74977_ (_24139_, _24138_, _24098_);
  or _74978_ (_24140_, _24139_, _06111_);
  and _74979_ (_24141_, _24140_, _07125_);
  and _74980_ (_24142_, _24141_, _24136_);
  and _74981_ (_24143_, _24142_, _24133_);
  and _74982_ (_24144_, _10295_, _07817_);
  or _74983_ (_24145_, _24144_, _24098_);
  and _74984_ (_24146_, _24145_, _06402_);
  or _74985_ (_24147_, _24146_, _24143_);
  and _74986_ (_24149_, _24147_, _07132_);
  or _74987_ (_24150_, _24098_, _08015_);
  and _74988_ (_24151_, _24139_, _06306_);
  and _74989_ (_24152_, _24151_, _24150_);
  or _74990_ (_24153_, _24152_, _24149_);
  and _74991_ (_24154_, _24153_, _07130_);
  and _74992_ (_24155_, _24103_, _06411_);
  and _74993_ (_24156_, _24155_, _24150_);
  or _74994_ (_24157_, _24156_, _06303_);
  or _74995_ (_24158_, _24157_, _24154_);
  and _74996_ (_24160_, _15410_, _07817_);
  or _74997_ (_24161_, _24098_, _08819_);
  or _74998_ (_24162_, _24161_, _24160_);
  and _74999_ (_24163_, _24162_, _08824_);
  and _75000_ (_24164_, _24163_, _24158_);
  nor _75001_ (_24165_, _10294_, _11740_);
  or _75002_ (_24166_, _24165_, _24098_);
  and _75003_ (_24167_, _24166_, _06396_);
  or _75004_ (_24168_, _24167_, _06433_);
  or _75005_ (_24169_, _24168_, _24164_);
  or _75006_ (_24171_, _24100_, _06829_);
  and _75007_ (_24172_, _24171_, _06444_);
  and _75008_ (_24173_, _24172_, _24169_);
  and _75009_ (_24174_, _15478_, _07817_);
  or _75010_ (_24175_, _24174_, _24098_);
  and _75011_ (_24176_, _24175_, _06440_);
  or _75012_ (_24177_, _24176_, _01321_);
  or _75013_ (_24178_, _24177_, _24173_);
  or _75014_ (_24179_, _01317_, \oc8051_golden_model_1.TH1 [6]);
  and _75015_ (_24180_, _24179_, _43100_);
  and _75016_ (_43676_, _24180_, _24178_);
  not _75017_ (_24182_, \oc8051_golden_model_1.TH0 [0]);
  nor _75018_ (_24183_, _01317_, _24182_);
  nand _75019_ (_24184_, _10276_, _07823_);
  nor _75020_ (_24185_, _07823_, _24182_);
  nor _75021_ (_24186_, _24185_, _07130_);
  nand _75022_ (_24187_, _24186_, _24184_);
  and _75023_ (_24188_, _07823_, \oc8051_golden_model_1.ACC [0]);
  or _75024_ (_24189_, _24188_, _24185_);
  and _75025_ (_24190_, _24189_, _06220_);
  or _75026_ (_24192_, _24190_, _09842_);
  nor _75027_ (_24193_, _08211_, _11817_);
  or _75028_ (_24194_, _24193_, _24185_);
  and _75029_ (_24195_, _24194_, _06160_);
  nor _75030_ (_24196_, _07056_, _24182_);
  and _75031_ (_24197_, _24189_, _07056_);
  or _75032_ (_24198_, _24197_, _24196_);
  and _75033_ (_24199_, _24198_, _06161_);
  or _75034_ (_24200_, _24199_, _06217_);
  or _75035_ (_24201_, _24200_, _24195_);
  and _75036_ (_24203_, _24201_, _06229_);
  or _75037_ (_24204_, _24203_, _24192_);
  and _75038_ (_24205_, _07823_, _07049_);
  and _75039_ (_24206_, _06132_, _07075_);
  or _75040_ (_24207_, _24185_, _24206_);
  or _75041_ (_24208_, _24207_, _24205_);
  and _75042_ (_24209_, _24208_, _24204_);
  or _75043_ (_24210_, _24209_, _06116_);
  and _75044_ (_24211_, _09160_, _07823_);
  or _75045_ (_24212_, _24185_, _06117_);
  or _75046_ (_24214_, _24212_, _24211_);
  and _75047_ (_24215_, _24214_, _24210_);
  or _75048_ (_24216_, _24215_, _05787_);
  and _75049_ (_24217_, _14260_, _07823_);
  or _75050_ (_24218_, _24217_, _24185_);
  or _75051_ (_24219_, _24218_, _06114_);
  and _75052_ (_24220_, _24219_, _06111_);
  and _75053_ (_24221_, _24220_, _24216_);
  and _75054_ (_24222_, _07823_, _08708_);
  or _75055_ (_24223_, _24222_, _24185_);
  and _75056_ (_24225_, _24223_, _06110_);
  or _75057_ (_24226_, _24225_, _06297_);
  or _75058_ (_24227_, _24226_, _24221_);
  and _75059_ (_24228_, _14275_, _07823_);
  or _75060_ (_24229_, _24228_, _24185_);
  or _75061_ (_24230_, _24229_, _07127_);
  and _75062_ (_24231_, _24230_, _07125_);
  and _75063_ (_24232_, _24231_, _24227_);
  nor _75064_ (_24233_, _12321_, _11817_);
  or _75065_ (_24234_, _24233_, _24185_);
  and _75066_ (_24236_, _24184_, _06402_);
  and _75067_ (_24237_, _24236_, _24234_);
  or _75068_ (_24238_, _24237_, _24232_);
  and _75069_ (_24239_, _24238_, _07132_);
  nand _75070_ (_24240_, _24223_, _06306_);
  nor _75071_ (_24241_, _24240_, _24193_);
  or _75072_ (_24242_, _24241_, _06411_);
  or _75073_ (_24243_, _24242_, _24239_);
  and _75074_ (_24244_, _24243_, _24187_);
  or _75075_ (_24245_, _24244_, _06303_);
  and _75076_ (_24247_, _14167_, _07823_);
  or _75077_ (_24248_, _24185_, _08819_);
  or _75078_ (_24249_, _24248_, _24247_);
  and _75079_ (_24250_, _24249_, _08824_);
  and _75080_ (_24251_, _24250_, _24245_);
  and _75081_ (_24252_, _24234_, _06396_);
  or _75082_ (_24253_, _24252_, _19287_);
  or _75083_ (_24254_, _24253_, _24251_);
  or _75084_ (_24255_, _24194_, _06630_);
  and _75085_ (_24256_, _24255_, _01317_);
  and _75086_ (_24258_, _24256_, _24254_);
  or _75087_ (_24259_, _24258_, _24183_);
  and _75088_ (_43678_, _24259_, _43100_);
  not _75089_ (_24260_, \oc8051_golden_model_1.TH0 [1]);
  nor _75090_ (_24261_, _01317_, _24260_);
  or _75091_ (_24262_, _14442_, _11817_);
  or _75092_ (_24263_, _07823_, \oc8051_golden_model_1.TH0 [1]);
  and _75093_ (_24264_, _24263_, _05787_);
  and _75094_ (_24265_, _24264_, _24262_);
  and _75095_ (_24266_, _09115_, _07823_);
  nor _75096_ (_24268_, _07823_, _24260_);
  or _75097_ (_24269_, _24268_, _06117_);
  or _75098_ (_24270_, _24269_, _24266_);
  and _75099_ (_24271_, _14363_, _07823_);
  not _75100_ (_24272_, _24271_);
  and _75101_ (_24273_, _24272_, _24263_);
  or _75102_ (_24274_, _24273_, _06161_);
  and _75103_ (_24275_, _07823_, \oc8051_golden_model_1.ACC [1]);
  or _75104_ (_24276_, _24275_, _24268_);
  and _75105_ (_24277_, _24276_, _07056_);
  nor _75106_ (_24279_, _07056_, _24260_);
  or _75107_ (_24280_, _24279_, _06160_);
  or _75108_ (_24281_, _24280_, _24277_);
  and _75109_ (_24282_, _24281_, _07075_);
  and _75110_ (_24283_, _24282_, _24274_);
  and _75111_ (_24284_, _07823_, _07306_);
  or _75112_ (_24285_, _24284_, _24268_);
  and _75113_ (_24286_, _24285_, _06217_);
  or _75114_ (_24287_, _24286_, _24283_);
  and _75115_ (_24288_, _24287_, _06229_);
  and _75116_ (_24290_, _24276_, _06220_);
  or _75117_ (_24291_, _24290_, _09842_);
  or _75118_ (_24292_, _24291_, _24288_);
  or _75119_ (_24293_, _24285_, _06132_);
  and _75120_ (_24294_, _24293_, _24292_);
  or _75121_ (_24295_, _24294_, _06116_);
  and _75122_ (_24296_, _24295_, _06114_);
  and _75123_ (_24297_, _24296_, _24270_);
  or _75124_ (_24298_, _24297_, _24265_);
  and _75125_ (_24299_, _24298_, _06298_);
  or _75126_ (_24301_, _14346_, _11817_);
  and _75127_ (_24302_, _24301_, _06297_);
  nand _75128_ (_24303_, _07823_, _06945_);
  and _75129_ (_24304_, _24303_, _06110_);
  or _75130_ (_24305_, _24304_, _24302_);
  and _75131_ (_24306_, _24305_, _24263_);
  or _75132_ (_24307_, _24306_, _06402_);
  or _75133_ (_24308_, _24307_, _24299_);
  nor _75134_ (_24309_, _10277_, _11817_);
  or _75135_ (_24310_, _24309_, _24268_);
  nand _75136_ (_24312_, _10275_, _07823_);
  and _75137_ (_24313_, _24312_, _24310_);
  or _75138_ (_24314_, _24313_, _07125_);
  and _75139_ (_24315_, _24314_, _07132_);
  and _75140_ (_24316_, _24315_, _24308_);
  or _75141_ (_24317_, _14344_, _11817_);
  and _75142_ (_24318_, _24263_, _06306_);
  and _75143_ (_24319_, _24318_, _24317_);
  or _75144_ (_24320_, _24319_, _06411_);
  or _75145_ (_24321_, _24320_, _24316_);
  nor _75146_ (_24323_, _24268_, _07130_);
  nand _75147_ (_24324_, _24323_, _24312_);
  and _75148_ (_24325_, _24324_, _08819_);
  and _75149_ (_24326_, _24325_, _24321_);
  or _75150_ (_24327_, _24303_, _08176_);
  and _75151_ (_24328_, _24263_, _06303_);
  and _75152_ (_24329_, _24328_, _24327_);
  or _75153_ (_24330_, _24329_, _06396_);
  or _75154_ (_24331_, _24330_, _24326_);
  or _75155_ (_24332_, _24310_, _08824_);
  and _75156_ (_24334_, _24332_, _06829_);
  and _75157_ (_24335_, _24334_, _24331_);
  and _75158_ (_24336_, _24273_, _06433_);
  or _75159_ (_24337_, _24336_, _06440_);
  or _75160_ (_24338_, _24337_, _24335_);
  or _75161_ (_24339_, _24268_, _06444_);
  or _75162_ (_24340_, _24339_, _24271_);
  and _75163_ (_24341_, _24340_, _01317_);
  and _75164_ (_24342_, _24341_, _24338_);
  or _75165_ (_24343_, _24342_, _24261_);
  and _75166_ (_43679_, _24343_, _43100_);
  and _75167_ (_24345_, _01321_, \oc8051_golden_model_1.TH0 [2]);
  and _75168_ (_24346_, _11817_, \oc8051_golden_model_1.TH0 [2]);
  and _75169_ (_24347_, _09211_, _07823_);
  or _75170_ (_24348_, _24347_, _24346_);
  and _75171_ (_24349_, _24348_, _06116_);
  and _75172_ (_24350_, _14542_, _07823_);
  or _75173_ (_24351_, _24350_, _24346_);
  or _75174_ (_24352_, _24351_, _06161_);
  and _75175_ (_24353_, _07823_, \oc8051_golden_model_1.ACC [2]);
  or _75176_ (_24355_, _24353_, _24346_);
  and _75177_ (_24356_, _24355_, _07056_);
  and _75178_ (_24357_, _07057_, \oc8051_golden_model_1.TH0 [2]);
  or _75179_ (_24358_, _24357_, _06160_);
  or _75180_ (_24359_, _24358_, _24356_);
  and _75181_ (_24360_, _24359_, _07075_);
  and _75182_ (_24361_, _24360_, _24352_);
  and _75183_ (_24362_, _07823_, _07708_);
  or _75184_ (_24363_, _24362_, _24346_);
  and _75185_ (_24364_, _24363_, _06217_);
  or _75186_ (_24366_, _24364_, _24361_);
  and _75187_ (_24367_, _24366_, _06229_);
  and _75188_ (_24368_, _24355_, _06220_);
  or _75189_ (_24369_, _24368_, _09842_);
  or _75190_ (_24370_, _24369_, _24367_);
  or _75191_ (_24371_, _24363_, _06132_);
  and _75192_ (_24372_, _24371_, _06117_);
  and _75193_ (_24373_, _24372_, _24370_);
  or _75194_ (_24374_, _24373_, _05787_);
  or _75195_ (_24375_, _24374_, _24349_);
  and _75196_ (_24378_, _14630_, _07823_);
  or _75197_ (_24379_, _24346_, _06114_);
  or _75198_ (_24380_, _24379_, _24378_);
  and _75199_ (_24381_, _24380_, _06111_);
  and _75200_ (_24382_, _24381_, _24375_);
  and _75201_ (_24383_, _07823_, _08768_);
  or _75202_ (_24384_, _24383_, _24346_);
  and _75203_ (_24385_, _24384_, _06110_);
  or _75204_ (_24386_, _24385_, _06297_);
  or _75205_ (_24387_, _24386_, _24382_);
  and _75206_ (_24389_, _14646_, _07823_);
  or _75207_ (_24390_, _24346_, _07127_);
  or _75208_ (_24391_, _24390_, _24389_);
  and _75209_ (_24392_, _24391_, _07125_);
  and _75210_ (_24393_, _24392_, _24387_);
  and _75211_ (_24394_, _10282_, _07823_);
  or _75212_ (_24395_, _24394_, _24346_);
  and _75213_ (_24396_, _24395_, _06402_);
  or _75214_ (_24397_, _24396_, _24393_);
  and _75215_ (_24398_, _24397_, _07132_);
  or _75216_ (_24400_, _24346_, _08248_);
  and _75217_ (_24401_, _24384_, _06306_);
  and _75218_ (_24402_, _24401_, _24400_);
  or _75219_ (_24403_, _24402_, _24398_);
  and _75220_ (_24404_, _24403_, _07130_);
  and _75221_ (_24405_, _24355_, _06411_);
  and _75222_ (_24406_, _24405_, _24400_);
  or _75223_ (_24407_, _24406_, _06303_);
  or _75224_ (_24408_, _24407_, _24404_);
  and _75225_ (_24409_, _14643_, _07823_);
  or _75226_ (_24411_, _24346_, _08819_);
  or _75227_ (_24412_, _24411_, _24409_);
  and _75228_ (_24413_, _24412_, _08824_);
  and _75229_ (_24414_, _24413_, _24408_);
  nor _75230_ (_24415_, _10281_, _11817_);
  or _75231_ (_24416_, _24415_, _24346_);
  and _75232_ (_24417_, _24416_, _06396_);
  or _75233_ (_24418_, _24417_, _24414_);
  and _75234_ (_24419_, _24418_, _06829_);
  and _75235_ (_24420_, _24351_, _06433_);
  or _75236_ (_24422_, _24420_, _06440_);
  or _75237_ (_24423_, _24422_, _24419_);
  and _75238_ (_24424_, _14710_, _07823_);
  or _75239_ (_24425_, _24346_, _06444_);
  or _75240_ (_24426_, _24425_, _24424_);
  and _75241_ (_24427_, _24426_, _01317_);
  and _75242_ (_24428_, _24427_, _24423_);
  or _75243_ (_24429_, _24428_, _24345_);
  and _75244_ (_43680_, _24429_, _43100_);
  and _75245_ (_24430_, _11817_, \oc8051_golden_model_1.TH0 [3]);
  and _75246_ (_24432_, _14738_, _07823_);
  or _75247_ (_24433_, _24432_, _24430_);
  or _75248_ (_24434_, _24433_, _06161_);
  and _75249_ (_24435_, _07823_, \oc8051_golden_model_1.ACC [3]);
  or _75250_ (_24436_, _24435_, _24430_);
  and _75251_ (_24437_, _24436_, _07056_);
  and _75252_ (_24438_, _07057_, \oc8051_golden_model_1.TH0 [3]);
  or _75253_ (_24439_, _24438_, _06160_);
  or _75254_ (_24440_, _24439_, _24437_);
  and _75255_ (_24441_, _24440_, _07075_);
  and _75256_ (_24443_, _24441_, _24434_);
  and _75257_ (_24444_, _07823_, _07544_);
  or _75258_ (_24445_, _24444_, _24430_);
  and _75259_ (_24446_, _24445_, _06217_);
  or _75260_ (_24447_, _24446_, _24443_);
  and _75261_ (_24448_, _24447_, _06229_);
  and _75262_ (_24449_, _24436_, _06220_);
  or _75263_ (_24450_, _24449_, _09842_);
  or _75264_ (_24451_, _24450_, _24448_);
  or _75265_ (_24452_, _24445_, _06132_);
  and _75266_ (_24454_, _24452_, _24451_);
  or _75267_ (_24455_, _24454_, _06116_);
  and _75268_ (_24456_, _09210_, _07823_);
  or _75269_ (_24457_, _24430_, _06117_);
  or _75270_ (_24458_, _24457_, _24456_);
  and _75271_ (_24459_, _24458_, _06114_);
  and _75272_ (_24460_, _24459_, _24455_);
  and _75273_ (_24461_, _14825_, _07823_);
  or _75274_ (_24462_, _24461_, _24430_);
  and _75275_ (_24463_, _24462_, _05787_);
  or _75276_ (_24465_, _24463_, _11136_);
  or _75277_ (_24466_, _24465_, _24460_);
  and _75278_ (_24467_, _14727_, _07823_);
  or _75279_ (_24468_, _24430_, _07127_);
  or _75280_ (_24469_, _24468_, _24467_);
  and _75281_ (_24470_, _07823_, _08712_);
  or _75282_ (_24471_, _24470_, _24430_);
  or _75283_ (_24472_, _24471_, _06111_);
  and _75284_ (_24473_, _24472_, _07125_);
  and _75285_ (_24474_, _24473_, _24469_);
  and _75286_ (_24476_, _24474_, _24466_);
  and _75287_ (_24477_, _12318_, _07823_);
  or _75288_ (_24478_, _24477_, _24430_);
  and _75289_ (_24479_, _24478_, _06402_);
  or _75290_ (_24480_, _24479_, _24476_);
  and _75291_ (_24481_, _24480_, _07132_);
  or _75292_ (_24482_, _24430_, _08140_);
  and _75293_ (_24483_, _24471_, _06306_);
  and _75294_ (_24484_, _24483_, _24482_);
  or _75295_ (_24485_, _24484_, _24481_);
  and _75296_ (_24487_, _24485_, _07130_);
  and _75297_ (_24488_, _24436_, _06411_);
  and _75298_ (_24489_, _24488_, _24482_);
  or _75299_ (_24490_, _24489_, _06303_);
  or _75300_ (_24491_, _24490_, _24487_);
  and _75301_ (_24492_, _14724_, _07823_);
  or _75302_ (_24493_, _24430_, _08819_);
  or _75303_ (_24494_, _24493_, _24492_);
  and _75304_ (_24495_, _24494_, _08824_);
  and _75305_ (_24496_, _24495_, _24491_);
  nor _75306_ (_24498_, _10273_, _11817_);
  or _75307_ (_24499_, _24498_, _24430_);
  and _75308_ (_24500_, _24499_, _06396_);
  or _75309_ (_24501_, _24500_, _06433_);
  or _75310_ (_24502_, _24501_, _24496_);
  or _75311_ (_24503_, _24433_, _06829_);
  and _75312_ (_24504_, _24503_, _06444_);
  and _75313_ (_24505_, _24504_, _24502_);
  and _75314_ (_24506_, _14897_, _07823_);
  or _75315_ (_24507_, _24506_, _24430_);
  and _75316_ (_24509_, _24507_, _06440_);
  or _75317_ (_24510_, _24509_, _01321_);
  or _75318_ (_24511_, _24510_, _24505_);
  or _75319_ (_24512_, _01317_, \oc8051_golden_model_1.TH0 [3]);
  and _75320_ (_24513_, _24512_, _43100_);
  and _75321_ (_43682_, _24513_, _24511_);
  and _75322_ (_24514_, _11817_, \oc8051_golden_model_1.TH0 [4]);
  and _75323_ (_24515_, _08336_, _07823_);
  or _75324_ (_24516_, _24515_, _24514_);
  or _75325_ (_24517_, _24516_, _06132_);
  and _75326_ (_24519_, _14928_, _07823_);
  or _75327_ (_24520_, _24519_, _24514_);
  or _75328_ (_24521_, _24520_, _06161_);
  and _75329_ (_24522_, _07823_, \oc8051_golden_model_1.ACC [4]);
  or _75330_ (_24523_, _24522_, _24514_);
  and _75331_ (_24524_, _24523_, _07056_);
  and _75332_ (_24525_, _07057_, \oc8051_golden_model_1.TH0 [4]);
  or _75333_ (_24526_, _24525_, _06160_);
  or _75334_ (_24527_, _24526_, _24524_);
  and _75335_ (_24528_, _24527_, _07075_);
  and _75336_ (_24530_, _24528_, _24521_);
  and _75337_ (_24531_, _24516_, _06217_);
  or _75338_ (_24532_, _24531_, _24530_);
  and _75339_ (_24533_, _24532_, _06229_);
  and _75340_ (_24534_, _24523_, _06220_);
  or _75341_ (_24535_, _24534_, _09842_);
  or _75342_ (_24536_, _24535_, _24533_);
  and _75343_ (_24537_, _24536_, _24517_);
  or _75344_ (_24538_, _24537_, _06116_);
  and _75345_ (_24539_, _09209_, _07823_);
  or _75346_ (_24541_, _24514_, _06117_);
  or _75347_ (_24542_, _24541_, _24539_);
  and _75348_ (_24543_, _24542_, _06114_);
  and _75349_ (_24544_, _24543_, _24538_);
  and _75350_ (_24545_, _15013_, _07823_);
  or _75351_ (_24546_, _24545_, _24514_);
  and _75352_ (_24547_, _24546_, _05787_);
  or _75353_ (_24548_, _24547_, _24544_);
  or _75354_ (_24549_, _24548_, _11136_);
  and _75355_ (_24550_, _15029_, _07823_);
  or _75356_ (_24552_, _24514_, _07127_);
  or _75357_ (_24553_, _24552_, _24550_);
  and _75358_ (_24554_, _08715_, _07823_);
  or _75359_ (_24555_, _24554_, _24514_);
  or _75360_ (_24556_, _24555_, _06111_);
  and _75361_ (_24557_, _24556_, _07125_);
  and _75362_ (_24558_, _24557_, _24553_);
  and _75363_ (_24559_, _24558_, _24549_);
  and _75364_ (_24560_, _10289_, _07823_);
  or _75365_ (_24561_, _24560_, _24514_);
  and _75366_ (_24563_, _24561_, _06402_);
  or _75367_ (_24564_, _24563_, _24559_);
  and _75368_ (_24565_, _24564_, _07132_);
  or _75369_ (_24566_, _24514_, _08339_);
  and _75370_ (_24567_, _24555_, _06306_);
  and _75371_ (_24568_, _24567_, _24566_);
  or _75372_ (_24569_, _24568_, _24565_);
  and _75373_ (_24570_, _24569_, _07130_);
  and _75374_ (_24571_, _24523_, _06411_);
  and _75375_ (_24572_, _24571_, _24566_);
  or _75376_ (_24574_, _24572_, _06303_);
  or _75377_ (_24575_, _24574_, _24570_);
  and _75378_ (_24576_, _15026_, _07823_);
  or _75379_ (_24577_, _24514_, _08819_);
  or _75380_ (_24578_, _24577_, _24576_);
  and _75381_ (_24579_, _24578_, _08824_);
  and _75382_ (_24580_, _24579_, _24575_);
  nor _75383_ (_24581_, _10288_, _11817_);
  or _75384_ (_24582_, _24581_, _24514_);
  and _75385_ (_24583_, _24582_, _06396_);
  or _75386_ (_24585_, _24583_, _06433_);
  or _75387_ (_24586_, _24585_, _24580_);
  or _75388_ (_24587_, _24520_, _06829_);
  and _75389_ (_24588_, _24587_, _06444_);
  and _75390_ (_24589_, _24588_, _24586_);
  and _75391_ (_24590_, _15087_, _07823_);
  or _75392_ (_24591_, _24590_, _24514_);
  and _75393_ (_24592_, _24591_, _06440_);
  or _75394_ (_24593_, _24592_, _01321_);
  or _75395_ (_24594_, _24593_, _24589_);
  or _75396_ (_24596_, _01317_, \oc8051_golden_model_1.TH0 [4]);
  and _75397_ (_24597_, _24596_, _43100_);
  and _75398_ (_43683_, _24597_, _24594_);
  and _75399_ (_24598_, _11817_, \oc8051_golden_model_1.TH0 [5]);
  and _75400_ (_24599_, _15119_, _07823_);
  or _75401_ (_24600_, _24599_, _24598_);
  or _75402_ (_24601_, _24600_, _06161_);
  and _75403_ (_24602_, _07823_, \oc8051_golden_model_1.ACC [5]);
  or _75404_ (_24603_, _24602_, _24598_);
  and _75405_ (_24604_, _24603_, _07056_);
  and _75406_ (_24605_, _07057_, \oc8051_golden_model_1.TH0 [5]);
  or _75407_ (_24606_, _24605_, _06160_);
  or _75408_ (_24607_, _24606_, _24604_);
  and _75409_ (_24608_, _24607_, _07075_);
  and _75410_ (_24609_, _24608_, _24601_);
  and _75411_ (_24610_, _08101_, _07823_);
  or _75412_ (_24611_, _24610_, _24598_);
  and _75413_ (_24612_, _24611_, _06217_);
  or _75414_ (_24613_, _24612_, _24609_);
  and _75415_ (_24614_, _24613_, _06229_);
  and _75416_ (_24617_, _24603_, _06220_);
  or _75417_ (_24618_, _24617_, _09842_);
  or _75418_ (_24619_, _24618_, _24614_);
  or _75419_ (_24620_, _24611_, _06132_);
  and _75420_ (_24621_, _24620_, _24619_);
  or _75421_ (_24622_, _24621_, _06116_);
  and _75422_ (_24623_, _09208_, _07823_);
  or _75423_ (_24624_, _24598_, _06117_);
  or _75424_ (_24625_, _24624_, _24623_);
  and _75425_ (_24626_, _24625_, _06114_);
  and _75426_ (_24628_, _24626_, _24622_);
  and _75427_ (_24629_, _15203_, _07823_);
  or _75428_ (_24630_, _24629_, _24598_);
  and _75429_ (_24631_, _24630_, _05787_);
  or _75430_ (_24632_, _24631_, _11136_);
  or _75431_ (_24633_, _24632_, _24628_);
  and _75432_ (_24634_, _15219_, _07823_);
  or _75433_ (_24635_, _24598_, _07127_);
  or _75434_ (_24636_, _24635_, _24634_);
  and _75435_ (_24637_, _08736_, _07823_);
  or _75436_ (_24639_, _24637_, _24598_);
  or _75437_ (_24640_, _24639_, _06111_);
  and _75438_ (_24641_, _24640_, _07125_);
  and _75439_ (_24642_, _24641_, _24636_);
  and _75440_ (_24643_, _24642_, _24633_);
  and _75441_ (_24644_, _12325_, _07823_);
  or _75442_ (_24645_, _24644_, _24598_);
  and _75443_ (_24646_, _24645_, _06402_);
  or _75444_ (_24647_, _24646_, _24643_);
  and _75445_ (_24648_, _24647_, _07132_);
  or _75446_ (_24650_, _24598_, _08104_);
  and _75447_ (_24651_, _24639_, _06306_);
  and _75448_ (_24652_, _24651_, _24650_);
  or _75449_ (_24653_, _24652_, _24648_);
  and _75450_ (_24654_, _24653_, _07130_);
  and _75451_ (_24655_, _24603_, _06411_);
  and _75452_ (_24656_, _24655_, _24650_);
  or _75453_ (_24657_, _24656_, _06303_);
  or _75454_ (_24658_, _24657_, _24654_);
  and _75455_ (_24659_, _15216_, _07823_);
  or _75456_ (_24661_, _24598_, _08819_);
  or _75457_ (_24662_, _24661_, _24659_);
  and _75458_ (_24663_, _24662_, _08824_);
  and _75459_ (_24664_, _24663_, _24658_);
  nor _75460_ (_24665_, _10269_, _11817_);
  or _75461_ (_24666_, _24665_, _24598_);
  and _75462_ (_24667_, _24666_, _06396_);
  or _75463_ (_24668_, _24667_, _06433_);
  or _75464_ (_24669_, _24668_, _24664_);
  or _75465_ (_24670_, _24600_, _06829_);
  and _75466_ (_24672_, _24670_, _06444_);
  and _75467_ (_24673_, _24672_, _24669_);
  and _75468_ (_24674_, _15275_, _07823_);
  or _75469_ (_24675_, _24674_, _24598_);
  and _75470_ (_24676_, _24675_, _06440_);
  or _75471_ (_24677_, _24676_, _01321_);
  or _75472_ (_24678_, _24677_, _24673_);
  or _75473_ (_24679_, _01317_, \oc8051_golden_model_1.TH0 [5]);
  and _75474_ (_24680_, _24679_, _43100_);
  and _75475_ (_43684_, _24680_, _24678_);
  and _75476_ (_24682_, _11817_, \oc8051_golden_model_1.TH0 [6]);
  or _75477_ (_24683_, _24682_, _08015_);
  and _75478_ (_24684_, _15402_, _07823_);
  or _75479_ (_24685_, _24684_, _24682_);
  and _75480_ (_24686_, _24685_, _06306_);
  and _75481_ (_24687_, _24686_, _24683_);
  and _75482_ (_24688_, _15300_, _07823_);
  or _75483_ (_24689_, _24688_, _24682_);
  or _75484_ (_24690_, _24689_, _06161_);
  and _75485_ (_24691_, _07823_, \oc8051_golden_model_1.ACC [6]);
  or _75486_ (_24693_, _24691_, _24682_);
  and _75487_ (_24694_, _24693_, _07056_);
  and _75488_ (_24695_, _07057_, \oc8051_golden_model_1.TH0 [6]);
  or _75489_ (_24696_, _24695_, _06160_);
  or _75490_ (_24697_, _24696_, _24694_);
  and _75491_ (_24698_, _24697_, _07075_);
  and _75492_ (_24699_, _24698_, _24690_);
  and _75493_ (_24700_, _08012_, _07823_);
  or _75494_ (_24701_, _24700_, _24682_);
  and _75495_ (_24702_, _24701_, _06217_);
  or _75496_ (_24704_, _24702_, _24699_);
  and _75497_ (_24705_, _24704_, _06229_);
  and _75498_ (_24706_, _24693_, _06220_);
  or _75499_ (_24707_, _24706_, _09842_);
  or _75500_ (_24708_, _24707_, _24705_);
  or _75501_ (_24709_, _24701_, _06132_);
  and _75502_ (_24710_, _24709_, _24708_);
  or _75503_ (_24711_, _24710_, _06116_);
  and _75504_ (_24712_, _09207_, _07823_);
  or _75505_ (_24713_, _24682_, _06117_);
  or _75506_ (_24715_, _24713_, _24712_);
  and _75507_ (_24716_, _24715_, _06114_);
  and _75508_ (_24717_, _24716_, _24711_);
  and _75509_ (_24718_, _15395_, _07823_);
  or _75510_ (_24719_, _24718_, _24682_);
  and _75511_ (_24720_, _24719_, _05787_);
  or _75512_ (_24721_, _24720_, _11136_);
  or _75513_ (_24722_, _24721_, _24717_);
  and _75514_ (_24723_, _15413_, _07823_);
  or _75515_ (_24724_, _24682_, _07127_);
  or _75516_ (_24726_, _24724_, _24723_);
  or _75517_ (_24727_, _24685_, _06111_);
  and _75518_ (_24728_, _24727_, _07125_);
  and _75519_ (_24729_, _24728_, _24726_);
  and _75520_ (_24730_, _24729_, _24722_);
  and _75521_ (_24731_, _10295_, _07823_);
  or _75522_ (_24732_, _24731_, _24682_);
  and _75523_ (_24733_, _24732_, _06402_);
  or _75524_ (_24734_, _24733_, _24730_);
  and _75525_ (_24735_, _24734_, _07132_);
  or _75526_ (_24737_, _24735_, _24687_);
  and _75527_ (_24738_, _24737_, _07130_);
  and _75528_ (_24739_, _24693_, _06411_);
  and _75529_ (_24740_, _24739_, _24683_);
  or _75530_ (_24741_, _24740_, _06303_);
  or _75531_ (_24742_, _24741_, _24738_);
  and _75532_ (_24743_, _15410_, _07823_);
  or _75533_ (_24744_, _24682_, _08819_);
  or _75534_ (_24745_, _24744_, _24743_);
  and _75535_ (_24746_, _24745_, _08824_);
  and _75536_ (_24748_, _24746_, _24742_);
  nor _75537_ (_24749_, _10294_, _11817_);
  or _75538_ (_24750_, _24749_, _24682_);
  and _75539_ (_24751_, _24750_, _06396_);
  or _75540_ (_24752_, _24751_, _06433_);
  or _75541_ (_24753_, _24752_, _24748_);
  or _75542_ (_24754_, _24689_, _06829_);
  and _75543_ (_24755_, _24754_, _06444_);
  and _75544_ (_24756_, _24755_, _24753_);
  and _75545_ (_24757_, _15478_, _07823_);
  or _75546_ (_24759_, _24757_, _24682_);
  and _75547_ (_24760_, _24759_, _06440_);
  or _75548_ (_24761_, _24760_, _01321_);
  or _75549_ (_24762_, _24761_, _24756_);
  or _75550_ (_24763_, _01317_, \oc8051_golden_model_1.TH0 [6]);
  and _75551_ (_24764_, _24763_, _43100_);
  and _75552_ (_43685_, _24764_, _24762_);
  and _75553_ (_24765_, _12744_, _12735_);
  nor _75554_ (_24766_, _24765_, _05444_);
  and _75555_ (_24767_, _12682_, \oc8051_golden_model_1.PC [0]);
  and _75556_ (_24769_, _06758_, \oc8051_golden_model_1.PC [0]);
  nor _75557_ (_24770_, _24769_, _12032_);
  nor _75558_ (_24771_, _24770_, _12682_);
  nor _75559_ (_24772_, _24771_, _24767_);
  and _75560_ (_24773_, _24772_, _05748_);
  and _75561_ (_24774_, _12711_, _12719_);
  nor _75562_ (_24775_, _24774_, _05444_);
  and _75563_ (_24776_, _11905_, _12693_);
  nor _75564_ (_24777_, _24776_, _05444_);
  nor _75565_ (_24778_, _10694_, _05444_);
  and _75566_ (_24780_, _10694_, _05444_);
  nor _75567_ (_24781_, _24780_, _24778_);
  nor _75568_ (_24782_, _24781_, _12539_);
  and _75569_ (_24783_, _11912_, _08819_);
  nor _75570_ (_24784_, _24783_, _05444_);
  and _75571_ (_24785_, _11914_, _07132_);
  nor _75572_ (_24786_, _24785_, _05444_);
  and _75573_ (_24787_, _11919_, _07127_);
  nor _75574_ (_24788_, _24787_, _05444_);
  and _75575_ (_24789_, _06110_, _05444_);
  not _75576_ (_24791_, _05791_);
  nor _75577_ (_24792_, _06758_, _24791_);
  nor _75578_ (_24793_, _06758_, _05769_);
  and _75579_ (_24794_, _06758_, _06581_);
  nor _75580_ (_24795_, _12263_, _05444_);
  nor _75581_ (_24796_, _12266_, _05444_);
  and _75582_ (_24797_, _12266_, _05444_);
  nor _75583_ (_24798_, _24797_, _24796_);
  and _75584_ (_24799_, _12263_, _06582_);
  not _75585_ (_24800_, _24799_);
  nor _75586_ (_24802_, _24800_, _24798_);
  nor _75587_ (_24803_, _24802_, _24795_);
  not _75588_ (_24804_, _24803_);
  nor _75589_ (_24805_, _24804_, _24794_);
  nor _75590_ (_24806_, _24805_, _08445_);
  and _75591_ (_24807_, _12258_, \oc8051_golden_model_1.PC [0]);
  and _75592_ (_24808_, _06107_, _05444_);
  nor _75593_ (_24809_, _24808_, _12200_);
  and _75594_ (_24810_, _24809_, _12256_);
  or _75595_ (_24811_, _24810_, _24807_);
  nor _75596_ (_24813_, _24811_, _08443_);
  nor _75597_ (_24814_, _24813_, _24806_);
  nor _75598_ (_24815_, _24814_, _07064_);
  and _75599_ (_24816_, _07064_, \oc8051_golden_model_1.PC [0]);
  nor _75600_ (_24817_, _24816_, _06160_);
  not _75601_ (_24818_, _24817_);
  nor _75602_ (_24819_, _24818_, _24815_);
  not _75603_ (_24820_, _24819_);
  not _75604_ (_24821_, _12134_);
  not _75605_ (_24822_, _24770_);
  and _75606_ (_24824_, _24822_, _12139_);
  and _75607_ (_24825_, _12141_, \oc8051_golden_model_1.PC [0]);
  or _75608_ (_24826_, _24825_, _06161_);
  nor _75609_ (_24827_, _24826_, _24824_);
  nor _75610_ (_24828_, _24827_, _24821_);
  and _75611_ (_24829_, _24828_, _24820_);
  nor _75612_ (_24830_, _12134_, _05444_);
  nor _75613_ (_24831_, _24830_, _07485_);
  not _75614_ (_24832_, _24831_);
  nor _75615_ (_24833_, _24832_, _24829_);
  nor _75616_ (_24835_, _06758_, _05764_);
  and _75617_ (_24836_, _12300_, _12292_);
  not _75618_ (_24837_, _24836_);
  nor _75619_ (_24838_, _24837_, _24835_);
  not _75620_ (_24839_, _24838_);
  nor _75621_ (_24840_, _24839_, _24833_);
  nor _75622_ (_24841_, _24836_, _05444_);
  nor _75623_ (_24842_, _24841_, _12304_);
  not _75624_ (_24843_, _24842_);
  nor _75625_ (_24844_, _24843_, _24840_);
  nor _75626_ (_24846_, _24844_, _24793_);
  or _75627_ (_24847_, _24846_, _12126_);
  and _75628_ (_24848_, _12120_, \oc8051_golden_model_1.PC [0]);
  nor _75629_ (_24849_, _24770_, _12120_);
  or _75630_ (_24850_, _24849_, _12125_);
  or _75631_ (_24851_, _24850_, _24848_);
  and _75632_ (_24852_, _24851_, _12089_);
  and _75633_ (_24853_, _24852_, _24847_);
  nor _75634_ (_24854_, _24853_, _06236_);
  nor _75635_ (_24855_, _11956_, \oc8051_golden_model_1.PC [0]);
  and _75636_ (_24857_, _24770_, _11956_);
  or _75637_ (_24858_, _24857_, _12089_);
  or _75638_ (_24859_, _24858_, _24855_);
  and _75639_ (_24860_, _24859_, _24854_);
  and _75640_ (_24861_, _12329_, _05444_);
  nor _75641_ (_24862_, _24822_, _12329_);
  nor _75642_ (_24863_, _24862_, _24861_);
  nor _75643_ (_24864_, _24863_, _06643_);
  nor _75644_ (_24865_, _24864_, _24860_);
  nor _75645_ (_24866_, _24865_, _06295_);
  and _75646_ (_24868_, _12346_, _05444_);
  nor _75647_ (_24869_, _24822_, _12346_);
  or _75648_ (_24870_, _24869_, _24868_);
  and _75649_ (_24871_, _24870_, _06295_);
  or _75650_ (_24872_, _24871_, _24866_);
  and _75651_ (_24873_, _24872_, _11925_);
  and _75652_ (_24874_, _11924_, _05444_);
  or _75653_ (_24875_, _24874_, _24873_);
  and _75654_ (_24876_, _24875_, _05760_);
  nor _75655_ (_24877_, _06758_, _05760_);
  nor _75656_ (_24879_, _24877_, _12373_);
  not _75657_ (_24880_, _24879_);
  nor _75658_ (_24881_, _24880_, _24876_);
  not _75659_ (_24882_, _05775_);
  nor _75660_ (_24883_, _12369_, _05444_);
  nor _75661_ (_24884_, _24883_, _24882_);
  not _75662_ (_24885_, _24884_);
  nor _75663_ (_24886_, _24885_, _24881_);
  nor _75664_ (_24887_, _06758_, _05775_);
  and _75665_ (_24888_, _12381_, _05805_);
  not _75666_ (_24890_, _24888_);
  nor _75667_ (_24891_, _24890_, _24887_);
  not _75668_ (_24892_, _24891_);
  nor _75669_ (_24893_, _24892_, _24886_);
  nor _75670_ (_24894_, _24888_, _05444_);
  nor _75671_ (_24895_, _24894_, _05791_);
  not _75672_ (_24896_, _24895_);
  nor _75673_ (_24897_, _24896_, _24893_);
  nor _75674_ (_24898_, _06293_, _05787_);
  and _75675_ (_24899_, _24898_, _11922_);
  not _75676_ (_24901_, _24899_);
  or _75677_ (_24902_, _24901_, _24897_);
  nor _75678_ (_24903_, _24902_, _24792_);
  nor _75679_ (_24904_, _24899_, _05444_);
  nor _75680_ (_24905_, _24904_, _05829_);
  not _75681_ (_24906_, _24905_);
  nor _75682_ (_24907_, _24906_, _24903_);
  nor _75683_ (_24908_, _06758_, _05830_);
  or _75684_ (_24909_, _24908_, _12416_);
  nor _75685_ (_24910_, _24909_, _24907_);
  nor _75686_ (_24912_, _24809_, _12417_);
  nor _75687_ (_24913_, _24912_, _24910_);
  and _75688_ (_24914_, _24913_, _06111_);
  or _75689_ (_24915_, _24914_, _24789_);
  and _75690_ (_24916_, _24915_, _12432_);
  and _75691_ (_24917_, _12431_, _05809_);
  or _75692_ (_24918_, _24917_, _24916_);
  and _75693_ (_24919_, _24918_, _05836_);
  nor _75694_ (_24920_, _06758_, _05836_);
  or _75695_ (_24921_, _24920_, _24919_);
  and _75696_ (_24923_, _24921_, _12474_);
  not _75697_ (_24924_, _24787_);
  nor _75698_ (_24925_, _24809_, _11101_);
  and _75699_ (_24926_, _11101_, _05444_);
  nor _75700_ (_24927_, _24926_, _12474_);
  not _75701_ (_24928_, _24927_);
  nor _75702_ (_24929_, _24928_, _24925_);
  nor _75703_ (_24930_, _24929_, _24924_);
  not _75704_ (_24931_, _24930_);
  nor _75705_ (_24932_, _24931_, _24923_);
  nor _75706_ (_24934_, _24932_, _24788_);
  and _75707_ (_24935_, _24934_, _05834_);
  nor _75708_ (_24936_, _06758_, _05834_);
  or _75709_ (_24937_, _24936_, _24935_);
  and _75710_ (_24938_, _24937_, _12497_);
  not _75711_ (_24939_, _24785_);
  nor _75712_ (_24940_, _24809_, _12480_);
  nor _75713_ (_24941_, _11101_, \oc8051_golden_model_1.PC [0]);
  nor _75714_ (_24942_, _24941_, _12497_);
  not _75715_ (_24943_, _24942_);
  nor _75716_ (_24945_, _24943_, _24940_);
  nor _75717_ (_24946_, _24945_, _24939_);
  not _75718_ (_24947_, _24946_);
  nor _75719_ (_24948_, _24947_, _24938_);
  nor _75720_ (_24949_, _24948_, _24786_);
  and _75721_ (_24950_, _24949_, _05848_);
  nor _75722_ (_24951_, _06758_, _05848_);
  or _75723_ (_24952_, _24951_, _24950_);
  and _75724_ (_24953_, _24952_, _12518_);
  not _75725_ (_24954_, _24783_);
  nor _75726_ (_24956_, _24809_, \oc8051_golden_model_1.PSW [7]);
  and _75727_ (_24957_, \oc8051_golden_model_1.PSW [7], _05444_);
  nor _75728_ (_24958_, _24957_, _12518_);
  not _75729_ (_24959_, _24958_);
  nor _75730_ (_24960_, _24959_, _24956_);
  nor _75731_ (_24961_, _24960_, _24954_);
  not _75732_ (_24962_, _24961_);
  nor _75733_ (_24963_, _24962_, _24953_);
  nor _75734_ (_24964_, _24963_, _24784_);
  and _75735_ (_24965_, _24964_, _05843_);
  nor _75736_ (_24967_, _06758_, _05843_);
  or _75737_ (_24968_, _24967_, _24965_);
  and _75738_ (_24969_, _24968_, _12539_);
  and _75739_ (_24970_, _11907_, _10926_);
  not _75740_ (_24971_, _24970_);
  or _75741_ (_24972_, _24971_, _24969_);
  nor _75742_ (_24973_, _24972_, _24782_);
  nor _75743_ (_24974_, _24970_, _05444_);
  nor _75744_ (_24975_, _24974_, _06417_);
  not _75745_ (_24976_, _24975_);
  nor _75746_ (_24978_, _24976_, _24973_);
  and _75747_ (_24979_, _09160_, _06417_);
  or _75748_ (_24980_, _24979_, _24978_);
  and _75749_ (_24981_, _24980_, _05846_);
  nor _75750_ (_24982_, _06758_, _05846_);
  or _75751_ (_24983_, _24982_, _24981_);
  and _75752_ (_24984_, _24983_, _06421_);
  not _75753_ (_24985_, _24776_);
  and _75754_ (_24986_, _24822_, _12682_);
  nor _75755_ (_24987_, _12682_, _05444_);
  or _75756_ (_24989_, _24987_, _06421_);
  nor _75757_ (_24990_, _24989_, _24986_);
  nor _75758_ (_24991_, _24990_, _24985_);
  not _75759_ (_24992_, _24991_);
  nor _75760_ (_24993_, _24992_, _24984_);
  nor _75761_ (_24994_, _24993_, _24777_);
  and _75762_ (_24995_, _24994_, _06168_);
  and _75763_ (_24996_, _09160_, _06167_);
  or _75764_ (_24997_, _24996_, _24995_);
  and _75765_ (_24998_, _24997_, _12703_);
  nor _75766_ (_25000_, _06758_, _12703_);
  nor _75767_ (_25001_, _25000_, _24998_);
  nor _75768_ (_25002_, _25001_, _06165_);
  not _75769_ (_25003_, _24774_);
  and _75770_ (_25004_, _24772_, _06165_);
  nor _75771_ (_25005_, _25004_, _25003_);
  not _75772_ (_25006_, _25005_);
  nor _75773_ (_25007_, _25006_, _25002_);
  or _75774_ (_25008_, _25007_, _24775_);
  nand _75775_ (_25009_, _25008_, _07160_);
  and _75776_ (_25011_, _07577_, _06758_);
  nor _75777_ (_25012_, _25011_, _05748_);
  nand _75778_ (_25013_, _25012_, _25009_);
  nand _75779_ (_25014_, _25013_, _24765_);
  nor _75780_ (_25015_, _25014_, _24773_);
  or _75781_ (_25016_, _25015_, _24766_);
  nor _75782_ (_25017_, _06305_, _05821_);
  nand _75783_ (_25018_, _25017_, _25016_);
  not _75784_ (_25019_, _25017_);
  and _75785_ (_25020_, _25019_, _06758_);
  nor _75786_ (_25022_, _25020_, _12754_);
  and _75787_ (_25023_, _25022_, _25018_);
  and _75788_ (_25024_, _12754_, _05444_);
  or _75789_ (_25025_, _25024_, _25023_);
  or _75790_ (_25026_, _25025_, _01321_);
  or _75791_ (_25027_, _01317_, \oc8051_golden_model_1.PC [0]);
  and _75792_ (_25028_, _25027_, _43100_);
  and _75793_ (_43687_, _25028_, _25026_);
  and _75794_ (_25029_, _06440_, _05407_);
  and _75795_ (_25030_, _12682_, _05879_);
  nor _75796_ (_25032_, _12034_, _12032_);
  nor _75797_ (_25033_, _25032_, _12035_);
  nor _75798_ (_25034_, _25033_, _12682_);
  nor _75799_ (_25035_, _25034_, _25030_);
  and _75800_ (_25036_, _25035_, _05748_);
  and _75801_ (_25037_, _06433_, _05407_);
  nor _75802_ (_25038_, _08362_, _05879_);
  or _75803_ (_25039_, _11905_, _05879_);
  or _75804_ (_25040_, _11907_, _05879_);
  or _75805_ (_25041_, _11914_, _05879_);
  or _75806_ (_25043_, _11919_, _05879_);
  or _75807_ (_25044_, _08787_, _05407_);
  or _75808_ (_25045_, _12381_, _05879_);
  nor _75809_ (_25046_, _12202_, _12200_);
  nor _75810_ (_25047_, _25046_, _12203_);
  and _75811_ (_25048_, _25047_, _12256_);
  and _75812_ (_25049_, _12258_, _05407_);
  or _75813_ (_25050_, _25049_, _25048_);
  or _75814_ (_25051_, _25050_, _08443_);
  or _75815_ (_25052_, _12263_, _05879_);
  nor _75816_ (_25054_, _06945_, _06582_);
  not _75817_ (_25055_, _12263_);
  and _75818_ (_25056_, _06653_, _05444_);
  nor _75819_ (_25057_, _12265_, _05444_);
  nor _75820_ (_25058_, _25057_, _06545_);
  nor _75821_ (_25059_, _25058_, _25056_);
  or _75822_ (_25060_, _25059_, \oc8051_golden_model_1.PC [1]);
  nand _75823_ (_25061_, _25059_, \oc8051_golden_model_1.PC [1]);
  and _75824_ (_25062_, _25061_, _06582_);
  and _75825_ (_25063_, _25062_, _25060_);
  or _75826_ (_25065_, _25063_, _25055_);
  or _75827_ (_25066_, _25065_, _25054_);
  and _75828_ (_25067_, _25066_, _25052_);
  or _75829_ (_25068_, _25067_, _08445_);
  and _75830_ (_25069_, _25068_, _07065_);
  and _75831_ (_25070_, _25069_, _25051_);
  and _75832_ (_25071_, _07064_, _05879_);
  or _75833_ (_25072_, _25071_, _06160_);
  or _75834_ (_25073_, _25072_, _25070_);
  and _75835_ (_25074_, _25033_, _12139_);
  and _75836_ (_25076_, _12141_, _05878_);
  or _75837_ (_25077_, _25076_, _06161_);
  or _75838_ (_25078_, _25077_, _25074_);
  and _75839_ (_25079_, _25078_, _25073_);
  or _75840_ (_25080_, _25079_, _24821_);
  or _75841_ (_25081_, _12134_, _05879_);
  and _75842_ (_25082_, _25081_, _06157_);
  and _75843_ (_25083_, _25082_, _25080_);
  and _75844_ (_25084_, _06156_, _05407_);
  or _75845_ (_25085_, _25084_, _07485_);
  or _75846_ (_25087_, _25085_, _25083_);
  nand _75847_ (_25088_, _06945_, _07485_);
  and _75848_ (_25089_, _25088_, _07075_);
  and _75849_ (_25090_, _25089_, _25087_);
  nand _75850_ (_25091_, _06217_, _05407_);
  nand _75851_ (_25092_, _25091_, _12292_);
  or _75852_ (_25093_, _25092_, _25090_);
  or _75853_ (_25094_, _12292_, _05879_);
  and _75854_ (_25095_, _25094_, _06229_);
  and _75855_ (_25096_, _25095_, _25093_);
  nand _75856_ (_25098_, _06220_, _05407_);
  nand _75857_ (_25099_, _25098_, _12300_);
  or _75858_ (_25100_, _25099_, _25096_);
  or _75859_ (_25101_, _12300_, _05879_);
  and _75860_ (_25102_, _25101_, _06153_);
  and _75861_ (_25103_, _25102_, _25100_);
  and _75862_ (_25104_, _06152_, _05407_);
  or _75863_ (_25105_, _25104_, _12304_);
  or _75864_ (_25106_, _25105_, _25103_);
  nand _75865_ (_25107_, _06945_, _12304_);
  and _75866_ (_25109_, _25107_, _07191_);
  and _75867_ (_25110_, _25109_, _25106_);
  nand _75868_ (_25111_, _06151_, _05407_);
  nand _75869_ (_25112_, _25111_, _12125_);
  or _75870_ (_25113_, _25112_, _25110_);
  nor _75871_ (_25114_, _06687_, _06236_);
  or _75872_ (_25115_, _25033_, _12120_);
  nand _75873_ (_25116_, _12120_, _05879_);
  and _75874_ (_25117_, _25116_, _25115_);
  or _75875_ (_25118_, _25117_, _12125_);
  and _75876_ (_25120_, _25118_, _25114_);
  and _75877_ (_25121_, _25120_, _25113_);
  and _75878_ (_25122_, _12329_, _05878_);
  not _75879_ (_25123_, _12329_);
  and _75880_ (_25124_, _25033_, _25123_);
  or _75881_ (_25125_, _25124_, _25122_);
  and _75882_ (_25126_, _25125_, _06236_);
  and _75883_ (_25127_, _11958_, _05878_);
  and _75884_ (_25128_, _25033_, _11956_);
  or _75885_ (_25129_, _25128_, _25127_);
  and _75886_ (_25131_, _25129_, _06687_);
  or _75887_ (_25132_, _25131_, _25126_);
  or _75888_ (_25133_, _25132_, _25121_);
  and _75889_ (_25134_, _25133_, _12317_);
  or _75890_ (_25135_, _25033_, _12346_);
  nand _75891_ (_25136_, _12346_, _05879_);
  and _75892_ (_25137_, _25136_, _06295_);
  and _75893_ (_25138_, _25137_, _25135_);
  or _75894_ (_25139_, _25138_, _11924_);
  or _75895_ (_25140_, _25139_, _25134_);
  nand _75896_ (_25142_, _11924_, _05878_);
  and _75897_ (_25143_, _25142_, _25140_);
  or _75898_ (_25144_, _25143_, _06145_);
  nand _75899_ (_25145_, _06145_, \oc8051_golden_model_1.PC [1]);
  and _75900_ (_25146_, _25145_, _05760_);
  and _75901_ (_25147_, _25146_, _25144_);
  nor _75902_ (_25148_, _06945_, _05760_);
  nor _75903_ (_25149_, _07292_, _06701_);
  and _75904_ (_25150_, _25149_, _12359_);
  and _75905_ (_25151_, _25150_, _12356_);
  not _75906_ (_25152_, _25151_);
  or _75907_ (_25153_, _25152_, _25148_);
  or _75908_ (_25154_, _25153_, _25147_);
  or _75909_ (_25155_, _25151_, _05407_);
  and _75910_ (_25156_, _25155_, _12367_);
  and _75911_ (_25157_, _25156_, _25154_);
  nand _75912_ (_25158_, _12366_, _05879_);
  nand _75913_ (_25159_, _25158_, _12368_);
  or _75914_ (_25160_, _25159_, _25157_);
  or _75915_ (_25161_, _12368_, _05879_);
  and _75916_ (_25164_, _25161_, _13844_);
  and _75917_ (_25165_, _25164_, _25160_);
  and _75918_ (_25166_, _06255_, _05407_);
  or _75919_ (_25167_, _25166_, _24882_);
  or _75920_ (_25168_, _25167_, _25165_);
  nand _75921_ (_25169_, _06945_, _24882_);
  and _75922_ (_25170_, _25169_, _13843_);
  and _75923_ (_25171_, _25170_, _25168_);
  or _75924_ (_25172_, _12379_, _10545_);
  and _75925_ (_25173_, _06254_, _05407_);
  nor _75926_ (_25175_, _25173_, _25172_);
  nand _75927_ (_25176_, _25175_, _10553_);
  or _75928_ (_25177_, _25176_, _25171_);
  and _75929_ (_25178_, _25177_, _25045_);
  or _75930_ (_25179_, _25178_, _12386_);
  or _75931_ (_25180_, _12385_, _05407_);
  and _75932_ (_25181_, _25180_, _05805_);
  and _75933_ (_25182_, _25181_, _25179_);
  nor _75934_ (_25183_, _05878_, _05805_);
  or _75935_ (_25184_, _25183_, _06139_);
  or _75936_ (_25186_, _25184_, _25182_);
  nand _75937_ (_25187_, _06139_, \oc8051_golden_model_1.PC [1]);
  and _75938_ (_25188_, _25187_, _25186_);
  or _75939_ (_25189_, _25188_, _05791_);
  nand _75940_ (_25190_, _06945_, _05791_);
  and _75941_ (_25191_, _25190_, _11296_);
  and _75942_ (_25192_, _25191_, _25189_);
  nand _75943_ (_25193_, _06293_, _05878_);
  nand _75944_ (_25194_, _25193_, _06133_);
  or _75945_ (_25195_, _25194_, _25192_);
  or _75946_ (_25197_, _06133_, _05407_);
  and _75947_ (_25198_, _25197_, _06114_);
  and _75948_ (_25199_, _25198_, _25195_);
  nand _75949_ (_25200_, _05878_, _05787_);
  nand _75950_ (_25201_, _25200_, _11922_);
  or _75951_ (_25202_, _25201_, _25199_);
  or _75952_ (_25203_, _11922_, _05879_);
  and _75953_ (_25204_, _25203_, _06762_);
  and _75954_ (_25205_, _25204_, _25202_);
  and _75955_ (_25206_, _06209_, _05407_);
  or _75956_ (_25208_, _25206_, _05829_);
  or _75957_ (_25209_, _25208_, _25205_);
  nand _75958_ (_25210_, _06945_, _05829_);
  and _75959_ (_25211_, _25210_, _12417_);
  and _75960_ (_25212_, _25211_, _25209_);
  and _75961_ (_25213_, _25047_, _12416_);
  or _75962_ (_25214_, _25213_, _08788_);
  or _75963_ (_25215_, _25214_, _25212_);
  and _75964_ (_25216_, _25215_, _25044_);
  or _75965_ (_25217_, _25216_, _06110_);
  nand _75966_ (_25219_, _06110_, _05879_);
  and _75967_ (_25220_, _25219_, _10752_);
  and _75968_ (_25221_, _25220_, _25217_);
  and _75969_ (_25222_, _10751_, _05407_);
  or _75970_ (_25223_, _25222_, _12431_);
  or _75971_ (_25224_, _25223_, _25221_);
  or _75972_ (_25225_, _12432_, _05876_);
  and _75973_ (_25226_, _25225_, _06768_);
  and _75974_ (_25227_, _25226_, _25224_);
  and _75975_ (_25228_, _06208_, _05407_);
  or _75976_ (_25230_, _25228_, _06076_);
  or _75977_ (_25231_, _25230_, _25227_);
  nand _75978_ (_25232_, _06945_, _06076_);
  and _75979_ (_25233_, _25232_, _12474_);
  and _75980_ (_25234_, _25233_, _25231_);
  or _75981_ (_25235_, _25047_, _11101_);
  nand _75982_ (_25236_, _11101_, \oc8051_golden_model_1.PC [1]);
  and _75983_ (_25237_, _25236_, _12473_);
  and _75984_ (_25238_, _25237_, _25235_);
  or _75985_ (_25239_, _25238_, _12478_);
  or _75986_ (_25241_, _25239_, _25234_);
  and _75987_ (_25242_, _25241_, _25043_);
  or _75988_ (_25243_, _25242_, _11917_);
  or _75989_ (_25244_, _11916_, _05407_);
  and _75990_ (_25245_, _25244_, _07127_);
  and _75991_ (_25246_, _25245_, _25243_);
  and _75992_ (_25247_, _06297_, _05878_);
  or _75993_ (_25248_, _25247_, _06402_);
  or _75994_ (_25249_, _25248_, _25246_);
  nand _75995_ (_25250_, _06402_, \oc8051_golden_model_1.PC [1]);
  and _75996_ (_25252_, _25250_, _25249_);
  or _75997_ (_25253_, _25252_, _12492_);
  nand _75998_ (_25254_, _06945_, _12492_);
  and _75999_ (_25255_, _25254_, _12497_);
  and _76000_ (_25256_, _25255_, _25253_);
  or _76001_ (_25257_, _25047_, _12480_);
  or _76002_ (_25258_, _11101_, _05407_);
  and _76003_ (_25259_, _25258_, _12496_);
  and _76004_ (_25260_, _25259_, _25257_);
  or _76005_ (_25261_, _25260_, _12505_);
  or _76006_ (_25263_, _25261_, _25256_);
  and _76007_ (_25264_, _25263_, _25041_);
  or _76008_ (_25265_, _25264_, _10822_);
  or _76009_ (_25266_, _10821_, _05407_);
  and _76010_ (_25267_, _25266_, _07132_);
  and _76011_ (_25268_, _25267_, _25265_);
  and _76012_ (_25269_, _06306_, _05878_);
  or _76013_ (_25270_, _25269_, _06411_);
  or _76014_ (_25271_, _25270_, _25268_);
  nand _76015_ (_25272_, _06411_, \oc8051_golden_model_1.PC [1]);
  and _76016_ (_25274_, _25272_, _25271_);
  or _76017_ (_25275_, _25274_, _07124_);
  nand _76018_ (_25276_, _06945_, _07124_);
  and _76019_ (_25277_, _25276_, _12518_);
  and _76020_ (_25278_, _25277_, _25275_);
  or _76021_ (_25279_, _25047_, \oc8051_golden_model_1.PSW [7]);
  nand _76022_ (_25280_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and _76023_ (_25281_, _25280_, _12517_);
  and _76024_ (_25282_, _25281_, _25279_);
  or _76025_ (_25283_, _25282_, _25278_);
  and _76026_ (_25285_, _25283_, _11910_);
  nor _76027_ (_25286_, _10466_, _06783_);
  and _76028_ (_25287_, _11909_, _05879_);
  or _76029_ (_25288_, _25287_, _25286_);
  or _76030_ (_25289_, _25288_, _25285_);
  and _76031_ (_25290_, _06281_, _05840_);
  and _76032_ (_25291_, _25286_, _05878_);
  nor _76033_ (_25292_, _25291_, _25290_);
  and _76034_ (_25293_, _25292_, _25289_);
  nand _76035_ (_25294_, _25290_, _05879_);
  nand _76036_ (_25296_, _25294_, _10849_);
  or _76037_ (_25297_, _25296_, _25293_);
  or _76038_ (_25298_, _10849_, _05407_);
  and _76039_ (_25299_, _25298_, _08819_);
  and _76040_ (_25300_, _25299_, _25297_);
  nand _76041_ (_25301_, _06303_, _05878_);
  nand _76042_ (_25302_, _25301_, _12535_);
  or _76043_ (_25303_, _25302_, _25300_);
  nand _76044_ (_25304_, _06945_, _05842_);
  and _76045_ (_25305_, _25304_, _12539_);
  or _76046_ (_25307_, _05842_, _05407_);
  or _76047_ (_25308_, _25307_, _08824_);
  and _76048_ (_25309_, _25308_, _25305_);
  and _76049_ (_25310_, _25309_, _25303_);
  or _76050_ (_25311_, _25047_, _10693_);
  or _76051_ (_25312_, \oc8051_golden_model_1.PSW [7], _05407_);
  and _76052_ (_25313_, _25312_, _12538_);
  and _76053_ (_25314_, _25313_, _25311_);
  or _76054_ (_25315_, _25314_, _12547_);
  or _76055_ (_25316_, _25315_, _25310_);
  and _76056_ (_25318_, _25316_, _25040_);
  or _76057_ (_25319_, _25318_, _10897_);
  or _76058_ (_25320_, _10896_, _05407_);
  and _76059_ (_25321_, _25320_, _10926_);
  and _76060_ (_25322_, _25321_, _25319_);
  and _76061_ (_25323_, _10925_, _05879_);
  or _76062_ (_25324_, _25323_, _06417_);
  or _76063_ (_25325_, _25324_, _25322_);
  or _76064_ (_25326_, _09115_, _12558_);
  and _76065_ (_25327_, _25326_, _25325_);
  or _76066_ (_25329_, _25327_, _07142_);
  nand _76067_ (_25330_, _06945_, _07142_);
  and _76068_ (_25331_, _25330_, _06421_);
  and _76069_ (_25332_, _25331_, _25329_);
  not _76070_ (_25333_, _12682_);
  or _76071_ (_25334_, _25033_, _25333_);
  or _76072_ (_25335_, _12682_, _05878_);
  and _76073_ (_25336_, _25335_, _06301_);
  and _76074_ (_25337_, _25336_, _25334_);
  or _76075_ (_25338_, _25337_, _12565_);
  or _76076_ (_25340_, _25338_, _25332_);
  nand _76077_ (_25341_, _25340_, _25039_);
  nand _76078_ (_25342_, _25341_, _12690_);
  nor _76079_ (_25343_, _12690_, _05407_);
  nor _76080_ (_25344_, _25343_, _10262_);
  nand _76081_ (_25345_, _25344_, _25342_);
  and _76082_ (_25346_, _10262_, _05879_);
  nor _76083_ (_25347_, _25346_, _06167_);
  and _76084_ (_25348_, _25347_, _25345_);
  and _76085_ (_25349_, _11935_, _06167_);
  or _76086_ (_25351_, _25349_, _25348_);
  nand _76087_ (_25352_, _25351_, _12703_);
  and _76088_ (_25353_, _06945_, _05826_);
  nor _76089_ (_25354_, _25353_, _06165_);
  nand _76090_ (_25355_, _25354_, _25352_);
  not _76091_ (_25356_, _08362_);
  and _76092_ (_25357_, _25035_, _06165_);
  nor _76093_ (_25358_, _25357_, _25356_);
  and _76094_ (_25359_, _25358_, _25355_);
  or _76095_ (_25360_, _25359_, _25038_);
  nand _76096_ (_25362_, _25360_, _07154_);
  and _76097_ (_25363_, _07153_, _05878_);
  nor _76098_ (_25364_, _25363_, _06433_);
  and _76099_ (_25365_, _25364_, _25362_);
  or _76100_ (_25366_, _25365_, _25037_);
  nand _76101_ (_25367_, _25366_, _12719_);
  nor _76102_ (_25368_, _12719_, _05878_);
  nor _76103_ (_25369_, _25368_, _07577_);
  nand _76104_ (_25370_, _25369_, _25367_);
  and _76105_ (_25371_, _07577_, _06945_);
  nor _76106_ (_25373_, _25371_, _05748_);
  and _76107_ (_25374_, _25373_, _25370_);
  or _76108_ (_25375_, _25374_, _25036_);
  and _76109_ (_25376_, _25375_, _09193_);
  nor _76110_ (_25377_, _07168_, _05879_);
  nor _76111_ (_25378_, _25377_, _12735_);
  or _76112_ (_25379_, _25378_, _25376_);
  and _76113_ (_25380_, _07168_, _05878_);
  nor _76114_ (_25381_, _25380_, _06440_);
  and _76115_ (_25382_, _25381_, _25379_);
  or _76116_ (_25384_, _25382_, _25029_);
  nand _76117_ (_25385_, _25384_, _12744_);
  nor _76118_ (_25386_, _12744_, _05878_);
  nor _76119_ (_25387_, _25386_, _25019_);
  nand _76120_ (_25388_, _25387_, _25385_);
  and _76121_ (_25389_, _25019_, _06945_);
  nor _76122_ (_25390_, _25389_, _12754_);
  and _76123_ (_25391_, _25390_, _25388_);
  and _76124_ (_25392_, _12754_, _05879_);
  or _76125_ (_25393_, _25392_, _25391_);
  or _76126_ (_25395_, _25393_, _01321_);
  or _76127_ (_25396_, _01317_, \oc8051_golden_model_1.PC [1]);
  and _76128_ (_25397_, _25396_, _43100_);
  and _76129_ (_43689_, _25397_, _25395_);
  and _76130_ (_25398_, _06440_, _05921_);
  nor _76131_ (_25399_, _11905_, _05907_);
  and _76132_ (_25400_, _09070_, _06417_);
  nor _76133_ (_25401_, _11907_, _05907_);
  nor _76134_ (_25402_, _11912_, _05907_);
  nor _76135_ (_25403_, _11914_, _05907_);
  nor _76136_ (_25405_, _11919_, _05907_);
  nor _76137_ (_25406_, _11922_, _05907_);
  nor _76138_ (_25407_, _06131_, _05921_);
  not _76139_ (_25408_, _05907_);
  and _76140_ (_25409_, _11924_, _25408_);
  or _76141_ (_25410_, _12028_, _11956_);
  and _76142_ (_25411_, _12039_, _12036_);
  nor _76143_ (_25412_, _25411_, _12040_);
  or _76144_ (_25413_, _25412_, _11958_);
  nand _76145_ (_25414_, _25413_, _25410_);
  nand _76146_ (_25415_, _25414_, _06687_);
  and _76147_ (_25416_, _06581_, _06521_);
  nor _76148_ (_25417_, _12263_, _05907_);
  or _76149_ (_25418_, _12265_, _25408_);
  nand _76150_ (_25419_, _12266_, \oc8051_golden_model_1.PC [2]);
  and _76151_ (_25420_, _25419_, _25418_);
  or _76152_ (_25421_, _25420_, _07056_);
  and _76153_ (_25422_, _06653_, _05907_);
  and _76154_ (_25423_, _07056_, _05921_);
  nor _76155_ (_25424_, _25423_, _25422_);
  and _76156_ (_25427_, _25424_, _24799_);
  and _76157_ (_25428_, _25427_, _25421_);
  or _76158_ (_25429_, _25428_, _25417_);
  nor _76159_ (_25430_, _25429_, _25416_);
  nor _76160_ (_25431_, _25430_, _08445_);
  and _76161_ (_25432_, _12207_, _12204_);
  nor _76162_ (_25433_, _25432_, _12208_);
  nand _76163_ (_25434_, _25433_, _12256_);
  or _76164_ (_25435_, _12256_, _05923_);
  and _76165_ (_25436_, _25435_, _08445_);
  and _76166_ (_25438_, _25436_, _25434_);
  or _76167_ (_25439_, _25438_, _25431_);
  nand _76168_ (_25440_, _25439_, _07065_);
  and _76169_ (_25441_, _07064_, _25408_);
  nor _76170_ (_25442_, _25441_, _06160_);
  nand _76171_ (_25443_, _25442_, _25440_);
  or _76172_ (_25444_, _25412_, _12141_);
  or _76173_ (_25445_, _12139_, _12028_);
  and _76174_ (_25446_, _25445_, _06160_);
  nand _76175_ (_25447_, _25446_, _25444_);
  and _76176_ (_25449_, _25447_, _12134_);
  nand _76177_ (_25450_, _25449_, _25443_);
  nor _76178_ (_25451_, _12134_, _05907_);
  nor _76179_ (_25452_, _25451_, _06156_);
  nand _76180_ (_25453_, _25452_, _25450_);
  and _76181_ (_25454_, _06156_, _05921_);
  nor _76182_ (_25455_, _25454_, _07485_);
  nand _76183_ (_25456_, _25455_, _25453_);
  and _76184_ (_25457_, _06521_, _07485_);
  nor _76185_ (_25458_, _25457_, _06217_);
  nand _76186_ (_25460_, _25458_, _25456_);
  and _76187_ (_25461_, _06217_, _05921_);
  nor _76188_ (_25462_, _25461_, _12293_);
  nand _76189_ (_25463_, _25462_, _25460_);
  nor _76190_ (_25464_, _12292_, _05907_);
  nor _76191_ (_25465_, _25464_, _06220_);
  nand _76192_ (_25466_, _25465_, _25463_);
  and _76193_ (_25467_, _06220_, _05921_);
  nor _76194_ (_25468_, _25467_, _12302_);
  nand _76195_ (_25469_, _25468_, _25466_);
  nor _76196_ (_25471_, _12300_, _05907_);
  nor _76197_ (_25472_, _25471_, _06152_);
  nand _76198_ (_25473_, _25472_, _25469_);
  and _76199_ (_25474_, _06152_, _05921_);
  nor _76200_ (_25475_, _25474_, _12304_);
  nand _76201_ (_25476_, _25475_, _25473_);
  and _76202_ (_25477_, _06521_, _12304_);
  nor _76203_ (_25478_, _25477_, _06151_);
  nand _76204_ (_25479_, _25478_, _25476_);
  and _76205_ (_25480_, _06151_, _05921_);
  nor _76206_ (_25482_, _25480_, _12126_);
  and _76207_ (_25483_, _25482_, _25479_);
  not _76208_ (_25484_, _25412_);
  nor _76209_ (_25485_, _25484_, _12120_);
  not _76210_ (_25486_, _25485_);
  and _76211_ (_25487_, _12120_, _12028_);
  nor _76212_ (_25488_, _25487_, _12125_);
  and _76213_ (_25489_, _25488_, _25486_);
  or _76214_ (_25490_, _25489_, _25483_);
  nand _76215_ (_25491_, _25490_, _12089_);
  nand _76216_ (_25493_, _25491_, _25415_);
  nand _76217_ (_25494_, _25493_, _06643_);
  and _76218_ (_25495_, _12329_, _12028_);
  not _76219_ (_25496_, _25495_);
  nor _76220_ (_25497_, _25484_, _12329_);
  nor _76221_ (_25498_, _25497_, _06643_);
  and _76222_ (_25499_, _25498_, _25496_);
  nor _76223_ (_25500_, _25499_, _06295_);
  nand _76224_ (_25501_, _25500_, _25494_);
  nor _76225_ (_25502_, _25412_, _12346_);
  and _76226_ (_25504_, _12346_, _12029_);
  or _76227_ (_25505_, _25504_, _12317_);
  or _76228_ (_25506_, _25505_, _25502_);
  and _76229_ (_25507_, _25506_, _11925_);
  and _76230_ (_25508_, _25507_, _25501_);
  or _76231_ (_25509_, _25508_, _25409_);
  nand _76232_ (_25510_, _25509_, _06146_);
  and _76233_ (_25511_, _06145_, _05923_);
  nor _76234_ (_25512_, _25511_, _07388_);
  nand _76235_ (_25513_, _25512_, _25510_);
  nor _76236_ (_25515_, _06521_, _05760_);
  nor _76237_ (_25516_, _25515_, _25152_);
  and _76238_ (_25517_, _25516_, _25513_);
  nor _76239_ (_25518_, _25151_, _05921_);
  or _76240_ (_25519_, _25518_, _25517_);
  nand _76241_ (_25520_, _25519_, _12369_);
  nor _76242_ (_25521_, _12369_, _05907_);
  nor _76243_ (_25522_, _25521_, _06255_);
  nand _76244_ (_25523_, _25522_, _25520_);
  and _76245_ (_25524_, _06255_, _05921_);
  nor _76246_ (_25526_, _25524_, _24882_);
  nand _76247_ (_25527_, _25526_, _25523_);
  and _76248_ (_25528_, _06521_, _24882_);
  nor _76249_ (_25529_, _25528_, _06254_);
  nand _76250_ (_25530_, _25529_, _25527_);
  and _76251_ (_25531_, _06254_, _05921_);
  nor _76252_ (_25532_, _25531_, _12387_);
  and _76253_ (_25533_, _25532_, _25530_);
  nor _76254_ (_25534_, _12381_, _05907_);
  or _76255_ (_25535_, _25534_, _25533_);
  nand _76256_ (_25537_, _25535_, _12385_);
  nor _76257_ (_25538_, _12385_, _05921_);
  nor _76258_ (_25539_, _25538_, _05870_);
  nand _76259_ (_25540_, _25539_, _25537_);
  nor _76260_ (_25541_, _25408_, _05805_);
  nor _76261_ (_25542_, _25541_, _06139_);
  and _76262_ (_25543_, _25542_, _25540_);
  and _76263_ (_25544_, _06139_, _05923_);
  or _76264_ (_25545_, _25544_, _25543_);
  nand _76265_ (_25546_, _25545_, _24791_);
  and _76266_ (_25548_, _06521_, _05791_);
  nor _76267_ (_25549_, _25548_, _06293_);
  nand _76268_ (_25550_, _25549_, _25546_);
  and _76269_ (_25551_, _12028_, _06293_);
  not _76270_ (_25552_, _25551_);
  and _76271_ (_25553_, _25552_, _06131_);
  and _76272_ (_25554_, _25553_, _25550_);
  nor _76273_ (_25555_, _25554_, _25407_);
  nor _76274_ (_25556_, _07365_, _05797_);
  or _76275_ (_25557_, _25556_, _25555_);
  and _76276_ (_25559_, _25556_, _05923_);
  nor _76277_ (_25560_, _25559_, _05787_);
  nand _76278_ (_25561_, _25560_, _25557_);
  and _76279_ (_25562_, _12028_, _05787_);
  nor _76280_ (_25563_, _25562_, _12412_);
  and _76281_ (_25564_, _25563_, _25561_);
  or _76282_ (_25565_, _25564_, _25406_);
  and _76283_ (_25566_, _25565_, _06762_);
  and _76284_ (_25567_, _06209_, _05923_);
  or _76285_ (_25568_, _25567_, _05829_);
  or _76286_ (_25570_, _25568_, _25566_);
  nor _76287_ (_25571_, _06521_, _05830_);
  nor _76288_ (_25572_, _25571_, _12416_);
  and _76289_ (_25573_, _25572_, _25570_);
  nor _76290_ (_25574_, _25433_, _12417_);
  or _76291_ (_25575_, _25574_, _25573_);
  nand _76292_ (_25576_, _25575_, _07352_);
  and _76293_ (_25577_, _07351_, _05923_);
  not _76294_ (_25578_, _25577_);
  and _76295_ (_25579_, _25578_, _08786_);
  nand _76296_ (_25581_, _25579_, _25576_);
  nor _76297_ (_25582_, _08786_, _05923_);
  nor _76298_ (_25583_, _25582_, _06110_);
  nand _76299_ (_25584_, _25583_, _25581_);
  and _76300_ (_25585_, _12029_, _06110_);
  nor _76301_ (_25586_, _25585_, _10751_);
  nand _76302_ (_25587_, _25586_, _25584_);
  and _76303_ (_25588_, _10751_, _05921_);
  nor _76304_ (_25589_, _25588_, _12431_);
  nand _76305_ (_25590_, _25589_, _25587_);
  and _76306_ (_25592_, _12431_, _05936_);
  nor _76307_ (_25593_, _25592_, _06208_);
  nand _76308_ (_25594_, _25593_, _25590_);
  and _76309_ (_25595_, _06208_, _05921_);
  nor _76310_ (_25596_, _25595_, _06076_);
  nand _76311_ (_25597_, _25596_, _25594_);
  and _76312_ (_25598_, _06521_, _06076_);
  nor _76313_ (_25599_, _25598_, _12473_);
  nand _76314_ (_25600_, _25599_, _25597_);
  and _76315_ (_25601_, _11101_, _05923_);
  nor _76316_ (_25603_, _25433_, _11101_);
  or _76317_ (_25604_, _25603_, _12474_);
  or _76318_ (_25605_, _25604_, _25601_);
  and _76319_ (_25606_, _25605_, _11919_);
  and _76320_ (_25607_, _25606_, _25600_);
  or _76321_ (_25608_, _25607_, _25405_);
  nand _76322_ (_25609_, _25608_, _11916_);
  nor _76323_ (_25610_, _11916_, _05921_);
  nor _76324_ (_25611_, _25610_, _06297_);
  nand _76325_ (_25612_, _25611_, _25609_);
  and _76326_ (_25614_, _12028_, _06297_);
  nor _76327_ (_25615_, _25614_, _06402_);
  and _76328_ (_25616_, _25615_, _25612_);
  and _76329_ (_25617_, _06402_, _05923_);
  or _76330_ (_25618_, _25617_, _25616_);
  nand _76331_ (_25619_, _25618_, _05834_);
  and _76332_ (_25620_, _06521_, _12492_);
  nor _76333_ (_25621_, _25620_, _12496_);
  nand _76334_ (_25622_, _25621_, _25619_);
  nor _76335_ (_25623_, _11101_, _05921_);
  nor _76336_ (_25625_, _25433_, _12480_);
  or _76337_ (_25626_, _25625_, _12497_);
  or _76338_ (_25627_, _25626_, _25623_);
  and _76339_ (_25628_, _25627_, _11914_);
  and _76340_ (_25629_, _25628_, _25622_);
  or _76341_ (_25630_, _25629_, _25403_);
  nand _76342_ (_25631_, _25630_, _10821_);
  nor _76343_ (_25632_, _10821_, _05921_);
  nor _76344_ (_25633_, _25632_, _06306_);
  nand _76345_ (_25634_, _25633_, _25631_);
  and _76346_ (_25636_, _12028_, _06306_);
  nor _76347_ (_25637_, _25636_, _06411_);
  and _76348_ (_25638_, _25637_, _25634_);
  and _76349_ (_25639_, _06411_, _05923_);
  or _76350_ (_25640_, _25639_, _25638_);
  nand _76351_ (_25641_, _25640_, _05848_);
  and _76352_ (_25642_, _06521_, _07124_);
  nor _76353_ (_25643_, _25642_, _12517_);
  nand _76354_ (_25644_, _25643_, _25641_);
  nor _76355_ (_25645_, _25433_, \oc8051_golden_model_1.PSW [7]);
  nor _76356_ (_25647_, _05921_, _10693_);
  nor _76357_ (_25648_, _25647_, _12518_);
  not _76358_ (_25649_, _25648_);
  nor _76359_ (_25650_, _25649_, _25645_);
  nor _76360_ (_25651_, _25650_, _12522_);
  and _76361_ (_25652_, _25651_, _25644_);
  or _76362_ (_25653_, _25652_, _25402_);
  nand _76363_ (_25654_, _25653_, _10849_);
  nor _76364_ (_25655_, _10849_, _05921_);
  nor _76365_ (_25656_, _25655_, _06303_);
  and _76366_ (_25658_, _25656_, _25654_);
  and _76367_ (_25659_, _12028_, _06303_);
  or _76368_ (_25660_, _25659_, _06396_);
  nor _76369_ (_25661_, _25660_, _25658_);
  and _76370_ (_25662_, _06396_, _05923_);
  or _76371_ (_25663_, _25662_, _25661_);
  nand _76372_ (_25664_, _25663_, _05843_);
  and _76373_ (_25665_, _06521_, _05842_);
  nor _76374_ (_25666_, _25665_, _12538_);
  nand _76375_ (_25667_, _25666_, _25664_);
  or _76376_ (_25669_, _25433_, _10693_);
  or _76377_ (_25670_, _05921_, \oc8051_golden_model_1.PSW [7]);
  and _76378_ (_25671_, _25670_, _12538_);
  and _76379_ (_25672_, _25671_, _25669_);
  nor _76380_ (_25673_, _25672_, _12547_);
  and _76381_ (_25674_, _25673_, _25667_);
  or _76382_ (_25675_, _25674_, _25401_);
  nand _76383_ (_25676_, _25675_, _10896_);
  nor _76384_ (_25677_, _10896_, _05921_);
  nor _76385_ (_25678_, _25677_, _10925_);
  nand _76386_ (_25680_, _25678_, _25676_);
  and _76387_ (_25681_, _10925_, _05907_);
  nor _76388_ (_25682_, _25681_, _06417_);
  and _76389_ (_25683_, _25682_, _25680_);
  or _76390_ (_25684_, _25683_, _25400_);
  nand _76391_ (_25685_, _25684_, _05846_);
  and _76392_ (_25686_, _06521_, _07142_);
  nor _76393_ (_25687_, _25686_, _06301_);
  nand _76394_ (_25688_, _25687_, _25685_);
  nor _76395_ (_25689_, _12028_, _12682_);
  and _76396_ (_25691_, _25484_, _12682_);
  or _76397_ (_25692_, _25691_, _06421_);
  nor _76398_ (_25693_, _25692_, _25689_);
  nor _76399_ (_25694_, _25693_, _12565_);
  and _76400_ (_25695_, _25694_, _25688_);
  or _76401_ (_25696_, _25695_, _25399_);
  nand _76402_ (_25697_, _25696_, _12690_);
  nor _76403_ (_25698_, _12690_, _05921_);
  nor _76404_ (_25699_, _25698_, _10262_);
  nand _76405_ (_25700_, _25699_, _25697_);
  and _76406_ (_25702_, _10262_, _05907_);
  nor _76407_ (_25703_, _25702_, _06167_);
  and _76408_ (_25704_, _25703_, _25700_);
  and _76409_ (_25705_, _09070_, _06167_);
  or _76410_ (_25706_, _25705_, _25704_);
  nand _76411_ (_25707_, _25706_, _12703_);
  and _76412_ (_25708_, _06521_, _05826_);
  nor _76413_ (_25709_, _25708_, _06165_);
  nand _76414_ (_25710_, _25709_, _25707_);
  nor _76415_ (_25711_, _25412_, _12682_);
  and _76416_ (_25713_, _12029_, _12682_);
  nor _76417_ (_25714_, _25713_, _25711_);
  and _76418_ (_25715_, _25714_, _06165_);
  nor _76419_ (_25716_, _25715_, _12712_);
  nand _76420_ (_25717_, _25716_, _25710_);
  nor _76421_ (_25718_, _12711_, _05907_);
  nor _76422_ (_25719_, _25718_, _06433_);
  nand _76423_ (_25720_, _25719_, _25717_);
  not _76424_ (_25721_, _12719_);
  and _76425_ (_25722_, _06433_, _05921_);
  nor _76426_ (_25723_, _25722_, _25721_);
  and _76427_ (_25724_, _25723_, _25720_);
  nor _76428_ (_25725_, _12719_, _05907_);
  or _76429_ (_25726_, _25725_, _25724_);
  nand _76430_ (_25727_, _25726_, _07160_);
  and _76431_ (_25728_, _07577_, _06521_);
  nor _76432_ (_25729_, _25728_, _05748_);
  nand _76433_ (_25730_, _25729_, _25727_);
  and _76434_ (_25731_, _25714_, _05748_);
  nor _76435_ (_25732_, _25731_, _12737_);
  nand _76436_ (_25735_, _25732_, _25730_);
  nor _76437_ (_25736_, _12735_, _05907_);
  nor _76438_ (_25737_, _25736_, _06440_);
  and _76439_ (_25738_, _25737_, _25735_);
  or _76440_ (_25739_, _25738_, _25398_);
  nand _76441_ (_25740_, _25739_, _12744_);
  nor _76442_ (_25741_, _12744_, _25408_);
  nor _76443_ (_25742_, _25741_, _25019_);
  nand _76444_ (_25743_, _25742_, _25740_);
  and _76445_ (_25744_, _25019_, _06521_);
  nor _76446_ (_25746_, _25744_, _12754_);
  and _76447_ (_25747_, _25746_, _25743_);
  and _76448_ (_25748_, _12754_, _05907_);
  or _76449_ (_25749_, _25748_, _25747_);
  or _76450_ (_25750_, _25749_, _01321_);
  or _76451_ (_25751_, _01317_, \oc8051_golden_model_1.PC [2]);
  and _76452_ (_25752_, _25751_, _43100_);
  and _76453_ (_43690_, _25752_, _25750_);
  and _76454_ (_25753_, _06440_, _05974_);
  and _76455_ (_25754_, _06433_, _05974_);
  or _76456_ (_25756_, _11905_, _06324_);
  or _76457_ (_25757_, _11907_, _06324_);
  or _76458_ (_25758_, _11912_, _06324_);
  or _76459_ (_25759_, _11914_, _06324_);
  or _76460_ (_25760_, _11919_, _06324_);
  or _76461_ (_25761_, _08787_, _05974_);
  or _76462_ (_25762_, _25151_, _05974_);
  nand _76463_ (_25763_, _11924_, _05951_);
  nor _76464_ (_25764_, _06582_, _06389_);
  nand _76465_ (_25765_, _07056_, _06322_);
  and _76466_ (_25767_, _25765_, _12264_);
  and _76467_ (_25768_, _12265_, \oc8051_golden_model_1.PC [3]);
  or _76468_ (_25769_, _25768_, _07056_);
  and _76469_ (_25770_, _25769_, _25767_);
  or _76470_ (_25771_, _12266_, _05951_);
  nand _76471_ (_25772_, _25771_, _12263_);
  or _76472_ (_25773_, _25772_, _25770_);
  and _76473_ (_25774_, _25773_, _06582_);
  or _76474_ (_25775_, _25774_, _25764_);
  or _76475_ (_25776_, _12263_, _06324_);
  and _76476_ (_25778_, _25776_, _25775_);
  or _76477_ (_25779_, _25778_, _08445_);
  or _76478_ (_25780_, _12197_, _12196_);
  nand _76479_ (_25781_, _25780_, _12209_);
  or _76480_ (_25782_, _25780_, _12209_);
  and _76481_ (_25783_, _25782_, _25781_);
  and _76482_ (_25784_, _25783_, _12256_);
  and _76483_ (_25785_, _12258_, _05974_);
  or _76484_ (_25786_, _25785_, _08443_);
  or _76485_ (_25787_, _25786_, _25784_);
  and _76486_ (_25789_, _25787_, _25779_);
  or _76487_ (_25790_, _25789_, _07064_);
  nand _76488_ (_25791_, _07064_, _05951_);
  and _76489_ (_25792_, _25791_, _06161_);
  and _76490_ (_25793_, _25792_, _25790_);
  or _76491_ (_25794_, _12139_, _12023_);
  or _76492_ (_25795_, _12026_, _12025_);
  and _76493_ (_25796_, _25795_, _12041_);
  nor _76494_ (_25797_, _25795_, _12041_);
  nor _76495_ (_25798_, _25797_, _25796_);
  or _76496_ (_25800_, _25798_, _12141_);
  and _76497_ (_25801_, _25800_, _06160_);
  and _76498_ (_25802_, _25801_, _25794_);
  or _76499_ (_25803_, _25802_, _24821_);
  or _76500_ (_25804_, _25803_, _25793_);
  or _76501_ (_25805_, _12134_, _06324_);
  and _76502_ (_25806_, _25805_, _06157_);
  and _76503_ (_25807_, _25806_, _25804_);
  and _76504_ (_25808_, _06156_, _05974_);
  or _76505_ (_25809_, _25808_, _07485_);
  or _76506_ (_25811_, _25809_, _25807_);
  nand _76507_ (_25812_, _06389_, _07485_);
  and _76508_ (_25813_, _25812_, _07075_);
  and _76509_ (_25814_, _25813_, _25811_);
  nand _76510_ (_25815_, _06217_, _05974_);
  nand _76511_ (_25816_, _25815_, _12292_);
  or _76512_ (_25817_, _25816_, _25814_);
  or _76513_ (_25818_, _12292_, _06324_);
  and _76514_ (_25819_, _25818_, _06229_);
  and _76515_ (_25820_, _25819_, _25817_);
  nand _76516_ (_25822_, _06220_, _05974_);
  nand _76517_ (_25823_, _25822_, _12300_);
  or _76518_ (_25824_, _25823_, _25820_);
  or _76519_ (_25825_, _12300_, _06324_);
  and _76520_ (_25826_, _25825_, _06153_);
  and _76521_ (_25827_, _25826_, _25824_);
  and _76522_ (_25828_, _06152_, _05974_);
  or _76523_ (_25829_, _25828_, _12304_);
  or _76524_ (_25830_, _25829_, _25827_);
  nand _76525_ (_25831_, _06389_, _12304_);
  and _76526_ (_25833_, _25831_, _07191_);
  and _76527_ (_25834_, _25833_, _25830_);
  nand _76528_ (_25835_, _06151_, _05974_);
  nand _76529_ (_25836_, _25835_, _12125_);
  or _76530_ (_25837_, _25836_, _25834_);
  not _76531_ (_25838_, _25798_);
  nor _76532_ (_25839_, _25838_, _12120_);
  and _76533_ (_25840_, _12120_, _12023_);
  or _76534_ (_25841_, _25840_, _12125_);
  or _76535_ (_25842_, _25841_, _25839_);
  and _76536_ (_25844_, _25842_, _25114_);
  and _76537_ (_25845_, _25844_, _25837_);
  and _76538_ (_25846_, _12329_, _12023_);
  nor _76539_ (_25847_, _25838_, _12329_);
  or _76540_ (_25848_, _25847_, _25846_);
  and _76541_ (_25849_, _25848_, _06236_);
  or _76542_ (_25850_, _12023_, _11956_);
  or _76543_ (_25851_, _25798_, _11958_);
  and _76544_ (_25852_, _25851_, _06687_);
  and _76545_ (_25853_, _25852_, _25850_);
  or _76546_ (_25855_, _25853_, _25849_);
  or _76547_ (_25856_, _25855_, _25845_);
  and _76548_ (_25857_, _25856_, _12317_);
  nand _76549_ (_25858_, _12346_, _12024_);
  or _76550_ (_25859_, _25798_, _12346_);
  and _76551_ (_25860_, _25859_, _06295_);
  and _76552_ (_25861_, _25860_, _25858_);
  or _76553_ (_25862_, _25861_, _11924_);
  or _76554_ (_25863_, _25862_, _25857_);
  and _76555_ (_25864_, _25863_, _25763_);
  or _76556_ (_25866_, _25864_, _06145_);
  nand _76557_ (_25867_, _06145_, _06322_);
  and _76558_ (_25868_, _25867_, _05760_);
  and _76559_ (_25869_, _25868_, _25866_);
  nor _76560_ (_25870_, _06389_, _05760_);
  or _76561_ (_25871_, _25870_, _25152_);
  or _76562_ (_25872_, _25871_, _25869_);
  and _76563_ (_25873_, _25872_, _25762_);
  or _76564_ (_25874_, _25873_, _12373_);
  or _76565_ (_25875_, _12369_, _06324_);
  and _76566_ (_25876_, _25875_, _13844_);
  and _76567_ (_25877_, _25876_, _25874_);
  and _76568_ (_25878_, _06255_, _05974_);
  or _76569_ (_25879_, _25878_, _24882_);
  or _76570_ (_25880_, _25879_, _25877_);
  nand _76571_ (_25881_, _06389_, _24882_);
  and _76572_ (_25882_, _25881_, _13843_);
  and _76573_ (_25883_, _25882_, _25880_);
  nand _76574_ (_25884_, _06254_, _05974_);
  nand _76575_ (_25885_, _25884_, _12381_);
  or _76576_ (_25887_, _25885_, _25883_);
  or _76577_ (_25888_, _12381_, _06324_);
  and _76578_ (_25889_, _25888_, _25887_);
  or _76579_ (_25890_, _25889_, _12386_);
  or _76580_ (_25891_, _12385_, _05974_);
  and _76581_ (_25892_, _25891_, _05805_);
  and _76582_ (_25893_, _25892_, _25890_);
  nor _76583_ (_25894_, _05805_, _05951_);
  or _76584_ (_25895_, _25894_, _06139_);
  or _76585_ (_25896_, _25895_, _25893_);
  nand _76586_ (_25898_, _06139_, _06322_);
  and _76587_ (_25899_, _25898_, _25896_);
  or _76588_ (_25900_, _25899_, _05791_);
  nand _76589_ (_25901_, _06389_, _05791_);
  and _76590_ (_25902_, _25901_, _11296_);
  and _76591_ (_25903_, _25902_, _25900_);
  nand _76592_ (_25904_, _12023_, _06293_);
  nand _76593_ (_25905_, _25904_, _06133_);
  or _76594_ (_25906_, _25905_, _25903_);
  or _76595_ (_25907_, _06133_, _05974_);
  and _76596_ (_25908_, _25907_, _06114_);
  and _76597_ (_25909_, _25908_, _25906_);
  nand _76598_ (_25910_, _12023_, _05787_);
  nand _76599_ (_25911_, _25910_, _11922_);
  or _76600_ (_25912_, _25911_, _25909_);
  or _76601_ (_25913_, _11922_, _06324_);
  and _76602_ (_25914_, _25913_, _06762_);
  and _76603_ (_25915_, _25914_, _25912_);
  and _76604_ (_25916_, _06209_, _05974_);
  or _76605_ (_25917_, _25916_, _05829_);
  or _76606_ (_25918_, _25917_, _25915_);
  nand _76607_ (_25919_, _06389_, _05829_);
  and _76608_ (_25920_, _25919_, _12417_);
  and _76609_ (_25921_, _25920_, _25918_);
  and _76610_ (_25922_, _25783_, _12416_);
  or _76611_ (_25923_, _25922_, _08788_);
  or _76612_ (_25924_, _25923_, _25921_);
  and _76613_ (_25925_, _25924_, _25761_);
  or _76614_ (_25926_, _25925_, _06110_);
  nand _76615_ (_25927_, _12024_, _06110_);
  and _76616_ (_25928_, _25927_, _10752_);
  and _76617_ (_25929_, _25928_, _25926_);
  and _76618_ (_25930_, _10751_, _05974_);
  or _76619_ (_25931_, _25930_, _12431_);
  or _76620_ (_25932_, _25931_, _25929_);
  or _76621_ (_25933_, _12432_, _05968_);
  and _76622_ (_25934_, _25933_, _06768_);
  and _76623_ (_25935_, _25934_, _25932_);
  and _76624_ (_25936_, _06208_, _05974_);
  or _76625_ (_25937_, _25936_, _06076_);
  or _76626_ (_25938_, _25937_, _25935_);
  nand _76627_ (_25939_, _06389_, _06076_);
  and _76628_ (_25940_, _25939_, _12474_);
  and _76629_ (_25941_, _25940_, _25938_);
  or _76630_ (_25942_, _25783_, _11101_);
  nand _76631_ (_25943_, _11101_, _06322_);
  and _76632_ (_25944_, _25943_, _12473_);
  and _76633_ (_25945_, _25944_, _25942_);
  or _76634_ (_25946_, _25945_, _12478_);
  or _76635_ (_25947_, _25946_, _25941_);
  and _76636_ (_25948_, _25947_, _25760_);
  or _76637_ (_25949_, _25948_, _11917_);
  or _76638_ (_25950_, _11916_, _05974_);
  and _76639_ (_25951_, _25950_, _07127_);
  and _76640_ (_25952_, _25951_, _25949_);
  and _76641_ (_25953_, _12023_, _06297_);
  or _76642_ (_25954_, _25953_, _06402_);
  or _76643_ (_25955_, _25954_, _25952_);
  nand _76644_ (_25956_, _06402_, _06322_);
  and _76645_ (_25957_, _25956_, _25955_);
  or _76646_ (_25959_, _25957_, _12492_);
  nand _76647_ (_25960_, _06389_, _12492_);
  and _76648_ (_25961_, _25960_, _12497_);
  and _76649_ (_25962_, _25961_, _25959_);
  or _76650_ (_25963_, _25783_, _12480_);
  or _76651_ (_25964_, _11101_, _05974_);
  and _76652_ (_25965_, _25964_, _12496_);
  and _76653_ (_25966_, _25965_, _25963_);
  or _76654_ (_25967_, _25966_, _12505_);
  or _76655_ (_25968_, _25967_, _25962_);
  and _76656_ (_25970_, _25968_, _25759_);
  or _76657_ (_25971_, _25970_, _10822_);
  or _76658_ (_25972_, _10821_, _05974_);
  and _76659_ (_25973_, _25972_, _07132_);
  and _76660_ (_25974_, _25973_, _25971_);
  and _76661_ (_25975_, _12023_, _06306_);
  or _76662_ (_25976_, _25975_, _06411_);
  or _76663_ (_25977_, _25976_, _25974_);
  nand _76664_ (_25978_, _06411_, _06322_);
  and _76665_ (_25979_, _25978_, _25977_);
  or _76666_ (_25980_, _25979_, _07124_);
  nand _76667_ (_25981_, _06389_, _07124_);
  and _76668_ (_25982_, _25981_, _12518_);
  and _76669_ (_25983_, _25982_, _25980_);
  or _76670_ (_25984_, _25783_, \oc8051_golden_model_1.PSW [7]);
  or _76671_ (_25985_, _05974_, _10693_);
  and _76672_ (_25986_, _25985_, _12517_);
  and _76673_ (_25987_, _25986_, _25984_);
  or _76674_ (_25988_, _25987_, _12522_);
  or _76675_ (_25989_, _25988_, _25983_);
  and _76676_ (_25991_, _25989_, _25758_);
  or _76677_ (_25992_, _25991_, _10850_);
  or _76678_ (_25993_, _10849_, _05974_);
  and _76679_ (_25994_, _25993_, _08819_);
  and _76680_ (_25995_, _25994_, _25992_);
  and _76681_ (_25996_, _12023_, _06303_);
  or _76682_ (_25997_, _25996_, _06396_);
  or _76683_ (_25998_, _25997_, _25995_);
  nand _76684_ (_25999_, _06396_, _06322_);
  and _76685_ (_26000_, _25999_, _25998_);
  or _76686_ (_26002_, _26000_, _05842_);
  nand _76687_ (_26003_, _06389_, _05842_);
  and _76688_ (_26004_, _26003_, _12539_);
  and _76689_ (_26005_, _26004_, _26002_);
  or _76690_ (_26006_, _25783_, _10693_);
  or _76691_ (_26007_, _05974_, \oc8051_golden_model_1.PSW [7]);
  and _76692_ (_26008_, _26007_, _12538_);
  and _76693_ (_26009_, _26008_, _26006_);
  or _76694_ (_26010_, _26009_, _12547_);
  or _76695_ (_26011_, _26010_, _26005_);
  and _76696_ (_26013_, _26011_, _25757_);
  or _76697_ (_26014_, _26013_, _10897_);
  or _76698_ (_26015_, _10896_, _05974_);
  and _76699_ (_26016_, _26015_, _10926_);
  and _76700_ (_26017_, _26016_, _26014_);
  and _76701_ (_26018_, _10925_, _06324_);
  or _76702_ (_26019_, _26018_, _06417_);
  or _76703_ (_26020_, _26019_, _26017_);
  or _76704_ (_26021_, _09210_, _12558_);
  and _76705_ (_26022_, _26021_, _26020_);
  or _76706_ (_26024_, _26022_, _07142_);
  nand _76707_ (_26025_, _06389_, _07142_);
  and _76708_ (_26026_, _26025_, _06421_);
  and _76709_ (_26027_, _26026_, _26024_);
  or _76710_ (_26028_, _12023_, _12682_);
  nand _76711_ (_26029_, _25838_, _12682_);
  and _76712_ (_26030_, _26029_, _06301_);
  and _76713_ (_26031_, _26030_, _26028_);
  or _76714_ (_26032_, _26031_, _12565_);
  or _76715_ (_26033_, _26032_, _26027_);
  and _76716_ (_26034_, _26033_, _25756_);
  or _76717_ (_26035_, _26034_, _12691_);
  or _76718_ (_26036_, _12690_, _05974_);
  and _76719_ (_26037_, _26036_, _12693_);
  and _76720_ (_26038_, _26037_, _26035_);
  and _76721_ (_26039_, _10262_, _06324_);
  or _76722_ (_26040_, _26039_, _06167_);
  or _76723_ (_26041_, _26040_, _26038_);
  or _76724_ (_26042_, _09210_, _06168_);
  and _76725_ (_26043_, _26042_, _26041_);
  or _76726_ (_26044_, _26043_, _05826_);
  nand _76727_ (_26045_, _06389_, _05826_);
  and _76728_ (_26046_, _26045_, _06166_);
  and _76729_ (_26047_, _26046_, _26044_);
  nor _76730_ (_26048_, _25798_, _12682_);
  and _76731_ (_26049_, _12024_, _12682_);
  nor _76732_ (_26050_, _26049_, _26048_);
  and _76733_ (_26051_, _26050_, _06165_);
  or _76734_ (_26052_, _26051_, _12712_);
  or _76735_ (_26053_, _26052_, _26047_);
  or _76736_ (_26056_, _12711_, _06324_);
  and _76737_ (_26057_, _26056_, _06829_);
  and _76738_ (_26058_, _26057_, _26053_);
  or _76739_ (_26059_, _26058_, _25754_);
  nand _76740_ (_26060_, _26059_, _12719_);
  nor _76741_ (_26061_, _12719_, _05951_);
  nor _76742_ (_26062_, _26061_, _07577_);
  nand _76743_ (_26063_, _26062_, _26060_);
  and _76744_ (_26064_, _07577_, _06389_);
  nor _76745_ (_26065_, _26064_, _05748_);
  nand _76746_ (_26067_, _26065_, _26063_);
  and _76747_ (_26068_, _26050_, _05748_);
  nor _76748_ (_26069_, _26068_, _12737_);
  nand _76749_ (_26070_, _26069_, _26067_);
  nor _76750_ (_26071_, _12735_, _06324_);
  nor _76751_ (_26072_, _26071_, _06440_);
  and _76752_ (_26073_, _26072_, _26070_);
  or _76753_ (_26074_, _26073_, _25753_);
  nand _76754_ (_26075_, _26074_, _12744_);
  nor _76755_ (_26076_, _12744_, _05951_);
  nor _76756_ (_26078_, _26076_, _25019_);
  nand _76757_ (_26079_, _26078_, _26075_);
  and _76758_ (_26080_, _25019_, _06389_);
  nor _76759_ (_26081_, _26080_, _12754_);
  and _76760_ (_26082_, _26081_, _26079_);
  and _76761_ (_26083_, _12754_, _06324_);
  or _76762_ (_26084_, _26083_, _26082_);
  or _76763_ (_26085_, _26084_, _01321_);
  or _76764_ (_26086_, _01317_, \oc8051_golden_model_1.PC [3]);
  and _76765_ (_26087_, _26086_, _43100_);
  and _76766_ (_43691_, _26087_, _26085_);
  and _76767_ (_26089_, _08670_, _07577_);
  nor _76768_ (_26090_, _12194_, _11101_);
  and _76769_ (_26091_, _12214_, _12211_);
  nor _76770_ (_26092_, _26091_, _12215_);
  and _76771_ (_26093_, _26092_, _11101_);
  or _76772_ (_26094_, _26093_, _26090_);
  and _76773_ (_26095_, _26094_, _12496_);
  and _76774_ (_26096_, _12193_, _11101_);
  and _76775_ (_26097_, _26092_, _12480_);
  or _76776_ (_26098_, _26097_, _26096_);
  and _76777_ (_26099_, _26098_, _12473_);
  nor _76778_ (_26100_, _12193_, _08787_);
  nor _76779_ (_26101_, _25151_, _12193_);
  and _76780_ (_26102_, _05426_, \oc8051_golden_model_1.PC [4]);
  nor _76781_ (_26103_, _05426_, \oc8051_golden_model_1.PC [4]);
  nor _76782_ (_26104_, _26103_, _26102_);
  not _76783_ (_26105_, _26104_);
  and _76784_ (_26106_, _26105_, _11924_);
  nand _76785_ (_26107_, _26105_, _12287_);
  and _76786_ (_26109_, _12046_, _12043_);
  nor _76787_ (_26110_, _26109_, _12047_);
  or _76788_ (_26111_, _26110_, _12141_);
  or _76789_ (_26112_, _12139_, _12018_);
  and _76790_ (_26113_, _26112_, _26111_);
  or _76791_ (_26114_, _26113_, _06161_);
  and _76792_ (_26115_, _08670_, _06581_);
  and _76793_ (_26116_, _12194_, _07056_);
  or _76794_ (_26117_, _26116_, _06653_);
  nand _76795_ (_26118_, _12265_, \oc8051_golden_model_1.PC [4]);
  and _76796_ (_26120_, _26118_, _07057_);
  or _76797_ (_26121_, _26120_, _26117_);
  or _76798_ (_26122_, _26105_, _12266_);
  and _76799_ (_26123_, _26122_, _06582_);
  and _76800_ (_26124_, _26123_, _26121_);
  or _76801_ (_26125_, _26124_, _25055_);
  or _76802_ (_26126_, _26125_, _26115_);
  or _76803_ (_26127_, _26105_, _12263_);
  and _76804_ (_26128_, _26127_, _08443_);
  and _76805_ (_26129_, _26128_, _26126_);
  or _76806_ (_26131_, _12256_, _12194_);
  nand _76807_ (_26132_, _26092_, _12256_);
  and _76808_ (_26133_, _26132_, _08445_);
  and _76809_ (_26134_, _26133_, _26131_);
  or _76810_ (_26135_, _26134_, _26129_);
  nand _76811_ (_26136_, _26135_, _12281_);
  and _76812_ (_26137_, _26136_, _26114_);
  or _76813_ (_26138_, _26137_, _24821_);
  nand _76814_ (_26139_, _26138_, _26107_);
  nand _76815_ (_26140_, _26139_, _06157_);
  and _76816_ (_26142_, _12194_, _06156_);
  nor _76817_ (_26143_, _26142_, _07485_);
  nand _76818_ (_26144_, _26143_, _26140_);
  nor _76819_ (_26145_, _08670_, _05764_);
  nor _76820_ (_26146_, _26145_, _06217_);
  and _76821_ (_26147_, _26146_, _26144_);
  and _76822_ (_26148_, _12194_, _06217_);
  or _76823_ (_26149_, _26148_, _26147_);
  and _76824_ (_26150_, _26149_, _12292_);
  nor _76825_ (_26151_, _26104_, _12292_);
  or _76826_ (_26153_, _26151_, _26150_);
  nand _76827_ (_26154_, _26153_, _06229_);
  and _76828_ (_26155_, _12194_, _06220_);
  nor _76829_ (_26156_, _26155_, _12302_);
  nand _76830_ (_26157_, _26156_, _26154_);
  nor _76831_ (_26158_, _26105_, _12300_);
  nor _76832_ (_26159_, _26158_, _06152_);
  and _76833_ (_26160_, _26159_, _26157_);
  and _76834_ (_26161_, _12194_, _06152_);
  or _76835_ (_26162_, _26161_, _26160_);
  nand _76836_ (_26163_, _26162_, _05769_);
  and _76837_ (_26164_, _08670_, _12304_);
  nor _76838_ (_26165_, _26164_, _06151_);
  nand _76839_ (_26166_, _26165_, _26163_);
  and _76840_ (_26167_, _12193_, _06151_);
  nor _76841_ (_26168_, _26167_, _12126_);
  nand _76842_ (_26169_, _26168_, _26166_);
  and _76843_ (_26170_, _12120_, _12018_);
  not _76844_ (_26171_, _26110_);
  nor _76845_ (_26172_, _26171_, _12120_);
  or _76846_ (_26174_, _26172_, _12125_);
  nor _76847_ (_26175_, _26174_, _26170_);
  not _76848_ (_26176_, _26175_);
  and _76849_ (_26177_, _26176_, _26169_);
  or _76850_ (_26178_, _26177_, _06687_);
  and _76851_ (_26179_, _26110_, _11956_);
  and _76852_ (_26180_, _12018_, _11958_);
  or _76853_ (_26181_, _26180_, _12089_);
  or _76854_ (_26182_, _26181_, _26179_);
  nand _76855_ (_26183_, _26182_, _26178_);
  nand _76856_ (_26185_, _26183_, _06643_);
  nor _76857_ (_26186_, _26171_, _12329_);
  not _76858_ (_26187_, _26186_);
  and _76859_ (_26188_, _12329_, _12018_);
  nor _76860_ (_26189_, _26188_, _06643_);
  and _76861_ (_26190_, _26189_, _26187_);
  nor _76862_ (_26191_, _26190_, _06295_);
  nand _76863_ (_26192_, _26191_, _26185_);
  nor _76864_ (_26193_, _26110_, _12346_);
  and _76865_ (_26194_, _12346_, _12019_);
  nor _76866_ (_26196_, _26194_, _12317_);
  not _76867_ (_26197_, _26196_);
  nor _76868_ (_26198_, _26197_, _26193_);
  nor _76869_ (_26199_, _26198_, _11924_);
  and _76870_ (_26200_, _26199_, _26192_);
  or _76871_ (_26201_, _26200_, _26106_);
  nand _76872_ (_26202_, _26201_, _06146_);
  and _76873_ (_26203_, _12194_, _06145_);
  nor _76874_ (_26204_, _26203_, _07388_);
  nand _76875_ (_26205_, _26204_, _26202_);
  nor _76876_ (_26207_, _08670_, _05760_);
  nor _76877_ (_26208_, _26207_, _25152_);
  and _76878_ (_26209_, _26208_, _26205_);
  or _76879_ (_26210_, _26209_, _26101_);
  nand _76880_ (_26211_, _26210_, _12369_);
  nor _76881_ (_26212_, _26104_, _12369_);
  nor _76882_ (_26213_, _26212_, _06255_);
  nand _76883_ (_26214_, _26213_, _26211_);
  and _76884_ (_26215_, _12193_, _06255_);
  nor _76885_ (_26216_, _26215_, _24882_);
  nand _76886_ (_26218_, _26216_, _26214_);
  and _76887_ (_26219_, _08670_, _24882_);
  nor _76888_ (_26220_, _26219_, _06254_);
  and _76889_ (_26221_, _26220_, _26218_);
  and _76890_ (_26222_, _12193_, _06254_);
  or _76891_ (_26223_, _26222_, _26221_);
  nand _76892_ (_26224_, _26223_, _12381_);
  nor _76893_ (_26225_, _26105_, _12381_);
  nor _76894_ (_26226_, _26225_, _12386_);
  nand _76895_ (_26227_, _26226_, _26224_);
  nor _76896_ (_26228_, _12193_, _12385_);
  nor _76897_ (_26229_, _26228_, _05870_);
  nand _76898_ (_26230_, _26229_, _26227_);
  nor _76899_ (_26231_, _26105_, _05805_);
  nor _76900_ (_26232_, _26231_, _06139_);
  and _76901_ (_26233_, _26232_, _26230_);
  and _76902_ (_26234_, _12194_, _06139_);
  or _76903_ (_26235_, _26234_, _26233_);
  nand _76904_ (_26236_, _26235_, _24791_);
  and _76905_ (_26237_, _08670_, _05791_);
  nor _76906_ (_26239_, _26237_, _06293_);
  nand _76907_ (_26240_, _26239_, _26236_);
  and _76908_ (_26241_, _12018_, _06293_);
  nor _76909_ (_26242_, _26241_, _13620_);
  nand _76910_ (_26243_, _26242_, _26240_);
  nor _76911_ (_26244_, _12193_, _06133_);
  nor _76912_ (_26245_, _26244_, _05787_);
  nand _76913_ (_26246_, _26245_, _26243_);
  and _76914_ (_26247_, _12018_, _05787_);
  nor _76915_ (_26248_, _26247_, _12412_);
  nand _76916_ (_26250_, _26248_, _26246_);
  nor _76917_ (_26251_, _26104_, _11922_);
  nor _76918_ (_26252_, _26251_, _06209_);
  nand _76919_ (_26253_, _26252_, _26250_);
  and _76920_ (_26254_, _12193_, _06209_);
  nor _76921_ (_26255_, _26254_, _05829_);
  nand _76922_ (_26256_, _26255_, _26253_);
  and _76923_ (_26257_, _08670_, _05829_);
  nor _76924_ (_26258_, _26257_, _12416_);
  nand _76925_ (_26259_, _26258_, _26256_);
  and _76926_ (_26261_, _26092_, _12416_);
  nor _76927_ (_26262_, _26261_, _08788_);
  and _76928_ (_26263_, _26262_, _26259_);
  or _76929_ (_26264_, _26263_, _26100_);
  nand _76930_ (_26265_, _26264_, _06111_);
  and _76931_ (_26266_, _12019_, _06110_);
  nor _76932_ (_26267_, _26266_, _10751_);
  nand _76933_ (_26268_, _26267_, _26265_);
  and _76934_ (_26269_, _12193_, _10751_);
  nor _76935_ (_26270_, _26269_, _12431_);
  nand _76936_ (_26272_, _26270_, _26268_);
  and _76937_ (_26273_, _12449_, _12446_);
  nor _76938_ (_26274_, _26273_, _12450_);
  nor _76939_ (_26275_, _26274_, _12432_);
  nor _76940_ (_26276_, _26275_, _06208_);
  nand _76941_ (_26277_, _26276_, _26272_);
  and _76942_ (_26278_, _12193_, _06208_);
  nor _76943_ (_26279_, _26278_, _06076_);
  nand _76944_ (_26280_, _26279_, _26277_);
  and _76945_ (_26281_, _08670_, _06076_);
  nor _76946_ (_26283_, _26281_, _12473_);
  and _76947_ (_26284_, _26283_, _26280_);
  or _76948_ (_26285_, _26284_, _26099_);
  nand _76949_ (_26286_, _26285_, _11919_);
  nor _76950_ (_26287_, _26105_, _11919_);
  nor _76951_ (_26288_, _26287_, _11917_);
  nand _76952_ (_26289_, _26288_, _26286_);
  nor _76953_ (_26290_, _12193_, _11916_);
  nor _76954_ (_26291_, _26290_, _06297_);
  nand _76955_ (_26292_, _26291_, _26289_);
  and _76956_ (_26293_, _12018_, _06297_);
  nor _76957_ (_26294_, _26293_, _06402_);
  and _76958_ (_26295_, _26294_, _26292_);
  and _76959_ (_26296_, _12194_, _06402_);
  or _76960_ (_26297_, _26296_, _26295_);
  nand _76961_ (_26298_, _26297_, _05834_);
  and _76962_ (_26299_, _08670_, _12492_);
  nor _76963_ (_26300_, _26299_, _12496_);
  and _76964_ (_26301_, _26300_, _26298_);
  or _76965_ (_26302_, _26301_, _26095_);
  nand _76966_ (_26304_, _26302_, _11914_);
  nor _76967_ (_26305_, _26105_, _11914_);
  nor _76968_ (_26306_, _26305_, _10822_);
  nand _76969_ (_26307_, _26306_, _26304_);
  nor _76970_ (_26308_, _12193_, _10821_);
  nor _76971_ (_26309_, _26308_, _06306_);
  nand _76972_ (_26310_, _26309_, _26307_);
  and _76973_ (_26311_, _12018_, _06306_);
  nor _76974_ (_26312_, _26311_, _06411_);
  and _76975_ (_26313_, _26312_, _26310_);
  and _76976_ (_26315_, _12194_, _06411_);
  or _76977_ (_26316_, _26315_, _26313_);
  nand _76978_ (_26317_, _26316_, _05848_);
  and _76979_ (_26318_, _08670_, _07124_);
  nor _76980_ (_26319_, _26318_, _12517_);
  and _76981_ (_26320_, _26319_, _26317_);
  and _76982_ (_26321_, _12193_, \oc8051_golden_model_1.PSW [7]);
  and _76983_ (_26322_, _26092_, _10693_);
  or _76984_ (_26323_, _26322_, _26321_);
  and _76985_ (_26324_, _26323_, _12517_);
  or _76986_ (_26326_, _26324_, _26320_);
  nand _76987_ (_26327_, _26326_, _11912_);
  nor _76988_ (_26328_, _26105_, _11912_);
  nor _76989_ (_26329_, _26328_, _10850_);
  nand _76990_ (_26330_, _26329_, _26327_);
  nor _76991_ (_26331_, _12193_, _10849_);
  nor _76992_ (_26332_, _26331_, _06303_);
  nand _76993_ (_26333_, _26332_, _26330_);
  and _76994_ (_26334_, _12018_, _06303_);
  nor _76995_ (_26335_, _26334_, _06396_);
  and _76996_ (_26337_, _26335_, _26333_);
  and _76997_ (_26338_, _12194_, _06396_);
  or _76998_ (_26339_, _26338_, _26337_);
  nand _76999_ (_26340_, _26339_, _05843_);
  and _77000_ (_26341_, _08670_, _05842_);
  nor _77001_ (_26342_, _26341_, _12538_);
  and _77002_ (_26343_, _26342_, _26340_);
  and _77003_ (_26344_, _12193_, _10693_);
  and _77004_ (_26345_, _26092_, \oc8051_golden_model_1.PSW [7]);
  or _77005_ (_26346_, _26345_, _26344_);
  and _77006_ (_26348_, _26346_, _12538_);
  or _77007_ (_26349_, _26348_, _26343_);
  nand _77008_ (_26350_, _26349_, _11907_);
  nor _77009_ (_26351_, _26105_, _11907_);
  nor _77010_ (_26352_, _26351_, _10897_);
  nand _77011_ (_26353_, _26352_, _26350_);
  nor _77012_ (_26354_, _12193_, _10896_);
  nor _77013_ (_26355_, _26354_, _10925_);
  nand _77014_ (_26356_, _26355_, _26353_);
  and _77015_ (_26357_, _26104_, _10925_);
  nor _77016_ (_26359_, _26357_, _06417_);
  and _77017_ (_26360_, _26359_, _26356_);
  and _77018_ (_26361_, _08980_, _06417_);
  or _77019_ (_26362_, _26361_, _26360_);
  nand _77020_ (_26363_, _26362_, _05846_);
  and _77021_ (_26364_, _08670_, _07142_);
  nor _77022_ (_26365_, _26364_, _06301_);
  and _77023_ (_26366_, _26365_, _26363_);
  nor _77024_ (_26367_, _12019_, _12682_);
  and _77025_ (_26368_, _26110_, _12682_);
  nor _77026_ (_26370_, _26368_, _26367_);
  nor _77027_ (_26371_, _26370_, _06421_);
  or _77028_ (_26372_, _26371_, _26366_);
  nand _77029_ (_26373_, _26372_, _11905_);
  nor _77030_ (_26374_, _26105_, _11905_);
  nor _77031_ (_26375_, _26374_, _12691_);
  nand _77032_ (_26376_, _26375_, _26373_);
  nor _77033_ (_26377_, _12690_, _12193_);
  nor _77034_ (_26378_, _26377_, _10262_);
  nand _77035_ (_26379_, _26378_, _26376_);
  and _77036_ (_26380_, _26104_, _10262_);
  nor _77037_ (_26381_, _26380_, _06167_);
  nand _77038_ (_26382_, _26381_, _26379_);
  and _77039_ (_26383_, _08980_, _06167_);
  nor _77040_ (_26384_, _26383_, _05826_);
  nand _77041_ (_26385_, _26384_, _26382_);
  nor _77042_ (_26386_, _08670_, _12703_);
  nor _77043_ (_26387_, _26386_, _06165_);
  nand _77044_ (_26388_, _26387_, _26385_);
  and _77045_ (_26389_, _12019_, _12682_);
  nor _77046_ (_26391_, _26110_, _12682_);
  nor _77047_ (_26392_, _26391_, _26389_);
  nor _77048_ (_26393_, _26392_, _06166_);
  nor _77049_ (_26394_, _26393_, _12712_);
  nand _77050_ (_26395_, _26394_, _26388_);
  nor _77051_ (_26396_, _26105_, _12711_);
  nor _77052_ (_26397_, _26396_, _06433_);
  nand _77053_ (_26398_, _26397_, _26395_);
  and _77054_ (_26399_, _12194_, _06433_);
  nor _77055_ (_26400_, _26399_, _25721_);
  nand _77056_ (_26402_, _26400_, _26398_);
  nor _77057_ (_26403_, _26105_, _12719_);
  nor _77058_ (_26404_, _26403_, _07577_);
  and _77059_ (_26405_, _26404_, _26402_);
  or _77060_ (_26406_, _26405_, _26089_);
  nand _77061_ (_26407_, _26406_, _05749_);
  nor _77062_ (_26408_, _26392_, _05749_);
  nor _77063_ (_26409_, _26408_, _12737_);
  nand _77064_ (_26410_, _26409_, _26407_);
  nor _77065_ (_26411_, _26105_, _12735_);
  nor _77066_ (_26413_, _26411_, _06440_);
  nand _77067_ (_26414_, _26413_, _26410_);
  not _77068_ (_26415_, _12744_);
  and _77069_ (_26416_, _12194_, _06440_);
  nor _77070_ (_26417_, _26416_, _26415_);
  nand _77071_ (_26418_, _26417_, _26414_);
  nor _77072_ (_26419_, _26105_, _12744_);
  nor _77073_ (_26420_, _26419_, _25019_);
  nand _77074_ (_26421_, _26420_, _26418_);
  and _77075_ (_26422_, _25019_, _08670_);
  nor _77076_ (_26424_, _26422_, _12754_);
  and _77077_ (_26425_, _26424_, _26421_);
  and _77078_ (_26426_, _26104_, _12754_);
  or _77079_ (_26427_, _26426_, _26425_);
  or _77080_ (_26428_, _26427_, _01321_);
  or _77081_ (_26429_, _01317_, \oc8051_golden_model_1.PC [4]);
  and _77082_ (_26430_, _26429_, _43100_);
  and _77083_ (_43692_, _26430_, _26428_);
  and _77084_ (_26431_, _12188_, _06440_);
  and _77085_ (_26432_, _12188_, _06433_);
  nor _77086_ (_26434_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor _77087_ (_26435_, _12188_, _05444_);
  nor _77088_ (_26436_, _26435_, _26434_);
  nor _77089_ (_26437_, _26436_, _11905_);
  and _77090_ (_26438_, _08931_, _06417_);
  nor _77091_ (_26439_, _26436_, _11907_);
  nor _77092_ (_26440_, _26436_, _11912_);
  nor _77093_ (_26441_, _26436_, _11914_);
  nor _77094_ (_26442_, _26436_, _11919_);
  nor _77095_ (_26443_, _12188_, _08787_);
  nor _77096_ (_26444_, _25151_, _12188_);
  not _77097_ (_26445_, _26436_);
  and _77098_ (_26446_, _26445_, _11924_);
  nor _77099_ (_26447_, _08701_, _06582_);
  and _77100_ (_26448_, _12189_, _07056_);
  nor _77101_ (_26449_, _26448_, _06653_);
  and _77102_ (_26450_, _12265_, \oc8051_golden_model_1.PC [5]);
  or _77103_ (_26451_, _26450_, _07056_);
  and _77104_ (_26452_, _26451_, _26449_);
  or _77105_ (_26453_, _26445_, _12266_);
  nand _77106_ (_26455_, _26453_, _12263_);
  or _77107_ (_26456_, _26455_, _26452_);
  and _77108_ (_26457_, _26456_, _06582_);
  nor _77109_ (_26458_, _26457_, _26447_);
  nor _77110_ (_26459_, _26436_, _12263_);
  nor _77111_ (_26460_, _26459_, _26458_);
  nor _77112_ (_26461_, _26460_, _08445_);
  or _77113_ (_26462_, _12256_, _12189_);
  or _77114_ (_26463_, _12191_, _12190_);
  and _77115_ (_26464_, _26463_, _12216_);
  nor _77116_ (_26466_, _26463_, _12216_);
  or _77117_ (_26467_, _26466_, _26464_);
  or _77118_ (_26468_, _26467_, _12258_);
  and _77119_ (_26469_, _26468_, _08445_);
  and _77120_ (_26470_, _26469_, _26462_);
  or _77121_ (_26471_, _26470_, _26461_);
  nand _77122_ (_26472_, _26471_, _07065_);
  and _77123_ (_26473_, _26445_, _07064_);
  nor _77124_ (_26474_, _26473_, _06160_);
  and _77125_ (_26475_, _26474_, _26472_);
  or _77126_ (_26477_, _12139_, _12014_);
  or _77127_ (_26478_, _12016_, _12015_);
  not _77128_ (_26479_, _26478_);
  nor _77129_ (_26480_, _26479_, _12048_);
  and _77130_ (_26481_, _26479_, _12048_);
  nor _77131_ (_26482_, _26481_, _26480_);
  or _77132_ (_26483_, _26482_, _12141_);
  nand _77133_ (_26484_, _26483_, _26477_);
  and _77134_ (_26485_, _26484_, _06160_);
  or _77135_ (_26486_, _26485_, _24821_);
  or _77136_ (_26488_, _26486_, _26475_);
  nor _77137_ (_26489_, _26436_, _12134_);
  nor _77138_ (_26490_, _26489_, _06156_);
  nand _77139_ (_26491_, _26490_, _26488_);
  and _77140_ (_26492_, _12188_, _06156_);
  nor _77141_ (_26493_, _26492_, _07485_);
  nand _77142_ (_26494_, _26493_, _26491_);
  and _77143_ (_26495_, _08701_, _07485_);
  nor _77144_ (_26496_, _26495_, _06217_);
  nand _77145_ (_26497_, _26496_, _26494_);
  and _77146_ (_26499_, _12188_, _06217_);
  nor _77147_ (_26500_, _26499_, _12293_);
  nand _77148_ (_26501_, _26500_, _26497_);
  nor _77149_ (_26502_, _26436_, _12292_);
  nor _77150_ (_26503_, _26502_, _06220_);
  nand _77151_ (_26504_, _26503_, _26501_);
  and _77152_ (_26505_, _12188_, _06220_);
  nor _77153_ (_26506_, _26505_, _12302_);
  nand _77154_ (_26507_, _26506_, _26504_);
  nor _77155_ (_26508_, _26436_, _12300_);
  nor _77156_ (_26510_, _26508_, _06152_);
  nand _77157_ (_26511_, _26510_, _26507_);
  and _77158_ (_26512_, _12188_, _06152_);
  nor _77159_ (_26513_, _26512_, _12304_);
  nand _77160_ (_26514_, _26513_, _26511_);
  and _77161_ (_26515_, _08701_, _12304_);
  nor _77162_ (_26516_, _26515_, _06151_);
  nand _77163_ (_26517_, _26516_, _26514_);
  and _77164_ (_26518_, _12188_, _06151_);
  nor _77165_ (_26519_, _26518_, _12126_);
  nand _77166_ (_26520_, _26519_, _26517_);
  and _77167_ (_26521_, _12120_, _12013_);
  nor _77168_ (_26522_, _26482_, _12120_);
  or _77169_ (_26523_, _26522_, _12125_);
  nor _77170_ (_26524_, _26523_, _26521_);
  not _77171_ (_26525_, _26524_);
  and _77172_ (_26526_, _26525_, _26520_);
  or _77173_ (_26527_, _26526_, _06687_);
  and _77174_ (_26528_, _12013_, _11958_);
  not _77175_ (_26529_, _26482_);
  and _77176_ (_26532_, _26529_, _11956_);
  or _77177_ (_26533_, _26532_, _12089_);
  or _77178_ (_26534_, _26533_, _26528_);
  nand _77179_ (_26535_, _26534_, _26527_);
  or _77180_ (_26536_, _26535_, _06236_);
  nor _77181_ (_26537_, _26482_, _12329_);
  and _77182_ (_26538_, _12329_, _12013_);
  nor _77183_ (_26539_, _26538_, _26537_);
  or _77184_ (_26540_, _26539_, _06643_);
  and _77185_ (_26541_, _26540_, _26536_);
  or _77186_ (_26543_, _26541_, _06295_);
  and _77187_ (_26544_, _12346_, _12013_);
  nor _77188_ (_26545_, _26482_, _12346_);
  nor _77189_ (_26546_, _26545_, _26544_);
  nor _77190_ (_26547_, _26546_, _12317_);
  nor _77191_ (_26548_, _26547_, _11924_);
  and _77192_ (_26549_, _26548_, _26543_);
  or _77193_ (_26550_, _26549_, _26446_);
  nand _77194_ (_26551_, _26550_, _06146_);
  and _77195_ (_26552_, _12189_, _06145_);
  nor _77196_ (_26554_, _26552_, _07388_);
  nand _77197_ (_26555_, _26554_, _26551_);
  nor _77198_ (_26556_, _08701_, _05760_);
  nor _77199_ (_26557_, _26556_, _25152_);
  and _77200_ (_26558_, _26557_, _26555_);
  or _77201_ (_26559_, _26558_, _26444_);
  nand _77202_ (_26560_, _26559_, _12369_);
  nor _77203_ (_26561_, _26436_, _12369_);
  nor _77204_ (_26562_, _26561_, _06255_);
  nand _77205_ (_26563_, _26562_, _26560_);
  and _77206_ (_26565_, _12188_, _06255_);
  nor _77207_ (_26566_, _26565_, _24882_);
  nand _77208_ (_26567_, _26566_, _26563_);
  and _77209_ (_26568_, _08701_, _24882_);
  nor _77210_ (_26569_, _26568_, _06254_);
  nand _77211_ (_26570_, _26569_, _26567_);
  and _77212_ (_26571_, _12188_, _06254_);
  nor _77213_ (_26572_, _26571_, _12387_);
  and _77214_ (_26573_, _26572_, _26570_);
  nor _77215_ (_26574_, _26436_, _12381_);
  or _77216_ (_26576_, _26574_, _26573_);
  nand _77217_ (_26577_, _26576_, _12385_);
  nor _77218_ (_26578_, _12188_, _12385_);
  nor _77219_ (_26579_, _26578_, _05870_);
  nand _77220_ (_26580_, _26579_, _26577_);
  nor _77221_ (_26581_, _26445_, _05805_);
  nor _77222_ (_26582_, _26581_, _06139_);
  and _77223_ (_26583_, _26582_, _26580_);
  and _77224_ (_26584_, _12189_, _06139_);
  or _77225_ (_26585_, _26584_, _26583_);
  nand _77226_ (_26587_, _26585_, _24791_);
  and _77227_ (_26588_, _08701_, _05791_);
  nor _77228_ (_26589_, _26588_, _06293_);
  nand _77229_ (_26590_, _26589_, _26587_);
  and _77230_ (_26591_, _12013_, _06293_);
  nor _77231_ (_26592_, _26591_, _13620_);
  nand _77232_ (_26593_, _26592_, _26590_);
  nor _77233_ (_26594_, _12188_, _06133_);
  nor _77234_ (_26595_, _26594_, _05787_);
  nand _77235_ (_26596_, _26595_, _26593_);
  and _77236_ (_26598_, _12013_, _05787_);
  nor _77237_ (_26599_, _26598_, _12412_);
  nand _77238_ (_26600_, _26599_, _26596_);
  nor _77239_ (_26601_, _26436_, _11922_);
  nor _77240_ (_26602_, _26601_, _06209_);
  nand _77241_ (_26603_, _26602_, _26600_);
  and _77242_ (_26604_, _12188_, _06209_);
  nor _77243_ (_26605_, _26604_, _05829_);
  nand _77244_ (_26606_, _26605_, _26603_);
  and _77245_ (_26607_, _08701_, _05829_);
  nor _77246_ (_26609_, _26607_, _12416_);
  nand _77247_ (_26610_, _26609_, _26606_);
  nor _77248_ (_26611_, _26467_, _12417_);
  nor _77249_ (_26612_, _26611_, _08788_);
  and _77250_ (_26613_, _26612_, _26610_);
  or _77251_ (_26614_, _26613_, _26443_);
  nand _77252_ (_26615_, _26614_, _06111_);
  and _77253_ (_26616_, _12014_, _06110_);
  nor _77254_ (_26617_, _26616_, _10751_);
  nand _77255_ (_26618_, _26617_, _26615_);
  and _77256_ (_26620_, _12188_, _10751_);
  nor _77257_ (_26621_, _26620_, _12431_);
  nand _77258_ (_26622_, _26621_, _26618_);
  and _77259_ (_26623_, _12451_, _12444_);
  nor _77260_ (_26624_, _26623_, _12452_);
  nor _77261_ (_26625_, _26624_, _12432_);
  nor _77262_ (_26626_, _26625_, _06208_);
  nand _77263_ (_26627_, _26626_, _26622_);
  and _77264_ (_26628_, _12188_, _06208_);
  nor _77265_ (_26629_, _26628_, _06076_);
  nand _77266_ (_26631_, _26629_, _26627_);
  and _77267_ (_26632_, _08701_, _06076_);
  nor _77268_ (_26633_, _26632_, _12473_);
  nand _77269_ (_26634_, _26633_, _26631_);
  and _77270_ (_26635_, _12188_, _11101_);
  nor _77271_ (_26636_, _26467_, _11101_);
  or _77272_ (_26637_, _26636_, _26635_);
  and _77273_ (_26638_, _26637_, _12473_);
  nor _77274_ (_26639_, _26638_, _12478_);
  and _77275_ (_26640_, _26639_, _26634_);
  or _77276_ (_26642_, _26640_, _26442_);
  nand _77277_ (_26643_, _26642_, _11916_);
  nor _77278_ (_26644_, _12188_, _11916_);
  nor _77279_ (_26645_, _26644_, _06297_);
  nand _77280_ (_26646_, _26645_, _26643_);
  and _77281_ (_26647_, _12013_, _06297_);
  nor _77282_ (_26648_, _26647_, _06402_);
  and _77283_ (_26649_, _26648_, _26646_);
  and _77284_ (_26650_, _12189_, _06402_);
  or _77285_ (_26651_, _26650_, _26649_);
  nand _77286_ (_26653_, _26651_, _05834_);
  and _77287_ (_26654_, _08701_, _12492_);
  nor _77288_ (_26655_, _26654_, _12496_);
  nand _77289_ (_26656_, _26655_, _26653_);
  and _77290_ (_26657_, _26467_, _11101_);
  nor _77291_ (_26658_, _12188_, _11101_);
  nor _77292_ (_26659_, _26658_, _12497_);
  not _77293_ (_26660_, _26659_);
  nor _77294_ (_26661_, _26660_, _26657_);
  nor _77295_ (_26662_, _26661_, _12505_);
  and _77296_ (_26664_, _26662_, _26656_);
  or _77297_ (_26665_, _26664_, _26441_);
  nand _77298_ (_26666_, _26665_, _10821_);
  nor _77299_ (_26667_, _12188_, _10821_);
  nor _77300_ (_26668_, _26667_, _06306_);
  nand _77301_ (_26669_, _26668_, _26666_);
  and _77302_ (_26670_, _12013_, _06306_);
  nor _77303_ (_26671_, _26670_, _06411_);
  and _77304_ (_26672_, _26671_, _26669_);
  and _77305_ (_26673_, _12189_, _06411_);
  or _77306_ (_26675_, _26673_, _26672_);
  nand _77307_ (_26676_, _26675_, _05848_);
  and _77308_ (_26677_, _08701_, _07124_);
  nor _77309_ (_26678_, _26677_, _12517_);
  nand _77310_ (_26679_, _26678_, _26676_);
  and _77311_ (_26680_, _12188_, \oc8051_golden_model_1.PSW [7]);
  nor _77312_ (_26681_, _26467_, \oc8051_golden_model_1.PSW [7]);
  or _77313_ (_26682_, _26681_, _26680_);
  and _77314_ (_26683_, _26682_, _12517_);
  nor _77315_ (_26684_, _26683_, _12522_);
  and _77316_ (_26686_, _26684_, _26679_);
  or _77317_ (_26687_, _26686_, _26440_);
  nand _77318_ (_26688_, _26687_, _10849_);
  nor _77319_ (_26689_, _12188_, _10849_);
  nor _77320_ (_26690_, _26689_, _06303_);
  nand _77321_ (_26691_, _26690_, _26688_);
  and _77322_ (_26692_, _12013_, _06303_);
  nor _77323_ (_26693_, _26692_, _06396_);
  and _77324_ (_26694_, _26693_, _26691_);
  and _77325_ (_26695_, _12189_, _06396_);
  or _77326_ (_26697_, _26695_, _26694_);
  nand _77327_ (_26698_, _26697_, _05843_);
  and _77328_ (_26699_, _08701_, _05842_);
  nor _77329_ (_26700_, _26699_, _12538_);
  nand _77330_ (_26701_, _26700_, _26698_);
  nand _77331_ (_26702_, _26467_, \oc8051_golden_model_1.PSW [7]);
  or _77332_ (_26703_, _12188_, \oc8051_golden_model_1.PSW [7]);
  and _77333_ (_26704_, _26703_, _12538_);
  and _77334_ (_26705_, _26704_, _26702_);
  nor _77335_ (_26706_, _26705_, _12547_);
  and _77336_ (_26708_, _26706_, _26701_);
  or _77337_ (_26709_, _26708_, _26439_);
  nand _77338_ (_26710_, _26709_, _10896_);
  nor _77339_ (_26711_, _12188_, _10896_);
  nor _77340_ (_26712_, _26711_, _10925_);
  nand _77341_ (_26713_, _26712_, _26710_);
  and _77342_ (_26714_, _26436_, _10925_);
  nor _77343_ (_26715_, _26714_, _06417_);
  and _77344_ (_26716_, _26715_, _26713_);
  or _77345_ (_26717_, _26716_, _26438_);
  nand _77346_ (_26719_, _26717_, _05846_);
  and _77347_ (_26720_, _08701_, _07142_);
  nor _77348_ (_26721_, _26720_, _06301_);
  nand _77349_ (_26722_, _26721_, _26719_);
  and _77350_ (_26723_, _26482_, _12682_);
  nor _77351_ (_26724_, _12013_, _12682_);
  or _77352_ (_26725_, _26724_, _06421_);
  nor _77353_ (_26726_, _26725_, _26723_);
  nor _77354_ (_26727_, _26726_, _12565_);
  and _77355_ (_26728_, _26727_, _26722_);
  or _77356_ (_26730_, _26728_, _26437_);
  nand _77357_ (_26731_, _26730_, _12690_);
  nor _77358_ (_26732_, _12690_, _12188_);
  nor _77359_ (_26733_, _26732_, _10262_);
  nand _77360_ (_26734_, _26733_, _26731_);
  and _77361_ (_26735_, _26436_, _10262_);
  nor _77362_ (_26736_, _26735_, _06167_);
  and _77363_ (_26737_, _26736_, _26734_);
  and _77364_ (_26738_, _08931_, _06167_);
  or _77365_ (_26739_, _26738_, _26737_);
  nand _77366_ (_26741_, _26739_, _12703_);
  and _77367_ (_26742_, _08701_, _05826_);
  nor _77368_ (_26743_, _26742_, _06165_);
  nand _77369_ (_26744_, _26743_, _26741_);
  nor _77370_ (_26745_, _26529_, _12682_);
  and _77371_ (_26746_, _12014_, _12682_);
  nor _77372_ (_26747_, _26746_, _26745_);
  and _77373_ (_26748_, _26747_, _06165_);
  nor _77374_ (_26749_, _26748_, _12712_);
  nand _77375_ (_26750_, _26749_, _26744_);
  nor _77376_ (_26751_, _26436_, _12711_);
  nor _77377_ (_26752_, _26751_, _06433_);
  and _77378_ (_26753_, _26752_, _26750_);
  or _77379_ (_26754_, _26753_, _26432_);
  nand _77380_ (_26755_, _26754_, _12719_);
  nor _77381_ (_26756_, _26445_, _12719_);
  nor _77382_ (_26757_, _26756_, _07577_);
  nand _77383_ (_26758_, _26757_, _26755_);
  and _77384_ (_26759_, _08701_, _07577_);
  nor _77385_ (_26760_, _26759_, _05748_);
  nand _77386_ (_26763_, _26760_, _26758_);
  and _77387_ (_26764_, _26747_, _05748_);
  nor _77388_ (_26765_, _26764_, _12737_);
  nand _77389_ (_26766_, _26765_, _26763_);
  nor _77390_ (_26767_, _26436_, _12735_);
  nor _77391_ (_26768_, _26767_, _06440_);
  and _77392_ (_26769_, _26768_, _26766_);
  or _77393_ (_26770_, _26769_, _26431_);
  nand _77394_ (_26771_, _26770_, _12744_);
  nor _77395_ (_26772_, _26445_, _12744_);
  nor _77396_ (_26774_, _26772_, _25019_);
  nand _77397_ (_26775_, _26774_, _26771_);
  and _77398_ (_26776_, _25019_, _08701_);
  nor _77399_ (_26777_, _26776_, _12754_);
  and _77400_ (_26778_, _26777_, _26775_);
  and _77401_ (_26779_, _26436_, _12754_);
  or _77402_ (_26780_, _26779_, _26778_);
  or _77403_ (_26781_, _26780_, _01321_);
  or _77404_ (_26782_, _01317_, \oc8051_golden_model_1.PC [5]);
  and _77405_ (_26783_, _26782_, _43100_);
  and _77406_ (_43693_, _26783_, _26781_);
  and _77407_ (_26785_, _08432_, _05426_);
  nor _77408_ (_26786_, _26785_, \oc8051_golden_model_1.PC [6]);
  nor _77409_ (_26787_, _26786_, _11894_);
  and _77410_ (_26788_, _26787_, _12754_);
  and _77411_ (_26789_, _08638_, _07577_);
  not _77412_ (_26790_, _26787_);
  and _77413_ (_26791_, _26790_, _10262_);
  and _77414_ (_26792_, _12181_, _06209_);
  or _77415_ (_26793_, _26792_, _05829_);
  nor _77416_ (_26795_, _25151_, _12180_);
  and _77417_ (_26796_, _12050_, _12010_);
  nor _77418_ (_26797_, _26796_, _12051_);
  or _77419_ (_26798_, _26797_, _12141_);
  or _77420_ (_26799_, _12139_, _12005_);
  and _77421_ (_26800_, _26799_, _06160_);
  nand _77422_ (_26801_, _26800_, _26798_);
  or _77423_ (_26802_, _12256_, _12181_);
  and _77424_ (_26803_, _12218_, _12185_);
  nor _77425_ (_26804_, _26803_, _12219_);
  nand _77426_ (_26806_, _26804_, _12256_);
  and _77427_ (_26807_, _26806_, _08445_);
  nand _77428_ (_26808_, _26807_, _26802_);
  and _77429_ (_26809_, _08638_, _06581_);
  and _77430_ (_26810_, _12181_, _07056_);
  or _77431_ (_26811_, _26810_, _06653_);
  nand _77432_ (_26812_, _12265_, \oc8051_golden_model_1.PC [6]);
  and _77433_ (_26813_, _26812_, _07057_);
  or _77434_ (_26814_, _26813_, _26811_);
  or _77435_ (_26815_, _26790_, _12266_);
  and _77436_ (_26817_, _26815_, _06582_);
  and _77437_ (_26818_, _26817_, _26814_);
  or _77438_ (_26819_, _26818_, _25055_);
  or _77439_ (_26820_, _26819_, _26809_);
  or _77440_ (_26821_, _26790_, _12263_);
  and _77441_ (_26822_, _26821_, _08443_);
  nand _77442_ (_26823_, _26822_, _26820_);
  and _77443_ (_26824_, _26823_, _12281_);
  nand _77444_ (_26825_, _26824_, _26808_);
  nand _77445_ (_26826_, _26825_, _26801_);
  and _77446_ (_26828_, _26826_, _12134_);
  and _77447_ (_26829_, _26787_, _12287_);
  or _77448_ (_26830_, _26829_, _06156_);
  or _77449_ (_26831_, _26830_, _26828_);
  and _77450_ (_26832_, _12181_, _06156_);
  nor _77451_ (_26833_, _26832_, _07485_);
  nand _77452_ (_26834_, _26833_, _26831_);
  nor _77453_ (_26835_, _08638_, _05764_);
  nor _77454_ (_26836_, _26835_, _06217_);
  nand _77455_ (_26837_, _26836_, _26834_);
  and _77456_ (_26839_, _12181_, _06217_);
  nor _77457_ (_26840_, _26839_, _12293_);
  nand _77458_ (_26841_, _26840_, _26837_);
  nor _77459_ (_26842_, _26790_, _12292_);
  nor _77460_ (_26843_, _26842_, _06220_);
  nand _77461_ (_26844_, _26843_, _26841_);
  and _77462_ (_26845_, _12181_, _06220_);
  nor _77463_ (_26846_, _26845_, _12302_);
  nand _77464_ (_26847_, _26846_, _26844_);
  nor _77465_ (_26848_, _26790_, _12300_);
  nor _77466_ (_26850_, _26848_, _06152_);
  and _77467_ (_26851_, _26850_, _26847_);
  and _77468_ (_26852_, _12181_, _06152_);
  or _77469_ (_26853_, _26852_, _26851_);
  nand _77470_ (_26854_, _26853_, _05769_);
  and _77471_ (_26855_, _08638_, _12304_);
  nor _77472_ (_26856_, _26855_, _06151_);
  nand _77473_ (_26857_, _26856_, _26854_);
  and _77474_ (_26858_, _12180_, _06151_);
  nor _77475_ (_26859_, _26858_, _12126_);
  nand _77476_ (_26861_, _26859_, _26857_);
  not _77477_ (_26862_, _25114_);
  and _77478_ (_26863_, _12120_, _12005_);
  not _77479_ (_26864_, _26797_);
  nor _77480_ (_26865_, _26864_, _12120_);
  or _77481_ (_26866_, _26865_, _26863_);
  nor _77482_ (_26867_, _26866_, _12125_);
  nor _77483_ (_26868_, _26867_, _26862_);
  nand _77484_ (_26869_, _26868_, _26861_);
  nor _77485_ (_26870_, _26864_, _12329_);
  and _77486_ (_26872_, _12329_, _12005_);
  nor _77487_ (_26873_, _26872_, _26870_);
  nor _77488_ (_26874_, _26873_, _06643_);
  or _77489_ (_26875_, _12005_, _11956_);
  or _77490_ (_26876_, _26797_, _11958_);
  and _77491_ (_26877_, _26876_, _06687_);
  and _77492_ (_26878_, _26877_, _26875_);
  nor _77493_ (_26879_, _26878_, _26874_);
  nand _77494_ (_26880_, _26879_, _26869_);
  nand _77495_ (_26881_, _26880_, _12317_);
  nand _77496_ (_26883_, _12346_, _12005_);
  nand _77497_ (_26884_, _26797_, _12347_);
  and _77498_ (_26885_, _26884_, _26883_);
  or _77499_ (_26886_, _26885_, _12317_);
  and _77500_ (_26887_, _26886_, _26881_);
  or _77501_ (_26888_, _26887_, _11924_);
  nand _77502_ (_26889_, _26787_, _11924_);
  and _77503_ (_26890_, _26889_, _26888_);
  nand _77504_ (_26891_, _26890_, _06146_);
  and _77505_ (_26892_, _12181_, _06145_);
  nor _77506_ (_26894_, _26892_, _07388_);
  nand _77507_ (_26895_, _26894_, _26891_);
  nor _77508_ (_26896_, _08638_, _05760_);
  nor _77509_ (_26897_, _26896_, _25152_);
  and _77510_ (_26898_, _26897_, _26895_);
  or _77511_ (_26899_, _26898_, _26795_);
  nand _77512_ (_26900_, _26899_, _12369_);
  nor _77513_ (_26901_, _26787_, _12369_);
  nor _77514_ (_26902_, _26901_, _06255_);
  nand _77515_ (_26903_, _26902_, _26900_);
  and _77516_ (_26905_, _12180_, _06255_);
  nor _77517_ (_26906_, _26905_, _24882_);
  nand _77518_ (_26907_, _26906_, _26903_);
  and _77519_ (_26908_, _08638_, _24882_);
  nor _77520_ (_26909_, _26908_, _06254_);
  nand _77521_ (_26910_, _26909_, _26907_);
  and _77522_ (_26911_, _12180_, _06254_);
  nor _77523_ (_26912_, _26911_, _12387_);
  nand _77524_ (_26913_, _26912_, _26910_);
  nor _77525_ (_26914_, _26787_, _12381_);
  nor _77526_ (_26916_, _26914_, _12386_);
  nand _77527_ (_26917_, _26916_, _26913_);
  nor _77528_ (_26918_, _12181_, _12385_);
  nor _77529_ (_26919_, _26918_, _05870_);
  and _77530_ (_26920_, _26919_, _26917_);
  nor _77531_ (_26921_, _26787_, _05805_);
  or _77532_ (_26922_, _26921_, _26920_);
  nand _77533_ (_26923_, _26922_, _06140_);
  and _77534_ (_26924_, _12181_, _06139_);
  nor _77535_ (_26925_, _26924_, _05791_);
  nand _77536_ (_26927_, _26925_, _26923_);
  nor _77537_ (_26928_, _08638_, _24791_);
  nor _77538_ (_26929_, _26928_, _06293_);
  and _77539_ (_26930_, _26929_, _26927_);
  and _77540_ (_26931_, _12006_, _06293_);
  or _77541_ (_26932_, _26931_, _26930_);
  and _77542_ (_26933_, _26932_, _06133_);
  nor _77543_ (_26934_, _12180_, _06133_);
  or _77544_ (_26935_, _26934_, _26933_);
  nand _77545_ (_26936_, _26935_, _06114_);
  and _77546_ (_26938_, _12006_, _05787_);
  nor _77547_ (_26939_, _26938_, _12412_);
  nand _77548_ (_26940_, _26939_, _26936_);
  nor _77549_ (_26941_, _26790_, _11922_);
  nor _77550_ (_26942_, _26941_, _06209_);
  and _77551_ (_26943_, _26942_, _26940_);
  or _77552_ (_26944_, _26943_, _26793_);
  nor _77553_ (_26945_, _08638_, _05830_);
  nor _77554_ (_26946_, _26945_, _12416_);
  and _77555_ (_26947_, _26946_, _26944_);
  nor _77556_ (_26949_, _26804_, _12417_);
  nor _77557_ (_26950_, _26949_, _26947_);
  nand _77558_ (_26951_, _26950_, _08787_);
  nor _77559_ (_26952_, _12181_, _08787_);
  nor _77560_ (_26953_, _26952_, _06110_);
  nand _77561_ (_26954_, _26953_, _26951_);
  and _77562_ (_26955_, _12006_, _06110_);
  nor _77563_ (_26956_, _26955_, _10751_);
  nand _77564_ (_26957_, _26956_, _26954_);
  and _77565_ (_26958_, _12180_, _10751_);
  nor _77566_ (_26960_, _26958_, _12431_);
  nand _77567_ (_26961_, _26960_, _26957_);
  and _77568_ (_26962_, _12453_, _12440_);
  nor _77569_ (_26963_, _26962_, _12454_);
  nor _77570_ (_26964_, _26963_, _12432_);
  nor _77571_ (_26965_, _26964_, _06208_);
  nand _77572_ (_26966_, _26965_, _26961_);
  and _77573_ (_26967_, _12180_, _06208_);
  nor _77574_ (_26968_, _26967_, _06076_);
  nand _77575_ (_26969_, _26968_, _26966_);
  and _77576_ (_26971_, _08638_, _06076_);
  nor _77577_ (_26972_, _26971_, _12473_);
  nand _77578_ (_26973_, _26972_, _26969_);
  and _77579_ (_26974_, _12180_, _11101_);
  and _77580_ (_26975_, _26804_, _12480_);
  or _77581_ (_26976_, _26975_, _26974_);
  and _77582_ (_26977_, _26976_, _12473_);
  nor _77583_ (_26978_, _26977_, _12478_);
  nand _77584_ (_26979_, _26978_, _26973_);
  nor _77585_ (_26980_, _26787_, _11919_);
  nor _77586_ (_26982_, _26980_, _11917_);
  nand _77587_ (_26983_, _26982_, _26979_);
  nor _77588_ (_26984_, _12181_, _11916_);
  nor _77589_ (_26985_, _26984_, _06297_);
  and _77590_ (_26986_, _26985_, _26983_);
  and _77591_ (_26987_, _12006_, _06297_);
  or _77592_ (_26988_, _26987_, _26986_);
  nand _77593_ (_26989_, _26988_, _07125_);
  and _77594_ (_26990_, _12181_, _06402_);
  nor _77595_ (_26991_, _26990_, _12492_);
  and _77596_ (_26993_, _26991_, _26989_);
  nor _77597_ (_26994_, _08638_, _05834_);
  or _77598_ (_26995_, _26994_, _26993_);
  nand _77599_ (_26996_, _26995_, _12497_);
  nor _77600_ (_26997_, _12181_, _11101_);
  and _77601_ (_26998_, _26804_, _11101_);
  or _77602_ (_26999_, _26998_, _26997_);
  and _77603_ (_27000_, _26999_, _12496_);
  nor _77604_ (_27001_, _27000_, _12505_);
  nand _77605_ (_27002_, _27001_, _26996_);
  nor _77606_ (_27004_, _26787_, _11914_);
  nor _77607_ (_27005_, _27004_, _10822_);
  nand _77608_ (_27006_, _27005_, _27002_);
  nor _77609_ (_27007_, _12181_, _10821_);
  nor _77610_ (_27008_, _27007_, _06306_);
  and _77611_ (_27009_, _27008_, _27006_);
  and _77612_ (_27010_, _12006_, _06306_);
  or _77613_ (_27011_, _27010_, _27009_);
  nand _77614_ (_27012_, _27011_, _07130_);
  and _77615_ (_27013_, _12181_, _06411_);
  nor _77616_ (_27015_, _27013_, _07124_);
  and _77617_ (_27016_, _27015_, _27012_);
  nor _77618_ (_27017_, _08638_, _05848_);
  or _77619_ (_27018_, _27017_, _27016_);
  nand _77620_ (_27019_, _27018_, _12518_);
  and _77621_ (_27020_, _12180_, \oc8051_golden_model_1.PSW [7]);
  and _77622_ (_27021_, _26804_, _10693_);
  or _77623_ (_27022_, _27021_, _27020_);
  and _77624_ (_27023_, _27022_, _12517_);
  nor _77625_ (_27024_, _27023_, _12522_);
  nand _77626_ (_27026_, _27024_, _27019_);
  nor _77627_ (_27027_, _26787_, _11912_);
  nor _77628_ (_27028_, _27027_, _10850_);
  nand _77629_ (_27029_, _27028_, _27026_);
  nor _77630_ (_27030_, _12181_, _10849_);
  nor _77631_ (_27031_, _27030_, _06303_);
  and _77632_ (_27032_, _27031_, _27029_);
  and _77633_ (_27033_, _12006_, _06303_);
  or _77634_ (_27034_, _27033_, _27032_);
  nand _77635_ (_27035_, _27034_, _08824_);
  and _77636_ (_27037_, _12181_, _06396_);
  nor _77637_ (_27038_, _27037_, _05842_);
  and _77638_ (_27039_, _27038_, _27035_);
  nor _77639_ (_27040_, _08638_, _05843_);
  or _77640_ (_27041_, _27040_, _27039_);
  nand _77641_ (_27042_, _27041_, _12539_);
  or _77642_ (_27043_, _26804_, _10693_);
  or _77643_ (_27044_, _12180_, \oc8051_golden_model_1.PSW [7]);
  and _77644_ (_27045_, _27044_, _12538_);
  and _77645_ (_27046_, _27045_, _27043_);
  nor _77646_ (_27048_, _27046_, _12547_);
  nand _77647_ (_27049_, _27048_, _27042_);
  nor _77648_ (_27050_, _26787_, _11907_);
  nor _77649_ (_27051_, _27050_, _10897_);
  nand _77650_ (_27052_, _27051_, _27049_);
  nor _77651_ (_27053_, _12181_, _10896_);
  nor _77652_ (_27054_, _27053_, _10925_);
  nand _77653_ (_27055_, _27054_, _27052_);
  and _77654_ (_27056_, _26790_, _10925_);
  nor _77655_ (_27057_, _27056_, _06417_);
  nand _77656_ (_27059_, _27057_, _27055_);
  and _77657_ (_27060_, _09207_, _06417_);
  nor _77658_ (_27061_, _27060_, _07142_);
  nand _77659_ (_27062_, _27061_, _27059_);
  and _77660_ (_27063_, _08638_, _07142_);
  nor _77661_ (_27064_, _27063_, _06301_);
  nand _77662_ (_27065_, _27064_, _27062_);
  and _77663_ (_27066_, _26864_, _12682_);
  nor _77664_ (_27067_, _12005_, _12682_);
  or _77665_ (_27068_, _27067_, _06421_);
  nor _77666_ (_27070_, _27068_, _27066_);
  nor _77667_ (_27071_, _27070_, _12565_);
  nand _77668_ (_27072_, _27071_, _27065_);
  nor _77669_ (_27073_, _26787_, _11905_);
  nor _77670_ (_27074_, _27073_, _12691_);
  nand _77671_ (_27075_, _27074_, _27072_);
  nor _77672_ (_27076_, _12690_, _12181_);
  nor _77673_ (_27077_, _27076_, _10262_);
  and _77674_ (_27078_, _27077_, _27075_);
  or _77675_ (_27079_, _27078_, _26791_);
  nand _77676_ (_27081_, _27079_, _06168_);
  and _77677_ (_27082_, _08883_, _06167_);
  nor _77678_ (_27083_, _27082_, _05826_);
  nand _77679_ (_27084_, _27083_, _27081_);
  nor _77680_ (_27085_, _08638_, _12703_);
  nor _77681_ (_27086_, _27085_, _06165_);
  and _77682_ (_27087_, _27086_, _27084_);
  and _77683_ (_27088_, _12006_, _12682_);
  nor _77684_ (_27089_, _26797_, _12682_);
  nor _77685_ (_27090_, _27089_, _27088_);
  nor _77686_ (_27092_, _27090_, _06166_);
  or _77687_ (_27093_, _27092_, _27087_);
  and _77688_ (_27094_, _27093_, _12711_);
  nor _77689_ (_27095_, _26787_, _12711_);
  or _77690_ (_27096_, _27095_, _27094_);
  nand _77691_ (_27097_, _27096_, _06829_);
  and _77692_ (_27098_, _12181_, _06433_);
  nor _77693_ (_27099_, _27098_, _25721_);
  nand _77694_ (_27100_, _27099_, _27097_);
  nor _77695_ (_27101_, _26790_, _12719_);
  nor _77696_ (_27103_, _27101_, _07577_);
  and _77697_ (_27104_, _27103_, _27100_);
  or _77698_ (_27105_, _27104_, _26789_);
  nand _77699_ (_27106_, _27105_, _05749_);
  nor _77700_ (_27107_, _27090_, _05749_);
  nor _77701_ (_27108_, _27107_, _12737_);
  nand _77702_ (_27109_, _27108_, _27106_);
  nor _77703_ (_27110_, _26790_, _12735_);
  nor _77704_ (_27111_, _27110_, _06440_);
  nand _77705_ (_27112_, _27111_, _27109_);
  and _77706_ (_27114_, _12181_, _06440_);
  nor _77707_ (_27115_, _27114_, _26415_);
  nand _77708_ (_27116_, _27115_, _27112_);
  nor _77709_ (_27117_, _26790_, _12744_);
  nor _77710_ (_27118_, _27117_, _25019_);
  nand _77711_ (_27119_, _27118_, _27116_);
  and _77712_ (_27120_, _25019_, _08638_);
  nor _77713_ (_27121_, _27120_, _12754_);
  and _77714_ (_27122_, _27121_, _27119_);
  or _77715_ (_27123_, _27122_, _26788_);
  or _77716_ (_27125_, _27123_, _01321_);
  or _77717_ (_27126_, _01317_, \oc8051_golden_model_1.PC [6]);
  and _77718_ (_27127_, _27126_, _43100_);
  and _77719_ (_43694_, _27127_, _27125_);
  and _77720_ (_27128_, _08437_, _06440_);
  nor _77721_ (_27129_, _11894_, \oc8051_golden_model_1.PC [7]);
  nor _77722_ (_27130_, _27129_, _11895_);
  nor _77723_ (_27131_, _27130_, _11905_);
  nor _77724_ (_27132_, _27130_, _11907_);
  nor _77725_ (_27133_, _27130_, _11912_);
  nor _77726_ (_27135_, _27130_, _11914_);
  nor _77727_ (_27136_, _27130_, _11919_);
  nor _77728_ (_27137_, _08787_, _08437_);
  nor _77729_ (_27138_, _25151_, _08437_);
  not _77730_ (_27139_, _27130_);
  nand _77731_ (_27140_, _27139_, _11924_);
  and _77732_ (_27141_, _12141_, _09180_);
  or _77733_ (_27142_, _12001_, _12002_);
  and _77734_ (_27143_, _27142_, _12052_);
  nor _77735_ (_27144_, _27142_, _12052_);
  nor _77736_ (_27146_, _27144_, _27143_);
  and _77737_ (_27147_, _27146_, _12139_);
  or _77738_ (_27148_, _27147_, _27141_);
  and _77739_ (_27149_, _27148_, _06160_);
  or _77740_ (_27150_, _12176_, _12177_);
  and _77741_ (_27151_, _27150_, _12220_);
  nor _77742_ (_27152_, _27150_, _12220_);
  nor _77743_ (_27153_, _27152_, _27151_);
  and _77744_ (_27154_, _27153_, _12256_);
  and _77745_ (_27155_, _12258_, _08437_);
  or _77746_ (_27157_, _27155_, _27154_);
  and _77747_ (_27158_, _27157_, _08445_);
  nor _77748_ (_27159_, _08395_, _06582_);
  nand _77749_ (_27160_, _08573_, _07056_);
  and _77750_ (_27161_, _27160_, _12264_);
  and _77751_ (_27162_, _12265_, \oc8051_golden_model_1.PC [7]);
  or _77752_ (_27163_, _27162_, _07056_);
  and _77753_ (_27164_, _27163_, _27161_);
  or _77754_ (_27165_, _27139_, _12266_);
  nand _77755_ (_27166_, _27165_, _12263_);
  or _77756_ (_27168_, _27166_, _27164_);
  and _77757_ (_27169_, _27168_, _06582_);
  or _77758_ (_27170_, _27169_, _27159_);
  or _77759_ (_27171_, _27130_, _12263_);
  and _77760_ (_27172_, _27171_, _08443_);
  and _77761_ (_27173_, _27172_, _27170_);
  or _77762_ (_27174_, _27173_, _07064_);
  or _77763_ (_27175_, _27174_, _27158_);
  nand _77764_ (_27176_, _27139_, _07064_);
  and _77765_ (_27177_, _27176_, _06161_);
  and _77766_ (_27179_, _27177_, _27175_);
  or _77767_ (_27180_, _27179_, _27149_);
  or _77768_ (_27181_, _27180_, _24821_);
  or _77769_ (_27182_, _27130_, _12134_);
  and _77770_ (_27183_, _27182_, _06157_);
  and _77771_ (_27184_, _27183_, _27181_);
  and _77772_ (_27185_, _08437_, _06156_);
  or _77773_ (_27186_, _27185_, _07485_);
  or _77774_ (_27187_, _27186_, _27184_);
  nand _77775_ (_27188_, _08395_, _07485_);
  and _77776_ (_27190_, _27188_, _07075_);
  and _77777_ (_27191_, _27190_, _27187_);
  nand _77778_ (_27192_, _08437_, _06217_);
  nand _77779_ (_27193_, _27192_, _12292_);
  or _77780_ (_27194_, _27193_, _27191_);
  or _77781_ (_27195_, _27130_, _12292_);
  and _77782_ (_27196_, _27195_, _06229_);
  and _77783_ (_27197_, _27196_, _27194_);
  nand _77784_ (_27198_, _08437_, _06220_);
  nand _77785_ (_27199_, _27198_, _12300_);
  or _77786_ (_27201_, _27199_, _27197_);
  or _77787_ (_27202_, _27130_, _12300_);
  and _77788_ (_27203_, _27202_, _06153_);
  and _77789_ (_27204_, _27203_, _27201_);
  and _77790_ (_27205_, _08437_, _06152_);
  or _77791_ (_27206_, _27205_, _12304_);
  or _77792_ (_27207_, _27206_, _27204_);
  nand _77793_ (_27208_, _08395_, _12304_);
  and _77794_ (_27209_, _27208_, _07191_);
  and _77795_ (_27210_, _27209_, _27207_);
  nand _77796_ (_27212_, _08437_, _06151_);
  nand _77797_ (_27213_, _27212_, _12125_);
  or _77798_ (_27214_, _27213_, _27210_);
  not _77799_ (_27215_, _27146_);
  nor _77800_ (_27216_, _27215_, _12120_);
  and _77801_ (_27217_, _12120_, _09180_);
  or _77802_ (_27218_, _27217_, _12125_);
  or _77803_ (_27219_, _27218_, _27216_);
  and _77804_ (_27220_, _27219_, _12089_);
  and _77805_ (_27221_, _27220_, _27214_);
  and _77806_ (_27223_, _27146_, _11956_);
  and _77807_ (_27224_, _11958_, _09180_);
  or _77808_ (_27225_, _27224_, _27223_);
  and _77809_ (_27226_, _27225_, _06687_);
  or _77810_ (_27227_, _27226_, _06236_);
  or _77811_ (_27228_, _27227_, _27221_);
  and _77812_ (_27229_, _12329_, _09180_);
  nor _77813_ (_27230_, _27215_, _12329_);
  or _77814_ (_27231_, _27230_, _06643_);
  or _77815_ (_27232_, _27231_, _27229_);
  and _77816_ (_27234_, _27232_, _12317_);
  and _77817_ (_27235_, _27234_, _27228_);
  or _77818_ (_27236_, _27146_, _12346_);
  nand _77819_ (_27237_, _12346_, _09181_);
  and _77820_ (_27238_, _27237_, _06295_);
  and _77821_ (_27239_, _27238_, _27236_);
  or _77822_ (_27240_, _27239_, _11924_);
  or _77823_ (_27241_, _27240_, _27235_);
  nand _77824_ (_27242_, _27241_, _27140_);
  nand _77825_ (_27243_, _27242_, _06146_);
  and _77826_ (_27245_, _08573_, _06145_);
  nor _77827_ (_27246_, _27245_, _07388_);
  nand _77828_ (_27247_, _27246_, _27243_);
  nor _77829_ (_27248_, _08395_, _05760_);
  nor _77830_ (_27249_, _27248_, _25152_);
  and _77831_ (_27250_, _27249_, _27247_);
  or _77832_ (_27251_, _27250_, _27138_);
  nand _77833_ (_27252_, _27251_, _12369_);
  nor _77834_ (_27253_, _27130_, _12369_);
  nor _77835_ (_27254_, _27253_, _06255_);
  nand _77836_ (_27256_, _27254_, _27252_);
  and _77837_ (_27257_, _08437_, _06255_);
  nor _77838_ (_27258_, _27257_, _24882_);
  nand _77839_ (_27259_, _27258_, _27256_);
  and _77840_ (_27260_, _08395_, _24882_);
  nor _77841_ (_27261_, _27260_, _06254_);
  nand _77842_ (_27262_, _27261_, _27259_);
  and _77843_ (_27263_, _08437_, _06254_);
  nor _77844_ (_27264_, _27263_, _12387_);
  and _77845_ (_27265_, _27264_, _27262_);
  nor _77846_ (_27267_, _27130_, _12381_);
  or _77847_ (_27268_, _27267_, _27265_);
  nand _77848_ (_27269_, _27268_, _12385_);
  nor _77849_ (_27270_, _12385_, _08437_);
  nor _77850_ (_27271_, _27270_, _05870_);
  nand _77851_ (_27272_, _27271_, _27269_);
  nor _77852_ (_27273_, _27139_, _05805_);
  nor _77853_ (_27274_, _27273_, _06139_);
  and _77854_ (_27275_, _27274_, _27272_);
  and _77855_ (_27276_, _08573_, _06139_);
  or _77856_ (_27278_, _27276_, _27275_);
  nand _77857_ (_27279_, _27278_, _24791_);
  and _77858_ (_27280_, _08395_, _05791_);
  nor _77859_ (_27281_, _27280_, _06293_);
  nand _77860_ (_27282_, _27281_, _27279_);
  and _77861_ (_27283_, _09180_, _06293_);
  nor _77862_ (_27284_, _27283_, _13620_);
  nand _77863_ (_27285_, _27284_, _27282_);
  nor _77864_ (_27286_, _08437_, _06133_);
  nor _77865_ (_27287_, _27286_, _05787_);
  nand _77866_ (_27289_, _27287_, _27285_);
  and _77867_ (_27290_, _09180_, _05787_);
  nor _77868_ (_27291_, _27290_, _12412_);
  nand _77869_ (_27292_, _27291_, _27289_);
  nor _77870_ (_27293_, _27130_, _11922_);
  nor _77871_ (_27294_, _27293_, _06209_);
  nand _77872_ (_27295_, _27294_, _27292_);
  and _77873_ (_27296_, _08437_, _06209_);
  nor _77874_ (_27297_, _27296_, _05829_);
  nand _77875_ (_27298_, _27297_, _27295_);
  and _77876_ (_27300_, _08395_, _05829_);
  nor _77877_ (_27301_, _27300_, _12416_);
  nand _77878_ (_27302_, _27301_, _27298_);
  and _77879_ (_27303_, _27153_, _12416_);
  nor _77880_ (_27304_, _27303_, _08788_);
  and _77881_ (_27305_, _27304_, _27302_);
  or _77882_ (_27306_, _27305_, _27137_);
  nand _77883_ (_27307_, _27306_, _06111_);
  and _77884_ (_27308_, _09181_, _06110_);
  nor _77885_ (_27309_, _27308_, _10751_);
  and _77886_ (_27311_, _27309_, _27307_);
  and _77887_ (_27312_, _10751_, _08437_);
  or _77888_ (_27313_, _27312_, _27311_);
  nand _77889_ (_27314_, _27313_, _12432_);
  or _77890_ (_27315_, _12436_, _12435_);
  nor _77891_ (_27316_, _27315_, _12455_);
  not _77892_ (_27317_, _27316_);
  and _77893_ (_27318_, _27315_, _12455_);
  nor _77894_ (_27319_, _27318_, _12432_);
  and _77895_ (_27320_, _27319_, _27317_);
  nor _77896_ (_27322_, _27320_, _06208_);
  and _77897_ (_27323_, _27322_, _27314_);
  and _77898_ (_27324_, _08573_, _06208_);
  or _77899_ (_27325_, _27324_, _27323_);
  nand _77900_ (_27326_, _27325_, _05836_);
  and _77901_ (_27327_, _08395_, _06076_);
  nor _77902_ (_27328_, _27327_, _12473_);
  nand _77903_ (_27329_, _27328_, _27326_);
  and _77904_ (_27330_, _11101_, _08437_);
  and _77905_ (_27331_, _27153_, _12480_);
  or _77906_ (_27332_, _27331_, _27330_);
  and _77907_ (_27333_, _27332_, _12473_);
  nor _77908_ (_27334_, _27333_, _12478_);
  and _77909_ (_27335_, _27334_, _27329_);
  or _77910_ (_27336_, _27335_, _27136_);
  nand _77911_ (_27337_, _27336_, _11916_);
  nor _77912_ (_27338_, _11916_, _08437_);
  nor _77913_ (_27339_, _27338_, _06297_);
  nand _77914_ (_27340_, _27339_, _27337_);
  and _77915_ (_27341_, _09180_, _06297_);
  nor _77916_ (_27344_, _27341_, _06402_);
  and _77917_ (_27345_, _27344_, _27340_);
  and _77918_ (_27346_, _08573_, _06402_);
  or _77919_ (_27347_, _27346_, _27345_);
  nand _77920_ (_27348_, _27347_, _05834_);
  and _77921_ (_27349_, _08395_, _12492_);
  nor _77922_ (_27350_, _27349_, _12496_);
  nand _77923_ (_27351_, _27350_, _27348_);
  nor _77924_ (_27352_, _27153_, _12480_);
  nor _77925_ (_27353_, _11101_, _08437_);
  nor _77926_ (_27355_, _27353_, _12497_);
  not _77927_ (_27356_, _27355_);
  nor _77928_ (_27357_, _27356_, _27352_);
  nor _77929_ (_27358_, _27357_, _12505_);
  and _77930_ (_27359_, _27358_, _27351_);
  or _77931_ (_27360_, _27359_, _27135_);
  nand _77932_ (_27361_, _27360_, _10821_);
  nor _77933_ (_27362_, _10821_, _08437_);
  nor _77934_ (_27363_, _27362_, _06306_);
  nand _77935_ (_27364_, _27363_, _27361_);
  and _77936_ (_27366_, _09180_, _06306_);
  nor _77937_ (_27367_, _27366_, _06411_);
  and _77938_ (_27368_, _27367_, _27364_);
  and _77939_ (_27369_, _08573_, _06411_);
  or _77940_ (_27370_, _27369_, _27368_);
  nand _77941_ (_27371_, _27370_, _05848_);
  and _77942_ (_27372_, _08395_, _07124_);
  nor _77943_ (_27373_, _27372_, _12517_);
  nand _77944_ (_27374_, _27373_, _27371_);
  and _77945_ (_27375_, _08437_, \oc8051_golden_model_1.PSW [7]);
  and _77946_ (_27377_, _27153_, _10693_);
  or _77947_ (_27378_, _27377_, _27375_);
  and _77948_ (_27379_, _27378_, _12517_);
  nor _77949_ (_27380_, _27379_, _12522_);
  and _77950_ (_27381_, _27380_, _27374_);
  or _77951_ (_27382_, _27381_, _27133_);
  nand _77952_ (_27383_, _27382_, _10849_);
  nor _77953_ (_27384_, _10849_, _08437_);
  nor _77954_ (_27385_, _27384_, _06303_);
  nand _77955_ (_27386_, _27385_, _27383_);
  and _77956_ (_27388_, _09180_, _06303_);
  nor _77957_ (_27389_, _27388_, _06396_);
  and _77958_ (_27390_, _27389_, _27386_);
  and _77959_ (_27391_, _08573_, _06396_);
  or _77960_ (_27392_, _27391_, _27390_);
  nand _77961_ (_27393_, _27392_, _05843_);
  and _77962_ (_27394_, _08395_, _05842_);
  nor _77963_ (_27395_, _27394_, _12538_);
  nand _77964_ (_27396_, _27395_, _27393_);
  and _77965_ (_27397_, _08437_, _10693_);
  and _77966_ (_27399_, _27153_, \oc8051_golden_model_1.PSW [7]);
  or _77967_ (_27400_, _27399_, _27397_);
  and _77968_ (_27401_, _27400_, _12538_);
  nor _77969_ (_27402_, _27401_, _12547_);
  and _77970_ (_27403_, _27402_, _27396_);
  or _77971_ (_27404_, _27403_, _27132_);
  nand _77972_ (_27405_, _27404_, _10896_);
  nor _77973_ (_27406_, _10896_, _08437_);
  nor _77974_ (_27407_, _27406_, _10925_);
  nand _77975_ (_27408_, _27407_, _27405_);
  and _77976_ (_27410_, _27130_, _10925_);
  nor _77977_ (_27411_, _27410_, _06417_);
  and _77978_ (_27412_, _27411_, _27408_);
  and _77979_ (_27413_, _08838_, _06417_);
  or _77980_ (_27414_, _27413_, _27412_);
  nand _77981_ (_27415_, _27414_, _05846_);
  and _77982_ (_27416_, _08395_, _07142_);
  nor _77983_ (_27417_, _27416_, _06301_);
  nand _77984_ (_27418_, _27417_, _27415_);
  and _77985_ (_27419_, _27215_, _12682_);
  nor _77986_ (_27421_, _09180_, _12682_);
  or _77987_ (_27422_, _27421_, _06421_);
  nor _77988_ (_27423_, _27422_, _27419_);
  nor _77989_ (_27424_, _27423_, _12565_);
  and _77990_ (_27425_, _27424_, _27418_);
  or _77991_ (_27426_, _27425_, _27131_);
  nand _77992_ (_27427_, _27426_, _12690_);
  nor _77993_ (_27428_, _12690_, _08437_);
  nor _77994_ (_27429_, _27428_, _10262_);
  nand _77995_ (_27430_, _27429_, _27427_);
  and _77996_ (_27432_, _27130_, _10262_);
  nor _77997_ (_27433_, _27432_, _06167_);
  and _77998_ (_27434_, _27433_, _27430_);
  and _77999_ (_27435_, _08838_, _06167_);
  or _78000_ (_27436_, _27435_, _27434_);
  nand _78001_ (_27437_, _27436_, _12703_);
  and _78002_ (_27438_, _08395_, _05826_);
  nor _78003_ (_27439_, _27438_, _06165_);
  nand _78004_ (_27440_, _27439_, _27437_);
  nor _78005_ (_27441_, _27146_, _12682_);
  and _78006_ (_27443_, _09181_, _12682_);
  nor _78007_ (_27444_, _27443_, _27441_);
  and _78008_ (_27445_, _27444_, _06165_);
  nor _78009_ (_27446_, _27445_, _12712_);
  nand _78010_ (_27447_, _27446_, _27440_);
  nor _78011_ (_27448_, _27130_, _12711_);
  nor _78012_ (_27449_, _27448_, _06433_);
  nand _78013_ (_27450_, _27449_, _27447_);
  and _78014_ (_27451_, _08437_, _06433_);
  nor _78015_ (_27452_, _27451_, _25721_);
  and _78016_ (_27454_, _27452_, _27450_);
  nor _78017_ (_27455_, _27130_, _12719_);
  or _78018_ (_27456_, _27455_, _27454_);
  nand _78019_ (_27457_, _27456_, _07160_);
  and _78020_ (_27458_, _08395_, _07577_);
  nor _78021_ (_27459_, _27458_, _05748_);
  nand _78022_ (_27460_, _27459_, _27457_);
  and _78023_ (_27461_, _27444_, _05748_);
  nor _78024_ (_27462_, _27461_, _12737_);
  nand _78025_ (_27463_, _27462_, _27460_);
  nor _78026_ (_27465_, _27130_, _12735_);
  nor _78027_ (_27466_, _27465_, _06440_);
  and _78028_ (_27467_, _27466_, _27463_);
  or _78029_ (_27468_, _27467_, _27128_);
  nand _78030_ (_27469_, _27468_, _12744_);
  nor _78031_ (_27470_, _27139_, _12744_);
  nor _78032_ (_27471_, _27470_, _25019_);
  nand _78033_ (_27472_, _27471_, _27469_);
  and _78034_ (_27473_, _25019_, _08395_);
  nor _78035_ (_27474_, _27473_, _12754_);
  and _78036_ (_27476_, _27474_, _27472_);
  and _78037_ (_27477_, _27130_, _12754_);
  or _78038_ (_27478_, _27477_, _27476_);
  or _78039_ (_27479_, _27478_, _01321_);
  or _78040_ (_27480_, _01317_, \oc8051_golden_model_1.PC [7]);
  and _78041_ (_27481_, _27480_, _43100_);
  and _78042_ (_43695_, _27481_, _27479_);
  nor _78043_ (_27482_, _12747_, _06107_);
  nor _78044_ (_27483_, _12723_, _06107_);
  nor _78045_ (_27484_, _12538_, _05842_);
  nor _78046_ (_27486_, _12416_, _05829_);
  and _78047_ (_27487_, _12224_, _06209_);
  and _78048_ (_27488_, _12224_, _06152_);
  nor _78049_ (_27489_, _06217_, _07485_);
  and _78050_ (_27490_, _12224_, _06156_);
  and _78051_ (_27491_, _11895_, \oc8051_golden_model_1.PC [8]);
  nor _78052_ (_27492_, _11895_, \oc8051_golden_model_1.PC [8]);
  nor _78053_ (_27493_, _27492_, _27491_);
  nor _78054_ (_27494_, _27493_, _12266_);
  not _78055_ (_27495_, _12224_);
  and _78056_ (_27497_, _27495_, _07056_);
  nor _78057_ (_27498_, _07056_, \oc8051_golden_model_1.PC [8]);
  and _78058_ (_27499_, _27498_, _12265_);
  or _78059_ (_27500_, _27499_, _27497_);
  and _78060_ (_27501_, _27500_, _12264_);
  nor _78061_ (_27502_, _27501_, _27494_);
  nor _78062_ (_27503_, _27502_, _24800_);
  nor _78063_ (_27504_, _27493_, _12263_);
  nor _78064_ (_27505_, _27504_, _27503_);
  nor _78065_ (_27506_, _27505_, _08445_);
  or _78066_ (_27508_, _12256_, _27495_);
  nor _78067_ (_27509_, _12227_, _12222_);
  nor _78068_ (_27510_, _27509_, _12228_);
  nand _78069_ (_27511_, _27510_, _12256_);
  and _78070_ (_27512_, _27511_, _08445_);
  and _78071_ (_27513_, _27512_, _27508_);
  or _78072_ (_27514_, _27513_, _27506_);
  nand _78073_ (_27515_, _27514_, _07065_);
  not _78074_ (_27516_, _27493_);
  and _78075_ (_27517_, _27516_, _07064_);
  nor _78076_ (_27519_, _27517_, _06160_);
  nand _78077_ (_27520_, _27519_, _27515_);
  or _78078_ (_27521_, _12139_, _12056_);
  nor _78079_ (_27522_, _12060_, _12054_);
  nor _78080_ (_27523_, _27522_, _12061_);
  or _78081_ (_27524_, _27523_, _12141_);
  and _78082_ (_27525_, _27524_, _06160_);
  nand _78083_ (_27526_, _27525_, _27521_);
  and _78084_ (_27527_, _27526_, _12134_);
  nand _78085_ (_27528_, _27527_, _27520_);
  nor _78086_ (_27530_, _27493_, _12134_);
  nor _78087_ (_27531_, _27530_, _06156_);
  and _78088_ (_27532_, _27531_, _27528_);
  or _78089_ (_27533_, _27532_, _27490_);
  nand _78090_ (_27534_, _27533_, _27489_);
  and _78091_ (_27535_, _12224_, _06217_);
  nor _78092_ (_27536_, _27535_, _12293_);
  nand _78093_ (_27537_, _27536_, _27534_);
  nor _78094_ (_27538_, _27493_, _12292_);
  nor _78095_ (_27539_, _27538_, _06220_);
  nand _78096_ (_27541_, _27539_, _27537_);
  and _78097_ (_27542_, _12224_, _06220_);
  nor _78098_ (_27543_, _27542_, _12302_);
  nand _78099_ (_27544_, _27543_, _27541_);
  nor _78100_ (_27545_, _27493_, _12300_);
  nor _78101_ (_27546_, _27545_, _06152_);
  and _78102_ (_27547_, _27546_, _27544_);
  or _78103_ (_27548_, _27547_, _27488_);
  nand _78104_ (_27549_, _27548_, _12305_);
  and _78105_ (_27550_, _12224_, _06151_);
  nor _78106_ (_27552_, _27550_, _12126_);
  nand _78107_ (_27553_, _27552_, _27549_);
  and _78108_ (_27554_, _12120_, _12056_);
  not _78109_ (_27555_, _27523_);
  nor _78110_ (_27556_, _27555_, _12120_);
  or _78111_ (_27557_, _27556_, _27554_);
  nor _78112_ (_27558_, _27557_, _12125_);
  nor _78113_ (_27559_, _27558_, _26862_);
  nand _78114_ (_27560_, _27559_, _27553_);
  nor _78115_ (_27561_, _27555_, _12329_);
  and _78116_ (_27563_, _12329_, _12056_);
  nor _78117_ (_27564_, _27563_, _27561_);
  nor _78118_ (_27565_, _27564_, _06643_);
  or _78119_ (_27566_, _12056_, _11956_);
  nand _78120_ (_27567_, _27555_, _11956_);
  and _78121_ (_27568_, _27567_, _06687_);
  and _78122_ (_27569_, _27568_, _27566_);
  nor _78123_ (_27570_, _27569_, _27565_);
  nand _78124_ (_27571_, _27570_, _27560_);
  nand _78125_ (_27572_, _27571_, _12317_);
  nor _78126_ (_27574_, _27523_, _12346_);
  and _78127_ (_27575_, _12346_, _12057_);
  nor _78128_ (_27576_, _27575_, _12317_);
  not _78129_ (_27577_, _27576_);
  nor _78130_ (_27578_, _27577_, _27574_);
  nor _78131_ (_27579_, _27578_, _11924_);
  nand _78132_ (_27580_, _27579_, _27572_);
  and _78133_ (_27581_, _27516_, _11924_);
  nor _78134_ (_27582_, _27581_, _06145_);
  nand _78135_ (_27583_, _27582_, _27580_);
  and _78136_ (_27585_, _12224_, _06145_);
  nor _78137_ (_27586_, _27585_, _07388_);
  nand _78138_ (_27587_, _27586_, _27583_);
  nand _78139_ (_27588_, _27587_, _25151_);
  nor _78140_ (_27589_, _25151_, _27495_);
  nor _78141_ (_27590_, _27589_, _12373_);
  nand _78142_ (_27591_, _27590_, _27588_);
  nor _78143_ (_27592_, _27493_, _12369_);
  nor _78144_ (_27593_, _27592_, _06255_);
  nand _78145_ (_27594_, _27593_, _27591_);
  and _78146_ (_27596_, _12224_, _06255_);
  nor _78147_ (_27597_, _27596_, _24882_);
  nand _78148_ (_27598_, _27597_, _27594_);
  nand _78149_ (_27599_, _27598_, _13843_);
  and _78150_ (_27600_, _12224_, _06254_);
  nor _78151_ (_27601_, _27600_, _12387_);
  nand _78152_ (_27602_, _27601_, _27599_);
  nor _78153_ (_27603_, _27493_, _12381_);
  nor _78154_ (_27604_, _27603_, _12386_);
  and _78155_ (_27605_, _27604_, _27602_);
  nor _78156_ (_27607_, _27495_, _12385_);
  or _78157_ (_27608_, _27607_, _05870_);
  nor _78158_ (_27609_, _27608_, _27605_);
  nor _78159_ (_27610_, _27493_, _05805_);
  or _78160_ (_27611_, _27610_, _27609_);
  nand _78161_ (_27612_, _27611_, _06140_);
  and _78162_ (_27613_, _27495_, _06139_);
  nor _78163_ (_27614_, _06293_, _05791_);
  not _78164_ (_27615_, _27614_);
  nor _78165_ (_27616_, _27615_, _27613_);
  nand _78166_ (_27618_, _27616_, _27612_);
  and _78167_ (_27619_, _12056_, _06293_);
  nor _78168_ (_27620_, _27619_, _13620_);
  nand _78169_ (_27621_, _27620_, _27618_);
  nor _78170_ (_27622_, _12224_, _06133_);
  nor _78171_ (_27623_, _27622_, _05787_);
  nand _78172_ (_27624_, _27623_, _27621_);
  and _78173_ (_27625_, _12056_, _05787_);
  nor _78174_ (_27626_, _27625_, _12412_);
  nand _78175_ (_27627_, _27626_, _27624_);
  nor _78176_ (_27629_, _27493_, _11922_);
  nor _78177_ (_27630_, _27629_, _06209_);
  and _78178_ (_27631_, _27630_, _27627_);
  or _78179_ (_27632_, _27631_, _27487_);
  nand _78180_ (_27633_, _27632_, _27486_);
  and _78181_ (_27634_, _27510_, _12416_);
  nor _78182_ (_27635_, _27634_, _08788_);
  and _78183_ (_27636_, _27635_, _27633_);
  nor _78184_ (_27637_, _12224_, _08787_);
  or _78185_ (_27638_, _27637_, _27636_);
  nand _78186_ (_27640_, _27638_, _06111_);
  and _78187_ (_27641_, _12057_, _06110_);
  nor _78188_ (_27642_, _27641_, _10751_);
  nand _78189_ (_27643_, _27642_, _27640_);
  and _78190_ (_27644_, _12224_, _10751_);
  nor _78191_ (_27645_, _27644_, _12431_);
  nand _78192_ (_27646_, _27645_, _27643_);
  and _78193_ (_27647_, _12457_, _12434_);
  nor _78194_ (_27648_, _27647_, _12458_);
  nor _78195_ (_27649_, _27648_, _12432_);
  nor _78196_ (_27651_, _27649_, _06208_);
  nand _78197_ (_27652_, _27651_, _27646_);
  and _78198_ (_27653_, _12224_, _06208_);
  nor _78199_ (_27654_, _27653_, _06076_);
  nand _78200_ (_27655_, _27654_, _27652_);
  nand _78201_ (_27656_, _27655_, _12474_);
  and _78202_ (_27657_, _12224_, _11101_);
  and _78203_ (_27658_, _27510_, _12480_);
  or _78204_ (_27659_, _27658_, _27657_);
  and _78205_ (_27660_, _27659_, _12473_);
  nor _78206_ (_27662_, _27660_, _12478_);
  nand _78207_ (_27663_, _27662_, _27656_);
  nor _78208_ (_27664_, _27493_, _11919_);
  nor _78209_ (_27665_, _27664_, _11917_);
  nand _78210_ (_27666_, _27665_, _27663_);
  nor _78211_ (_27667_, _27495_, _11916_);
  nor _78212_ (_27668_, _27667_, _06297_);
  nand _78213_ (_27669_, _27668_, _27666_);
  and _78214_ (_27670_, _12057_, _06297_);
  nor _78215_ (_27671_, _27670_, _06402_);
  nand _78216_ (_27673_, _27671_, _27669_);
  and _78217_ (_27674_, _12224_, _06402_);
  nor _78218_ (_27675_, _27674_, _12492_);
  nand _78219_ (_27676_, _27675_, _27673_);
  nand _78220_ (_27677_, _27676_, _12497_);
  nor _78221_ (_27678_, _27510_, _12480_);
  nor _78222_ (_27679_, _12224_, _11101_);
  nor _78223_ (_27680_, _27679_, _12497_);
  not _78224_ (_27681_, _27680_);
  nor _78225_ (_27682_, _27681_, _27678_);
  nor _78226_ (_27684_, _27682_, _12505_);
  nand _78227_ (_27685_, _27684_, _27677_);
  nor _78228_ (_27686_, _27493_, _11914_);
  nor _78229_ (_27687_, _27686_, _10822_);
  nand _78230_ (_27688_, _27687_, _27685_);
  nor _78231_ (_27689_, _27495_, _10821_);
  nor _78232_ (_27690_, _27689_, _06306_);
  and _78233_ (_27691_, _27690_, _27688_);
  and _78234_ (_27692_, _12057_, _06306_);
  or _78235_ (_27693_, _27692_, _27691_);
  nand _78236_ (_27695_, _27693_, _07130_);
  nor _78237_ (_27696_, _12517_, _07124_);
  and _78238_ (_27697_, _27495_, _06411_);
  not _78239_ (_27698_, _27697_);
  and _78240_ (_27699_, _27698_, _27696_);
  nand _78241_ (_27700_, _27699_, _27695_);
  and _78242_ (_27701_, _12224_, \oc8051_golden_model_1.PSW [7]);
  and _78243_ (_27702_, _27510_, _10693_);
  or _78244_ (_27703_, _27702_, _27701_);
  and _78245_ (_27704_, _27703_, _12517_);
  nor _78246_ (_27706_, _27704_, _12522_);
  nand _78247_ (_27707_, _27706_, _27700_);
  nor _78248_ (_27708_, _27493_, _11912_);
  nor _78249_ (_27709_, _27708_, _10850_);
  and _78250_ (_27710_, _27709_, _27707_);
  nor _78251_ (_27711_, _27495_, _10849_);
  or _78252_ (_27712_, _27711_, _06303_);
  or _78253_ (_27713_, _27712_, _27710_);
  and _78254_ (_27714_, _12057_, _06303_);
  nor _78255_ (_27715_, _27714_, _06396_);
  and _78256_ (_27717_, _27715_, _27713_);
  and _78257_ (_27718_, _12224_, _06396_);
  or _78258_ (_27719_, _27718_, _27717_);
  nand _78259_ (_27720_, _27719_, _27484_);
  and _78260_ (_27721_, _12224_, _10693_);
  and _78261_ (_27722_, _27510_, \oc8051_golden_model_1.PSW [7]);
  or _78262_ (_27723_, _27722_, _27721_);
  and _78263_ (_27724_, _27723_, _12538_);
  nor _78264_ (_27725_, _27724_, _12547_);
  nand _78265_ (_27726_, _27725_, _27720_);
  nor _78266_ (_27728_, _27493_, _11907_);
  nor _78267_ (_27729_, _27728_, _10897_);
  nand _78268_ (_27730_, _27729_, _27726_);
  nor _78269_ (_27731_, _27495_, _10896_);
  nor _78270_ (_27732_, _27731_, _10925_);
  nand _78271_ (_27733_, _27732_, _27730_);
  and _78272_ (_27734_, _27516_, _10925_);
  nor _78273_ (_27735_, _27734_, _06417_);
  nand _78274_ (_27736_, _27735_, _27733_);
  and _78275_ (_27737_, _07049_, _06417_);
  nor _78276_ (_27739_, _27737_, _07142_);
  nand _78277_ (_27740_, _27739_, _27736_);
  nand _78278_ (_27741_, _27740_, _06421_);
  and _78279_ (_27742_, _27555_, _12682_);
  nor _78280_ (_27743_, _12056_, _12682_);
  or _78281_ (_27744_, _27743_, _06421_);
  nor _78282_ (_27745_, _27744_, _27742_);
  nor _78283_ (_27746_, _27745_, _12565_);
  nand _78284_ (_27747_, _27746_, _27741_);
  nor _78285_ (_27748_, _27493_, _11905_);
  nor _78286_ (_27750_, _27748_, _12691_);
  nand _78287_ (_27751_, _27750_, _27747_);
  nor _78288_ (_27752_, _12690_, _27495_);
  nor _78289_ (_27753_, _27752_, _10262_);
  nand _78290_ (_27754_, _27753_, _27751_);
  and _78291_ (_27755_, _27516_, _10262_);
  nor _78292_ (_27756_, _27755_, _06167_);
  nand _78293_ (_27757_, _27756_, _27754_);
  and _78294_ (_27758_, _07049_, _06167_);
  nor _78295_ (_27759_, _27758_, _05826_);
  nand _78296_ (_27761_, _27759_, _27757_);
  nand _78297_ (_27762_, _27761_, _06166_);
  nor _78298_ (_27763_, _27523_, _12682_);
  and _78299_ (_27764_, _12057_, _12682_);
  nor _78300_ (_27765_, _27764_, _27763_);
  and _78301_ (_27766_, _27765_, _06165_);
  nor _78302_ (_27767_, _27766_, _12712_);
  nand _78303_ (_27768_, _27767_, _27762_);
  nor _78304_ (_27769_, _27493_, _12711_);
  nor _78305_ (_27770_, _27769_, _06433_);
  nand _78306_ (_27772_, _27770_, _27768_);
  and _78307_ (_27773_, _12224_, _06433_);
  nor _78308_ (_27774_, _27773_, _25721_);
  nand _78309_ (_27775_, _27774_, _27772_);
  nor _78310_ (_27776_, _27493_, _12719_);
  nor _78311_ (_27777_, _27776_, _06310_);
  and _78312_ (_27778_, _27777_, _27775_);
  or _78313_ (_27779_, _27778_, _27483_);
  nor _78314_ (_27780_, _05823_, _05748_);
  nand _78315_ (_27781_, _27780_, _27779_);
  and _78316_ (_27783_, _27765_, _05748_);
  nor _78317_ (_27784_, _27783_, _12737_);
  nand _78318_ (_27785_, _27784_, _27781_);
  nor _78319_ (_27786_, _27493_, _12735_);
  nor _78320_ (_27787_, _27786_, _06440_);
  nand _78321_ (_27788_, _27787_, _27785_);
  and _78322_ (_27789_, _12224_, _06440_);
  nor _78323_ (_27790_, _27789_, _26415_);
  nand _78324_ (_27791_, _27790_, _27788_);
  nor _78325_ (_27792_, _27493_, _12744_);
  nor _78326_ (_27794_, _27792_, _06305_);
  and _78327_ (_27795_, _27794_, _27791_);
  or _78328_ (_27796_, _27795_, _27482_);
  nor _78329_ (_27797_, _12754_, _05821_);
  and _78330_ (_27798_, _27797_, _27796_);
  and _78331_ (_27799_, _27493_, _12754_);
  or _78332_ (_27800_, _27799_, _27798_);
  or _78333_ (_27801_, _27800_, _01321_);
  or _78334_ (_27802_, _01317_, \oc8051_golden_model_1.PC [8]);
  and _78335_ (_27803_, _27802_, _43100_);
  and _78336_ (_43696_, _27803_, _27801_);
  nor _78337_ (_27805_, _06912_, _12747_);
  nor _78338_ (_27806_, _06912_, _12723_);
  nor _78339_ (_27807_, _27491_, \oc8051_golden_model_1.PC [9]);
  nor _78340_ (_27808_, _27807_, _11896_);
  nor _78341_ (_27809_, _27808_, _11905_);
  nor _78342_ (_27810_, _27808_, _11907_);
  and _78343_ (_27811_, _11996_, _06303_);
  nor _78344_ (_27812_, _27808_, _11912_);
  and _78345_ (_27813_, _11996_, _06306_);
  nor _78346_ (_27815_, _27808_, _11914_);
  and _78347_ (_27816_, _11996_, _06297_);
  nor _78348_ (_27817_, _27808_, _11919_);
  nor _78349_ (_27818_, _12172_, _08787_);
  and _78350_ (_27819_, _12172_, _06209_);
  and _78351_ (_27820_, _12172_, _06254_);
  nor _78352_ (_27821_, _06254_, _24882_);
  and _78353_ (_27822_, _12172_, _06255_);
  or _78354_ (_27823_, _12139_, _11996_);
  nor _78355_ (_27824_, _12061_, _12058_);
  and _78356_ (_27826_, _27824_, _12000_);
  nor _78357_ (_27827_, _27824_, _12000_);
  nor _78358_ (_27828_, _27827_, _27826_);
  not _78359_ (_27829_, _27828_);
  or _78360_ (_27830_, _27829_, _12141_);
  and _78361_ (_27831_, _27830_, _27823_);
  or _78362_ (_27832_, _27831_, _06161_);
  nor _78363_ (_27833_, _12228_, _12225_);
  and _78364_ (_27834_, _27833_, _12175_);
  nor _78365_ (_27835_, _27833_, _12175_);
  nor _78366_ (_27837_, _27835_, _27834_);
  or _78367_ (_27838_, _27837_, _12258_);
  not _78368_ (_27839_, _12172_);
  or _78369_ (_27840_, _12256_, _27839_);
  and _78370_ (_27841_, _27840_, _08445_);
  nand _78371_ (_27842_, _27841_, _27838_);
  and _78372_ (_27843_, _12265_, _12263_);
  or _78373_ (_27844_, _27843_, _27808_);
  and _78374_ (_27845_, _27839_, _07056_);
  nor _78375_ (_27846_, _27845_, _06653_);
  nor _78376_ (_27848_, _07056_, \oc8051_golden_model_1.PC [9]);
  nand _78377_ (_27849_, _27848_, _12265_);
  nand _78378_ (_27850_, _27849_, _27846_);
  nand _78379_ (_27851_, _27850_, _24799_);
  and _78380_ (_27852_, _27851_, _27844_);
  and _78381_ (_27853_, _27808_, _06653_);
  nor _78382_ (_27854_, _27853_, _08445_);
  not _78383_ (_27855_, _27854_);
  nor _78384_ (_27856_, _27855_, _27852_);
  nor _78385_ (_27857_, _27856_, _07064_);
  and _78386_ (_27859_, _27857_, _27842_);
  and _78387_ (_27860_, _27808_, _07064_);
  or _78388_ (_27861_, _27860_, _06160_);
  or _78389_ (_27862_, _27861_, _27859_);
  nand _78390_ (_27863_, _27862_, _27832_);
  nand _78391_ (_27864_, _27863_, _12134_);
  nor _78392_ (_27865_, _27808_, _12134_);
  nor _78393_ (_27866_, _27865_, _06156_);
  nand _78394_ (_27867_, _27866_, _27864_);
  and _78395_ (_27868_, _12172_, _06156_);
  nor _78396_ (_27870_, _27868_, _07485_);
  nand _78397_ (_27871_, _27870_, _27867_);
  nand _78398_ (_27872_, _27871_, _07075_);
  and _78399_ (_27873_, _12172_, _06217_);
  nor _78400_ (_27874_, _27873_, _12293_);
  nand _78401_ (_27875_, _27874_, _27872_);
  nor _78402_ (_27876_, _27808_, _12292_);
  nor _78403_ (_27877_, _27876_, _06220_);
  nand _78404_ (_27878_, _27877_, _27875_);
  and _78405_ (_27879_, _12172_, _06220_);
  nor _78406_ (_27881_, _27879_, _12302_);
  nand _78407_ (_27882_, _27881_, _27878_);
  nor _78408_ (_27883_, _27808_, _12300_);
  nor _78409_ (_27884_, _27883_, _06152_);
  nand _78410_ (_27885_, _27884_, _27882_);
  and _78411_ (_27886_, _12172_, _06152_);
  nor _78412_ (_27887_, _27886_, _12304_);
  nand _78413_ (_27888_, _27887_, _27885_);
  nand _78414_ (_27889_, _27888_, _07191_);
  and _78415_ (_27890_, _12172_, _06151_);
  nor _78416_ (_27892_, _27890_, _12126_);
  nand _78417_ (_27893_, _27892_, _27889_);
  and _78418_ (_27894_, _12120_, _11996_);
  nor _78419_ (_27895_, _27828_, _12120_);
  or _78420_ (_27896_, _27895_, _27894_);
  nor _78421_ (_27897_, _27896_, _12125_);
  nor _78422_ (_27898_, _27897_, _06687_);
  and _78423_ (_27899_, _27898_, _27893_);
  and _78424_ (_27900_, _27829_, _11956_);
  and _78425_ (_27901_, _11996_, _11958_);
  or _78426_ (_27903_, _27901_, _27900_);
  and _78427_ (_27904_, _27903_, _06687_);
  or _78428_ (_27905_, _27904_, _06236_);
  or _78429_ (_27906_, _27905_, _27899_);
  nor _78430_ (_27907_, _27828_, _12329_);
  not _78431_ (_27908_, _27907_);
  and _78432_ (_27909_, _12329_, _11996_);
  nor _78433_ (_27910_, _27909_, _06643_);
  and _78434_ (_27911_, _27910_, _27908_);
  nor _78435_ (_27912_, _27911_, _06295_);
  nand _78436_ (_27914_, _27912_, _27906_);
  nand _78437_ (_27915_, _12346_, _11996_);
  or _78438_ (_27916_, _27828_, _12346_);
  and _78439_ (_27917_, _27916_, _27915_);
  or _78440_ (_27918_, _27917_, _12317_);
  and _78441_ (_27919_, _27918_, _27914_);
  or _78442_ (_27920_, _27919_, _11924_);
  nand _78443_ (_27921_, _27808_, _11924_);
  and _78444_ (_27922_, _27921_, _27920_);
  nand _78445_ (_27923_, _27922_, _06146_);
  and _78446_ (_27925_, _27839_, _06145_);
  nor _78447_ (_27926_, _27925_, _07388_);
  and _78448_ (_27927_, _27926_, _25151_);
  nand _78449_ (_27928_, _27927_, _27923_);
  nor _78450_ (_27929_, _25151_, _27839_);
  nor _78451_ (_27930_, _27929_, _12373_);
  nand _78452_ (_27931_, _27930_, _27928_);
  nor _78453_ (_27932_, _27808_, _12369_);
  nor _78454_ (_27933_, _27932_, _06255_);
  and _78455_ (_27934_, _27933_, _27931_);
  or _78456_ (_27936_, _27934_, _27822_);
  and _78457_ (_27937_, _27936_, _27821_);
  or _78458_ (_27938_, _27937_, _27820_);
  nand _78459_ (_27939_, _27938_, _12381_);
  and _78460_ (_27940_, _27808_, _12387_);
  nor _78461_ (_27941_, _27940_, _12386_);
  nand _78462_ (_27942_, _27941_, _27939_);
  nor _78463_ (_27943_, _12172_, _12385_);
  nor _78464_ (_27944_, _27943_, _05870_);
  nand _78465_ (_27945_, _27944_, _27942_);
  and _78466_ (_27947_, _27808_, _05870_);
  nor _78467_ (_27948_, _27947_, _06139_);
  nand _78468_ (_27949_, _27948_, _27945_);
  and _78469_ (_27950_, _27839_, _06139_);
  nor _78470_ (_27951_, _27950_, _27615_);
  nand _78471_ (_27952_, _27951_, _27949_);
  and _78472_ (_27953_, _11996_, _06293_);
  nor _78473_ (_27954_, _27953_, _13620_);
  nand _78474_ (_27955_, _27954_, _27952_);
  nor _78475_ (_27956_, _12172_, _06133_);
  nor _78476_ (_27958_, _27956_, _05787_);
  nand _78477_ (_27959_, _27958_, _27955_);
  and _78478_ (_27960_, _11996_, _05787_);
  nor _78479_ (_27961_, _27960_, _12412_);
  nand _78480_ (_27962_, _27961_, _27959_);
  nor _78481_ (_27963_, _27808_, _11922_);
  nor _78482_ (_27964_, _27963_, _06209_);
  and _78483_ (_27965_, _27964_, _27962_);
  or _78484_ (_27966_, _27965_, _27819_);
  nand _78485_ (_27967_, _27966_, _27486_);
  nor _78486_ (_27968_, _27837_, _12417_);
  nor _78487_ (_27969_, _27968_, _08788_);
  and _78488_ (_27970_, _27969_, _27967_);
  or _78489_ (_27971_, _27970_, _27818_);
  nand _78490_ (_27972_, _27971_, _06111_);
  and _78491_ (_27973_, _11997_, _06110_);
  nor _78492_ (_27974_, _27973_, _10751_);
  nand _78493_ (_27975_, _27974_, _27972_);
  and _78494_ (_27976_, _12172_, _10751_);
  nor _78495_ (_27977_, _27976_, _12431_);
  nand _78496_ (_27980_, _27977_, _27975_);
  nor _78497_ (_27981_, _12458_, \oc8051_golden_model_1.DPH [1]);
  nor _78498_ (_27982_, _27981_, _12459_);
  nor _78499_ (_27983_, _27982_, _12432_);
  nor _78500_ (_27984_, _27983_, _06208_);
  nand _78501_ (_27985_, _27984_, _27980_);
  and _78502_ (_27986_, _12172_, _06208_);
  nor _78503_ (_27987_, _27986_, _06076_);
  nand _78504_ (_27988_, _27987_, _27985_);
  nand _78505_ (_27989_, _27988_, _12474_);
  and _78506_ (_27991_, _12172_, _11101_);
  nor _78507_ (_27992_, _27837_, _11101_);
  or _78508_ (_27993_, _27992_, _27991_);
  and _78509_ (_27994_, _27993_, _12473_);
  nor _78510_ (_27995_, _27994_, _12478_);
  and _78511_ (_27996_, _27995_, _27989_);
  or _78512_ (_27997_, _27996_, _27817_);
  nand _78513_ (_27998_, _27997_, _11916_);
  nor _78514_ (_27999_, _12172_, _11916_);
  nor _78515_ (_28000_, _27999_, _06297_);
  and _78516_ (_28002_, _28000_, _27998_);
  or _78517_ (_28003_, _28002_, _27816_);
  nand _78518_ (_28004_, _28003_, _07125_);
  and _78519_ (_28005_, _12172_, _06402_);
  nor _78520_ (_28006_, _28005_, _12492_);
  nand _78521_ (_28007_, _28006_, _28004_);
  nand _78522_ (_28008_, _28007_, _12497_);
  and _78523_ (_28009_, _12172_, _12480_);
  nor _78524_ (_28010_, _27837_, _12480_);
  or _78525_ (_28011_, _28010_, _28009_);
  and _78526_ (_28013_, _28011_, _12496_);
  nor _78527_ (_28014_, _28013_, _12505_);
  and _78528_ (_28015_, _28014_, _28008_);
  or _78529_ (_28016_, _28015_, _27815_);
  nand _78530_ (_28017_, _28016_, _10821_);
  nor _78531_ (_28018_, _12172_, _10821_);
  nor _78532_ (_28019_, _28018_, _06306_);
  and _78533_ (_28020_, _28019_, _28017_);
  or _78534_ (_28021_, _28020_, _27813_);
  nand _78535_ (_28022_, _28021_, _07130_);
  and _78536_ (_28024_, _12172_, _06411_);
  nor _78537_ (_28025_, _28024_, _07124_);
  nand _78538_ (_28026_, _28025_, _28022_);
  nand _78539_ (_28027_, _28026_, _12518_);
  and _78540_ (_28028_, _12172_, \oc8051_golden_model_1.PSW [7]);
  nor _78541_ (_28029_, _27837_, \oc8051_golden_model_1.PSW [7]);
  or _78542_ (_28030_, _28029_, _28028_);
  and _78543_ (_28031_, _28030_, _12517_);
  nor _78544_ (_28032_, _28031_, _12522_);
  and _78545_ (_28033_, _28032_, _28027_);
  or _78546_ (_28035_, _28033_, _27812_);
  nand _78547_ (_28036_, _28035_, _10849_);
  nor _78548_ (_28037_, _12172_, _10849_);
  nor _78549_ (_28038_, _28037_, _06303_);
  and _78550_ (_28039_, _28038_, _28036_);
  or _78551_ (_28040_, _28039_, _27811_);
  nand _78552_ (_28041_, _28040_, _08824_);
  and _78553_ (_28042_, _12172_, _06396_);
  nor _78554_ (_28043_, _28042_, _05842_);
  nand _78555_ (_28044_, _28043_, _28041_);
  nand _78556_ (_28046_, _28044_, _12539_);
  nand _78557_ (_28047_, _27837_, \oc8051_golden_model_1.PSW [7]);
  or _78558_ (_28048_, _12172_, \oc8051_golden_model_1.PSW [7]);
  and _78559_ (_28049_, _28048_, _12538_);
  and _78560_ (_28050_, _28049_, _28047_);
  nor _78561_ (_28051_, _28050_, _12547_);
  and _78562_ (_28052_, _28051_, _28046_);
  or _78563_ (_28053_, _28052_, _27810_);
  nand _78564_ (_28054_, _28053_, _10896_);
  nor _78565_ (_28055_, _12172_, _10896_);
  nor _78566_ (_28057_, _28055_, _10925_);
  nand _78567_ (_28058_, _28057_, _28054_);
  and _78568_ (_28059_, _27808_, _10925_);
  nor _78569_ (_28060_, _28059_, _06417_);
  nand _78570_ (_28061_, _28060_, _28058_);
  nor _78571_ (_28062_, _06301_, _07142_);
  not _78572_ (_28063_, _28062_);
  and _78573_ (_28064_, _07252_, _06417_);
  nor _78574_ (_28065_, _28064_, _28063_);
  nand _78575_ (_28066_, _28065_, _28061_);
  nor _78576_ (_28068_, _11996_, _12682_);
  and _78577_ (_28069_, _27828_, _12682_);
  or _78578_ (_28070_, _28069_, _06421_);
  nor _78579_ (_28071_, _28070_, _28068_);
  nor _78580_ (_28072_, _28071_, _12565_);
  and _78581_ (_28073_, _28072_, _28066_);
  or _78582_ (_28074_, _28073_, _27809_);
  nand _78583_ (_28075_, _28074_, _12690_);
  nor _78584_ (_28076_, _12690_, _12172_);
  nor _78585_ (_28077_, _28076_, _10262_);
  nand _78586_ (_28079_, _28077_, _28075_);
  and _78587_ (_28080_, _27808_, _10262_);
  nor _78588_ (_28081_, _28080_, _06167_);
  nand _78589_ (_28082_, _28081_, _28079_);
  nor _78590_ (_28083_, _06165_, _05826_);
  not _78591_ (_28084_, _28083_);
  and _78592_ (_28085_, _07252_, _06167_);
  nor _78593_ (_28086_, _28085_, _28084_);
  nand _78594_ (_28087_, _28086_, _28082_);
  nor _78595_ (_28088_, _27829_, _12682_);
  and _78596_ (_28090_, _11997_, _12682_);
  nor _78597_ (_28091_, _28090_, _28088_);
  and _78598_ (_28092_, _28091_, _06165_);
  nor _78599_ (_28093_, _28092_, _12712_);
  nand _78600_ (_28094_, _28093_, _28087_);
  nor _78601_ (_28095_, _27808_, _12711_);
  nor _78602_ (_28096_, _28095_, _06433_);
  nand _78603_ (_28097_, _28096_, _28094_);
  and _78604_ (_28098_, _12172_, _06433_);
  nor _78605_ (_28099_, _28098_, _25721_);
  nand _78606_ (_28101_, _28099_, _28097_);
  nor _78607_ (_28102_, _27808_, _12719_);
  nor _78608_ (_28103_, _28102_, _06310_);
  and _78609_ (_28104_, _28103_, _28101_);
  or _78610_ (_28105_, _28104_, _27806_);
  nand _78611_ (_28106_, _28105_, _27780_);
  and _78612_ (_28107_, _28091_, _05748_);
  nor _78613_ (_28108_, _28107_, _12737_);
  nand _78614_ (_28109_, _28108_, _28106_);
  nor _78615_ (_28110_, _27808_, _12735_);
  nor _78616_ (_28112_, _28110_, _06440_);
  nand _78617_ (_28113_, _28112_, _28109_);
  and _78618_ (_28114_, _12172_, _06440_);
  nor _78619_ (_28115_, _28114_, _26415_);
  nand _78620_ (_28116_, _28115_, _28113_);
  nor _78621_ (_28117_, _27808_, _12744_);
  nor _78622_ (_28118_, _28117_, _06305_);
  and _78623_ (_28119_, _28118_, _28116_);
  or _78624_ (_28120_, _28119_, _27805_);
  and _78625_ (_28121_, _28120_, _27797_);
  and _78626_ (_28123_, _27808_, _12754_);
  or _78627_ (_28124_, _28123_, _28121_);
  or _78628_ (_28125_, _28124_, _01321_);
  or _78629_ (_28126_, _01317_, \oc8051_golden_model_1.PC [9]);
  and _78630_ (_28127_, _28126_, _43100_);
  and _78631_ (_43697_, _28127_, _28125_);
  nor _78632_ (_28128_, _11896_, \oc8051_golden_model_1.PC [10]);
  nor _78633_ (_28129_, _28128_, _11897_);
  not _78634_ (_28130_, _28129_);
  nand _78635_ (_28131_, _28130_, _10925_);
  nand _78636_ (_28133_, _11989_, _06303_);
  nand _78637_ (_28134_, _11989_, _06306_);
  nand _78638_ (_28135_, _11989_, _06297_);
  nor _78639_ (_28136_, _12473_, _06076_);
  not _78640_ (_28137_, _06286_);
  or _78641_ (_28138_, _28129_, _12292_);
  and _78642_ (_28139_, _12159_, _07056_);
  and _78643_ (_28140_, _07057_, \oc8051_golden_model_1.PC [10]);
  and _78644_ (_28141_, _28140_, _12265_);
  or _78645_ (_28142_, _28141_, _28139_);
  and _78646_ (_28144_, _28142_, _12264_);
  or _78647_ (_28145_, _28144_, _06581_);
  and _78648_ (_28146_, _28145_, _12263_);
  nor _78649_ (_28147_, _28130_, _12267_);
  or _78650_ (_28148_, _28147_, _08445_);
  or _78651_ (_28149_, _28148_, _28146_);
  and _78652_ (_28150_, _12258_, _12159_);
  nor _78653_ (_28151_, _12232_, _12229_);
  not _78654_ (_28152_, _28151_);
  and _78655_ (_28153_, _28152_, _12168_);
  nor _78656_ (_28155_, _28152_, _12168_);
  nor _78657_ (_28156_, _28155_, _28153_);
  and _78658_ (_28157_, _28156_, _12256_);
  or _78659_ (_28158_, _28157_, _28150_);
  or _78660_ (_28159_, _28158_, _08443_);
  and _78661_ (_28160_, _28159_, _28149_);
  or _78662_ (_28161_, _28160_, _07064_);
  nand _78663_ (_28162_, _28130_, _07064_);
  and _78664_ (_28163_, _28162_, _06161_);
  and _78665_ (_28164_, _28163_, _28161_);
  not _78666_ (_28166_, _11992_);
  nor _78667_ (_28167_, _12065_, _12062_);
  nor _78668_ (_28168_, _28167_, _28166_);
  and _78669_ (_28169_, _28167_, _28166_);
  nor _78670_ (_28170_, _28169_, _28168_);
  or _78671_ (_28171_, _28170_, _12141_);
  or _78672_ (_28172_, _12139_, _11988_);
  and _78673_ (_28173_, _28172_, _06160_);
  and _78674_ (_28174_, _28173_, _28171_);
  or _78675_ (_28175_, _28174_, _24821_);
  or _78676_ (_28177_, _28175_, _28164_);
  or _78677_ (_28178_, _28129_, _12134_);
  and _78678_ (_28179_, _28178_, _06157_);
  and _78679_ (_28180_, _28179_, _28177_);
  or _78680_ (_28181_, _28180_, _07485_);
  and _78681_ (_28182_, _28181_, _07075_);
  not _78682_ (_28183_, _12159_);
  or _78683_ (_28184_, _28183_, _06221_);
  nand _78684_ (_28185_, _28184_, _12292_);
  or _78685_ (_28186_, _28185_, _28182_);
  and _78686_ (_28188_, _28186_, _28138_);
  or _78687_ (_28189_, _28188_, _06220_);
  nand _78688_ (_28190_, _28183_, _06220_);
  and _78689_ (_28191_, _28190_, _12300_);
  and _78690_ (_28192_, _28191_, _28189_);
  nor _78691_ (_28193_, _28130_, _12300_);
  or _78692_ (_28194_, _28193_, _28192_);
  and _78693_ (_28195_, _28194_, _06153_);
  and _78694_ (_28196_, _12159_, _06152_);
  or _78695_ (_28197_, _28196_, _12304_);
  or _78696_ (_28199_, _28197_, _28195_);
  and _78697_ (_28200_, _28199_, _07191_);
  nand _78698_ (_28201_, _12159_, _06151_);
  nand _78699_ (_28202_, _28201_, _12125_);
  or _78700_ (_28203_, _28202_, _28200_);
  or _78701_ (_28204_, _28170_, _12120_);
  nand _78702_ (_28205_, _12120_, _11989_);
  and _78703_ (_28206_, _28205_, _28204_);
  or _78704_ (_28207_, _28206_, _12125_);
  and _78705_ (_28208_, _28207_, _28203_);
  or _78706_ (_28210_, _28208_, _28137_);
  and _78707_ (_28211_, _11988_, _11958_);
  and _78708_ (_28212_, _28170_, _11956_);
  or _78709_ (_28213_, _28212_, _28211_);
  or _78710_ (_28214_, _28213_, _12089_);
  and _78711_ (_28215_, _28214_, _28210_);
  or _78712_ (_28216_, _28215_, _06236_);
  and _78713_ (_28217_, _12329_, _11988_);
  and _78714_ (_28218_, _28170_, _25123_);
  or _78715_ (_28219_, _28218_, _06643_);
  or _78716_ (_28221_, _28219_, _28217_);
  and _78717_ (_28222_, _28221_, _12317_);
  and _78718_ (_28223_, _28222_, _28216_);
  or _78719_ (_28224_, _28170_, _12346_);
  nand _78720_ (_28225_, _12346_, _11989_);
  and _78721_ (_28226_, _28225_, _06295_);
  and _78722_ (_28227_, _28226_, _28224_);
  or _78723_ (_28228_, _28227_, _11924_);
  or _78724_ (_28229_, _28228_, _28223_);
  nand _78725_ (_28230_, _28130_, _11924_);
  and _78726_ (_28232_, _25151_, _06146_);
  and _78727_ (_28233_, _28232_, _28230_);
  and _78728_ (_28234_, _28233_, _28229_);
  nor _78729_ (_28235_, _28232_, _28183_);
  nand _78730_ (_28236_, _12369_, _05760_);
  or _78731_ (_28237_, _28236_, _28235_);
  or _78732_ (_28238_, _28237_, _28234_);
  or _78733_ (_28239_, _28129_, _12369_);
  and _78734_ (_28240_, _28239_, _13844_);
  and _78735_ (_28241_, _28240_, _28238_);
  or _78736_ (_28243_, _28241_, _24882_);
  and _78737_ (_28244_, _28243_, _13843_);
  or _78738_ (_28245_, _28183_, _06256_);
  nand _78739_ (_28246_, _28245_, _12381_);
  or _78740_ (_28247_, _28246_, _28244_);
  or _78741_ (_28248_, _28129_, _12381_);
  and _78742_ (_28249_, _28248_, _12385_);
  and _78743_ (_28250_, _28249_, _28247_);
  nor _78744_ (_28251_, _28183_, _12385_);
  or _78745_ (_28252_, _28251_, _05870_);
  or _78746_ (_28254_, _28252_, _28250_);
  or _78747_ (_28255_, _28129_, _05805_);
  and _78748_ (_28256_, _28255_, _06140_);
  and _78749_ (_28257_, _28256_, _28254_);
  nand _78750_ (_28258_, _12159_, _06139_);
  nand _78751_ (_28259_, _28258_, _27614_);
  or _78752_ (_28260_, _28259_, _28257_);
  nand _78753_ (_28261_, _11989_, _06293_);
  and _78754_ (_28262_, _28261_, _06133_);
  and _78755_ (_28263_, _28262_, _28260_);
  nor _78756_ (_28265_, _28183_, _06133_);
  or _78757_ (_28266_, _28265_, _05787_);
  or _78758_ (_28267_, _28266_, _28263_);
  nand _78759_ (_28268_, _11989_, _05787_);
  and _78760_ (_28269_, _28268_, _11922_);
  and _78761_ (_28270_, _28269_, _28267_);
  nor _78762_ (_28271_, _28130_, _11922_);
  or _78763_ (_28272_, _28271_, _28270_);
  and _78764_ (_28273_, _28272_, _06762_);
  nand _78765_ (_28274_, _12159_, _06209_);
  nand _78766_ (_28275_, _28274_, _27486_);
  or _78767_ (_28276_, _28275_, _28273_);
  or _78768_ (_28277_, _28156_, _12417_);
  and _78769_ (_28278_, _28277_, _08787_);
  and _78770_ (_28279_, _28278_, _28276_);
  nor _78771_ (_28280_, _28183_, _08787_);
  or _78772_ (_28281_, _28280_, _06110_);
  or _78773_ (_28282_, _28281_, _28279_);
  nand _78774_ (_28283_, _11989_, _06110_);
  and _78775_ (_28284_, _28283_, _10752_);
  and _78776_ (_28287_, _28284_, _28282_);
  and _78777_ (_28288_, _12159_, _10751_);
  or _78778_ (_28289_, _28288_, _12431_);
  or _78779_ (_28290_, _28289_, _28287_);
  nor _78780_ (_28291_, _12459_, \oc8051_golden_model_1.DPH [2]);
  nor _78781_ (_28292_, _28291_, _12460_);
  or _78782_ (_28293_, _28292_, _12432_);
  and _78783_ (_28294_, _28293_, _06768_);
  and _78784_ (_28295_, _28294_, _28290_);
  and _78785_ (_28296_, _12159_, _06208_);
  or _78786_ (_28298_, _28296_, _28295_);
  and _78787_ (_28299_, _28298_, _28136_);
  or _78788_ (_28300_, _28156_, _11101_);
  or _78789_ (_28301_, _12159_, _12480_);
  and _78790_ (_28302_, _28301_, _12473_);
  and _78791_ (_28303_, _28302_, _28300_);
  or _78792_ (_28304_, _28303_, _12478_);
  or _78793_ (_28305_, _28304_, _28299_);
  or _78794_ (_28306_, _28129_, _11919_);
  and _78795_ (_28307_, _28306_, _11916_);
  and _78796_ (_28309_, _28307_, _28305_);
  nor _78797_ (_28310_, _28183_, _11916_);
  or _78798_ (_28311_, _28310_, _06297_);
  or _78799_ (_28312_, _28311_, _28309_);
  and _78800_ (_28313_, _28312_, _28135_);
  or _78801_ (_28314_, _28313_, _06402_);
  nand _78802_ (_28315_, _28183_, _06402_);
  nor _78803_ (_28316_, _12496_, _12492_);
  and _78804_ (_28317_, _28316_, _28315_);
  and _78805_ (_28318_, _28317_, _28314_);
  or _78806_ (_28320_, _28156_, _12480_);
  or _78807_ (_28321_, _12159_, _11101_);
  and _78808_ (_28322_, _28321_, _12496_);
  and _78809_ (_28323_, _28322_, _28320_);
  or _78810_ (_28324_, _28323_, _12505_);
  or _78811_ (_28325_, _28324_, _28318_);
  or _78812_ (_28326_, _28129_, _11914_);
  and _78813_ (_28327_, _28326_, _10821_);
  and _78814_ (_28328_, _28327_, _28325_);
  nor _78815_ (_28329_, _28183_, _10821_);
  or _78816_ (_28331_, _28329_, _06306_);
  or _78817_ (_28332_, _28331_, _28328_);
  and _78818_ (_28333_, _28332_, _28134_);
  or _78819_ (_28334_, _28333_, _06411_);
  nand _78820_ (_28335_, _28183_, _06411_);
  and _78821_ (_28336_, _28335_, _27696_);
  and _78822_ (_28337_, _28336_, _28334_);
  or _78823_ (_28338_, _28156_, \oc8051_golden_model_1.PSW [7]);
  or _78824_ (_28339_, _12159_, _10693_);
  and _78825_ (_28340_, _28339_, _12517_);
  and _78826_ (_28342_, _28340_, _28338_);
  or _78827_ (_28343_, _28342_, _12522_);
  or _78828_ (_28344_, _28343_, _28337_);
  or _78829_ (_28345_, _28129_, _11912_);
  and _78830_ (_28346_, _28345_, _10849_);
  and _78831_ (_28347_, _28346_, _28344_);
  nor _78832_ (_28348_, _28183_, _10849_);
  or _78833_ (_28349_, _28348_, _06303_);
  or _78834_ (_28350_, _28349_, _28347_);
  and _78835_ (_28351_, _28350_, _28133_);
  or _78836_ (_28353_, _28351_, _06396_);
  nand _78837_ (_28354_, _28183_, _06396_);
  and _78838_ (_28355_, _28354_, _27484_);
  and _78839_ (_28356_, _28355_, _28353_);
  or _78840_ (_28357_, _28156_, _10693_);
  or _78841_ (_28358_, _12159_, \oc8051_golden_model_1.PSW [7]);
  and _78842_ (_28359_, _28358_, _12538_);
  and _78843_ (_28360_, _28359_, _28357_);
  or _78844_ (_28361_, _28360_, _12547_);
  or _78845_ (_28362_, _28361_, _28356_);
  or _78846_ (_28364_, _28129_, _11907_);
  and _78847_ (_28365_, _28364_, _10896_);
  and _78848_ (_28366_, _28365_, _28362_);
  nor _78849_ (_28367_, _28183_, _10896_);
  or _78850_ (_28368_, _28367_, _10925_);
  or _78851_ (_28369_, _28368_, _28366_);
  and _78852_ (_28370_, _28369_, _28131_);
  or _78853_ (_28371_, _28370_, _06417_);
  or _78854_ (_28372_, _07708_, _12558_);
  and _78855_ (_28373_, _28372_, _28062_);
  and _78856_ (_28375_, _28373_, _28371_);
  or _78857_ (_28376_, _28170_, _25333_);
  or _78858_ (_28377_, _11988_, _12682_);
  and _78859_ (_28378_, _28377_, _06301_);
  and _78860_ (_28379_, _28378_, _28376_);
  or _78861_ (_28380_, _28379_, _12565_);
  or _78862_ (_28381_, _28380_, _28375_);
  or _78863_ (_28382_, _28129_, _11905_);
  and _78864_ (_28383_, _28382_, _12690_);
  and _78865_ (_28384_, _28383_, _28381_);
  nor _78866_ (_28386_, _12690_, _28183_);
  or _78867_ (_28387_, _28386_, _10262_);
  or _78868_ (_28388_, _28387_, _28384_);
  nand _78869_ (_28389_, _28130_, _10262_);
  and _78870_ (_28390_, _28389_, _28388_);
  or _78871_ (_28391_, _28390_, _06167_);
  or _78872_ (_28392_, _07708_, _06168_);
  and _78873_ (_28393_, _28392_, _28083_);
  and _78874_ (_28394_, _28393_, _28391_);
  nor _78875_ (_28395_, _28170_, _12682_);
  and _78876_ (_28397_, _11989_, _12682_);
  nor _78877_ (_28398_, _28397_, _28395_);
  and _78878_ (_28399_, _28398_, _06165_);
  or _78879_ (_28400_, _28399_, _12712_);
  or _78880_ (_28401_, _28400_, _28394_);
  or _78881_ (_28402_, _28129_, _12711_);
  and _78882_ (_28403_, _28402_, _28401_);
  nor _78883_ (_28404_, _28403_, _06433_);
  and _78884_ (_28405_, _28183_, _06433_);
  nor _78885_ (_28406_, _28405_, _25721_);
  not _78886_ (_28408_, _28406_);
  nor _78887_ (_28409_, _28408_, _28404_);
  nor _78888_ (_28410_, _28130_, _12719_);
  nor _78889_ (_28411_, _28410_, _06310_);
  not _78890_ (_28412_, _28411_);
  nor _78891_ (_28413_, _28412_, _28409_);
  not _78892_ (_28414_, _27780_);
  and _78893_ (_28415_, _06625_, _06310_);
  nor _78894_ (_28416_, _28415_, _28414_);
  not _78895_ (_28417_, _28416_);
  nor _78896_ (_28419_, _28417_, _28413_);
  and _78897_ (_28420_, _28398_, _05748_);
  nor _78898_ (_28421_, _28420_, _12737_);
  not _78899_ (_28422_, _28421_);
  nor _78900_ (_28423_, _28422_, _28419_);
  nor _78901_ (_28424_, _28129_, _12735_);
  or _78902_ (_28425_, _28424_, _28423_);
  nand _78903_ (_28426_, _28425_, _06444_);
  and _78904_ (_28427_, _28183_, _06440_);
  nor _78905_ (_28428_, _28427_, _26415_);
  and _78906_ (_28430_, _28428_, _28426_);
  nor _78907_ (_28431_, _28130_, _12744_);
  or _78908_ (_28432_, _28431_, _06305_);
  or _78909_ (_28433_, _28432_, _28430_);
  not _78910_ (_28434_, _27797_);
  and _78911_ (_28435_, _06625_, _06305_);
  nor _78912_ (_28436_, _28435_, _28434_);
  and _78913_ (_28437_, _28436_, _28433_);
  and _78914_ (_28438_, _28129_, _12754_);
  or _78915_ (_28439_, _28438_, _28437_);
  or _78916_ (_28441_, _28439_, _01321_);
  or _78917_ (_28442_, _01317_, \oc8051_golden_model_1.PC [10]);
  and _78918_ (_28443_, _28442_, _43100_);
  and _78919_ (_43698_, _28443_, _28441_);
  nor _78920_ (_28444_, _11897_, \oc8051_golden_model_1.PC [11]);
  nor _78921_ (_28445_, _28444_, _11898_);
  or _78922_ (_28446_, _28445_, _11905_);
  nor _78923_ (_28447_, _28153_, _12160_);
  nor _78924_ (_28448_, _28447_, _12166_);
  and _78925_ (_28449_, _28447_, _12166_);
  or _78926_ (_28451_, _28449_, _28448_);
  or _78927_ (_28452_, _28451_, _10693_);
  or _78928_ (_28453_, _12163_, \oc8051_golden_model_1.PSW [7]);
  and _78929_ (_28454_, _28453_, _12538_);
  and _78930_ (_28455_, _28454_, _28452_);
  or _78931_ (_28456_, _28451_, \oc8051_golden_model_1.PSW [7]);
  or _78932_ (_28457_, _12163_, _10693_);
  and _78933_ (_28458_, _28457_, _12517_);
  and _78934_ (_28459_, _28458_, _28456_);
  or _78935_ (_28460_, _28445_, _11914_);
  or _78936_ (_28462_, _28445_, _11919_);
  or _78937_ (_28463_, _12163_, _08787_);
  and _78938_ (_28464_, _11981_, _05787_);
  or _78939_ (_28465_, _11981_, _11956_);
  nor _78940_ (_28466_, _28168_, _11990_);
  and _78941_ (_28467_, _28466_, _11985_);
  nor _78942_ (_28468_, _28466_, _11985_);
  nor _78943_ (_28469_, _28468_, _28467_);
  not _78944_ (_28470_, _28469_);
  or _78945_ (_28471_, _28470_, _11958_);
  and _78946_ (_28473_, _28471_, _06687_);
  and _78947_ (_28474_, _28473_, _28465_);
  nand _78948_ (_28475_, _12120_, _11982_);
  or _78949_ (_28476_, _28470_, _12120_);
  and _78950_ (_28477_, _28476_, _12126_);
  and _78951_ (_28478_, _28477_, _28475_);
  and _78952_ (_28479_, _12163_, _06220_);
  or _78953_ (_28480_, _12131_, _12163_);
  or _78954_ (_28481_, _12139_, _11981_);
  or _78955_ (_28482_, _28470_, _12141_);
  and _78956_ (_28484_, _28482_, _06160_);
  and _78957_ (_28485_, _28484_, _28481_);
  and _78958_ (_28486_, _12258_, _12163_);
  and _78959_ (_28487_, _28451_, _12256_);
  or _78960_ (_28488_, _28487_, _08443_);
  or _78961_ (_28489_, _28488_, _28486_);
  or _78962_ (_28490_, _28445_, _12267_);
  or _78963_ (_28491_, _12163_, _06582_);
  or _78964_ (_28492_, _12163_, _07057_);
  nor _78965_ (_28493_, _07056_, \oc8051_golden_model_1.PC [11]);
  nand _78966_ (_28495_, _28493_, _12265_);
  and _78967_ (_28496_, _28495_, _28492_);
  nor _78968_ (_28497_, _28496_, _06653_);
  nand _78969_ (_28498_, _28497_, _24799_);
  and _78970_ (_28499_, _28498_, _28491_);
  and _78971_ (_28500_, _28499_, _28490_);
  or _78972_ (_28501_, _28500_, _08445_);
  and _78973_ (_28502_, _28501_, _12281_);
  and _78974_ (_28503_, _28502_, _28489_);
  or _78975_ (_28504_, _28503_, _28485_);
  and _78976_ (_28506_, _28504_, _12134_);
  and _78977_ (_28507_, _28445_, _12287_);
  or _78978_ (_28508_, _28507_, _12286_);
  or _78979_ (_28509_, _28508_, _28506_);
  and _78980_ (_28510_, _28509_, _28480_);
  or _78981_ (_28511_, _28510_, _12293_);
  or _78982_ (_28512_, _28445_, _12292_);
  and _78983_ (_28513_, _28512_, _06229_);
  and _78984_ (_28514_, _28513_, _28511_);
  or _78985_ (_28515_, _28514_, _28479_);
  and _78986_ (_28517_, _28515_, _12300_);
  and _78987_ (_28518_, _28445_, _12302_);
  or _78988_ (_28519_, _28518_, _12307_);
  or _78989_ (_28520_, _28519_, _28517_);
  or _78990_ (_28521_, _12306_, _12163_);
  and _78991_ (_28522_, _28521_, _12125_);
  and _78992_ (_28523_, _28522_, _28520_);
  or _78993_ (_28524_, _28523_, _28478_);
  and _78994_ (_28525_, _28524_, _12089_);
  or _78995_ (_28526_, _28525_, _06236_);
  or _78996_ (_28528_, _28526_, _28474_);
  and _78997_ (_28529_, _12329_, _11981_);
  nor _78998_ (_28530_, _28469_, _12329_);
  or _78999_ (_28531_, _28530_, _06643_);
  or _79000_ (_28532_, _28531_, _28529_);
  and _79001_ (_28533_, _28532_, _12317_);
  and _79002_ (_28534_, _28533_, _28528_);
  nand _79003_ (_28535_, _28469_, _12347_);
  nand _79004_ (_28536_, _12346_, _11982_);
  and _79005_ (_28537_, _28536_, _06295_);
  and _79006_ (_28539_, _28537_, _28535_);
  or _79007_ (_28540_, _28539_, _28534_);
  and _79008_ (_28541_, _28540_, _11925_);
  nand _79009_ (_28542_, _28445_, _11924_);
  nand _79010_ (_28543_, _28542_, _12363_);
  or _79011_ (_28544_, _28543_, _28541_);
  or _79012_ (_28545_, _12363_, _12163_);
  and _79013_ (_28546_, _28545_, _12369_);
  and _79014_ (_28547_, _28546_, _28544_);
  and _79015_ (_28548_, _28445_, _12373_);
  or _79016_ (_28550_, _28548_, _12376_);
  or _79017_ (_28551_, _28550_, _28547_);
  or _79018_ (_28552_, _12375_, _12163_);
  and _79019_ (_28553_, _28552_, _12381_);
  and _79020_ (_28554_, _28553_, _28551_);
  and _79021_ (_28555_, _28445_, _12387_);
  or _79022_ (_28556_, _28555_, _12386_);
  or _79023_ (_28557_, _28556_, _28554_);
  or _79024_ (_28558_, _12163_, _12385_);
  and _79025_ (_28559_, _28558_, _05805_);
  and _79026_ (_28561_, _28559_, _28557_);
  nand _79027_ (_28562_, _28445_, _05870_);
  nand _79028_ (_28563_, _28562_, _12395_);
  or _79029_ (_28564_, _28563_, _28561_);
  or _79030_ (_28565_, _12395_, _12163_);
  and _79031_ (_28566_, _28565_, _11296_);
  and _79032_ (_28567_, _28566_, _28564_);
  nand _79033_ (_28568_, _11981_, _06293_);
  nand _79034_ (_28569_, _28568_, _06133_);
  or _79035_ (_28570_, _28569_, _28567_);
  or _79036_ (_28572_, _12163_, _06133_);
  and _79037_ (_28573_, _28572_, _06114_);
  and _79038_ (_28574_, _28573_, _28570_);
  or _79039_ (_28575_, _28574_, _28464_);
  and _79040_ (_28576_, _28575_, _11922_);
  and _79041_ (_28577_, _28445_, _12412_);
  or _79042_ (_28578_, _28577_, _12411_);
  or _79043_ (_28579_, _28578_, _28576_);
  or _79044_ (_28580_, _12410_, _12163_);
  and _79045_ (_28581_, _28580_, _12417_);
  and _79046_ (_28583_, _28581_, _28579_);
  and _79047_ (_28584_, _28451_, _12416_);
  or _79048_ (_28585_, _28584_, _08788_);
  or _79049_ (_28586_, _28585_, _28583_);
  and _79050_ (_28587_, _28586_, _28463_);
  or _79051_ (_28588_, _28587_, _06110_);
  nand _79052_ (_28589_, _11982_, _06110_);
  and _79053_ (_28590_, _28589_, _10752_);
  and _79054_ (_28591_, _28590_, _28588_);
  and _79055_ (_28592_, _12163_, _10751_);
  or _79056_ (_28594_, _28592_, _28591_);
  and _79057_ (_28595_, _28594_, _12432_);
  or _79058_ (_28596_, _12460_, \oc8051_golden_model_1.DPH [3]);
  nor _79059_ (_28597_, _12461_, _12432_);
  and _79060_ (_28598_, _28597_, _28596_);
  or _79061_ (_28599_, _28598_, _12470_);
  or _79062_ (_28600_, _28599_, _28595_);
  or _79063_ (_28601_, _12469_, _12163_);
  and _79064_ (_28602_, _28601_, _12474_);
  and _79065_ (_28603_, _28602_, _28600_);
  or _79066_ (_28605_, _28451_, _11101_);
  or _79067_ (_28606_, _12163_, _12480_);
  and _79068_ (_28607_, _28606_, _12473_);
  and _79069_ (_28608_, _28607_, _28605_);
  or _79070_ (_28609_, _28608_, _12478_);
  or _79071_ (_28610_, _28609_, _28603_);
  and _79072_ (_28611_, _28610_, _28462_);
  or _79073_ (_28612_, _28611_, _11917_);
  or _79074_ (_28613_, _12163_, _11916_);
  and _79075_ (_28614_, _28613_, _07127_);
  and _79076_ (_28616_, _28614_, _28612_);
  nand _79077_ (_28617_, _11981_, _06297_);
  nand _79078_ (_28618_, _28617_, _12493_);
  or _79079_ (_28619_, _28618_, _28616_);
  or _79080_ (_28620_, _12493_, _12163_);
  and _79081_ (_28621_, _28620_, _12497_);
  and _79082_ (_28622_, _28621_, _28619_);
  or _79083_ (_28623_, _28451_, _12480_);
  or _79084_ (_28624_, _12163_, _11101_);
  and _79085_ (_28625_, _28624_, _12496_);
  and _79086_ (_28626_, _28625_, _28623_);
  or _79087_ (_28627_, _28626_, _12505_);
  or _79088_ (_28628_, _28627_, _28622_);
  and _79089_ (_28629_, _28628_, _28460_);
  or _79090_ (_28630_, _28629_, _10822_);
  or _79091_ (_28631_, _12163_, _10821_);
  and _79092_ (_28632_, _28631_, _07132_);
  and _79093_ (_28633_, _28632_, _28630_);
  nand _79094_ (_28634_, _11981_, _06306_);
  nand _79095_ (_28635_, _28634_, _12514_);
  or _79096_ (_28638_, _28635_, _28633_);
  or _79097_ (_28639_, _12514_, _12163_);
  and _79098_ (_28640_, _28639_, _12518_);
  and _79099_ (_28641_, _28640_, _28638_);
  or _79100_ (_28642_, _28641_, _28459_);
  and _79101_ (_28643_, _28642_, _11912_);
  and _79102_ (_28644_, _28445_, _12522_);
  or _79103_ (_28645_, _28644_, _10850_);
  or _79104_ (_28646_, _28645_, _28643_);
  or _79105_ (_28647_, _12163_, _10849_);
  and _79106_ (_28649_, _28647_, _08819_);
  and _79107_ (_28650_, _28649_, _28646_);
  nand _79108_ (_28651_, _11981_, _06303_);
  nand _79109_ (_28652_, _28651_, _12535_);
  or _79110_ (_28653_, _28652_, _28650_);
  or _79111_ (_28654_, _12535_, _12163_);
  and _79112_ (_28655_, _28654_, _12539_);
  and _79113_ (_28656_, _28655_, _28653_);
  or _79114_ (_28657_, _28656_, _28455_);
  and _79115_ (_28658_, _28657_, _11907_);
  and _79116_ (_28660_, _28445_, _12547_);
  or _79117_ (_28661_, _28660_, _10897_);
  or _79118_ (_28662_, _28661_, _28658_);
  or _79119_ (_28663_, _12163_, _10896_);
  and _79120_ (_28664_, _28663_, _10926_);
  and _79121_ (_28665_, _28664_, _28662_);
  and _79122_ (_28666_, _28445_, _10925_);
  or _79123_ (_28667_, _28666_, _06417_);
  or _79124_ (_28668_, _28667_, _28665_);
  or _79125_ (_28669_, _07544_, _12558_);
  and _79126_ (_28671_, _28669_, _28668_);
  or _79127_ (_28672_, _28671_, _07142_);
  nor _79128_ (_28673_, _12163_, _05846_);
  nor _79129_ (_28674_, _28673_, _06301_);
  and _79130_ (_28675_, _28674_, _28672_);
  nand _79131_ (_28676_, _28469_, _12682_);
  or _79132_ (_28677_, _11981_, _12682_);
  and _79133_ (_28678_, _28677_, _06301_);
  and _79134_ (_28679_, _28678_, _28676_);
  or _79135_ (_28680_, _28679_, _12565_);
  or _79136_ (_28682_, _28680_, _28675_);
  and _79137_ (_28683_, _28682_, _28446_);
  or _79138_ (_28684_, _28683_, _12691_);
  or _79139_ (_28685_, _12690_, _12163_);
  and _79140_ (_28686_, _28685_, _12693_);
  and _79141_ (_28687_, _28686_, _28684_);
  and _79142_ (_28688_, _28445_, _10262_);
  or _79143_ (_28689_, _28688_, _06167_);
  or _79144_ (_28690_, _28689_, _28687_);
  or _79145_ (_28691_, _07544_, _06168_);
  and _79146_ (_28693_, _28691_, _28690_);
  or _79147_ (_28694_, _28693_, _05826_);
  or _79148_ (_28695_, _12163_, _12703_);
  and _79149_ (_28696_, _28695_, _06166_);
  and _79150_ (_28697_, _28696_, _28694_);
  or _79151_ (_28698_, _28470_, _12682_);
  nand _79152_ (_28699_, _11982_, _12682_);
  and _79153_ (_28700_, _28699_, _28698_);
  and _79154_ (_28701_, _28700_, _06165_);
  or _79155_ (_28702_, _28701_, _12712_);
  or _79156_ (_28704_, _28702_, _28697_);
  or _79157_ (_28705_, _28445_, _12711_);
  and _79158_ (_28706_, _28705_, _06829_);
  and _79159_ (_28707_, _28706_, _28704_);
  nand _79160_ (_28708_, _12163_, _06433_);
  nand _79161_ (_28709_, _28708_, _12719_);
  or _79162_ (_28710_, _28709_, _28707_);
  or _79163_ (_28711_, _28445_, _12719_);
  and _79164_ (_28712_, _28711_, _12723_);
  and _79165_ (_28713_, _28712_, _28710_);
  nor _79166_ (_28715_, _12723_, _06070_);
  or _79167_ (_28716_, _28715_, _05823_);
  or _79168_ (_28717_, _28716_, _28713_);
  or _79169_ (_28718_, _12163_, _12730_);
  and _79170_ (_28719_, _28718_, _05749_);
  and _79171_ (_28720_, _28719_, _28717_);
  and _79172_ (_28721_, _28700_, _05748_);
  or _79173_ (_28722_, _28721_, _12737_);
  or _79174_ (_28723_, _28722_, _28720_);
  or _79175_ (_28724_, _28445_, _12735_);
  and _79176_ (_28726_, _28724_, _06444_);
  and _79177_ (_28727_, _28726_, _28723_);
  nand _79178_ (_28728_, _12163_, _06440_);
  nand _79179_ (_28729_, _28728_, _12744_);
  or _79180_ (_28730_, _28729_, _28727_);
  or _79181_ (_28731_, _28445_, _12744_);
  and _79182_ (_28732_, _28731_, _12747_);
  and _79183_ (_28733_, _28732_, _28730_);
  nor _79184_ (_28734_, _12747_, _06070_);
  or _79185_ (_28735_, _28734_, _05821_);
  or _79186_ (_28737_, _28735_, _28733_);
  or _79187_ (_28738_, _12163_, _05822_);
  and _79188_ (_28739_, _28738_, _12755_);
  and _79189_ (_28740_, _28739_, _28737_);
  and _79190_ (_28741_, _28445_, _12754_);
  or _79191_ (_28742_, _28741_, _28740_);
  or _79192_ (_28743_, _28742_, _01321_);
  or _79193_ (_28744_, _01317_, \oc8051_golden_model_1.PC [11]);
  and _79194_ (_28745_, _28744_, _43100_);
  and _79195_ (_43700_, _28745_, _28743_);
  and _79196_ (_28747_, _11895_, _09242_);
  and _79197_ (_28748_, _28747_, \oc8051_golden_model_1.PC [11]);
  and _79198_ (_28749_, _28748_, \oc8051_golden_model_1.PC [12]);
  nor _79199_ (_28750_, _28748_, \oc8051_golden_model_1.PC [12]);
  nor _79200_ (_28751_, _28750_, _28749_);
  not _79201_ (_28752_, _28751_);
  and _79202_ (_28753_, _28752_, _12754_);
  and _79203_ (_28754_, _06876_, _06305_);
  or _79204_ (_28755_, _28754_, _05821_);
  and _79205_ (_28756_, _12156_, _10693_);
  and _79206_ (_28758_, _12239_, _12236_);
  nor _79207_ (_28759_, _28758_, _12240_);
  and _79208_ (_28760_, _28759_, \oc8051_golden_model_1.PSW [7]);
  or _79209_ (_28761_, _28760_, _28756_);
  and _79210_ (_28762_, _28761_, _12538_);
  and _79211_ (_28763_, _12156_, \oc8051_golden_model_1.PSW [7]);
  and _79212_ (_28764_, _28759_, _10693_);
  or _79213_ (_28765_, _28764_, _28763_);
  and _79214_ (_28766_, _28765_, _12517_);
  and _79215_ (_28767_, _12156_, _11101_);
  and _79216_ (_28769_, _28759_, _12480_);
  or _79217_ (_28770_, _28769_, _28767_);
  and _79218_ (_28771_, _28770_, _12473_);
  nor _79219_ (_28772_, _12156_, _08787_);
  and _79220_ (_28773_, _11977_, _05787_);
  and _79221_ (_28774_, _28751_, _11924_);
  and _79222_ (_28775_, _12072_, _12069_);
  nor _79223_ (_28776_, _28775_, _12073_);
  not _79224_ (_28777_, _28776_);
  and _79225_ (_28778_, _28777_, _11956_);
  nor _79226_ (_28780_, _11977_, _11956_);
  or _79227_ (_28781_, _28780_, _12089_);
  or _79228_ (_28782_, _28781_, _28778_);
  and _79229_ (_28783_, _12329_, _11977_);
  nor _79230_ (_28784_, _28777_, _12329_);
  nor _79231_ (_28785_, _28784_, _28783_);
  nor _79232_ (_28786_, _28785_, _06643_);
  not _79233_ (_28787_, _28786_);
  nand _79234_ (_28788_, _12120_, _11978_);
  or _79235_ (_28789_, _28776_, _12120_);
  and _79236_ (_28791_, _28789_, _12126_);
  and _79237_ (_28792_, _28791_, _28788_);
  or _79238_ (_28793_, _12139_, _11977_);
  or _79239_ (_28794_, _28776_, _12141_);
  and _79240_ (_28795_, _28794_, _06160_);
  nand _79241_ (_28796_, _28795_, _28793_);
  nand _79242_ (_28797_, _28759_, _12256_);
  not _79243_ (_28798_, _12156_);
  or _79244_ (_28799_, _12256_, _28798_);
  and _79245_ (_28800_, _28799_, _28797_);
  nand _79246_ (_28802_, _28800_, _08445_);
  and _79247_ (_28803_, _12263_, _28798_);
  nor _79248_ (_28804_, _28751_, _12263_);
  nor _79249_ (_28805_, _28804_, _28803_);
  nor _79250_ (_28806_, _28805_, _24799_);
  nor _79251_ (_28807_, _28752_, _12267_);
  not _79252_ (_28808_, _28807_);
  and _79253_ (_28809_, _28798_, _07056_);
  nor _79254_ (_28810_, _28809_, _06653_);
  not _79255_ (_28811_, _28810_);
  and _79256_ (_28813_, _12265_, \oc8051_golden_model_1.PC [12]);
  nor _79257_ (_28814_, _28813_, _07056_);
  nor _79258_ (_28815_, _28814_, _28811_);
  nor _79259_ (_28816_, _28815_, _06581_);
  and _79260_ (_28817_, _28816_, _28808_);
  nor _79261_ (_28818_, _28817_, _28806_);
  nor _79262_ (_28819_, _28818_, _08445_);
  not _79263_ (_28820_, _28819_);
  and _79264_ (_28821_, _28820_, _12281_);
  nand _79265_ (_28822_, _28821_, _28802_);
  nand _79266_ (_28824_, _28822_, _28796_);
  and _79267_ (_28825_, _28824_, _12134_);
  and _79268_ (_28826_, _28751_, _12287_);
  or _79269_ (_28827_, _28826_, _12286_);
  or _79270_ (_28828_, _28827_, _28825_);
  nor _79271_ (_28829_, _12131_, _12156_);
  nor _79272_ (_28830_, _28829_, _12293_);
  nand _79273_ (_28831_, _28830_, _28828_);
  nor _79274_ (_28832_, _28752_, _12292_);
  nor _79275_ (_28833_, _28832_, _06220_);
  nand _79276_ (_28835_, _28833_, _28831_);
  and _79277_ (_28836_, _28798_, _06220_);
  nor _79278_ (_28837_, _28836_, _12302_);
  nand _79279_ (_28838_, _28837_, _28835_);
  nor _79280_ (_28839_, _28752_, _12300_);
  nor _79281_ (_28840_, _28839_, _12307_);
  nand _79282_ (_28841_, _28840_, _28838_);
  nor _79283_ (_28842_, _12306_, _12156_);
  not _79284_ (_28843_, _28842_);
  and _79285_ (_28844_, _28843_, _12125_);
  and _79286_ (_28846_, _28844_, _28841_);
  nor _79287_ (_28847_, _28846_, _28792_);
  or _79288_ (_28848_, _28847_, _26862_);
  and _79289_ (_28849_, _28848_, _28787_);
  nand _79290_ (_28850_, _28849_, _28782_);
  nand _79291_ (_28851_, _28850_, _12317_);
  nand _79292_ (_28852_, _12346_, _11977_);
  nand _79293_ (_28853_, _28776_, _12347_);
  and _79294_ (_28854_, _28853_, _28852_);
  or _79295_ (_28855_, _28854_, _12317_);
  nand _79296_ (_28857_, _28855_, _28851_);
  nand _79297_ (_28858_, _28857_, _11925_);
  nand _79298_ (_28859_, _28858_, _12363_);
  or _79299_ (_28860_, _28859_, _28774_);
  nor _79300_ (_28861_, _12363_, _12156_);
  nor _79301_ (_28862_, _28861_, _12373_);
  nand _79302_ (_28863_, _28862_, _28860_);
  nor _79303_ (_28864_, _28752_, _12369_);
  nor _79304_ (_28865_, _28864_, _12376_);
  nand _79305_ (_28866_, _28865_, _28863_);
  nor _79306_ (_28868_, _12375_, _12156_);
  nor _79307_ (_28869_, _28868_, _12387_);
  nand _79308_ (_28870_, _28869_, _28866_);
  nor _79309_ (_28871_, _28752_, _12381_);
  nor _79310_ (_28872_, _28871_, _12386_);
  nand _79311_ (_28873_, _28872_, _28870_);
  nor _79312_ (_28874_, _12156_, _12385_);
  nor _79313_ (_28875_, _28874_, _05870_);
  nand _79314_ (_28876_, _28875_, _28873_);
  nor _79315_ (_28877_, _28752_, _05805_);
  nor _79316_ (_28879_, _28877_, _12396_);
  nand _79317_ (_28880_, _28879_, _28876_);
  nor _79318_ (_28881_, _12395_, _12156_);
  nor _79319_ (_28882_, _28881_, _06293_);
  nand _79320_ (_28883_, _28882_, _28880_);
  and _79321_ (_28884_, _11977_, _06293_);
  nor _79322_ (_28885_, _28884_, _13620_);
  nand _79323_ (_28886_, _28885_, _28883_);
  nor _79324_ (_28887_, _12156_, _06133_);
  nor _79325_ (_28888_, _28887_, _05787_);
  and _79326_ (_28890_, _28888_, _28886_);
  or _79327_ (_28891_, _28890_, _28773_);
  nand _79328_ (_28892_, _28891_, _11922_);
  nor _79329_ (_28893_, _28752_, _11922_);
  nor _79330_ (_28894_, _28893_, _12411_);
  nand _79331_ (_28895_, _28894_, _28892_);
  nor _79332_ (_28896_, _12410_, _12156_);
  nor _79333_ (_28897_, _28896_, _12416_);
  nand _79334_ (_28898_, _28897_, _28895_);
  and _79335_ (_28899_, _28759_, _12416_);
  nor _79336_ (_28901_, _28899_, _08788_);
  and _79337_ (_28902_, _28901_, _28898_);
  or _79338_ (_28903_, _28902_, _28772_);
  nand _79339_ (_28904_, _28903_, _06111_);
  and _79340_ (_28905_, _11978_, _06110_);
  nor _79341_ (_28906_, _28905_, _10751_);
  and _79342_ (_28907_, _28906_, _28904_);
  and _79343_ (_28908_, _12156_, _10751_);
  or _79344_ (_28909_, _28908_, _28907_);
  nand _79345_ (_28910_, _28909_, _12432_);
  nor _79346_ (_28912_, _12461_, \oc8051_golden_model_1.DPH [4]);
  nor _79347_ (_28913_, _28912_, _12462_);
  and _79348_ (_28914_, _28913_, _12431_);
  nor _79349_ (_28915_, _28914_, _12470_);
  nand _79350_ (_28916_, _28915_, _28910_);
  nor _79351_ (_28917_, _12469_, _12156_);
  nor _79352_ (_28918_, _28917_, _12473_);
  and _79353_ (_28919_, _28918_, _28916_);
  or _79354_ (_28920_, _28919_, _28771_);
  nand _79355_ (_28921_, _28920_, _11919_);
  nor _79356_ (_28923_, _28752_, _11919_);
  nor _79357_ (_28924_, _28923_, _11917_);
  nand _79358_ (_28925_, _28924_, _28921_);
  nor _79359_ (_28926_, _12156_, _11916_);
  nor _79360_ (_28927_, _28926_, _06297_);
  nand _79361_ (_28928_, _28927_, _28925_);
  and _79362_ (_28929_, _11977_, _06297_);
  not _79363_ (_28930_, _28929_);
  and _79364_ (_28931_, _28930_, _12493_);
  nand _79365_ (_28932_, _28931_, _28928_);
  nor _79366_ (_28934_, _12493_, _12156_);
  nor _79367_ (_28935_, _28934_, _12496_);
  and _79368_ (_28936_, _28935_, _28932_);
  and _79369_ (_28937_, _12156_, _12480_);
  and _79370_ (_28938_, _28759_, _11101_);
  or _79371_ (_28939_, _28938_, _28937_);
  and _79372_ (_28940_, _28939_, _12496_);
  or _79373_ (_28941_, _28940_, _28936_);
  nand _79374_ (_28942_, _28941_, _11914_);
  nor _79375_ (_28943_, _28752_, _11914_);
  nor _79376_ (_28945_, _28943_, _10822_);
  nand _79377_ (_28946_, _28945_, _28942_);
  nor _79378_ (_28947_, _12156_, _10821_);
  nor _79379_ (_28948_, _28947_, _06306_);
  nand _79380_ (_28949_, _28948_, _28946_);
  and _79381_ (_28950_, _11977_, _06306_);
  not _79382_ (_28951_, _28950_);
  and _79383_ (_28952_, _28951_, _12514_);
  nand _79384_ (_28953_, _28952_, _28949_);
  nor _79385_ (_28954_, _12514_, _12156_);
  nor _79386_ (_28956_, _28954_, _12517_);
  and _79387_ (_28957_, _28956_, _28953_);
  or _79388_ (_28958_, _28957_, _28766_);
  nand _79389_ (_28959_, _28958_, _11912_);
  nor _79390_ (_28960_, _28752_, _11912_);
  nor _79391_ (_28961_, _28960_, _10850_);
  nand _79392_ (_28962_, _28961_, _28959_);
  nor _79393_ (_28963_, _12156_, _10849_);
  nor _79394_ (_28964_, _28963_, _06303_);
  nand _79395_ (_28965_, _28964_, _28962_);
  not _79396_ (_28967_, _12535_);
  and _79397_ (_28968_, _11977_, _06303_);
  nor _79398_ (_28969_, _28968_, _28967_);
  nand _79399_ (_28970_, _28969_, _28965_);
  nor _79400_ (_28971_, _12535_, _12156_);
  nor _79401_ (_28972_, _28971_, _12538_);
  and _79402_ (_28973_, _28972_, _28970_);
  or _79403_ (_28974_, _28973_, _28762_);
  nand _79404_ (_28975_, _28974_, _11907_);
  nor _79405_ (_28976_, _28752_, _11907_);
  nor _79406_ (_28978_, _28976_, _10897_);
  nand _79407_ (_28979_, _28978_, _28975_);
  nor _79408_ (_28980_, _12156_, _10896_);
  nor _79409_ (_28981_, _28980_, _10925_);
  nand _79410_ (_28982_, _28981_, _28979_);
  and _79411_ (_28983_, _28751_, _10925_);
  nor _79412_ (_28984_, _28983_, _06417_);
  and _79413_ (_28985_, _28984_, _28982_);
  and _79414_ (_28986_, _08349_, _06417_);
  or _79415_ (_28987_, _28986_, _28985_);
  nand _79416_ (_28989_, _28987_, _05846_);
  nor _79417_ (_28990_, _12156_, _05846_);
  nor _79418_ (_28991_, _28990_, _06301_);
  and _79419_ (_28992_, _28991_, _28989_);
  nor _79420_ (_28993_, _11978_, _12682_);
  and _79421_ (_28994_, _28776_, _12682_);
  nor _79422_ (_28995_, _28994_, _28993_);
  nor _79423_ (_28996_, _28995_, _06421_);
  or _79424_ (_28997_, _28996_, _28992_);
  nand _79425_ (_28998_, _28997_, _11905_);
  nor _79426_ (_28999_, _28752_, _11905_);
  nor _79427_ (_29000_, _28999_, _12691_);
  nand _79428_ (_29001_, _29000_, _28998_);
  nor _79429_ (_29002_, _12690_, _12156_);
  nor _79430_ (_29003_, _29002_, _10262_);
  nand _79431_ (_29004_, _29003_, _29001_);
  and _79432_ (_29005_, _28751_, _10262_);
  nor _79433_ (_29006_, _29005_, _06167_);
  nand _79434_ (_29007_, _29006_, _29004_);
  and _79435_ (_29008_, _08349_, _06167_);
  nor _79436_ (_29011_, _29008_, _05826_);
  and _79437_ (_29012_, _29011_, _29007_);
  and _79438_ (_29013_, _12156_, _05826_);
  or _79439_ (_29014_, _29013_, _06165_);
  or _79440_ (_29015_, _29014_, _29012_);
  and _79441_ (_29016_, _11978_, _12682_);
  nor _79442_ (_29017_, _28776_, _12682_);
  nor _79443_ (_29018_, _29017_, _29016_);
  nor _79444_ (_29019_, _29018_, _06166_);
  nor _79445_ (_29020_, _29019_, _12712_);
  nand _79446_ (_29022_, _29020_, _29015_);
  nor _79447_ (_29023_, _28752_, _12711_);
  nor _79448_ (_29024_, _29023_, _06433_);
  nand _79449_ (_29025_, _29024_, _29022_);
  and _79450_ (_29026_, _28798_, _06433_);
  nor _79451_ (_29027_, _29026_, _25721_);
  nand _79452_ (_29028_, _29027_, _29025_);
  nor _79453_ (_29029_, _28752_, _12719_);
  nor _79454_ (_29030_, _29029_, _06310_);
  nand _79455_ (_29031_, _29030_, _29028_);
  and _79456_ (_29033_, _06876_, _06310_);
  nor _79457_ (_29034_, _29033_, _05823_);
  and _79458_ (_29035_, _29034_, _29031_);
  and _79459_ (_29036_, _12156_, _05823_);
  or _79460_ (_29037_, _29036_, _05748_);
  or _79461_ (_29038_, _29037_, _29035_);
  nor _79462_ (_29039_, _29018_, _05749_);
  nor _79463_ (_29040_, _29039_, _12737_);
  nand _79464_ (_29041_, _29040_, _29038_);
  nor _79465_ (_29042_, _28752_, _12735_);
  nor _79466_ (_29044_, _29042_, _06440_);
  nand _79467_ (_29045_, _29044_, _29041_);
  and _79468_ (_29046_, _28798_, _06440_);
  nor _79469_ (_29047_, _29046_, _26415_);
  nand _79470_ (_29048_, _29047_, _29045_);
  nor _79471_ (_29049_, _28752_, _12744_);
  nor _79472_ (_29050_, _29049_, _06305_);
  and _79473_ (_29051_, _29050_, _29048_);
  or _79474_ (_29052_, _29051_, _28755_);
  and _79475_ (_29053_, _12156_, _05821_);
  nor _79476_ (_29055_, _29053_, _12754_);
  and _79477_ (_29056_, _29055_, _29052_);
  nor _79478_ (_29057_, _29056_, _28753_);
  or _79479_ (_29058_, _29057_, _01321_);
  or _79480_ (_29059_, _01317_, \oc8051_golden_model_1.PC [12]);
  and _79481_ (_29060_, _29059_, _43100_);
  and _79482_ (_43701_, _29060_, _29058_);
  and _79483_ (_29061_, _12152_, _05823_);
  and _79484_ (_29062_, _28749_, \oc8051_golden_model_1.PC [13]);
  nor _79485_ (_29063_, _28749_, \oc8051_golden_model_1.PC [13]);
  nor _79486_ (_29065_, _29063_, _29062_);
  or _79487_ (_29066_, _29065_, _12719_);
  or _79488_ (_29067_, _29065_, _11905_);
  or _79489_ (_29068_, _29065_, _11912_);
  or _79490_ (_29069_, _29065_, _11919_);
  and _79491_ (_29070_, _11972_, _05787_);
  or _79492_ (_29071_, _11975_, _11974_);
  not _79493_ (_29072_, _29071_);
  nor _79494_ (_29073_, _29072_, _12074_);
  and _79495_ (_29074_, _29072_, _12074_);
  nor _79496_ (_29076_, _29074_, _29073_);
  not _79497_ (_29077_, _29076_);
  or _79498_ (_29078_, _29077_, _11958_);
  or _79499_ (_29079_, _11972_, _11956_);
  and _79500_ (_29080_, _29079_, _06687_);
  and _79501_ (_29081_, _29080_, _29078_);
  and _79502_ (_29082_, _12152_, _06220_);
  and _79503_ (_29083_, _29065_, _12287_);
  or _79504_ (_29084_, _29077_, _12141_);
  or _79505_ (_29085_, _12139_, _11972_);
  and _79506_ (_29087_, _29085_, _06160_);
  and _79507_ (_29088_, _29087_, _29084_);
  or _79508_ (_29089_, _29065_, _12267_);
  not _79509_ (_29090_, _12152_);
  nand _79510_ (_29091_, _29090_, _06581_);
  nand _79511_ (_29092_, _29090_, _07056_);
  nor _79512_ (_29093_, _07056_, \oc8051_golden_model_1.PC [13]);
  nand _79513_ (_29094_, _29093_, _12265_);
  nand _79514_ (_29095_, _29094_, _29092_);
  and _79515_ (_29096_, _29095_, _12264_);
  nand _79516_ (_29098_, _29096_, _24799_);
  and _79517_ (_29099_, _29098_, _08443_);
  and _79518_ (_29100_, _29099_, _29091_);
  and _79519_ (_29101_, _29100_, _29089_);
  or _79520_ (_29102_, _12256_, _12152_);
  or _79521_ (_29103_, _12154_, _12153_);
  not _79522_ (_29104_, _29103_);
  nor _79523_ (_29105_, _29104_, _12241_);
  and _79524_ (_29106_, _29104_, _12241_);
  or _79525_ (_29107_, _29106_, _29105_);
  or _79526_ (_29109_, _29107_, _12258_);
  and _79527_ (_29110_, _29109_, _08445_);
  and _79528_ (_29111_, _29110_, _29102_);
  or _79529_ (_29112_, _29111_, _29101_);
  and _79530_ (_29113_, _29112_, _12281_);
  or _79531_ (_29114_, _29113_, _29088_);
  and _79532_ (_29115_, _29114_, _12134_);
  or _79533_ (_29116_, _29115_, _29083_);
  and _79534_ (_29117_, _29116_, _12131_);
  or _79535_ (_29118_, _12131_, _29090_);
  nand _79536_ (_29120_, _29118_, _12292_);
  or _79537_ (_29121_, _29120_, _29117_);
  or _79538_ (_29122_, _29065_, _12292_);
  and _79539_ (_29123_, _29122_, _06229_);
  and _79540_ (_29124_, _29123_, _29121_);
  or _79541_ (_29125_, _29124_, _29082_);
  and _79542_ (_29126_, _29125_, _12300_);
  not _79543_ (_29127_, _29065_);
  or _79544_ (_29128_, _29127_, _12300_);
  nand _79545_ (_29129_, _29128_, _12306_);
  or _79546_ (_29131_, _29129_, _29126_);
  or _79547_ (_29132_, _12306_, _12152_);
  and _79548_ (_29133_, _29132_, _29131_);
  or _79549_ (_29134_, _29133_, _12126_);
  and _79550_ (_29135_, _12120_, _11972_);
  nor _79551_ (_29136_, _29076_, _12120_);
  or _79552_ (_29137_, _29136_, _29135_);
  or _79553_ (_29138_, _29137_, _12125_);
  and _79554_ (_29139_, _29138_, _12089_);
  and _79555_ (_29140_, _29139_, _29134_);
  or _79556_ (_29142_, _29140_, _06236_);
  or _79557_ (_29143_, _29142_, _29081_);
  and _79558_ (_29144_, _12329_, _11972_);
  nor _79559_ (_29145_, _29076_, _12329_);
  or _79560_ (_29146_, _29145_, _06643_);
  or _79561_ (_29147_, _29146_, _29144_);
  and _79562_ (_29148_, _29147_, _12317_);
  and _79563_ (_29149_, _29148_, _29143_);
  nand _79564_ (_29150_, _29076_, _12347_);
  nand _79565_ (_29151_, _12346_, _11973_);
  and _79566_ (_29153_, _29151_, _06295_);
  and _79567_ (_29154_, _29153_, _29150_);
  or _79568_ (_29155_, _29154_, _29149_);
  and _79569_ (_29156_, _29155_, _11925_);
  nand _79570_ (_29157_, _29065_, _11924_);
  nand _79571_ (_29158_, _29157_, _12363_);
  or _79572_ (_29159_, _29158_, _29156_);
  or _79573_ (_29160_, _12363_, _12152_);
  and _79574_ (_29161_, _29160_, _12369_);
  and _79575_ (_29162_, _29161_, _29159_);
  nor _79576_ (_29164_, _29127_, _12369_);
  or _79577_ (_29165_, _29164_, _12376_);
  or _79578_ (_29166_, _29165_, _29162_);
  or _79579_ (_29167_, _12375_, _12152_);
  and _79580_ (_29168_, _29167_, _12381_);
  and _79581_ (_29169_, _29168_, _29166_);
  nor _79582_ (_29170_, _29127_, _12381_);
  or _79583_ (_29171_, _29170_, _12386_);
  or _79584_ (_29172_, _29171_, _29169_);
  or _79585_ (_29173_, _12152_, _12385_);
  and _79586_ (_29175_, _29173_, _05805_);
  and _79587_ (_29176_, _29175_, _29172_);
  or _79588_ (_29177_, _29127_, _05805_);
  nand _79589_ (_29178_, _29177_, _12395_);
  or _79590_ (_29179_, _29178_, _29176_);
  or _79591_ (_29180_, _12395_, _12152_);
  and _79592_ (_29181_, _29180_, _11296_);
  and _79593_ (_29182_, _29181_, _29179_);
  nand _79594_ (_29183_, _11972_, _06293_);
  nand _79595_ (_29184_, _29183_, _06133_);
  or _79596_ (_29186_, _29184_, _29182_);
  or _79597_ (_29187_, _12152_, _06133_);
  and _79598_ (_29188_, _29187_, _06114_);
  and _79599_ (_29189_, _29188_, _29186_);
  or _79600_ (_29190_, _29189_, _29070_);
  and _79601_ (_29191_, _29190_, _11922_);
  nor _79602_ (_29192_, _29127_, _11922_);
  or _79603_ (_29193_, _29192_, _12411_);
  or _79604_ (_29194_, _29193_, _29191_);
  or _79605_ (_29195_, _12410_, _12152_);
  and _79606_ (_29197_, _29195_, _12417_);
  and _79607_ (_29198_, _29197_, _29194_);
  and _79608_ (_29199_, _29107_, _12416_);
  or _79609_ (_29200_, _29199_, _08788_);
  or _79610_ (_29201_, _29200_, _29198_);
  or _79611_ (_29202_, _12152_, _08787_);
  and _79612_ (_29203_, _29202_, _06111_);
  and _79613_ (_29204_, _29203_, _29201_);
  and _79614_ (_29205_, _11972_, _06110_);
  or _79615_ (_29206_, _29205_, _10751_);
  or _79616_ (_29208_, _29206_, _29204_);
  nand _79617_ (_29209_, _29090_, _10751_);
  and _79618_ (_29210_, _29209_, _12432_);
  and _79619_ (_29211_, _29210_, _29208_);
  or _79620_ (_29212_, _12462_, \oc8051_golden_model_1.DPH [5]);
  nor _79621_ (_29213_, _12463_, _12432_);
  and _79622_ (_29214_, _29213_, _29212_);
  or _79623_ (_29215_, _29214_, _12470_);
  or _79624_ (_29216_, _29215_, _29211_);
  or _79625_ (_29217_, _12469_, _12152_);
  and _79626_ (_29219_, _29217_, _12474_);
  and _79627_ (_29220_, _29219_, _29216_);
  or _79628_ (_29221_, _29107_, _11101_);
  or _79629_ (_29222_, _12152_, _12480_);
  and _79630_ (_29223_, _29222_, _12473_);
  and _79631_ (_29224_, _29223_, _29221_);
  or _79632_ (_29225_, _29224_, _12478_);
  or _79633_ (_29226_, _29225_, _29220_);
  and _79634_ (_29227_, _29226_, _29069_);
  or _79635_ (_29228_, _29227_, _11917_);
  or _79636_ (_29230_, _12152_, _11916_);
  and _79637_ (_29231_, _29230_, _07127_);
  and _79638_ (_29232_, _29231_, _29228_);
  nand _79639_ (_29233_, _11972_, _06297_);
  nand _79640_ (_29234_, _29233_, _12493_);
  or _79641_ (_29235_, _29234_, _29232_);
  or _79642_ (_29236_, _12493_, _12152_);
  and _79643_ (_29237_, _29236_, _12497_);
  and _79644_ (_29238_, _29237_, _29235_);
  or _79645_ (_29239_, _29107_, _12480_);
  or _79646_ (_29241_, _12152_, _11101_);
  and _79647_ (_29242_, _29241_, _12496_);
  and _79648_ (_29243_, _29242_, _29239_);
  or _79649_ (_29244_, _29243_, _29238_);
  and _79650_ (_29245_, _29244_, _11914_);
  nor _79651_ (_29246_, _29127_, _11914_);
  or _79652_ (_29247_, _29246_, _10822_);
  or _79653_ (_29248_, _29247_, _29245_);
  or _79654_ (_29249_, _12152_, _10821_);
  and _79655_ (_29250_, _29249_, _07132_);
  and _79656_ (_29252_, _29250_, _29248_);
  nand _79657_ (_29253_, _11972_, _06306_);
  nand _79658_ (_29254_, _29253_, _12514_);
  or _79659_ (_29255_, _29254_, _29252_);
  or _79660_ (_29256_, _12514_, _12152_);
  and _79661_ (_29257_, _29256_, _12518_);
  and _79662_ (_29258_, _29257_, _29255_);
  or _79663_ (_29259_, _29107_, \oc8051_golden_model_1.PSW [7]);
  or _79664_ (_29260_, _12152_, _10693_);
  and _79665_ (_29261_, _29260_, _12517_);
  and _79666_ (_29263_, _29261_, _29259_);
  or _79667_ (_29264_, _29263_, _12522_);
  or _79668_ (_29265_, _29264_, _29258_);
  and _79669_ (_29266_, _29265_, _29068_);
  or _79670_ (_29267_, _29266_, _10850_);
  or _79671_ (_29268_, _12152_, _10849_);
  and _79672_ (_29269_, _29268_, _08819_);
  and _79673_ (_29270_, _29269_, _29267_);
  nand _79674_ (_29271_, _11972_, _06303_);
  nand _79675_ (_29272_, _29271_, _12535_);
  or _79676_ (_29274_, _29272_, _29270_);
  or _79677_ (_29275_, _12535_, _12152_);
  and _79678_ (_29276_, _29275_, _12539_);
  and _79679_ (_29277_, _29276_, _29274_);
  or _79680_ (_29278_, _29107_, _10693_);
  or _79681_ (_29279_, _12152_, \oc8051_golden_model_1.PSW [7]);
  and _79682_ (_29280_, _29279_, _12538_);
  and _79683_ (_29281_, _29280_, _29278_);
  or _79684_ (_29282_, _29281_, _29277_);
  and _79685_ (_29283_, _29282_, _11907_);
  nor _79686_ (_29285_, _29127_, _11907_);
  or _79687_ (_29286_, _29285_, _10897_);
  or _79688_ (_29287_, _29286_, _29283_);
  or _79689_ (_29288_, _12152_, _10896_);
  and _79690_ (_29289_, _29288_, _10926_);
  and _79691_ (_29290_, _29289_, _29287_);
  and _79692_ (_29291_, _29065_, _10925_);
  or _79693_ (_29292_, _29291_, _06417_);
  or _79694_ (_29293_, _29292_, _29290_);
  or _79695_ (_29294_, _08101_, _12558_);
  and _79696_ (_29296_, _29294_, _29293_);
  or _79697_ (_29297_, _29296_, _07142_);
  nor _79698_ (_29298_, _12152_, _05846_);
  nor _79699_ (_29299_, _29298_, _06301_);
  and _79700_ (_29300_, _29299_, _29297_);
  or _79701_ (_29301_, _11972_, _12682_);
  nand _79702_ (_29302_, _29076_, _12682_);
  and _79703_ (_29303_, _29302_, _06301_);
  and _79704_ (_29304_, _29303_, _29301_);
  or _79705_ (_29305_, _29304_, _12565_);
  or _79706_ (_29307_, _29305_, _29300_);
  and _79707_ (_29308_, _29307_, _29067_);
  or _79708_ (_29309_, _29308_, _12691_);
  or _79709_ (_29310_, _12690_, _12152_);
  and _79710_ (_29311_, _29310_, _12693_);
  and _79711_ (_29312_, _29311_, _29309_);
  and _79712_ (_29313_, _29065_, _10262_);
  or _79713_ (_29314_, _29313_, _06167_);
  or _79714_ (_29315_, _29314_, _29312_);
  or _79715_ (_29316_, _08101_, _06168_);
  and _79716_ (_29318_, _29316_, _29315_);
  or _79717_ (_29319_, _29318_, _05826_);
  nand _79718_ (_29320_, _29090_, _05826_);
  and _79719_ (_29321_, _29320_, _06166_);
  and _79720_ (_29322_, _29321_, _29319_);
  or _79721_ (_29323_, _29077_, _12682_);
  nand _79722_ (_29324_, _11973_, _12682_);
  and _79723_ (_29325_, _29324_, _29323_);
  and _79724_ (_29326_, _29325_, _06165_);
  or _79725_ (_29327_, _29326_, _12712_);
  or _79726_ (_29329_, _29327_, _29322_);
  or _79727_ (_29330_, _29065_, _12711_);
  and _79728_ (_29331_, _29330_, _06829_);
  and _79729_ (_29332_, _29331_, _29329_);
  nand _79730_ (_29333_, _12152_, _06433_);
  nand _79731_ (_29334_, _29333_, _12719_);
  or _79732_ (_29335_, _29334_, _29332_);
  and _79733_ (_29336_, _29335_, _29066_);
  or _79734_ (_29337_, _29336_, _06310_);
  nand _79735_ (_29338_, _06477_, _06310_);
  and _79736_ (_29340_, _29338_, _12730_);
  and _79737_ (_29341_, _29340_, _29337_);
  or _79738_ (_29342_, _29341_, _29061_);
  and _79739_ (_29343_, _29342_, _05749_);
  and _79740_ (_29344_, _29325_, _05748_);
  or _79741_ (_29345_, _29344_, _12737_);
  or _79742_ (_29346_, _29345_, _29343_);
  or _79743_ (_29347_, _29065_, _12735_);
  and _79744_ (_29348_, _29347_, _06444_);
  and _79745_ (_29349_, _29348_, _29346_);
  nand _79746_ (_29351_, _12152_, _06440_);
  nand _79747_ (_29352_, _29351_, _12744_);
  or _79748_ (_29353_, _29352_, _29349_);
  or _79749_ (_29354_, _29065_, _12744_);
  and _79750_ (_29355_, _29354_, _12747_);
  and _79751_ (_29356_, _29355_, _29353_);
  nor _79752_ (_29357_, _06477_, _12747_);
  or _79753_ (_29358_, _29357_, _05821_);
  or _79754_ (_29359_, _29358_, _29356_);
  nand _79755_ (_29360_, _29090_, _05821_);
  and _79756_ (_29362_, _29360_, _12755_);
  and _79757_ (_29363_, _29362_, _29359_);
  and _79758_ (_29364_, _29065_, _12754_);
  or _79759_ (_29365_, _29364_, _29363_);
  or _79760_ (_29366_, _29365_, _01321_);
  or _79761_ (_29367_, _01317_, \oc8051_golden_model_1.PC [13]);
  and _79762_ (_29368_, _29367_, _43100_);
  and _79763_ (_43702_, _29368_, _29366_);
  and _79764_ (_29369_, _06305_, _06203_);
  or _79765_ (_29370_, _29369_, _05821_);
  nor _79766_ (_29372_, _29062_, \oc8051_golden_model_1.PC [14]);
  nor _79767_ (_29373_, _29372_, _11901_);
  not _79768_ (_29374_, _29373_);
  and _79769_ (_29375_, _29374_, _10262_);
  not _79770_ (_29376_, _12146_);
  or _79771_ (_29377_, _12535_, _29376_);
  or _79772_ (_29378_, _12514_, _29376_);
  or _79773_ (_29379_, _12493_, _29376_);
  nor _79774_ (_29380_, _12410_, _12146_);
  and _79775_ (_29381_, _12076_, _11970_);
  or _79776_ (_29383_, _29381_, _12077_);
  and _79777_ (_29384_, _29383_, _11956_);
  nor _79778_ (_29385_, _11965_, _11956_);
  or _79779_ (_29386_, _29385_, _12089_);
  or _79780_ (_29387_, _29386_, _29384_);
  or _79781_ (_29388_, _29383_, _12329_);
  nand _79782_ (_29389_, _12329_, _11965_);
  and _79783_ (_29390_, _29389_, _29388_);
  or _79784_ (_29391_, _29390_, _06643_);
  and _79785_ (_29392_, _29376_, _06220_);
  and _79786_ (_29394_, _29374_, _12287_);
  and _79787_ (_29395_, _29383_, _12139_);
  and _79788_ (_29396_, _12141_, _11966_);
  or _79789_ (_29397_, _29396_, _29395_);
  and _79790_ (_29398_, _29397_, _06160_);
  nor _79791_ (_29399_, _29373_, _12263_);
  and _79792_ (_29400_, _12263_, _29376_);
  or _79793_ (_29401_, _29400_, _29399_);
  and _79794_ (_29402_, _29401_, _24800_);
  or _79795_ (_29403_, _29374_, _12267_);
  and _79796_ (_29405_, _29376_, _07056_);
  or _79797_ (_29406_, _29405_, _06653_);
  nand _79798_ (_29407_, _12265_, \oc8051_golden_model_1.PC [14]);
  and _79799_ (_29408_, _29407_, _07057_);
  or _79800_ (_29409_, _29408_, _29406_);
  and _79801_ (_29410_, _29409_, _06582_);
  and _79802_ (_29411_, _29410_, _29403_);
  or _79803_ (_29412_, _29411_, _29402_);
  and _79804_ (_29413_, _29412_, _08443_);
  or _79805_ (_29414_, _12256_, _29376_);
  and _79806_ (_29416_, _12243_, _12150_);
  nor _79807_ (_29417_, _29416_, _12244_);
  nand _79808_ (_29418_, _29417_, _12256_);
  and _79809_ (_29419_, _29418_, _08445_);
  and _79810_ (_29420_, _29419_, _29414_);
  or _79811_ (_29421_, _29420_, _29413_);
  and _79812_ (_29422_, _29421_, _12281_);
  or _79813_ (_29423_, _29422_, _29398_);
  and _79814_ (_29424_, _29423_, _12134_);
  or _79815_ (_29425_, _29424_, _29394_);
  and _79816_ (_29427_, _29425_, _12131_);
  or _79817_ (_29428_, _12131_, _12146_);
  nand _79818_ (_29429_, _29428_, _12292_);
  or _79819_ (_29430_, _29429_, _29427_);
  or _79820_ (_29431_, _29374_, _12292_);
  and _79821_ (_29432_, _29431_, _06229_);
  and _79822_ (_29433_, _29432_, _29430_);
  or _79823_ (_29434_, _29433_, _29392_);
  and _79824_ (_29435_, _29434_, _12300_);
  or _79825_ (_29436_, _29373_, _12300_);
  nand _79826_ (_29438_, _29436_, _12306_);
  or _79827_ (_29439_, _29438_, _29435_);
  or _79828_ (_29440_, _12306_, _29376_);
  and _79829_ (_29441_, _29440_, _12125_);
  and _79830_ (_29442_, _29441_, _29439_);
  nand _79831_ (_29443_, _12120_, _11965_);
  or _79832_ (_29444_, _29383_, _12120_);
  and _79833_ (_29445_, _29444_, _29443_);
  and _79834_ (_29446_, _29445_, _12126_);
  or _79835_ (_29447_, _29446_, _26862_);
  or _79836_ (_29449_, _29447_, _29442_);
  and _79837_ (_29450_, _29449_, _29391_);
  and _79838_ (_29451_, _29450_, _29387_);
  or _79839_ (_29452_, _29451_, _06295_);
  and _79840_ (_29453_, _29383_, _12347_);
  and _79841_ (_29454_, _12346_, _11966_);
  or _79842_ (_29455_, _29454_, _12317_);
  or _79843_ (_29456_, _29455_, _29453_);
  and _79844_ (_29457_, _29456_, _11925_);
  and _79845_ (_29458_, _29457_, _29452_);
  and _79846_ (_29460_, _29374_, _11924_);
  or _79847_ (_29461_, _29460_, _29458_);
  and _79848_ (_29462_, _29461_, _12363_);
  nor _79849_ (_29463_, _12363_, _12146_);
  or _79850_ (_29464_, _29463_, _29462_);
  and _79851_ (_29465_, _29464_, _12369_);
  nor _79852_ (_29466_, _29373_, _12369_);
  or _79853_ (_29467_, _29466_, _12376_);
  or _79854_ (_29468_, _29467_, _29465_);
  or _79855_ (_29469_, _12375_, _29376_);
  and _79856_ (_29471_, _29469_, _12381_);
  and _79857_ (_29472_, _29471_, _29468_);
  nor _79858_ (_29473_, _29373_, _12381_);
  or _79859_ (_29474_, _29473_, _12386_);
  or _79860_ (_29475_, _29474_, _29472_);
  or _79861_ (_29476_, _29376_, _12385_);
  and _79862_ (_29477_, _29476_, _05805_);
  and _79863_ (_29478_, _29477_, _29475_);
  or _79864_ (_29479_, _29373_, _05805_);
  nand _79865_ (_29480_, _29479_, _12395_);
  or _79866_ (_29482_, _29480_, _29478_);
  or _79867_ (_29483_, _12395_, _29376_);
  and _79868_ (_29484_, _29483_, _11296_);
  and _79869_ (_29485_, _29484_, _29482_);
  nand _79870_ (_29486_, _11966_, _06293_);
  nand _79871_ (_29487_, _29486_, _06133_);
  or _79872_ (_29488_, _29487_, _29485_);
  or _79873_ (_29489_, _29376_, _06133_);
  and _79874_ (_29490_, _29489_, _06114_);
  and _79875_ (_29491_, _29490_, _29488_);
  nand _79876_ (_29493_, _11966_, _05787_);
  nand _79877_ (_29494_, _29493_, _11922_);
  or _79878_ (_29495_, _29494_, _29491_);
  or _79879_ (_29496_, _29374_, _11922_);
  and _79880_ (_29497_, _29496_, _12410_);
  and _79881_ (_29498_, _29497_, _29495_);
  or _79882_ (_29499_, _29498_, _29380_);
  and _79883_ (_29500_, _29499_, _12417_);
  nor _79884_ (_29501_, _29417_, _12417_);
  or _79885_ (_29502_, _29501_, _08788_);
  or _79886_ (_29504_, _29502_, _29500_);
  or _79887_ (_29505_, _29376_, _08787_);
  and _79888_ (_29506_, _29505_, _06111_);
  and _79889_ (_29507_, _29506_, _29504_);
  and _79890_ (_29508_, _11966_, _06110_);
  or _79891_ (_29509_, _29508_, _29507_);
  and _79892_ (_29510_, _29509_, _10752_);
  and _79893_ (_29511_, _29376_, _10751_);
  or _79894_ (_29512_, _29511_, _12431_);
  or _79895_ (_29513_, _29512_, _29510_);
  nor _79896_ (_29515_, _12463_, \oc8051_golden_model_1.DPH [6]);
  or _79897_ (_29516_, _12464_, _12432_);
  or _79898_ (_29517_, _29516_, _29515_);
  and _79899_ (_29518_, _29517_, _12469_);
  and _79900_ (_29519_, _29518_, _29513_);
  nor _79901_ (_29520_, _12469_, _12146_);
  or _79902_ (_29521_, _29520_, _12473_);
  or _79903_ (_29522_, _29521_, _29519_);
  nor _79904_ (_29523_, _29417_, _11101_);
  or _79905_ (_29524_, _12146_, _12480_);
  nand _79906_ (_29525_, _29524_, _12473_);
  or _79907_ (_29526_, _29525_, _29523_);
  and _79908_ (_29527_, _29526_, _11919_);
  and _79909_ (_29528_, _29527_, _29522_);
  nor _79910_ (_29529_, _29373_, _11919_);
  or _79911_ (_29530_, _29529_, _11917_);
  or _79912_ (_29531_, _29530_, _29528_);
  or _79913_ (_29532_, _29376_, _11916_);
  and _79914_ (_29533_, _29532_, _07127_);
  and _79915_ (_29534_, _29533_, _29531_);
  nand _79916_ (_29537_, _11966_, _06297_);
  nand _79917_ (_29538_, _29537_, _12493_);
  or _79918_ (_29539_, _29538_, _29534_);
  and _79919_ (_29540_, _29539_, _29379_);
  or _79920_ (_29541_, _29540_, _12496_);
  nor _79921_ (_29542_, _29417_, _12480_);
  or _79922_ (_29543_, _12146_, _11101_);
  nand _79923_ (_29544_, _29543_, _12496_);
  or _79924_ (_29545_, _29544_, _29542_);
  and _79925_ (_29546_, _29545_, _11914_);
  and _79926_ (_29548_, _29546_, _29541_);
  nor _79927_ (_29549_, _29373_, _11914_);
  or _79928_ (_29550_, _29549_, _10822_);
  or _79929_ (_29551_, _29550_, _29548_);
  or _79930_ (_29552_, _29376_, _10821_);
  and _79931_ (_29553_, _29552_, _07132_);
  and _79932_ (_29554_, _29553_, _29551_);
  nand _79933_ (_29555_, _11966_, _06306_);
  nand _79934_ (_29556_, _29555_, _12514_);
  or _79935_ (_29557_, _29556_, _29554_);
  and _79936_ (_29559_, _29557_, _29378_);
  or _79937_ (_29560_, _29559_, _12517_);
  nor _79938_ (_29561_, _29417_, \oc8051_golden_model_1.PSW [7]);
  or _79939_ (_29562_, _12146_, _10693_);
  nand _79940_ (_29563_, _29562_, _12517_);
  or _79941_ (_29564_, _29563_, _29561_);
  and _79942_ (_29565_, _29564_, _11912_);
  and _79943_ (_29566_, _29565_, _29560_);
  nor _79944_ (_29567_, _29373_, _11912_);
  or _79945_ (_29568_, _29567_, _10850_);
  or _79946_ (_29570_, _29568_, _29566_);
  or _79947_ (_29571_, _29376_, _10849_);
  and _79948_ (_29572_, _29571_, _08819_);
  and _79949_ (_29573_, _29572_, _29570_);
  nand _79950_ (_29574_, _11966_, _06303_);
  nand _79951_ (_29575_, _29574_, _12535_);
  or _79952_ (_29576_, _29575_, _29573_);
  and _79953_ (_29577_, _29576_, _29377_);
  or _79954_ (_29578_, _29577_, _12538_);
  or _79955_ (_29579_, _29417_, _10693_);
  or _79956_ (_29581_, _12146_, \oc8051_golden_model_1.PSW [7]);
  and _79957_ (_29582_, _29581_, _12538_);
  and _79958_ (_29583_, _29582_, _29579_);
  nor _79959_ (_29584_, _29583_, _12547_);
  and _79960_ (_29585_, _29584_, _29578_);
  nor _79961_ (_29586_, _29373_, _11907_);
  or _79962_ (_29587_, _29586_, _10897_);
  or _79963_ (_29588_, _29587_, _29585_);
  or _79964_ (_29589_, _29376_, _10896_);
  and _79965_ (_29590_, _29589_, _10926_);
  and _79966_ (_29592_, _29590_, _29588_);
  and _79967_ (_29593_, _29374_, _10925_);
  or _79968_ (_29594_, _29593_, _06417_);
  or _79969_ (_29595_, _29594_, _29592_);
  or _79970_ (_29596_, _08347_, _12558_);
  and _79971_ (_29597_, _29596_, _05846_);
  and _79972_ (_29598_, _29597_, _29595_);
  nor _79973_ (_29599_, _12146_, _05846_);
  or _79974_ (_29600_, _29599_, _06301_);
  or _79975_ (_29601_, _29600_, _29598_);
  nor _79976_ (_29603_, _11965_, _12682_);
  and _79977_ (_29604_, _29383_, _12682_);
  or _79978_ (_29605_, _29604_, _06421_);
  or _79979_ (_29606_, _29605_, _29603_);
  and _79980_ (_29607_, _29606_, _11905_);
  and _79981_ (_29608_, _29607_, _29601_);
  nor _79982_ (_29609_, _29373_, _11905_);
  or _79983_ (_29610_, _29609_, _12691_);
  or _79984_ (_29611_, _29610_, _29608_);
  or _79985_ (_29612_, _12690_, _29376_);
  and _79986_ (_29614_, _29612_, _12693_);
  and _79987_ (_29615_, _29614_, _29611_);
  or _79988_ (_29616_, _29615_, _29375_);
  and _79989_ (_29617_, _29616_, _06168_);
  and _79990_ (_29618_, _08347_, _06167_);
  or _79991_ (_29619_, _29618_, _05826_);
  or _79992_ (_29620_, _29619_, _29617_);
  nand _79993_ (_29621_, _12146_, _05826_);
  and _79994_ (_29622_, _29621_, _06166_);
  and _79995_ (_29623_, _29622_, _29620_);
  nand _79996_ (_29625_, _11965_, _12682_);
  or _79997_ (_29626_, _29383_, _12682_);
  and _79998_ (_29627_, _29626_, _29625_);
  and _79999_ (_29628_, _29627_, _06165_);
  or _80000_ (_29629_, _29628_, _29623_);
  and _80001_ (_29630_, _29629_, _12711_);
  nor _80002_ (_29631_, _29373_, _12711_);
  or _80003_ (_29632_, _29631_, _29630_);
  and _80004_ (_29633_, _29632_, _06829_);
  nand _80005_ (_29634_, _29376_, _06433_);
  nand _80006_ (_29636_, _29634_, _12719_);
  or _80007_ (_29637_, _29636_, _29633_);
  or _80008_ (_29638_, _29374_, _12719_);
  and _80009_ (_29639_, _29638_, _12723_);
  and _80010_ (_29640_, _29639_, _29637_);
  and _80011_ (_29641_, _06310_, _06203_);
  or _80012_ (_29642_, _29641_, _05823_);
  or _80013_ (_29643_, _29642_, _29640_);
  nand _80014_ (_29644_, _12146_, _05823_);
  and _80015_ (_29645_, _29644_, _05749_);
  and _80016_ (_29647_, _29645_, _29643_);
  and _80017_ (_29648_, _29627_, _05748_);
  or _80018_ (_29649_, _29648_, _12737_);
  or _80019_ (_29650_, _29649_, _29647_);
  or _80020_ (_29651_, _29374_, _12735_);
  and _80021_ (_29652_, _29651_, _06444_);
  and _80022_ (_29653_, _29652_, _29650_);
  nand _80023_ (_29654_, _29376_, _06440_);
  nand _80024_ (_29655_, _29654_, _12744_);
  or _80025_ (_29656_, _29655_, _29653_);
  or _80026_ (_29658_, _29374_, _12744_);
  and _80027_ (_29659_, _29658_, _12747_);
  and _80028_ (_29660_, _29659_, _29656_);
  nor _80029_ (_29661_, _29660_, _29370_);
  and _80030_ (_29662_, _12146_, _05821_);
  nor _80031_ (_29663_, _29662_, _29661_);
  or _80032_ (_29664_, _29663_, _12754_);
  nand _80033_ (_29665_, _29373_, _12754_);
  and _80034_ (_29666_, _29665_, _29664_);
  nand _80035_ (_29667_, _29666_, _01317_);
  or _80036_ (_29669_, _01317_, \oc8051_golden_model_1.PC [14]);
  and _80037_ (_29670_, _29669_, _43100_);
  and _80038_ (_43703_, _29670_, _29667_);
  not _80039_ (_29671_, _12768_);
  and _80040_ (_29672_, _29671_, \oc8051_golden_model_1.P2 [0]);
  or _80041_ (_29673_, _12858_, \oc8051_golden_model_1.ACC [0]);
  nand _80042_ (_29674_, _12858_, \oc8051_golden_model_1.ACC [0]);
  and _80043_ (_29675_, _29674_, _29673_);
  and _80044_ (_29676_, _29675_, _12768_);
  or _80045_ (_29677_, _29676_, _29672_);
  and _80046_ (_29679_, _29677_, _06402_);
  and _80047_ (_29680_, _12768_, _07049_);
  or _80048_ (_29681_, _29680_, _29672_);
  or _80049_ (_29682_, _29681_, _06132_);
  nor _80050_ (_29683_, _12858_, _29671_);
  or _80051_ (_29684_, _29683_, _29672_);
  or _80052_ (_29685_, _29684_, _06161_);
  and _80053_ (_29686_, _12768_, \oc8051_golden_model_1.ACC [0]);
  or _80054_ (_29687_, _29686_, _29672_);
  and _80055_ (_29688_, _29687_, _07056_);
  and _80056_ (_29690_, _07057_, \oc8051_golden_model_1.P2 [0]);
  or _80057_ (_29691_, _29690_, _06160_);
  or _80058_ (_29692_, _29691_, _29688_);
  and _80059_ (_29693_, _29692_, _06157_);
  and _80060_ (_29694_, _29693_, _29685_);
  not _80061_ (_29695_, _12773_);
  and _80062_ (_29696_, _29695_, \oc8051_golden_model_1.P2 [0]);
  and _80063_ (_29697_, _07847_, \oc8051_golden_model_1.P0 [0]);
  and _80064_ (_29698_, _12773_, \oc8051_golden_model_1.P2 [0]);
  or _80065_ (_29699_, _29698_, _29697_);
  and _80066_ (_29701_, _12778_, \oc8051_golden_model_1.P1 [0]);
  and _80067_ (_29702_, _12780_, \oc8051_golden_model_1.P3 [0]);
  or _80068_ (_29703_, _29702_, _29701_);
  or _80069_ (_29704_, _29703_, _29699_);
  or _80070_ (_29705_, _14169_, _29704_);
  and _80071_ (_29706_, _29705_, _12773_);
  or _80072_ (_29707_, _29706_, _29696_);
  and _80073_ (_29708_, _29707_, _06156_);
  or _80074_ (_29709_, _29708_, _29694_);
  and _80075_ (_29710_, _29709_, _07075_);
  and _80076_ (_29712_, _29681_, _06217_);
  or _80077_ (_29713_, _29712_, _06220_);
  or _80078_ (_29714_, _29713_, _29710_);
  or _80079_ (_29715_, _29687_, _06229_);
  and _80080_ (_29716_, _29715_, _06153_);
  and _80081_ (_29717_, _29716_, _29714_);
  and _80082_ (_29718_, _29672_, _06152_);
  or _80083_ (_29719_, _29718_, _06145_);
  or _80084_ (_29720_, _29719_, _29717_);
  or _80085_ (_29721_, _29684_, _06146_);
  and _80086_ (_29723_, _29721_, _06140_);
  and _80087_ (_29724_, _29723_, _29720_);
  or _80088_ (_29725_, _29696_, _14170_);
  and _80089_ (_29726_, _29725_, _06139_);
  and _80090_ (_29727_, _29726_, _29707_);
  or _80091_ (_29728_, _29727_, _09842_);
  or _80092_ (_29729_, _29728_, _29724_);
  and _80093_ (_29730_, _29729_, _29682_);
  or _80094_ (_29731_, _29730_, _06116_);
  and _80095_ (_29732_, _12768_, _09160_);
  or _80096_ (_29734_, _29672_, _06117_);
  or _80097_ (_29735_, _29734_, _29732_);
  and _80098_ (_29736_, _29735_, _06114_);
  and _80099_ (_29737_, _29736_, _29731_);
  and _80100_ (_29738_, _12918_, \oc8051_golden_model_1.P1 [0]);
  and _80101_ (_29739_, _12916_, \oc8051_golden_model_1.P0 [0]);
  and _80102_ (_29740_, _12920_, \oc8051_golden_model_1.P2 [0]);
  and _80103_ (_29741_, _12922_, \oc8051_golden_model_1.P3 [0]);
  or _80104_ (_29742_, _29741_, _29740_);
  or _80105_ (_29743_, _29742_, _29739_);
  or _80106_ (_29745_, _29743_, _29738_);
  or _80107_ (_29746_, _29745_, _14260_);
  and _80108_ (_29747_, _29746_, _12768_);
  or _80109_ (_29748_, _29747_, _29672_);
  and _80110_ (_29749_, _29748_, _05787_);
  or _80111_ (_29750_, _29749_, _29737_);
  or _80112_ (_29751_, _29750_, _11136_);
  or _80113_ (_29752_, _12858_, _08708_);
  and _80114_ (_29753_, _12858_, _08708_);
  not _80115_ (_29754_, _29753_);
  and _80116_ (_29756_, _29754_, _29752_);
  and _80117_ (_29757_, _29756_, _12768_);
  or _80118_ (_29758_, _29672_, _07127_);
  or _80119_ (_29759_, _29758_, _29757_);
  and _80120_ (_29760_, _12768_, _08708_);
  or _80121_ (_29761_, _29760_, _29672_);
  or _80122_ (_29762_, _29761_, _06111_);
  and _80123_ (_29763_, _29762_, _07125_);
  and _80124_ (_29764_, _29763_, _29759_);
  and _80125_ (_29765_, _29764_, _29751_);
  or _80126_ (_29767_, _29765_, _29679_);
  and _80127_ (_29768_, _29767_, _07132_);
  nand _80128_ (_29769_, _29761_, _06306_);
  nor _80129_ (_29770_, _29769_, _29683_);
  or _80130_ (_29771_, _29770_, _29768_);
  and _80131_ (_29772_, _29771_, _07130_);
  or _80132_ (_29773_, _29672_, _12858_);
  and _80133_ (_29774_, _29687_, _06411_);
  and _80134_ (_29775_, _29774_, _29773_);
  or _80135_ (_29776_, _29775_, _06303_);
  or _80136_ (_29778_, _29776_, _29772_);
  and _80137_ (_29779_, _29752_, _12768_);
  or _80138_ (_29780_, _29672_, _08819_);
  or _80139_ (_29781_, _29780_, _29779_);
  and _80140_ (_29782_, _29781_, _08824_);
  and _80141_ (_29783_, _29782_, _29778_);
  and _80142_ (_29784_, _29673_, _12768_);
  or _80143_ (_29785_, _29784_, _29672_);
  and _80144_ (_29786_, _29785_, _06396_);
  or _80145_ (_29787_, _29786_, _06433_);
  or _80146_ (_29789_, _29787_, _29783_);
  or _80147_ (_29790_, _29684_, _06829_);
  and _80148_ (_29791_, _29790_, _05749_);
  and _80149_ (_29792_, _29791_, _29789_);
  and _80150_ (_29793_, _29672_, _05748_);
  or _80151_ (_29794_, _29793_, _06440_);
  or _80152_ (_29795_, _29794_, _29792_);
  or _80153_ (_29796_, _29684_, _06444_);
  and _80154_ (_29797_, _29796_, _01317_);
  and _80155_ (_29798_, _29797_, _29795_);
  nor _80156_ (_29799_, \oc8051_golden_model_1.P2 [0], rst);
  nor _80157_ (_29800_, _29799_, _00000_);
  or _80158_ (_43705_, _29800_, _29798_);
  nor _80159_ (_29801_, \oc8051_golden_model_1.P2 [1], rst);
  nor _80160_ (_29802_, _29801_, _00000_);
  and _80161_ (_29803_, _07847_, \oc8051_golden_model_1.P0 [1]);
  and _80162_ (_29804_, _12778_, \oc8051_golden_model_1.P1 [1]);
  or _80163_ (_29805_, _29804_, _29803_);
  and _80164_ (_29806_, _12773_, \oc8051_golden_model_1.P2 [1]);
  and _80165_ (_29807_, _12780_, \oc8051_golden_model_1.P3 [1]);
  or _80166_ (_29810_, _29807_, _29806_);
  or _80167_ (_29811_, _29810_, _29805_);
  or _80168_ (_29812_, _29811_, _12627_);
  nand _80169_ (_29813_, _29812_, _07781_);
  or _80170_ (_29814_, _14367_, _29811_);
  and _80171_ (_29815_, _29814_, _12773_);
  and _80172_ (_29816_, _29815_, _29813_);
  and _80173_ (_29817_, _29695_, \oc8051_golden_model_1.P2 [1]);
  or _80174_ (_29818_, _29817_, _06146_);
  or _80175_ (_29819_, _29818_, _29816_);
  or _80176_ (_29821_, _12768_, \oc8051_golden_model_1.P2 [1]);
  not _80177_ (_29822_, _12977_);
  and _80178_ (_29823_, _29822_, _12859_);
  and _80179_ (_29824_, _29823_, _12768_);
  not _80180_ (_29825_, _29824_);
  and _80181_ (_29826_, _29825_, _29821_);
  or _80182_ (_29827_, _29826_, _06161_);
  nand _80183_ (_29828_, _12768_, _05887_);
  and _80184_ (_29829_, _29828_, _29821_);
  and _80185_ (_29830_, _29829_, _07056_);
  and _80186_ (_29832_, _07057_, \oc8051_golden_model_1.P2 [1]);
  or _80187_ (_29833_, _29832_, _06160_);
  or _80188_ (_29834_, _29833_, _29830_);
  and _80189_ (_29835_, _29834_, _06157_);
  and _80190_ (_29836_, _29835_, _29827_);
  or _80191_ (_29837_, _29817_, _06217_);
  or _80192_ (_29838_, _29837_, _29815_);
  and _80193_ (_29839_, _29838_, _13860_);
  or _80194_ (_29840_, _29839_, _29836_);
  and _80195_ (_29841_, _29671_, \oc8051_golden_model_1.P2 [1]);
  and _80196_ (_29843_, _12768_, _07306_);
  or _80197_ (_29844_, _29843_, _29841_);
  or _80198_ (_29845_, _29844_, _07075_);
  and _80199_ (_29846_, _29845_, _29840_);
  or _80200_ (_29847_, _29846_, _06220_);
  or _80201_ (_29848_, _29829_, _06229_);
  and _80202_ (_29849_, _29848_, _06153_);
  and _80203_ (_29850_, _29849_, _29847_);
  and _80204_ (_29851_, _29812_, _14348_);
  and _80205_ (_29852_, _29851_, _12773_);
  or _80206_ (_29854_, _29852_, _29817_);
  and _80207_ (_29855_, _29854_, _06152_);
  or _80208_ (_29856_, _29855_, _06145_);
  or _80209_ (_29857_, _29856_, _29850_);
  and _80210_ (_29858_, _29857_, _29819_);
  and _80211_ (_29859_, _29858_, _06140_);
  or _80212_ (_29860_, _29851_, _14350_);
  and _80213_ (_29861_, _29860_, _12773_);
  or _80214_ (_29862_, _29817_, _29861_);
  and _80215_ (_29863_, _29862_, _06139_);
  or _80216_ (_29865_, _29863_, _09842_);
  or _80217_ (_29866_, _29865_, _29859_);
  or _80218_ (_29867_, _29844_, _06132_);
  and _80219_ (_29868_, _29867_, _29866_);
  or _80220_ (_29869_, _29868_, _06116_);
  and _80221_ (_29870_, _12768_, _09115_);
  or _80222_ (_29871_, _29841_, _06117_);
  or _80223_ (_29872_, _29871_, _29870_);
  and _80224_ (_29873_, _29872_, _06114_);
  and _80225_ (_29874_, _29873_, _29869_);
  and _80226_ (_29876_, _12916_, \oc8051_golden_model_1.P0 [1]);
  and _80227_ (_29877_, _12918_, \oc8051_golden_model_1.P1 [1]);
  and _80228_ (_29878_, _12920_, \oc8051_golden_model_1.P2 [1]);
  and _80229_ (_29879_, _12922_, \oc8051_golden_model_1.P3 [1]);
  or _80230_ (_29880_, _29879_, _29878_);
  or _80231_ (_29881_, _29880_, _29877_);
  or _80232_ (_29882_, _29881_, _29876_);
  or _80233_ (_29883_, _29882_, _14442_);
  and _80234_ (_29884_, _29883_, _12768_);
  or _80235_ (_29885_, _29884_, _29841_);
  and _80236_ (_29887_, _29885_, _05787_);
  or _80237_ (_29888_, _29887_, _29874_);
  and _80238_ (_29889_, _29888_, _06298_);
  nand _80239_ (_29890_, _12768_, _06945_);
  and _80240_ (_29891_, _29821_, _06110_);
  and _80241_ (_29892_, _29891_, _29890_);
  or _80242_ (_29893_, _12850_, _08763_);
  and _80243_ (_29894_, _29893_, _12768_);
  or _80244_ (_29895_, _29894_, _29841_);
  and _80245_ (_29896_, _12850_, _08763_);
  not _80246_ (_29898_, _29896_);
  or _80247_ (_29899_, _29898_, _29841_);
  and _80248_ (_29900_, _29899_, _06297_);
  and _80249_ (_29901_, _29900_, _29895_);
  or _80250_ (_29902_, _29901_, _29892_);
  or _80251_ (_29903_, _29902_, _29889_);
  and _80252_ (_29904_, _29903_, _07125_);
  or _80253_ (_29905_, _12850_, \oc8051_golden_model_1.ACC [1]);
  and _80254_ (_29906_, _29905_, _12768_);
  or _80255_ (_29907_, _29906_, _29841_);
  nand _80256_ (_29909_, _12850_, \oc8051_golden_model_1.ACC [1]);
  or _80257_ (_29910_, _29909_, _29841_);
  and _80258_ (_29911_, _29910_, _06402_);
  and _80259_ (_29912_, _29911_, _29907_);
  or _80260_ (_29913_, _29912_, _29904_);
  and _80261_ (_29914_, _29913_, _07132_);
  or _80262_ (_29915_, _29896_, _29671_);
  and _80263_ (_29916_, _29821_, _06306_);
  and _80264_ (_29917_, _29916_, _29915_);
  or _80265_ (_29918_, _29917_, _29914_);
  and _80266_ (_29920_, _29918_, _07130_);
  or _80267_ (_29921_, _29841_, _12850_);
  and _80268_ (_29922_, _29829_, _06411_);
  and _80269_ (_29923_, _29922_, _29921_);
  or _80270_ (_29924_, _29923_, _06303_);
  or _80271_ (_29925_, _29924_, _29920_);
  or _80272_ (_29926_, _29895_, _08819_);
  and _80273_ (_29927_, _29926_, _08824_);
  and _80274_ (_29928_, _29927_, _29925_);
  and _80275_ (_29929_, _29907_, _06396_);
  or _80276_ (_29931_, _29929_, _06433_);
  or _80277_ (_29932_, _29931_, _29928_);
  or _80278_ (_29933_, _29826_, _06829_);
  and _80279_ (_29934_, _29933_, _05749_);
  and _80280_ (_29935_, _29934_, _29932_);
  and _80281_ (_29936_, _29854_, _05748_);
  or _80282_ (_29937_, _29936_, _06440_);
  or _80283_ (_29938_, _29937_, _29935_);
  or _80284_ (_29939_, _29841_, _06444_);
  or _80285_ (_29940_, _29939_, _29824_);
  and _80286_ (_29942_, _29940_, _01317_);
  and _80287_ (_29943_, _29942_, _29938_);
  or _80288_ (_43706_, _29943_, _29802_);
  and _80289_ (_29944_, _29671_, \oc8051_golden_model_1.P2 [2]);
  or _80290_ (_29945_, _12842_, _08768_);
  and _80291_ (_29946_, _29945_, _12768_);
  or _80292_ (_29947_, _29946_, _29944_);
  nand _80293_ (_29948_, _12842_, _08768_);
  or _80294_ (_29949_, _29948_, _29944_);
  and _80295_ (_29950_, _29949_, _06297_);
  and _80296_ (_29952_, _29950_, _29947_);
  and _80297_ (_29953_, _12859_, _12842_);
  or _80298_ (_29954_, _29953_, _12860_);
  and _80299_ (_29955_, _29954_, _12768_);
  or _80300_ (_29956_, _29955_, _29944_);
  or _80301_ (_29957_, _29956_, _06161_);
  and _80302_ (_29958_, _12768_, \oc8051_golden_model_1.ACC [2]);
  or _80303_ (_29959_, _29958_, _29944_);
  and _80304_ (_29960_, _29959_, _07056_);
  and _80305_ (_29961_, _07057_, \oc8051_golden_model_1.P2 [2]);
  or _80306_ (_29963_, _29961_, _06160_);
  or _80307_ (_29964_, _29963_, _29960_);
  and _80308_ (_29965_, _29964_, _06157_);
  and _80309_ (_29966_, _29965_, _29957_);
  and _80310_ (_29967_, _29695_, \oc8051_golden_model_1.P2 [2]);
  and _80311_ (_29968_, _07847_, \oc8051_golden_model_1.P0 [2]);
  and _80312_ (_29969_, _12773_, \oc8051_golden_model_1.P2 [2]);
  or _80313_ (_29970_, _29969_, _29968_);
  and _80314_ (_29971_, _12778_, \oc8051_golden_model_1.P1 [2]);
  and _80315_ (_29972_, _12780_, \oc8051_golden_model_1.P3 [2]);
  or _80316_ (_29974_, _29972_, _29971_);
  or _80317_ (_29975_, _29974_, _29970_);
  or _80318_ (_29976_, _14538_, _29975_);
  and _80319_ (_29977_, _29976_, _12773_);
  or _80320_ (_29978_, _29977_, _29967_);
  and _80321_ (_29979_, _29978_, _06156_);
  or _80322_ (_29980_, _29979_, _06217_);
  or _80323_ (_29981_, _29980_, _29966_);
  and _80324_ (_29982_, _12768_, _07708_);
  or _80325_ (_29983_, _29982_, _29944_);
  or _80326_ (_29985_, _29983_, _07075_);
  and _80327_ (_29986_, _29985_, _29981_);
  or _80328_ (_29987_, _29986_, _06220_);
  or _80329_ (_29988_, _29959_, _06229_);
  and _80330_ (_29989_, _29988_, _06153_);
  and _80331_ (_29990_, _29989_, _29987_);
  or _80332_ (_29991_, _29975_, _12644_);
  and _80333_ (_29992_, _29991_, _14535_);
  and _80334_ (_29993_, _29992_, _12773_);
  or _80335_ (_29994_, _29993_, _29967_);
  and _80336_ (_29996_, _29994_, _06152_);
  or _80337_ (_29997_, _29996_, _06145_);
  or _80338_ (_29998_, _29997_, _29990_);
  nand _80339_ (_29999_, _29991_, _07848_);
  or _80340_ (_30000_, _29967_, _29999_);
  and _80341_ (_30001_, _30000_, _29978_);
  or _80342_ (_30002_, _30001_, _06146_);
  and _80343_ (_30003_, _30002_, _06140_);
  and _80344_ (_30004_, _30003_, _29998_);
  or _80345_ (_30005_, _29992_, _14582_);
  and _80346_ (_30007_, _30005_, _12773_);
  or _80347_ (_30008_, _30007_, _29967_);
  and _80348_ (_30009_, _30008_, _06139_);
  or _80349_ (_30010_, _30009_, _09842_);
  or _80350_ (_30011_, _30010_, _30004_);
  or _80351_ (_30012_, _29983_, _06132_);
  and _80352_ (_30013_, _30012_, _30011_);
  or _80353_ (_30014_, _30013_, _06116_);
  and _80354_ (_30015_, _12768_, _09211_);
  or _80355_ (_30016_, _29944_, _06117_);
  or _80356_ (_30018_, _30016_, _30015_);
  and _80357_ (_30019_, _30018_, _06114_);
  and _80358_ (_30020_, _30019_, _30014_);
  and _80359_ (_30021_, _12916_, \oc8051_golden_model_1.P0 [2]);
  and _80360_ (_30022_, _12918_, \oc8051_golden_model_1.P1 [2]);
  and _80361_ (_30023_, _12920_, \oc8051_golden_model_1.P2 [2]);
  and _80362_ (_30024_, _12922_, \oc8051_golden_model_1.P3 [2]);
  or _80363_ (_30025_, _30024_, _30023_);
  or _80364_ (_30026_, _30025_, _30022_);
  or _80365_ (_30027_, _30026_, _30021_);
  or _80366_ (_30029_, _30027_, _14630_);
  and _80367_ (_30030_, _30029_, _12768_);
  or _80368_ (_30031_, _30030_, _29944_);
  and _80369_ (_30032_, _30031_, _05787_);
  or _80370_ (_30033_, _30032_, _06110_);
  or _80371_ (_30034_, _30033_, _30020_);
  and _80372_ (_30035_, _12768_, _08768_);
  or _80373_ (_30036_, _30035_, _29944_);
  or _80374_ (_30037_, _30036_, _06111_);
  and _80375_ (_30038_, _30037_, _07127_);
  and _80376_ (_30040_, _30038_, _30034_);
  or _80377_ (_30041_, _30040_, _29952_);
  and _80378_ (_30042_, _30041_, _07125_);
  or _80379_ (_30043_, _12842_, \oc8051_golden_model_1.ACC [2]);
  and _80380_ (_30044_, _30043_, _12768_);
  or _80381_ (_30045_, _30044_, _29944_);
  nand _80382_ (_30046_, _12842_, \oc8051_golden_model_1.ACC [2]);
  or _80383_ (_30047_, _30046_, _29944_);
  and _80384_ (_30048_, _30047_, _06402_);
  and _80385_ (_30049_, _30048_, _30045_);
  or _80386_ (_30051_, _30049_, _30042_);
  and _80387_ (_30052_, _30051_, _07132_);
  or _80388_ (_30053_, _29944_, _12842_);
  and _80389_ (_30054_, _30036_, _06306_);
  and _80390_ (_30055_, _30054_, _30053_);
  or _80391_ (_30056_, _30055_, _30052_);
  and _80392_ (_30057_, _30056_, _07130_);
  and _80393_ (_30058_, _29959_, _06411_);
  and _80394_ (_30059_, _30058_, _30053_);
  or _80395_ (_30060_, _30059_, _06303_);
  or _80396_ (_30062_, _30060_, _30057_);
  or _80397_ (_30063_, _29947_, _08819_);
  and _80398_ (_30064_, _30063_, _08824_);
  and _80399_ (_30065_, _30064_, _30062_);
  and _80400_ (_30066_, _30045_, _06396_);
  or _80401_ (_30067_, _30066_, _06433_);
  or _80402_ (_30068_, _30067_, _30065_);
  or _80403_ (_30069_, _29956_, _06829_);
  and _80404_ (_30070_, _30069_, _05749_);
  and _80405_ (_30071_, _30070_, _30068_);
  and _80406_ (_30073_, _29994_, _05748_);
  or _80407_ (_30074_, _30073_, _06440_);
  or _80408_ (_30075_, _30074_, _30071_);
  nor _80409_ (_30076_, _12977_, _12842_);
  nor _80410_ (_30077_, _30076_, _12978_);
  and _80411_ (_30078_, _30077_, _12768_);
  or _80412_ (_30079_, _29944_, _06444_);
  or _80413_ (_30080_, _30079_, _30078_);
  and _80414_ (_30081_, _30080_, _01317_);
  and _80415_ (_30082_, _30081_, _30075_);
  nor _80416_ (_30084_, \oc8051_golden_model_1.P2 [2], rst);
  nor _80417_ (_30085_, _30084_, _00000_);
  or _80418_ (_43707_, _30085_, _30082_);
  and _80419_ (_30086_, _29671_, \oc8051_golden_model_1.P2 [3]);
  and _80420_ (_30087_, _12768_, _07544_);
  or _80421_ (_30088_, _30087_, _30086_);
  or _80422_ (_30089_, _30088_, _06132_);
  and _80423_ (_30090_, _29695_, \oc8051_golden_model_1.P2 [3]);
  and _80424_ (_30091_, _07847_, \oc8051_golden_model_1.P0 [3]);
  and _80425_ (_30092_, _12778_, \oc8051_golden_model_1.P1 [3]);
  or _80426_ (_30094_, _30092_, _30091_);
  and _80427_ (_30095_, _12773_, \oc8051_golden_model_1.P2 [3]);
  and _80428_ (_30096_, _12780_, \oc8051_golden_model_1.P3 [3]);
  or _80429_ (_30097_, _30096_, _30095_);
  or _80430_ (_30098_, _30097_, _30094_);
  or _80431_ (_30099_, _30098_, _12595_);
  and _80432_ (_30100_, _30099_, _14730_);
  and _80433_ (_30101_, _30100_, _12773_);
  or _80434_ (_30102_, _30101_, _30090_);
  and _80435_ (_30103_, _30102_, _06152_);
  and _80436_ (_30105_, _12861_, _12834_);
  or _80437_ (_30106_, _30105_, _12862_);
  and _80438_ (_30107_, _30106_, _12768_);
  or _80439_ (_30108_, _30107_, _30086_);
  or _80440_ (_30109_, _30108_, _06161_);
  and _80441_ (_30110_, _12768_, \oc8051_golden_model_1.ACC [3]);
  or _80442_ (_30111_, _30110_, _30086_);
  and _80443_ (_30112_, _30111_, _07056_);
  and _80444_ (_30113_, _07057_, \oc8051_golden_model_1.P2 [3]);
  or _80445_ (_30114_, _30113_, _06160_);
  or _80446_ (_30116_, _30114_, _30112_);
  and _80447_ (_30117_, _30116_, _06157_);
  and _80448_ (_30118_, _30117_, _30109_);
  or _80449_ (_30119_, _14735_, _30098_);
  and _80450_ (_30120_, _30119_, _12773_);
  or _80451_ (_30121_, _30120_, _30090_);
  and _80452_ (_30122_, _30121_, _06156_);
  or _80453_ (_30123_, _30122_, _06217_);
  or _80454_ (_30124_, _30123_, _30118_);
  or _80455_ (_30125_, _30088_, _07075_);
  and _80456_ (_30127_, _30125_, _30124_);
  or _80457_ (_30128_, _30127_, _06220_);
  or _80458_ (_30129_, _30111_, _06229_);
  and _80459_ (_30130_, _30129_, _06153_);
  and _80460_ (_30131_, _30130_, _30128_);
  or _80461_ (_30132_, _30131_, _30103_);
  and _80462_ (_30133_, _30132_, _06146_);
  nand _80463_ (_30134_, _30099_, _07851_);
  or _80464_ (_30135_, _30090_, _30134_);
  and _80465_ (_30136_, _30121_, _06145_);
  and _80466_ (_30138_, _30136_, _30135_);
  or _80467_ (_30139_, _30138_, _30133_);
  and _80468_ (_30140_, _30139_, _06140_);
  or _80469_ (_30141_, _30100_, _14729_);
  and _80470_ (_30142_, _30141_, _12773_);
  or _80471_ (_30143_, _30142_, _30090_);
  and _80472_ (_30144_, _30143_, _06139_);
  or _80473_ (_30145_, _30144_, _09842_);
  or _80474_ (_30146_, _30145_, _30140_);
  and _80475_ (_30147_, _30146_, _30089_);
  or _80476_ (_30149_, _30147_, _06116_);
  and _80477_ (_30150_, _12768_, _09210_);
  or _80478_ (_30151_, _30086_, _06117_);
  or _80479_ (_30152_, _30151_, _30150_);
  and _80480_ (_30153_, _30152_, _06114_);
  and _80481_ (_30154_, _30153_, _30149_);
  and _80482_ (_30155_, _12916_, \oc8051_golden_model_1.P0 [3]);
  and _80483_ (_30156_, _12918_, \oc8051_golden_model_1.P1 [3]);
  and _80484_ (_30157_, _12920_, \oc8051_golden_model_1.P2 [3]);
  and _80485_ (_30158_, _12922_, \oc8051_golden_model_1.P3 [3]);
  or _80486_ (_30160_, _30158_, _30157_);
  or _80487_ (_30161_, _30160_, _30156_);
  or _80488_ (_30162_, _30161_, _30155_);
  or _80489_ (_30163_, _30162_, _14825_);
  and _80490_ (_30164_, _30163_, _12768_);
  or _80491_ (_30165_, _30164_, _30086_);
  and _80492_ (_30166_, _30165_, _05787_);
  or _80493_ (_30167_, _30166_, _06110_);
  or _80494_ (_30168_, _30167_, _30154_);
  and _80495_ (_30169_, _12768_, _08712_);
  or _80496_ (_30171_, _30169_, _30086_);
  or _80497_ (_30172_, _30171_, _06111_);
  and _80498_ (_30173_, _30172_, _07127_);
  and _80499_ (_30174_, _30173_, _30168_);
  or _80500_ (_30175_, _12834_, _08712_);
  and _80501_ (_30176_, _30175_, _12768_);
  or _80502_ (_30177_, _30176_, _30086_);
  nand _80503_ (_30178_, _12834_, _08712_);
  or _80504_ (_30179_, _30178_, _30086_);
  and _80505_ (_30180_, _30179_, _06297_);
  and _80506_ (_30182_, _30180_, _30177_);
  or _80507_ (_30183_, _30182_, _30174_);
  and _80508_ (_30184_, _30183_, _07125_);
  or _80509_ (_30185_, _12834_, \oc8051_golden_model_1.ACC [3]);
  and _80510_ (_30186_, _30185_, _12768_);
  or _80511_ (_30187_, _30186_, _30086_);
  nand _80512_ (_30188_, _12834_, \oc8051_golden_model_1.ACC [3]);
  or _80513_ (_30189_, _30188_, _30086_);
  and _80514_ (_30190_, _30189_, _06402_);
  and _80515_ (_30191_, _30190_, _30187_);
  or _80516_ (_30193_, _30191_, _30184_);
  and _80517_ (_30194_, _30193_, _07132_);
  or _80518_ (_30195_, _30086_, _12834_);
  and _80519_ (_30196_, _30171_, _06306_);
  and _80520_ (_30197_, _30196_, _30195_);
  or _80521_ (_30198_, _30197_, _30194_);
  and _80522_ (_30199_, _30198_, _07130_);
  and _80523_ (_30200_, _30111_, _06411_);
  and _80524_ (_30201_, _30200_, _30195_);
  or _80525_ (_30202_, _30201_, _06303_);
  or _80526_ (_30204_, _30202_, _30199_);
  or _80527_ (_30205_, _30177_, _08819_);
  and _80528_ (_30206_, _30205_, _08824_);
  and _80529_ (_30207_, _30206_, _30204_);
  and _80530_ (_30208_, _30187_, _06396_);
  or _80531_ (_30209_, _30208_, _06433_);
  or _80532_ (_30210_, _30209_, _30207_);
  or _80533_ (_30211_, _30108_, _06829_);
  and _80534_ (_30212_, _30211_, _05749_);
  and _80535_ (_30213_, _30212_, _30210_);
  and _80536_ (_30215_, _30102_, _05748_);
  or _80537_ (_30216_, _30215_, _06440_);
  or _80538_ (_30217_, _30216_, _30213_);
  nor _80539_ (_30218_, _12978_, _12834_);
  nor _80540_ (_30219_, _30218_, _12979_);
  and _80541_ (_30220_, _30219_, _12768_);
  or _80542_ (_30221_, _30086_, _06444_);
  or _80543_ (_30222_, _30221_, _30220_);
  and _80544_ (_30223_, _30222_, _01317_);
  and _80545_ (_30224_, _30223_, _30217_);
  nor _80546_ (_30226_, \oc8051_golden_model_1.P2 [3], rst);
  nor _80547_ (_30227_, _30226_, _00000_);
  or _80548_ (_43708_, _30227_, _30224_);
  and _80549_ (_30228_, _29671_, \oc8051_golden_model_1.P2 [4]);
  and _80550_ (_30229_, _12768_, _08336_);
  or _80551_ (_30230_, _30229_, _30228_);
  or _80552_ (_30231_, _30230_, _06132_);
  and _80553_ (_30232_, _29695_, \oc8051_golden_model_1.P2 [4]);
  and _80554_ (_30233_, _07847_, \oc8051_golden_model_1.P0 [4]);
  and _80555_ (_30234_, _12778_, \oc8051_golden_model_1.P1 [4]);
  or _80556_ (_30236_, _30234_, _30233_);
  and _80557_ (_30237_, _12773_, \oc8051_golden_model_1.P2 [4]);
  and _80558_ (_30238_, _12780_, \oc8051_golden_model_1.P3 [4]);
  or _80559_ (_30239_, _30238_, _30237_);
  nor _80560_ (_30240_, _30239_, _30236_);
  nand _80561_ (_30241_, _30240_, _12676_);
  and _80562_ (_30242_, _30241_, _12678_);
  and _80563_ (_30243_, _30242_, _12773_);
  or _80564_ (_30244_, _30243_, _30232_);
  and _80565_ (_30245_, _30244_, _06152_);
  and _80566_ (_30247_, _12863_, _12826_);
  or _80567_ (_30248_, _30247_, _12864_);
  and _80568_ (_30249_, _30248_, _12768_);
  or _80569_ (_30250_, _30249_, _30228_);
  or _80570_ (_30251_, _30250_, _06161_);
  and _80571_ (_30252_, _12768_, \oc8051_golden_model_1.ACC [4]);
  or _80572_ (_30253_, _30252_, _30228_);
  and _80573_ (_30254_, _30253_, _07056_);
  and _80574_ (_30255_, _07057_, \oc8051_golden_model_1.P2 [4]);
  or _80575_ (_30256_, _30255_, _06160_);
  or _80576_ (_30258_, _30256_, _30254_);
  and _80577_ (_30259_, _30258_, _06157_);
  and _80578_ (_30260_, _30259_, _30251_);
  or _80579_ (_30261_, _30241_, _12677_);
  and _80580_ (_30262_, _30261_, _12773_);
  or _80581_ (_30263_, _30262_, _30232_);
  and _80582_ (_30264_, _30263_, _06156_);
  or _80583_ (_30265_, _30264_, _06217_);
  or _80584_ (_30266_, _30265_, _30260_);
  or _80585_ (_30267_, _30230_, _07075_);
  and _80586_ (_30269_, _30267_, _30266_);
  or _80587_ (_30270_, _30269_, _06220_);
  or _80588_ (_30271_, _30253_, _06229_);
  and _80589_ (_30272_, _30271_, _06153_);
  and _80590_ (_30273_, _30272_, _30270_);
  or _80591_ (_30274_, _30273_, _30245_);
  and _80592_ (_30275_, _30274_, _06146_);
  nand _80593_ (_30276_, _30241_, _12677_);
  or _80594_ (_30277_, _30232_, _30276_);
  and _80595_ (_30278_, _30263_, _06145_);
  and _80596_ (_30280_, _30278_, _30277_);
  or _80597_ (_30281_, _30280_, _30275_);
  and _80598_ (_30282_, _30281_, _06140_);
  or _80599_ (_30283_, _30242_, _14965_);
  and _80600_ (_30284_, _30283_, _12773_);
  or _80601_ (_30285_, _30284_, _30232_);
  and _80602_ (_30286_, _30285_, _06139_);
  or _80603_ (_30287_, _30286_, _09842_);
  or _80604_ (_30288_, _30287_, _30282_);
  and _80605_ (_30289_, _30288_, _30231_);
  or _80606_ (_30291_, _30289_, _06116_);
  and _80607_ (_30292_, _12768_, _09209_);
  or _80608_ (_30293_, _30228_, _06117_);
  or _80609_ (_30294_, _30293_, _30292_);
  and _80610_ (_30295_, _30294_, _06114_);
  and _80611_ (_30296_, _30295_, _30291_);
  and _80612_ (_30297_, _12918_, \oc8051_golden_model_1.P1 [4]);
  and _80613_ (_30298_, _12916_, \oc8051_golden_model_1.P0 [4]);
  and _80614_ (_30299_, _12920_, \oc8051_golden_model_1.P2 [4]);
  and _80615_ (_30300_, _12922_, \oc8051_golden_model_1.P3 [4]);
  or _80616_ (_30302_, _30300_, _30299_);
  or _80617_ (_30303_, _30302_, _30298_);
  or _80618_ (_30304_, _30303_, _30297_);
  or _80619_ (_30305_, _30304_, _15013_);
  and _80620_ (_30306_, _30305_, _12768_);
  or _80621_ (_30307_, _30306_, _30228_);
  and _80622_ (_30308_, _30307_, _05787_);
  or _80623_ (_30309_, _30308_, _06110_);
  or _80624_ (_30310_, _30309_, _30296_);
  and _80625_ (_30311_, _12768_, _08715_);
  or _80626_ (_30313_, _30311_, _30228_);
  or _80627_ (_30314_, _30313_, _06111_);
  and _80628_ (_30315_, _30314_, _07127_);
  and _80629_ (_30316_, _30315_, _30310_);
  or _80630_ (_30317_, _12826_, _08715_);
  and _80631_ (_30318_, _30317_, _12768_);
  or _80632_ (_30319_, _30318_, _30228_);
  nand _80633_ (_30320_, _12826_, _08715_);
  or _80634_ (_30321_, _30320_, _30228_);
  and _80635_ (_30322_, _30321_, _06297_);
  and _80636_ (_30324_, _30322_, _30319_);
  or _80637_ (_30325_, _30324_, _30316_);
  and _80638_ (_30326_, _30325_, _07125_);
  or _80639_ (_30327_, _12826_, \oc8051_golden_model_1.ACC [4]);
  and _80640_ (_30328_, _30327_, _12768_);
  or _80641_ (_30329_, _30328_, _30228_);
  nand _80642_ (_30330_, _12826_, \oc8051_golden_model_1.ACC [4]);
  or _80643_ (_30331_, _30330_, _30228_);
  and _80644_ (_30332_, _30331_, _06402_);
  and _80645_ (_30333_, _30332_, _30329_);
  or _80646_ (_30335_, _30333_, _30326_);
  and _80647_ (_30336_, _30335_, _07132_);
  or _80648_ (_30337_, _30228_, _12826_);
  and _80649_ (_30338_, _30313_, _06306_);
  and _80650_ (_30339_, _30338_, _30337_);
  or _80651_ (_30340_, _30339_, _30336_);
  and _80652_ (_30341_, _30340_, _07130_);
  and _80653_ (_30342_, _30253_, _06411_);
  and _80654_ (_30343_, _30342_, _30337_);
  or _80655_ (_30344_, _30343_, _06303_);
  or _80656_ (_30346_, _30344_, _30341_);
  or _80657_ (_30347_, _30319_, _08819_);
  and _80658_ (_30348_, _30347_, _08824_);
  and _80659_ (_30349_, _30348_, _30346_);
  and _80660_ (_30350_, _30329_, _06396_);
  or _80661_ (_30351_, _30350_, _06433_);
  or _80662_ (_30352_, _30351_, _30349_);
  or _80663_ (_30353_, _30250_, _06829_);
  and _80664_ (_30354_, _30353_, _05749_);
  and _80665_ (_30355_, _30354_, _30352_);
  and _80666_ (_30357_, _30244_, _05748_);
  or _80667_ (_30358_, _30357_, _06440_);
  or _80668_ (_30359_, _30358_, _30355_);
  nor _80669_ (_30360_, _12979_, _12826_);
  nor _80670_ (_30361_, _30360_, _12980_);
  and _80671_ (_30362_, _30361_, _12768_);
  or _80672_ (_30363_, _30228_, _06444_);
  or _80673_ (_30364_, _30363_, _30362_);
  and _80674_ (_30365_, _30364_, _01317_);
  and _80675_ (_30366_, _30365_, _30359_);
  nor _80676_ (_30368_, \oc8051_golden_model_1.P2 [4], rst);
  nor _80677_ (_30369_, _30368_, _00000_);
  or _80678_ (_43709_, _30369_, _30366_);
  nor _80679_ (_30370_, \oc8051_golden_model_1.P2 [5], rst);
  nor _80680_ (_30371_, _30370_, _00000_);
  and _80681_ (_30372_, _29671_, \oc8051_golden_model_1.P2 [5]);
  and _80682_ (_30373_, _12768_, _08101_);
  or _80683_ (_30374_, _30373_, _30372_);
  or _80684_ (_30375_, _30374_, _06132_);
  and _80685_ (_30376_, _12865_, _12818_);
  or _80686_ (_30378_, _30376_, _12866_);
  and _80687_ (_30379_, _30378_, _12768_);
  or _80688_ (_30380_, _30379_, _30372_);
  or _80689_ (_30381_, _30380_, _06161_);
  and _80690_ (_30382_, _12768_, \oc8051_golden_model_1.ACC [5]);
  or _80691_ (_30383_, _30382_, _30372_);
  and _80692_ (_30384_, _30383_, _07056_);
  and _80693_ (_30385_, _07057_, \oc8051_golden_model_1.P2 [5]);
  or _80694_ (_30386_, _30385_, _06160_);
  or _80695_ (_30387_, _30386_, _30384_);
  and _80696_ (_30389_, _30387_, _06157_);
  and _80697_ (_30390_, _30389_, _30381_);
  and _80698_ (_30391_, _29695_, \oc8051_golden_model_1.P2 [5]);
  and _80699_ (_30392_, _07847_, \oc8051_golden_model_1.P0 [5]);
  and _80700_ (_30393_, _12773_, \oc8051_golden_model_1.P2 [5]);
  or _80701_ (_30394_, _30393_, _30392_);
  and _80702_ (_30395_, _12778_, \oc8051_golden_model_1.P1 [5]);
  and _80703_ (_30396_, _12780_, \oc8051_golden_model_1.P3 [5]);
  or _80704_ (_30397_, _30396_, _30395_);
  or _80705_ (_30398_, _30397_, _30394_);
  or _80706_ (_30400_, _15123_, _30398_);
  and _80707_ (_30401_, _30400_, _12773_);
  or _80708_ (_30402_, _30401_, _30391_);
  and _80709_ (_30403_, _30402_, _06156_);
  or _80710_ (_30404_, _30403_, _06217_);
  or _80711_ (_30405_, _30404_, _30390_);
  or _80712_ (_30406_, _30374_, _07075_);
  and _80713_ (_30407_, _30406_, _30405_);
  or _80714_ (_30408_, _30407_, _06220_);
  or _80715_ (_30409_, _30383_, _06229_);
  and _80716_ (_30411_, _30409_, _06153_);
  and _80717_ (_30412_, _30411_, _30408_);
  or _80718_ (_30413_, _30398_, _12611_);
  and _80719_ (_30414_, _30413_, _15103_);
  and _80720_ (_30415_, _30414_, _12773_);
  or _80721_ (_30416_, _30415_, _30391_);
  and _80722_ (_30417_, _30416_, _06152_);
  or _80723_ (_30418_, _30417_, _06145_);
  or _80724_ (_30419_, _30418_, _30412_);
  nand _80725_ (_30420_, _30413_, _12612_);
  or _80726_ (_30421_, _30391_, _30420_);
  and _80727_ (_30422_, _30421_, _30402_);
  or _80728_ (_30423_, _30422_, _06146_);
  and _80729_ (_30424_, _30423_, _06140_);
  and _80730_ (_30425_, _30424_, _30419_);
  or _80731_ (_30426_, _30414_, _15154_);
  and _80732_ (_30427_, _30426_, _12773_);
  or _80733_ (_30428_, _30427_, _30391_);
  and _80734_ (_30429_, _30428_, _06139_);
  or _80735_ (_30430_, _30429_, _09842_);
  or _80736_ (_30433_, _30430_, _30425_);
  and _80737_ (_30434_, _30433_, _30375_);
  or _80738_ (_30435_, _30434_, _06116_);
  and _80739_ (_30436_, _12768_, _09208_);
  or _80740_ (_30437_, _30372_, _06117_);
  or _80741_ (_30438_, _30437_, _30436_);
  and _80742_ (_30439_, _30438_, _06114_);
  and _80743_ (_30440_, _30439_, _30435_);
  and _80744_ (_30441_, _12918_, \oc8051_golden_model_1.P1 [5]);
  and _80745_ (_30442_, _12916_, \oc8051_golden_model_1.P0 [5]);
  and _80746_ (_30444_, _12920_, \oc8051_golden_model_1.P2 [5]);
  and _80747_ (_30445_, _12922_, \oc8051_golden_model_1.P3 [5]);
  or _80748_ (_30446_, _30445_, _30444_);
  or _80749_ (_30447_, _30446_, _30442_);
  or _80750_ (_30448_, _30447_, _30441_);
  or _80751_ (_30449_, _30448_, _15203_);
  and _80752_ (_30450_, _30449_, _12768_);
  or _80753_ (_30451_, _30450_, _30372_);
  and _80754_ (_30452_, _30451_, _05787_);
  or _80755_ (_30453_, _30452_, _06110_);
  or _80756_ (_30455_, _30453_, _30440_);
  and _80757_ (_30456_, _12768_, _08736_);
  or _80758_ (_30457_, _30456_, _30372_);
  or _80759_ (_30458_, _30457_, _06111_);
  and _80760_ (_30459_, _30458_, _07127_);
  and _80761_ (_30460_, _30459_, _30455_);
  or _80762_ (_30461_, _12818_, _08736_);
  and _80763_ (_30462_, _30461_, _12768_);
  or _80764_ (_30463_, _30462_, _30372_);
  nand _80765_ (_30464_, _12818_, _08736_);
  or _80766_ (_30466_, _30464_, _30372_);
  and _80767_ (_30467_, _30466_, _06297_);
  and _80768_ (_30468_, _30467_, _30463_);
  or _80769_ (_30469_, _30468_, _30460_);
  and _80770_ (_30470_, _30469_, _07125_);
  or _80771_ (_30471_, _12818_, \oc8051_golden_model_1.ACC [5]);
  and _80772_ (_30472_, _30471_, _12768_);
  or _80773_ (_30473_, _30472_, _30372_);
  nand _80774_ (_30474_, _12818_, \oc8051_golden_model_1.ACC [5]);
  or _80775_ (_30475_, _30474_, _30372_);
  and _80776_ (_30477_, _30475_, _06402_);
  and _80777_ (_30478_, _30477_, _30473_);
  or _80778_ (_30479_, _30478_, _30470_);
  and _80779_ (_30480_, _30479_, _07132_);
  or _80780_ (_30481_, _30372_, _12818_);
  and _80781_ (_30482_, _30457_, _06306_);
  and _80782_ (_30483_, _30482_, _30481_);
  or _80783_ (_30484_, _30483_, _30480_);
  and _80784_ (_30485_, _30484_, _07130_);
  and _80785_ (_30486_, _30383_, _06411_);
  and _80786_ (_30488_, _30486_, _30481_);
  or _80787_ (_30489_, _30488_, _06303_);
  or _80788_ (_30490_, _30489_, _30485_);
  or _80789_ (_30491_, _30463_, _08819_);
  and _80790_ (_30492_, _30491_, _08824_);
  and _80791_ (_30493_, _30492_, _30490_);
  and _80792_ (_30494_, _30473_, _06396_);
  or _80793_ (_30495_, _30494_, _06433_);
  or _80794_ (_30496_, _30495_, _30493_);
  or _80795_ (_30497_, _30380_, _06829_);
  and _80796_ (_30499_, _30497_, _05749_);
  and _80797_ (_30500_, _30499_, _30496_);
  and _80798_ (_30501_, _30416_, _05748_);
  or _80799_ (_30502_, _30501_, _06440_);
  or _80800_ (_30503_, _30502_, _30500_);
  nor _80801_ (_30504_, _12980_, _12818_);
  nor _80802_ (_30505_, _30504_, _12981_);
  and _80803_ (_30506_, _30505_, _12768_);
  or _80804_ (_30507_, _30372_, _06444_);
  or _80805_ (_30508_, _30507_, _30506_);
  and _80806_ (_30510_, _30508_, _01317_);
  and _80807_ (_30511_, _30510_, _30503_);
  or _80808_ (_43710_, _30511_, _30371_);
  and _80809_ (_30512_, _29671_, \oc8051_golden_model_1.P2 [6]);
  and _80810_ (_30513_, _12768_, _08012_);
  or _80811_ (_30514_, _30513_, _30512_);
  or _80812_ (_30515_, _30514_, _06132_);
  and _80813_ (_30516_, _29695_, \oc8051_golden_model_1.P2 [6]);
  and _80814_ (_30517_, _07847_, \oc8051_golden_model_1.P0 [6]);
  and _80815_ (_30518_, _12773_, \oc8051_golden_model_1.P2 [6]);
  or _80816_ (_30520_, _30518_, _30517_);
  and _80817_ (_30521_, _12778_, \oc8051_golden_model_1.P1 [6]);
  and _80818_ (_30522_, _12780_, \oc8051_golden_model_1.P3 [6]);
  or _80819_ (_30523_, _30522_, _30521_);
  or _80820_ (_30524_, _30523_, _30520_);
  or _80821_ (_30525_, _30524_, _12579_);
  and _80822_ (_30526_, _30525_, _15296_);
  and _80823_ (_30527_, _30526_, _12773_);
  or _80824_ (_30528_, _30527_, _30516_);
  and _80825_ (_30529_, _30528_, _06152_);
  and _80826_ (_30531_, _12867_, _12810_);
  or _80827_ (_30532_, _30531_, _12868_);
  and _80828_ (_30533_, _30532_, _12768_);
  or _80829_ (_30534_, _30533_, _30512_);
  or _80830_ (_30535_, _30534_, _06161_);
  and _80831_ (_30536_, _12768_, \oc8051_golden_model_1.ACC [6]);
  or _80832_ (_30537_, _30536_, _30512_);
  and _80833_ (_30538_, _30537_, _07056_);
  and _80834_ (_30539_, _07057_, \oc8051_golden_model_1.P2 [6]);
  or _80835_ (_30540_, _30539_, _06160_);
  or _80836_ (_30542_, _30540_, _30538_);
  and _80837_ (_30543_, _30542_, _06157_);
  and _80838_ (_30544_, _30543_, _30535_);
  or _80839_ (_30545_, _15316_, _30524_);
  and _80840_ (_30546_, _30545_, _12773_);
  or _80841_ (_30547_, _30546_, _30516_);
  and _80842_ (_30548_, _30547_, _06156_);
  or _80843_ (_30549_, _30548_, _06217_);
  or _80844_ (_30550_, _30549_, _30544_);
  or _80845_ (_30551_, _30514_, _07075_);
  and _80846_ (_30553_, _30551_, _30550_);
  or _80847_ (_30554_, _30553_, _06220_);
  or _80848_ (_30555_, _30537_, _06229_);
  and _80849_ (_30556_, _30555_, _06153_);
  and _80850_ (_30557_, _30556_, _30554_);
  or _80851_ (_30558_, _30557_, _30529_);
  and _80852_ (_30559_, _30558_, _06146_);
  nand _80853_ (_30560_, _30525_, _12580_);
  or _80854_ (_30561_, _30516_, _30560_);
  and _80855_ (_30562_, _30547_, _06145_);
  and _80856_ (_30564_, _30562_, _30561_);
  or _80857_ (_30565_, _30564_, _30559_);
  and _80858_ (_30566_, _30565_, _06140_);
  or _80859_ (_30567_, _30526_, _15347_);
  and _80860_ (_30568_, _30567_, _12773_);
  or _80861_ (_30569_, _30568_, _30516_);
  and _80862_ (_30570_, _30569_, _06139_);
  or _80863_ (_30571_, _30570_, _09842_);
  or _80864_ (_30572_, _30571_, _30566_);
  and _80865_ (_30573_, _30572_, _30515_);
  or _80866_ (_30575_, _30573_, _06116_);
  and _80867_ (_30576_, _12768_, _09207_);
  or _80868_ (_30577_, _30512_, _06117_);
  or _80869_ (_30578_, _30577_, _30576_);
  and _80870_ (_30579_, _30578_, _06114_);
  and _80871_ (_30580_, _30579_, _30575_);
  and _80872_ (_30581_, _12916_, \oc8051_golden_model_1.P0 [6]);
  and _80873_ (_30582_, _12918_, \oc8051_golden_model_1.P1 [6]);
  and _80874_ (_30583_, _12920_, \oc8051_golden_model_1.P2 [6]);
  and _80875_ (_30584_, _12922_, \oc8051_golden_model_1.P3 [6]);
  or _80876_ (_30586_, _30584_, _30583_);
  or _80877_ (_30587_, _30586_, _30582_);
  or _80878_ (_30588_, _30587_, _30581_);
  or _80879_ (_30589_, _30588_, _15395_);
  and _80880_ (_30590_, _30589_, _12768_);
  or _80881_ (_30591_, _30590_, _30512_);
  and _80882_ (_30592_, _30591_, _05787_);
  or _80883_ (_30593_, _30592_, _06110_);
  or _80884_ (_30594_, _30593_, _30580_);
  and _80885_ (_30595_, _12768_, _15402_);
  or _80886_ (_30597_, _30595_, _30512_);
  or _80887_ (_30598_, _30597_, _06111_);
  and _80888_ (_30599_, _30598_, _07127_);
  and _80889_ (_30600_, _30599_, _30594_);
  or _80890_ (_30601_, _12810_, _15402_);
  and _80891_ (_30602_, _30601_, _12768_);
  or _80892_ (_30603_, _30602_, _30512_);
  nand _80893_ (_30604_, _12810_, _15402_);
  or _80894_ (_30605_, _30604_, _30512_);
  and _80895_ (_30606_, _30605_, _06297_);
  and _80896_ (_30608_, _30606_, _30603_);
  or _80897_ (_30609_, _30608_, _06402_);
  or _80898_ (_30610_, _30609_, _30600_);
  or _80899_ (_30611_, _12810_, \oc8051_golden_model_1.ACC [6]);
  nand _80900_ (_30612_, _12810_, \oc8051_golden_model_1.ACC [6]);
  and _80901_ (_30613_, _30612_, _30611_);
  and _80902_ (_30614_, _30613_, _12768_);
  or _80903_ (_30615_, _30512_, _07125_);
  or _80904_ (_30616_, _30615_, _30614_);
  and _80905_ (_30617_, _30616_, _07132_);
  and _80906_ (_30619_, _30617_, _30610_);
  or _80907_ (_30620_, _30512_, _12810_);
  and _80908_ (_30621_, _30597_, _06306_);
  and _80909_ (_30622_, _30621_, _30620_);
  or _80910_ (_30623_, _30622_, _30619_);
  and _80911_ (_30624_, _30623_, _07130_);
  and _80912_ (_30625_, _30537_, _06411_);
  and _80913_ (_30626_, _30625_, _30620_);
  or _80914_ (_30627_, _30626_, _06303_);
  or _80915_ (_30628_, _30627_, _30624_);
  or _80916_ (_30630_, _30603_, _08819_);
  and _80917_ (_30631_, _30630_, _08824_);
  and _80918_ (_30632_, _30631_, _30628_);
  and _80919_ (_30633_, _30611_, _12768_);
  or _80920_ (_30634_, _30633_, _30512_);
  and _80921_ (_30635_, _30634_, _06396_);
  or _80922_ (_30636_, _30635_, _06433_);
  or _80923_ (_30637_, _30636_, _30632_);
  or _80924_ (_30638_, _30534_, _06829_);
  and _80925_ (_30639_, _30638_, _05749_);
  and _80926_ (_30641_, _30639_, _30637_);
  and _80927_ (_30642_, _30528_, _05748_);
  or _80928_ (_30643_, _30642_, _06440_);
  or _80929_ (_30644_, _30643_, _30641_);
  or _80930_ (_30645_, _12981_, _12810_);
  and _80931_ (_30646_, _30645_, _12982_);
  and _80932_ (_30647_, _30646_, _12768_);
  or _80933_ (_30648_, _30512_, _06444_);
  or _80934_ (_30649_, _30648_, _30647_);
  and _80935_ (_30650_, _30649_, _01317_);
  and _80936_ (_30652_, _30650_, _30644_);
  nor _80937_ (_30653_, \oc8051_golden_model_1.P2 [6], rst);
  nor _80938_ (_30654_, _30653_, _00000_);
  or _80939_ (_43711_, _30654_, _30652_);
  and _80940_ (_30655_, _12996_, \oc8051_golden_model_1.P3 [0]);
  and _80941_ (_30656_, _29705_, _12780_);
  or _80942_ (_30657_, _30656_, _30655_);
  or _80943_ (_30658_, _30657_, _06157_);
  and _80944_ (_30659_, _12991_, \oc8051_golden_model_1.P3 [0]);
  nor _80945_ (_30660_, _12858_, _12991_);
  or _80946_ (_30662_, _30660_, _30659_);
  and _80947_ (_30663_, _30662_, _06160_);
  and _80948_ (_30664_, _07057_, \oc8051_golden_model_1.P3 [0]);
  and _80949_ (_30665_, _12797_, \oc8051_golden_model_1.ACC [0]);
  or _80950_ (_30666_, _30665_, _30659_);
  and _80951_ (_30667_, _30666_, _07056_);
  or _80952_ (_30668_, _30667_, _30664_);
  and _80953_ (_30669_, _30668_, _06161_);
  or _80954_ (_30670_, _30669_, _06156_);
  or _80955_ (_30671_, _30670_, _30663_);
  and _80956_ (_30673_, _30671_, _30658_);
  and _80957_ (_30674_, _30673_, _07075_);
  and _80958_ (_30675_, _12797_, _07049_);
  or _80959_ (_30676_, _30675_, _30659_);
  and _80960_ (_30677_, _30676_, _06217_);
  or _80961_ (_30678_, _30677_, _06220_);
  or _80962_ (_30679_, _30678_, _30674_);
  or _80963_ (_30680_, _30666_, _06229_);
  and _80964_ (_30681_, _30680_, _06153_);
  and _80965_ (_30682_, _30681_, _30679_);
  and _80966_ (_30684_, _30659_, _06152_);
  or _80967_ (_30685_, _30684_, _06145_);
  or _80968_ (_30686_, _30685_, _30682_);
  or _80969_ (_30687_, _30662_, _06146_);
  and _80970_ (_30688_, _30687_, _06140_);
  and _80971_ (_30689_, _30688_, _30686_);
  or _80972_ (_30690_, _30655_, _14170_);
  and _80973_ (_30691_, _30690_, _06139_);
  and _80974_ (_30692_, _30691_, _30657_);
  or _80975_ (_30693_, _30692_, _09842_);
  or _80976_ (_30695_, _30693_, _30689_);
  or _80977_ (_30696_, _30676_, _06132_);
  and _80978_ (_30697_, _30696_, _30695_);
  or _80979_ (_30698_, _30697_, _06116_);
  and _80980_ (_30699_, _12797_, _09160_);
  or _80981_ (_30700_, _30659_, _06117_);
  or _80982_ (_30701_, _30700_, _30699_);
  and _80983_ (_30702_, _30701_, _06114_);
  and _80984_ (_30703_, _30702_, _30698_);
  and _80985_ (_30704_, _29746_, _12797_);
  or _80986_ (_30706_, _30704_, _30659_);
  and _80987_ (_30707_, _30706_, _05787_);
  or _80988_ (_30708_, _30707_, _06110_);
  or _80989_ (_30709_, _30708_, _30703_);
  and _80990_ (_30710_, _12797_, _08708_);
  or _80991_ (_30711_, _30710_, _30659_);
  or _80992_ (_30712_, _30711_, _06111_);
  and _80993_ (_30713_, _30712_, _07127_);
  and _80994_ (_30714_, _30713_, _30709_);
  and _80995_ (_30715_, _29752_, _12797_);
  or _80996_ (_30717_, _30715_, _30659_);
  or _80997_ (_30718_, _30659_, _29754_);
  and _80998_ (_30719_, _30718_, _06297_);
  and _80999_ (_30720_, _30719_, _30717_);
  or _81000_ (_30721_, _30720_, _06402_);
  or _81001_ (_30722_, _30721_, _30714_);
  and _81002_ (_30723_, _29675_, _12797_);
  or _81003_ (_30724_, _30659_, _07125_);
  or _81004_ (_30725_, _30724_, _30723_);
  and _81005_ (_30726_, _30725_, _07132_);
  and _81006_ (_30728_, _30726_, _30722_);
  nand _81007_ (_30729_, _30711_, _06306_);
  nor _81008_ (_30730_, _30729_, _30660_);
  or _81009_ (_30731_, _30730_, _30728_);
  and _81010_ (_30732_, _30731_, _07130_);
  or _81011_ (_30733_, _30659_, _12858_);
  and _81012_ (_30734_, _30666_, _06411_);
  and _81013_ (_30735_, _30734_, _30733_);
  or _81014_ (_30736_, _30735_, _06303_);
  or _81015_ (_30737_, _30736_, _30732_);
  or _81016_ (_30739_, _30717_, _08819_);
  and _81017_ (_30740_, _30739_, _08824_);
  and _81018_ (_30741_, _30740_, _30737_);
  and _81019_ (_30742_, _29673_, _12797_);
  or _81020_ (_30743_, _30742_, _30659_);
  and _81021_ (_30744_, _30743_, _06396_);
  or _81022_ (_30745_, _30744_, _06433_);
  or _81023_ (_30746_, _30745_, _30741_);
  or _81024_ (_30747_, _30662_, _06829_);
  and _81025_ (_30748_, _30747_, _05749_);
  and _81026_ (_30750_, _30748_, _30746_);
  and _81027_ (_30751_, _30659_, _05748_);
  or _81028_ (_30752_, _30751_, _06440_);
  or _81029_ (_30753_, _30752_, _30750_);
  or _81030_ (_30754_, _30662_, _06444_);
  and _81031_ (_30755_, _30754_, _01317_);
  and _81032_ (_30756_, _30755_, _30753_);
  nor _81033_ (_30757_, \oc8051_golden_model_1.P3 [0], rst);
  nor _81034_ (_30758_, _30757_, _00000_);
  or _81035_ (_43713_, _30758_, _30756_);
  nor _81036_ (_30760_, \oc8051_golden_model_1.P3 [1], rst);
  nor _81037_ (_30761_, _30760_, _00000_);
  or _81038_ (_30762_, _29883_, _12991_);
  or _81039_ (_30763_, _12797_, \oc8051_golden_model_1.P3 [1]);
  and _81040_ (_30764_, _30763_, _05787_);
  and _81041_ (_30765_, _30764_, _30762_);
  and _81042_ (_30766_, _29814_, _12780_);
  and _81043_ (_30767_, _30766_, _29813_);
  and _81044_ (_30768_, _12996_, \oc8051_golden_model_1.P3 [1]);
  or _81045_ (_30769_, _30768_, _06146_);
  or _81046_ (_30771_, _30769_, _30767_);
  and _81047_ (_30772_, _29823_, _12797_);
  not _81048_ (_30773_, _30772_);
  and _81049_ (_30774_, _30773_, _30763_);
  or _81050_ (_30775_, _30774_, _06161_);
  nand _81051_ (_30776_, _12797_, _05887_);
  and _81052_ (_30777_, _30776_, _30763_);
  and _81053_ (_30778_, _30777_, _07056_);
  and _81054_ (_30779_, _07057_, \oc8051_golden_model_1.P3 [1]);
  or _81055_ (_30780_, _30779_, _06160_);
  or _81056_ (_30782_, _30780_, _30778_);
  and _81057_ (_30783_, _30782_, _06157_);
  and _81058_ (_30784_, _30783_, _30775_);
  or _81059_ (_30785_, _30768_, _06217_);
  or _81060_ (_30786_, _30785_, _30766_);
  and _81061_ (_30787_, _30786_, _13860_);
  or _81062_ (_30788_, _30787_, _30784_);
  and _81063_ (_30789_, _12991_, \oc8051_golden_model_1.P3 [1]);
  and _81064_ (_30790_, _12797_, _07306_);
  or _81065_ (_30791_, _30790_, _30789_);
  or _81066_ (_30793_, _30791_, _07075_);
  and _81067_ (_30794_, _30793_, _30788_);
  or _81068_ (_30795_, _30794_, _06220_);
  or _81069_ (_30796_, _30777_, _06229_);
  and _81070_ (_30797_, _30796_, _06153_);
  and _81071_ (_30798_, _30797_, _30795_);
  and _81072_ (_30799_, _29851_, _12780_);
  or _81073_ (_30800_, _30799_, _30768_);
  and _81074_ (_30801_, _30800_, _06152_);
  or _81075_ (_30802_, _30801_, _06145_);
  or _81076_ (_30804_, _30802_, _30798_);
  and _81077_ (_30805_, _30804_, _30771_);
  and _81078_ (_30806_, _30805_, _06140_);
  and _81079_ (_30807_, _29860_, _12780_);
  or _81080_ (_30808_, _30768_, _30807_);
  and _81081_ (_30809_, _30808_, _06139_);
  or _81082_ (_30810_, _30809_, _09842_);
  or _81083_ (_30811_, _30810_, _30806_);
  or _81084_ (_30812_, _30791_, _06132_);
  and _81085_ (_30813_, _30812_, _30811_);
  or _81086_ (_30815_, _30813_, _06116_);
  and _81087_ (_30816_, _12797_, _09115_);
  or _81088_ (_30817_, _30789_, _06117_);
  or _81089_ (_30818_, _30817_, _30816_);
  and _81090_ (_30819_, _30818_, _06114_);
  and _81091_ (_30820_, _30819_, _30815_);
  or _81092_ (_30821_, _30820_, _30765_);
  and _81093_ (_30822_, _30821_, _06298_);
  and _81094_ (_30823_, _29898_, _29893_);
  or _81095_ (_30824_, _30823_, _12991_);
  and _81096_ (_30826_, _30824_, _06297_);
  nand _81097_ (_30827_, _12797_, _06945_);
  and _81098_ (_30828_, _30827_, _06110_);
  or _81099_ (_30829_, _30828_, _30826_);
  and _81100_ (_30830_, _30829_, _30763_);
  or _81101_ (_30831_, _30830_, _30822_);
  and _81102_ (_30832_, _30831_, _07125_);
  and _81103_ (_30833_, _29909_, _29905_);
  or _81104_ (_30834_, _30833_, _12991_);
  and _81105_ (_30835_, _30763_, _06402_);
  and _81106_ (_30837_, _30835_, _30834_);
  or _81107_ (_30838_, _30837_, _30832_);
  and _81108_ (_30839_, _30838_, _07132_);
  or _81109_ (_30840_, _29896_, _12991_);
  and _81110_ (_30841_, _30763_, _06306_);
  and _81111_ (_30842_, _30841_, _30840_);
  or _81112_ (_30843_, _30842_, _30839_);
  and _81113_ (_30844_, _30843_, _07130_);
  or _81114_ (_30845_, _30789_, _12850_);
  and _81115_ (_30846_, _30777_, _06411_);
  and _81116_ (_30848_, _30846_, _30845_);
  or _81117_ (_30849_, _30848_, _30844_);
  and _81118_ (_30850_, _30849_, _06397_);
  or _81119_ (_30851_, _30827_, _12850_);
  and _81120_ (_30852_, _30763_, _06303_);
  and _81121_ (_30853_, _30852_, _30851_);
  or _81122_ (_30854_, _30776_, _12850_);
  and _81123_ (_30855_, _30763_, _06396_);
  and _81124_ (_30856_, _30855_, _30854_);
  or _81125_ (_30857_, _30856_, _06433_);
  or _81126_ (_30859_, _30857_, _30853_);
  or _81127_ (_30860_, _30859_, _30850_);
  or _81128_ (_30861_, _30774_, _06829_);
  and _81129_ (_30862_, _30861_, _05749_);
  and _81130_ (_30863_, _30862_, _30860_);
  and _81131_ (_30864_, _30800_, _05748_);
  or _81132_ (_30865_, _30864_, _06440_);
  or _81133_ (_30866_, _30865_, _30863_);
  or _81134_ (_30867_, _30789_, _06444_);
  or _81135_ (_30868_, _30867_, _30772_);
  and _81136_ (_30870_, _30868_, _01317_);
  and _81137_ (_30871_, _30870_, _30866_);
  or _81138_ (_43714_, _30871_, _30761_);
  and _81139_ (_30872_, _12991_, \oc8051_golden_model_1.P3 [2]);
  and _81140_ (_30873_, _29954_, _12797_);
  or _81141_ (_30874_, _30873_, _30872_);
  or _81142_ (_30875_, _30874_, _06161_);
  and _81143_ (_30876_, _12797_, \oc8051_golden_model_1.ACC [2]);
  or _81144_ (_30877_, _30876_, _30872_);
  and _81145_ (_30878_, _30877_, _07056_);
  and _81146_ (_30880_, _07057_, \oc8051_golden_model_1.P3 [2]);
  or _81147_ (_30881_, _30880_, _06160_);
  or _81148_ (_30882_, _30881_, _30878_);
  and _81149_ (_30883_, _30882_, _06157_);
  and _81150_ (_30884_, _30883_, _30875_);
  and _81151_ (_30885_, _12996_, \oc8051_golden_model_1.P3 [2]);
  and _81152_ (_30886_, _29976_, _12780_);
  or _81153_ (_30887_, _30886_, _30885_);
  and _81154_ (_30888_, _30887_, _06156_);
  or _81155_ (_30889_, _30888_, _06217_);
  or _81156_ (_30891_, _30889_, _30884_);
  and _81157_ (_30892_, _12797_, _07708_);
  or _81158_ (_30893_, _30892_, _30872_);
  or _81159_ (_30894_, _30893_, _07075_);
  and _81160_ (_30895_, _30894_, _30891_);
  or _81161_ (_30896_, _30895_, _06220_);
  or _81162_ (_30897_, _30877_, _06229_);
  and _81163_ (_30898_, _30897_, _06153_);
  and _81164_ (_30899_, _30898_, _30896_);
  and _81165_ (_30900_, _29992_, _12780_);
  or _81166_ (_30902_, _30900_, _30885_);
  and _81167_ (_30903_, _30902_, _06152_);
  or _81168_ (_30904_, _30903_, _06145_);
  or _81169_ (_30905_, _30904_, _30899_);
  or _81170_ (_30906_, _30885_, _29999_);
  and _81171_ (_30907_, _30906_, _30887_);
  or _81172_ (_30908_, _30907_, _06146_);
  and _81173_ (_30909_, _30908_, _06140_);
  and _81174_ (_30910_, _30909_, _30905_);
  and _81175_ (_30911_, _30005_, _12780_);
  or _81176_ (_30913_, _30911_, _30885_);
  and _81177_ (_30914_, _30913_, _06139_);
  or _81178_ (_30915_, _30914_, _09842_);
  or _81179_ (_30916_, _30915_, _30910_);
  or _81180_ (_30917_, _30893_, _06132_);
  and _81181_ (_30918_, _30917_, _30916_);
  or _81182_ (_30919_, _30918_, _06116_);
  and _81183_ (_30920_, _12797_, _09211_);
  or _81184_ (_30921_, _30872_, _06117_);
  or _81185_ (_30922_, _30921_, _30920_);
  and _81186_ (_30924_, _30922_, _06114_);
  and _81187_ (_30925_, _30924_, _30919_);
  and _81188_ (_30926_, _30029_, _12797_);
  or _81189_ (_30927_, _30926_, _30872_);
  and _81190_ (_30928_, _30927_, _05787_);
  or _81191_ (_30929_, _30928_, _06110_);
  or _81192_ (_30930_, _30929_, _30925_);
  and _81193_ (_30931_, _12797_, _08768_);
  or _81194_ (_30932_, _30931_, _30872_);
  or _81195_ (_30933_, _30932_, _06111_);
  and _81196_ (_30935_, _30933_, _07127_);
  and _81197_ (_30936_, _30935_, _30930_);
  and _81198_ (_30937_, _29945_, _12797_);
  or _81199_ (_30938_, _30937_, _30872_);
  or _81200_ (_30939_, _30872_, _29948_);
  and _81201_ (_30940_, _30939_, _06297_);
  and _81202_ (_30941_, _30940_, _30938_);
  or _81203_ (_30942_, _30941_, _30936_);
  and _81204_ (_30943_, _30942_, _07125_);
  and _81205_ (_30944_, _30043_, _12797_);
  or _81206_ (_30946_, _30944_, _30872_);
  or _81207_ (_30947_, _30872_, _30046_);
  and _81208_ (_30948_, _30947_, _06402_);
  and _81209_ (_30949_, _30948_, _30946_);
  or _81210_ (_30950_, _30949_, _30943_);
  and _81211_ (_30951_, _30950_, _07132_);
  or _81212_ (_30952_, _30872_, _12842_);
  and _81213_ (_30953_, _30932_, _06306_);
  and _81214_ (_30954_, _30953_, _30952_);
  or _81215_ (_30955_, _30954_, _30951_);
  and _81216_ (_30957_, _30955_, _07130_);
  and _81217_ (_30958_, _30877_, _06411_);
  and _81218_ (_30959_, _30958_, _30952_);
  or _81219_ (_30960_, _30959_, _06303_);
  or _81220_ (_30961_, _30960_, _30957_);
  or _81221_ (_30962_, _30938_, _08819_);
  and _81222_ (_30963_, _30962_, _08824_);
  and _81223_ (_30964_, _30963_, _30961_);
  and _81224_ (_30965_, _30946_, _06396_);
  or _81225_ (_30966_, _30965_, _06433_);
  or _81226_ (_30968_, _30966_, _30964_);
  or _81227_ (_30969_, _30874_, _06829_);
  and _81228_ (_30970_, _30969_, _05749_);
  and _81229_ (_30971_, _30970_, _30968_);
  and _81230_ (_30972_, _30902_, _05748_);
  or _81231_ (_30973_, _30972_, _06440_);
  or _81232_ (_30974_, _30973_, _30971_);
  and _81233_ (_30975_, _30077_, _12797_);
  or _81234_ (_30976_, _30872_, _06444_);
  or _81235_ (_30977_, _30976_, _30975_);
  and _81236_ (_30979_, _30977_, _01317_);
  and _81237_ (_30980_, _30979_, _30974_);
  nor _81238_ (_30981_, \oc8051_golden_model_1.P3 [2], rst);
  nor _81239_ (_30982_, _30981_, _00000_);
  or _81240_ (_43715_, _30982_, _30980_);
  and _81241_ (_30983_, _12991_, \oc8051_golden_model_1.P3 [3]);
  and _81242_ (_30984_, _12797_, _07544_);
  or _81243_ (_30985_, _30984_, _30983_);
  or _81244_ (_30986_, _30985_, _06132_);
  and _81245_ (_30987_, _12996_, \oc8051_golden_model_1.P3 [3]);
  and _81246_ (_30989_, _30100_, _12780_);
  or _81247_ (_30990_, _30989_, _30987_);
  and _81248_ (_30991_, _30990_, _06152_);
  and _81249_ (_30992_, _30106_, _12797_);
  or _81250_ (_30993_, _30992_, _30983_);
  or _81251_ (_30994_, _30993_, _06161_);
  and _81252_ (_30995_, _12797_, \oc8051_golden_model_1.ACC [3]);
  or _81253_ (_30996_, _30995_, _30983_);
  and _81254_ (_30997_, _30996_, _07056_);
  and _81255_ (_30998_, _07057_, \oc8051_golden_model_1.P3 [3]);
  or _81256_ (_31000_, _30998_, _06160_);
  or _81257_ (_31001_, _31000_, _30997_);
  and _81258_ (_31002_, _31001_, _06157_);
  and _81259_ (_31003_, _31002_, _30994_);
  and _81260_ (_31004_, _30119_, _12780_);
  or _81261_ (_31005_, _31004_, _30987_);
  and _81262_ (_31006_, _31005_, _06156_);
  or _81263_ (_31007_, _31006_, _06217_);
  or _81264_ (_31008_, _31007_, _31003_);
  or _81265_ (_31009_, _30985_, _07075_);
  and _81266_ (_31011_, _31009_, _31008_);
  or _81267_ (_31012_, _31011_, _06220_);
  or _81268_ (_31013_, _30996_, _06229_);
  and _81269_ (_31014_, _31013_, _06153_);
  and _81270_ (_31015_, _31014_, _31012_);
  or _81271_ (_31016_, _31015_, _30991_);
  and _81272_ (_31017_, _31016_, _06146_);
  or _81273_ (_31018_, _30987_, _30134_);
  and _81274_ (_31019_, _31005_, _06145_);
  and _81275_ (_31020_, _31019_, _31018_);
  or _81276_ (_31022_, _31020_, _31017_);
  and _81277_ (_31023_, _31022_, _06140_);
  and _81278_ (_31024_, _30141_, _12780_);
  or _81279_ (_31025_, _31024_, _30987_);
  and _81280_ (_31026_, _31025_, _06139_);
  or _81281_ (_31027_, _31026_, _09842_);
  or _81282_ (_31028_, _31027_, _31023_);
  and _81283_ (_31029_, _31028_, _30986_);
  or _81284_ (_31030_, _31029_, _06116_);
  and _81285_ (_31031_, _12797_, _09210_);
  or _81286_ (_31033_, _30983_, _06117_);
  or _81287_ (_31034_, _31033_, _31031_);
  and _81288_ (_31035_, _31034_, _06114_);
  and _81289_ (_31036_, _31035_, _31030_);
  and _81290_ (_31037_, _30163_, _12797_);
  or _81291_ (_31038_, _31037_, _30983_);
  and _81292_ (_31039_, _31038_, _05787_);
  or _81293_ (_31040_, _31039_, _11136_);
  or _81294_ (_31041_, _31040_, _31036_);
  and _81295_ (_31042_, _30178_, _30175_);
  and _81296_ (_31044_, _31042_, _12797_);
  or _81297_ (_31045_, _30983_, _07127_);
  or _81298_ (_31046_, _31045_, _31044_);
  and _81299_ (_31047_, _12797_, _08712_);
  or _81300_ (_31048_, _31047_, _30983_);
  or _81301_ (_31049_, _31048_, _06111_);
  and _81302_ (_31050_, _31049_, _07125_);
  and _81303_ (_31051_, _31050_, _31046_);
  and _81304_ (_31052_, _31051_, _31041_);
  and _81305_ (_31053_, _30188_, _30185_);
  and _81306_ (_31055_, _31053_, _12797_);
  or _81307_ (_31056_, _31055_, _30983_);
  and _81308_ (_31057_, _31056_, _06402_);
  or _81309_ (_31058_, _31057_, _31052_);
  and _81310_ (_31059_, _31058_, _07132_);
  or _81311_ (_31060_, _30983_, _12834_);
  and _81312_ (_31061_, _31048_, _06306_);
  and _81313_ (_31062_, _31061_, _31060_);
  or _81314_ (_31063_, _31062_, _31059_);
  and _81315_ (_31064_, _31063_, _07130_);
  and _81316_ (_31066_, _30996_, _06411_);
  and _81317_ (_31067_, _31066_, _31060_);
  or _81318_ (_31068_, _31067_, _06303_);
  or _81319_ (_31069_, _31068_, _31064_);
  and _81320_ (_31070_, _30175_, _12797_);
  or _81321_ (_31071_, _30983_, _08819_);
  or _81322_ (_31072_, _31071_, _31070_);
  and _81323_ (_31073_, _31072_, _08824_);
  and _81324_ (_31074_, _31073_, _31069_);
  and _81325_ (_31075_, _30185_, _12797_);
  or _81326_ (_31077_, _31075_, _30983_);
  and _81327_ (_31078_, _31077_, _06396_);
  or _81328_ (_31079_, _31078_, _06433_);
  or _81329_ (_31080_, _31079_, _31074_);
  or _81330_ (_31081_, _30993_, _06829_);
  and _81331_ (_31082_, _31081_, _05749_);
  and _81332_ (_31083_, _31082_, _31080_);
  and _81333_ (_31084_, _30990_, _05748_);
  or _81334_ (_31085_, _31084_, _06440_);
  or _81335_ (_31086_, _31085_, _31083_);
  and _81336_ (_31088_, _30219_, _12797_);
  or _81337_ (_31089_, _30983_, _06444_);
  or _81338_ (_31090_, _31089_, _31088_);
  and _81339_ (_31091_, _31090_, _01317_);
  and _81340_ (_31092_, _31091_, _31086_);
  nor _81341_ (_31093_, \oc8051_golden_model_1.P3 [3], rst);
  nor _81342_ (_31094_, _31093_, _00000_);
  or _81343_ (_43716_, _31094_, _31092_);
  nor _81344_ (_31095_, \oc8051_golden_model_1.P3 [4], rst);
  nor _81345_ (_31096_, _31095_, _00000_);
  and _81346_ (_31098_, _12991_, \oc8051_golden_model_1.P3 [4]);
  and _81347_ (_31099_, _12797_, _08336_);
  or _81348_ (_31100_, _31099_, _31098_);
  or _81349_ (_31101_, _31100_, _06132_);
  and _81350_ (_31102_, _12996_, \oc8051_golden_model_1.P3 [4]);
  and _81351_ (_31103_, _30242_, _12780_);
  or _81352_ (_31104_, _31103_, _31102_);
  and _81353_ (_31105_, _31104_, _06152_);
  and _81354_ (_31106_, _30248_, _12797_);
  or _81355_ (_31107_, _31106_, _31098_);
  or _81356_ (_31109_, _31107_, _06161_);
  and _81357_ (_31110_, _12797_, \oc8051_golden_model_1.ACC [4]);
  or _81358_ (_31111_, _31110_, _31098_);
  and _81359_ (_31112_, _31111_, _07056_);
  and _81360_ (_31113_, _07057_, \oc8051_golden_model_1.P3 [4]);
  or _81361_ (_31114_, _31113_, _06160_);
  or _81362_ (_31115_, _31114_, _31112_);
  and _81363_ (_31116_, _31115_, _06157_);
  and _81364_ (_31117_, _31116_, _31109_);
  and _81365_ (_31118_, _30261_, _12780_);
  or _81366_ (_31120_, _31118_, _31102_);
  and _81367_ (_31121_, _31120_, _06156_);
  or _81368_ (_31122_, _31121_, _06217_);
  or _81369_ (_31123_, _31122_, _31117_);
  or _81370_ (_31124_, _31100_, _07075_);
  and _81371_ (_31125_, _31124_, _31123_);
  or _81372_ (_31126_, _31125_, _06220_);
  or _81373_ (_31127_, _31111_, _06229_);
  and _81374_ (_31128_, _31127_, _06153_);
  and _81375_ (_31129_, _31128_, _31126_);
  or _81376_ (_31131_, _31129_, _31105_);
  and _81377_ (_31132_, _31131_, _06146_);
  or _81378_ (_31133_, _31102_, _30276_);
  and _81379_ (_31134_, _31120_, _06145_);
  and _81380_ (_31135_, _31134_, _31133_);
  or _81381_ (_31136_, _31135_, _31132_);
  and _81382_ (_31137_, _31136_, _06140_);
  and _81383_ (_31138_, _30283_, _12780_);
  or _81384_ (_31139_, _31138_, _31102_);
  and _81385_ (_31140_, _31139_, _06139_);
  or _81386_ (_31143_, _31140_, _09842_);
  or _81387_ (_31144_, _31143_, _31137_);
  and _81388_ (_31145_, _31144_, _31101_);
  or _81389_ (_31146_, _31145_, _06116_);
  and _81390_ (_31147_, _12797_, _09209_);
  or _81391_ (_31148_, _31098_, _06117_);
  or _81392_ (_31149_, _31148_, _31147_);
  and _81393_ (_31150_, _31149_, _06114_);
  and _81394_ (_31151_, _31150_, _31146_);
  and _81395_ (_31152_, _30305_, _12797_);
  or _81396_ (_31154_, _31152_, _31098_);
  and _81397_ (_31155_, _31154_, _05787_);
  or _81398_ (_31156_, _31155_, _06110_);
  or _81399_ (_31157_, _31156_, _31151_);
  and _81400_ (_31158_, _12797_, _08715_);
  or _81401_ (_31159_, _31158_, _31098_);
  or _81402_ (_31160_, _31159_, _06111_);
  and _81403_ (_31161_, _31160_, _07127_);
  and _81404_ (_31162_, _31161_, _31157_);
  and _81405_ (_31163_, _30317_, _12797_);
  or _81406_ (_31166_, _31163_, _31098_);
  or _81407_ (_31167_, _31098_, _30320_);
  and _81408_ (_31168_, _31167_, _06297_);
  and _81409_ (_31169_, _31168_, _31166_);
  or _81410_ (_31170_, _31169_, _06402_);
  or _81411_ (_31171_, _31170_, _31162_);
  and _81412_ (_31172_, _30330_, _30327_);
  and _81413_ (_31173_, _31172_, _12797_);
  or _81414_ (_31174_, _31098_, _07125_);
  or _81415_ (_31175_, _31174_, _31173_);
  and _81416_ (_31177_, _31175_, _07132_);
  and _81417_ (_31178_, _31177_, _31171_);
  or _81418_ (_31179_, _31098_, _12826_);
  and _81419_ (_31180_, _31159_, _06306_);
  and _81420_ (_31181_, _31180_, _31179_);
  or _81421_ (_31182_, _31181_, _31178_);
  and _81422_ (_31183_, _31182_, _07130_);
  and _81423_ (_31184_, _31111_, _06411_);
  and _81424_ (_31185_, _31184_, _31179_);
  or _81425_ (_31186_, _31185_, _06303_);
  or _81426_ (_31189_, _31186_, _31183_);
  or _81427_ (_31190_, _31166_, _08819_);
  and _81428_ (_31191_, _31190_, _08824_);
  and _81429_ (_31192_, _31191_, _31189_);
  and _81430_ (_31193_, _30327_, _12797_);
  or _81431_ (_31194_, _31193_, _31098_);
  and _81432_ (_31195_, _31194_, _06396_);
  or _81433_ (_31196_, _31195_, _06433_);
  or _81434_ (_31197_, _31196_, _31192_);
  or _81435_ (_31198_, _31107_, _06829_);
  and _81436_ (_31200_, _31198_, _05749_);
  and _81437_ (_31201_, _31200_, _31197_);
  and _81438_ (_31202_, _31104_, _05748_);
  or _81439_ (_31203_, _31202_, _06440_);
  or _81440_ (_31204_, _31203_, _31201_);
  and _81441_ (_31205_, _30361_, _12797_);
  or _81442_ (_31206_, _31098_, _06444_);
  or _81443_ (_31207_, _31206_, _31205_);
  and _81444_ (_31208_, _31207_, _01317_);
  and _81445_ (_31209_, _31208_, _31204_);
  or _81446_ (_43717_, _31209_, _31096_);
  and _81447_ (_31212_, _12991_, \oc8051_golden_model_1.P3 [5]);
  and _81448_ (_31213_, _12797_, _08101_);
  or _81449_ (_31214_, _31213_, _31212_);
  or _81450_ (_31215_, _31214_, _06132_);
  and _81451_ (_31216_, _30378_, _12797_);
  or _81452_ (_31217_, _31216_, _31212_);
  or _81453_ (_31218_, _31217_, _06161_);
  and _81454_ (_31219_, _12797_, \oc8051_golden_model_1.ACC [5]);
  or _81455_ (_31220_, _31219_, _31212_);
  and _81456_ (_31222_, _31220_, _07056_);
  and _81457_ (_31223_, _07057_, \oc8051_golden_model_1.P3 [5]);
  or _81458_ (_31224_, _31223_, _06160_);
  or _81459_ (_31225_, _31224_, _31222_);
  and _81460_ (_31226_, _31225_, _06157_);
  and _81461_ (_31227_, _31226_, _31218_);
  and _81462_ (_31228_, _12996_, \oc8051_golden_model_1.P3 [5]);
  and _81463_ (_31229_, _30400_, _12780_);
  or _81464_ (_31230_, _31229_, _31228_);
  and _81465_ (_31231_, _31230_, _06156_);
  or _81466_ (_31233_, _31231_, _06217_);
  or _81467_ (_31234_, _31233_, _31227_);
  or _81468_ (_31235_, _31214_, _07075_);
  and _81469_ (_31236_, _31235_, _31234_);
  or _81470_ (_31237_, _31236_, _06220_);
  or _81471_ (_31238_, _31220_, _06229_);
  and _81472_ (_31239_, _31238_, _06153_);
  and _81473_ (_31240_, _31239_, _31237_);
  and _81474_ (_31241_, _30414_, _12780_);
  or _81475_ (_31242_, _31241_, _31228_);
  and _81476_ (_31244_, _31242_, _06152_);
  or _81477_ (_31245_, _31244_, _06145_);
  or _81478_ (_31246_, _31245_, _31240_);
  or _81479_ (_31247_, _31228_, _30420_);
  and _81480_ (_31248_, _31247_, _31230_);
  or _81481_ (_31249_, _31248_, _06146_);
  and _81482_ (_31250_, _31249_, _06140_);
  and _81483_ (_31251_, _31250_, _31246_);
  and _81484_ (_31252_, _30426_, _12780_);
  or _81485_ (_31253_, _31252_, _31228_);
  and _81486_ (_31254_, _31253_, _06139_);
  or _81487_ (_31255_, _31254_, _09842_);
  or _81488_ (_31256_, _31255_, _31251_);
  and _81489_ (_31257_, _31256_, _31215_);
  or _81490_ (_31258_, _31257_, _06116_);
  and _81491_ (_31259_, _12797_, _09208_);
  or _81492_ (_31260_, _31212_, _06117_);
  or _81493_ (_31261_, _31260_, _31259_);
  and _81494_ (_31262_, _31261_, _06114_);
  and _81495_ (_31263_, _31262_, _31258_);
  and _81496_ (_31266_, _30449_, _12797_);
  or _81497_ (_31267_, _31266_, _31212_);
  and _81498_ (_31268_, _31267_, _05787_);
  or _81499_ (_31269_, _31268_, _06110_);
  or _81500_ (_31270_, _31269_, _31263_);
  and _81501_ (_31271_, _12797_, _08736_);
  or _81502_ (_31272_, _31271_, _31212_);
  or _81503_ (_31273_, _31272_, _06111_);
  and _81504_ (_31274_, _31273_, _07127_);
  and _81505_ (_31275_, _31274_, _31270_);
  and _81506_ (_31276_, _30461_, _12797_);
  or _81507_ (_31277_, _31276_, _31212_);
  or _81508_ (_31278_, _31212_, _30464_);
  and _81509_ (_31279_, _31278_, _06297_);
  and _81510_ (_31280_, _31279_, _31277_);
  or _81511_ (_31281_, _31280_, _31275_);
  and _81512_ (_31282_, _31281_, _07125_);
  and _81513_ (_31283_, _30471_, _12797_);
  or _81514_ (_31284_, _31283_, _31212_);
  or _81515_ (_31285_, _31212_, _30474_);
  and _81516_ (_31288_, _31285_, _06402_);
  and _81517_ (_31289_, _31288_, _31284_);
  or _81518_ (_31290_, _31289_, _31282_);
  and _81519_ (_31291_, _31290_, _07132_);
  or _81520_ (_31292_, _31212_, _12818_);
  and _81521_ (_31293_, _31272_, _06306_);
  and _81522_ (_31294_, _31293_, _31292_);
  or _81523_ (_31295_, _31294_, _31291_);
  and _81524_ (_31296_, _31295_, _07130_);
  and _81525_ (_31297_, _31220_, _06411_);
  and _81526_ (_31298_, _31297_, _31292_);
  or _81527_ (_31299_, _31298_, _06303_);
  or _81528_ (_31300_, _31299_, _31296_);
  or _81529_ (_31301_, _31277_, _08819_);
  and _81530_ (_31302_, _31301_, _08824_);
  and _81531_ (_31303_, _31302_, _31300_);
  and _81532_ (_31304_, _31284_, _06396_);
  or _81533_ (_31305_, _31304_, _06433_);
  or _81534_ (_31306_, _31305_, _31303_);
  or _81535_ (_31307_, _31217_, _06829_);
  and _81536_ (_31310_, _31307_, _05749_);
  and _81537_ (_31311_, _31310_, _31306_);
  and _81538_ (_31312_, _31242_, _05748_);
  or _81539_ (_31313_, _31312_, _06440_);
  or _81540_ (_31314_, _31313_, _31311_);
  and _81541_ (_31315_, _30505_, _12797_);
  or _81542_ (_31316_, _31212_, _06444_);
  or _81543_ (_31317_, _31316_, _31315_);
  and _81544_ (_31318_, _31317_, _01317_);
  and _81545_ (_31319_, _31318_, _31314_);
  nor _81546_ (_31320_, \oc8051_golden_model_1.P3 [5], rst);
  nor _81547_ (_31321_, _31320_, _00000_);
  or _81548_ (_43719_, _31321_, _31319_);
  and _81549_ (_31322_, _12991_, \oc8051_golden_model_1.P3 [6]);
  and _81550_ (_31323_, _12797_, _08012_);
  or _81551_ (_31324_, _31323_, _31322_);
  or _81552_ (_31325_, _31324_, _06132_);
  and _81553_ (_31326_, _12996_, \oc8051_golden_model_1.P3 [6]);
  and _81554_ (_31327_, _30526_, _12780_);
  or _81555_ (_31328_, _31327_, _31326_);
  and _81556_ (_31331_, _31328_, _06152_);
  and _81557_ (_31332_, _30532_, _12797_);
  or _81558_ (_31333_, _31332_, _31322_);
  or _81559_ (_31334_, _31333_, _06161_);
  and _81560_ (_31335_, _12797_, \oc8051_golden_model_1.ACC [6]);
  or _81561_ (_31336_, _31335_, _31322_);
  and _81562_ (_31337_, _31336_, _07056_);
  and _81563_ (_31338_, _07057_, \oc8051_golden_model_1.P3 [6]);
  or _81564_ (_31339_, _31338_, _06160_);
  or _81565_ (_31340_, _31339_, _31337_);
  and _81566_ (_31341_, _31340_, _06157_);
  and _81567_ (_31342_, _31341_, _31334_);
  and _81568_ (_31343_, _30545_, _12780_);
  or _81569_ (_31344_, _31343_, _31326_);
  and _81570_ (_31345_, _31344_, _06156_);
  or _81571_ (_31346_, _31345_, _06217_);
  or _81572_ (_31347_, _31346_, _31342_);
  or _81573_ (_31348_, _31324_, _07075_);
  and _81574_ (_31349_, _31348_, _31347_);
  or _81575_ (_31350_, _31349_, _06220_);
  or _81576_ (_31353_, _31336_, _06229_);
  and _81577_ (_31354_, _31353_, _06153_);
  and _81578_ (_31355_, _31354_, _31350_);
  or _81579_ (_31356_, _31355_, _31331_);
  and _81580_ (_31357_, _31356_, _06146_);
  or _81581_ (_31358_, _31326_, _30560_);
  and _81582_ (_31359_, _31344_, _06145_);
  and _81583_ (_31360_, _31359_, _31358_);
  or _81584_ (_31361_, _31360_, _31357_);
  and _81585_ (_31362_, _31361_, _06140_);
  and _81586_ (_31363_, _30567_, _12780_);
  or _81587_ (_31364_, _31363_, _31326_);
  and _81588_ (_31365_, _31364_, _06139_);
  or _81589_ (_31366_, _31365_, _09842_);
  or _81590_ (_31367_, _31366_, _31362_);
  and _81591_ (_31368_, _31367_, _31325_);
  or _81592_ (_31369_, _31368_, _06116_);
  and _81593_ (_31370_, _12797_, _09207_);
  or _81594_ (_31371_, _31322_, _06117_);
  or _81595_ (_31372_, _31371_, _31370_);
  and _81596_ (_31375_, _31372_, _06114_);
  and _81597_ (_31376_, _31375_, _31369_);
  and _81598_ (_31377_, _30589_, _12797_);
  or _81599_ (_31378_, _31377_, _31322_);
  and _81600_ (_31379_, _31378_, _05787_);
  or _81601_ (_31380_, _31379_, _06110_);
  or _81602_ (_31381_, _31380_, _31376_);
  and _81603_ (_31382_, _12797_, _15402_);
  or _81604_ (_31383_, _31382_, _31322_);
  or _81605_ (_31384_, _31383_, _06111_);
  and _81606_ (_31385_, _31384_, _07127_);
  and _81607_ (_31386_, _31385_, _31381_);
  and _81608_ (_31387_, _30601_, _12797_);
  or _81609_ (_31388_, _31387_, _31322_);
  or _81610_ (_31389_, _31322_, _30604_);
  and _81611_ (_31390_, _31389_, _06297_);
  and _81612_ (_31391_, _31390_, _31388_);
  or _81613_ (_31392_, _31391_, _06402_);
  or _81614_ (_31393_, _31392_, _31386_);
  and _81615_ (_31394_, _30613_, _12797_);
  or _81616_ (_31396_, _31322_, _07125_);
  or _81617_ (_31397_, _31396_, _31394_);
  and _81618_ (_31398_, _31397_, _07132_);
  and _81619_ (_31399_, _31398_, _31393_);
  or _81620_ (_31400_, _31322_, _12810_);
  and _81621_ (_31401_, _31383_, _06306_);
  and _81622_ (_31402_, _31401_, _31400_);
  or _81623_ (_31403_, _31402_, _31399_);
  and _81624_ (_31404_, _31403_, _07130_);
  and _81625_ (_31405_, _31336_, _06411_);
  and _81626_ (_31406_, _31405_, _31400_);
  or _81627_ (_31407_, _31406_, _06303_);
  or _81628_ (_31408_, _31407_, _31404_);
  or _81629_ (_31409_, _31388_, _08819_);
  and _81630_ (_31410_, _31409_, _08824_);
  and _81631_ (_31411_, _31410_, _31408_);
  and _81632_ (_31412_, _30611_, _12797_);
  or _81633_ (_31413_, _31412_, _31322_);
  and _81634_ (_31414_, _31413_, _06396_);
  or _81635_ (_31415_, _31414_, _06433_);
  or _81636_ (_31418_, _31415_, _31411_);
  or _81637_ (_31419_, _31333_, _06829_);
  and _81638_ (_31420_, _31419_, _05749_);
  and _81639_ (_31421_, _31420_, _31418_);
  and _81640_ (_31422_, _31328_, _05748_);
  or _81641_ (_31423_, _31422_, _06440_);
  or _81642_ (_31424_, _31423_, _31421_);
  and _81643_ (_31425_, _30646_, _12797_);
  or _81644_ (_31426_, _31322_, _06444_);
  or _81645_ (_31427_, _31426_, _31425_);
  and _81646_ (_31428_, _31427_, _01317_);
  and _81647_ (_31429_, _31428_, _31424_);
  nor _81648_ (_31430_, \oc8051_golden_model_1.P3 [6], rst);
  nor _81649_ (_31431_, _31430_, _00000_);
  or _81650_ (_43720_, _31431_, _31429_);
  nor _81651_ (_31432_, \oc8051_golden_model_1.P0 [0], rst);
  nor _81652_ (_31433_, _31432_, _00000_);
  and _81653_ (_31434_, _13096_, \oc8051_golden_model_1.P0 [0]);
  and _81654_ (_31435_, _29675_, _12789_);
  or _81655_ (_31436_, _31435_, _31434_);
  and _81656_ (_31439_, _31436_, _06402_);
  and _81657_ (_31440_, _12789_, _07049_);
  or _81658_ (_31441_, _31440_, _31434_);
  or _81659_ (_31442_, _31441_, _06132_);
  and _81660_ (_31443_, _13101_, \oc8051_golden_model_1.P0 [0]);
  and _81661_ (_31444_, _29705_, _07847_);
  or _81662_ (_31445_, _31444_, _31443_);
  or _81663_ (_31446_, _31445_, _06157_);
  nor _81664_ (_31447_, _12858_, _13096_);
  or _81665_ (_31448_, _31447_, _31434_);
  and _81666_ (_31449_, _31448_, _06160_);
  and _81667_ (_31450_, _07057_, \oc8051_golden_model_1.P0 [0]);
  and _81668_ (_31451_, _12789_, \oc8051_golden_model_1.ACC [0]);
  or _81669_ (_31452_, _31451_, _31434_);
  and _81670_ (_31453_, _31452_, _07056_);
  or _81671_ (_31454_, _31453_, _31450_);
  and _81672_ (_31455_, _31454_, _06161_);
  or _81673_ (_31456_, _31455_, _06156_);
  or _81674_ (_31457_, _31456_, _31449_);
  and _81675_ (_31458_, _31457_, _31446_);
  and _81676_ (_31461_, _31458_, _07075_);
  and _81677_ (_31462_, _31441_, _06217_);
  or _81678_ (_31463_, _31462_, _06220_);
  or _81679_ (_31464_, _31463_, _31461_);
  or _81680_ (_31465_, _31452_, _06229_);
  and _81681_ (_31466_, _31465_, _06153_);
  and _81682_ (_31467_, _31466_, _31464_);
  and _81683_ (_31468_, _31434_, _06152_);
  or _81684_ (_31469_, _31468_, _06145_);
  or _81685_ (_31470_, _31469_, _31467_);
  or _81686_ (_31471_, _31448_, _06146_);
  and _81687_ (_31472_, _31471_, _06140_);
  and _81688_ (_31473_, _31472_, _31470_);
  or _81689_ (_31474_, _31443_, _14170_);
  and _81690_ (_31475_, _31474_, _06139_);
  and _81691_ (_31476_, _31475_, _31445_);
  or _81692_ (_31477_, _31476_, _09842_);
  or _81693_ (_31478_, _31477_, _31473_);
  and _81694_ (_31479_, _31478_, _31442_);
  or _81695_ (_31480_, _31479_, _06116_);
  and _81696_ (_31483_, _12789_, _09160_);
  or _81697_ (_31484_, _31434_, _06117_);
  or _81698_ (_31485_, _31484_, _31483_);
  and _81699_ (_31486_, _31485_, _06114_);
  and _81700_ (_31487_, _31486_, _31480_);
  and _81701_ (_31488_, _29746_, _12789_);
  or _81702_ (_31489_, _31488_, _31434_);
  and _81703_ (_31490_, _31489_, _05787_);
  or _81704_ (_31491_, _31490_, _31487_);
  or _81705_ (_31492_, _31491_, _11136_);
  and _81706_ (_31493_, _29756_, _12789_);
  or _81707_ (_31494_, _31434_, _07127_);
  or _81708_ (_31495_, _31494_, _31493_);
  and _81709_ (_31496_, _12789_, _08708_);
  or _81710_ (_31497_, _31496_, _31434_);
  or _81711_ (_31498_, _31497_, _06111_);
  and _81712_ (_31499_, _31498_, _07125_);
  and _81713_ (_31500_, _31499_, _31495_);
  and _81714_ (_31501_, _31500_, _31492_);
  or _81715_ (_31502_, _31501_, _31439_);
  and _81716_ (_31505_, _31502_, _07132_);
  nand _81717_ (_31506_, _31497_, _06306_);
  nor _81718_ (_31507_, _31506_, _31447_);
  or _81719_ (_31508_, _31507_, _31505_);
  and _81720_ (_31509_, _31508_, _07130_);
  or _81721_ (_31510_, _31434_, _12858_);
  and _81722_ (_31511_, _31452_, _06411_);
  and _81723_ (_31512_, _31511_, _31510_);
  or _81724_ (_31513_, _31512_, _06303_);
  or _81725_ (_31514_, _31513_, _31509_);
  and _81726_ (_31515_, _29752_, _12789_);
  or _81727_ (_31516_, _31434_, _08819_);
  or _81728_ (_31517_, _31516_, _31515_);
  and _81729_ (_31518_, _31517_, _08824_);
  and _81730_ (_31519_, _31518_, _31514_);
  and _81731_ (_31520_, _29673_, _12789_);
  or _81732_ (_31521_, _31520_, _31434_);
  and _81733_ (_31522_, _31521_, _06396_);
  or _81734_ (_31523_, _31522_, _06433_);
  or _81735_ (_31524_, _31523_, _31519_);
  or _81736_ (_31527_, _31448_, _06829_);
  and _81737_ (_31528_, _31527_, _05749_);
  and _81738_ (_31529_, _31528_, _31524_);
  and _81739_ (_31530_, _31434_, _05748_);
  or _81740_ (_31531_, _31530_, _06440_);
  or _81741_ (_31532_, _31531_, _31529_);
  or _81742_ (_31533_, _31448_, _06444_);
  and _81743_ (_31534_, _31533_, _01317_);
  and _81744_ (_31535_, _31534_, _31532_);
  or _81745_ (_43721_, _31535_, _31433_);
  nor _81746_ (_31536_, \oc8051_golden_model_1.P0 [1], rst);
  nor _81747_ (_31537_, _31536_, _00000_);
  or _81748_ (_31538_, _29883_, _13096_);
  or _81749_ (_31539_, _12789_, \oc8051_golden_model_1.P0 [1]);
  and _81750_ (_31540_, _31539_, _05787_);
  and _81751_ (_31541_, _31540_, _31538_);
  and _81752_ (_31542_, _29814_, _07847_);
  and _81753_ (_31543_, _31542_, _29813_);
  and _81754_ (_31544_, _13101_, \oc8051_golden_model_1.P0 [1]);
  or _81755_ (_31545_, _31544_, _06146_);
  or _81756_ (_31548_, _31545_, _31543_);
  and _81757_ (_31549_, _29823_, _12789_);
  not _81758_ (_31550_, _31549_);
  and _81759_ (_31551_, _31550_, _31539_);
  or _81760_ (_31552_, _31551_, _06161_);
  nand _81761_ (_31553_, _12789_, _05887_);
  and _81762_ (_31554_, _31553_, _31539_);
  and _81763_ (_31555_, _31554_, _07056_);
  and _81764_ (_31556_, _07057_, \oc8051_golden_model_1.P0 [1]);
  or _81765_ (_31557_, _31556_, _06160_);
  or _81766_ (_31558_, _31557_, _31555_);
  and _81767_ (_31559_, _31558_, _06157_);
  and _81768_ (_31560_, _31559_, _31552_);
  or _81769_ (_31561_, _31544_, _06217_);
  or _81770_ (_31562_, _31561_, _31542_);
  and _81771_ (_31563_, _31562_, _13860_);
  or _81772_ (_31564_, _31563_, _31560_);
  and _81773_ (_31565_, _13096_, \oc8051_golden_model_1.P0 [1]);
  and _81774_ (_31566_, _12789_, _07306_);
  or _81775_ (_31567_, _31566_, _31565_);
  or _81776_ (_31570_, _31567_, _07075_);
  and _81777_ (_31571_, _31570_, _31564_);
  or _81778_ (_31572_, _31571_, _06220_);
  or _81779_ (_31573_, _31554_, _06229_);
  and _81780_ (_31574_, _31573_, _06153_);
  and _81781_ (_31575_, _31574_, _31572_);
  and _81782_ (_31576_, _29851_, _07847_);
  or _81783_ (_31577_, _31576_, _31544_);
  and _81784_ (_31578_, _31577_, _06152_);
  or _81785_ (_31579_, _31578_, _06145_);
  or _81786_ (_31580_, _31579_, _31575_);
  and _81787_ (_31581_, _31580_, _31548_);
  and _81788_ (_31582_, _31581_, _06140_);
  and _81789_ (_31583_, _29860_, _07847_);
  or _81790_ (_31584_, _31544_, _31583_);
  and _81791_ (_31585_, _31584_, _06139_);
  or _81792_ (_31586_, _31585_, _09842_);
  or _81793_ (_31587_, _31586_, _31582_);
  or _81794_ (_31588_, _31567_, _06132_);
  and _81795_ (_31589_, _31588_, _31587_);
  or _81796_ (_31592_, _31589_, _06116_);
  and _81797_ (_31593_, _12789_, _09115_);
  or _81798_ (_31594_, _31565_, _06117_);
  or _81799_ (_31595_, _31594_, _31593_);
  and _81800_ (_31596_, _31595_, _06114_);
  and _81801_ (_31597_, _31596_, _31592_);
  or _81802_ (_31598_, _31597_, _31541_);
  and _81803_ (_31599_, _31598_, _06298_);
  or _81804_ (_31600_, _30823_, _13096_);
  and _81805_ (_31601_, _31600_, _06297_);
  nand _81806_ (_31602_, _12789_, _06945_);
  and _81807_ (_31603_, _31602_, _06110_);
  or _81808_ (_31604_, _31603_, _31601_);
  and _81809_ (_31605_, _31604_, _31539_);
  or _81810_ (_31606_, _31605_, _31599_);
  and _81811_ (_31607_, _31606_, _07125_);
  or _81812_ (_31608_, _30833_, _13096_);
  and _81813_ (_31609_, _31539_, _06402_);
  and _81814_ (_31610_, _31609_, _31608_);
  or _81815_ (_31611_, _31610_, _31607_);
  and _81816_ (_31614_, _31611_, _07132_);
  or _81817_ (_31615_, _29896_, _13096_);
  and _81818_ (_31616_, _31539_, _06306_);
  and _81819_ (_31617_, _31616_, _31615_);
  or _81820_ (_31618_, _31617_, _31614_);
  and _81821_ (_31619_, _31618_, _07130_);
  or _81822_ (_31620_, _31565_, _12850_);
  and _81823_ (_31621_, _31554_, _06411_);
  and _81824_ (_31622_, _31621_, _31620_);
  or _81825_ (_31623_, _31622_, _31619_);
  and _81826_ (_31624_, _31623_, _06397_);
  or _81827_ (_31625_, _31602_, _12850_);
  and _81828_ (_31626_, _31539_, _06303_);
  and _81829_ (_31627_, _31626_, _31625_);
  or _81830_ (_31628_, _31553_, _12850_);
  and _81831_ (_31629_, _31539_, _06396_);
  and _81832_ (_31630_, _31629_, _31628_);
  or _81833_ (_31631_, _31630_, _06433_);
  or _81834_ (_31632_, _31631_, _31627_);
  or _81835_ (_31633_, _31632_, _31624_);
  or _81836_ (_31636_, _31551_, _06829_);
  and _81837_ (_31637_, _31636_, _05749_);
  and _81838_ (_31638_, _31637_, _31633_);
  and _81839_ (_31639_, _31577_, _05748_);
  or _81840_ (_31640_, _31639_, _06440_);
  or _81841_ (_31641_, _31640_, _31638_);
  or _81842_ (_31642_, _31565_, _06444_);
  or _81843_ (_31643_, _31642_, _31549_);
  and _81844_ (_31644_, _31643_, _01317_);
  and _81845_ (_31645_, _31644_, _31641_);
  or _81846_ (_43723_, _31645_, _31537_);
  nor _81847_ (_31646_, \oc8051_golden_model_1.P0 [2], rst);
  nor _81848_ (_31647_, _31646_, _00000_);
  and _81849_ (_31648_, _13096_, \oc8051_golden_model_1.P0 [2]);
  and _81850_ (_31649_, _12789_, _07708_);
  or _81851_ (_31650_, _31649_, _31648_);
  or _81852_ (_31651_, _31650_, _06132_);
  and _81853_ (_31652_, _29954_, _12789_);
  or _81854_ (_31653_, _31652_, _31648_);
  or _81855_ (_31654_, _31653_, _06161_);
  and _81856_ (_31657_, _12789_, \oc8051_golden_model_1.ACC [2]);
  or _81857_ (_31658_, _31657_, _31648_);
  and _81858_ (_31659_, _31658_, _07056_);
  and _81859_ (_31660_, _07057_, \oc8051_golden_model_1.P0 [2]);
  or _81860_ (_31661_, _31660_, _06160_);
  or _81861_ (_31662_, _31661_, _31659_);
  and _81862_ (_31663_, _31662_, _06157_);
  and _81863_ (_31664_, _31663_, _31654_);
  and _81864_ (_31665_, _13101_, \oc8051_golden_model_1.P0 [2]);
  and _81865_ (_31666_, _29976_, _07847_);
  or _81866_ (_31667_, _31666_, _31665_);
  and _81867_ (_31668_, _31667_, _06156_);
  or _81868_ (_31669_, _31668_, _06217_);
  or _81869_ (_31670_, _31669_, _31664_);
  or _81870_ (_31671_, _31650_, _07075_);
  and _81871_ (_31672_, _31671_, _31670_);
  or _81872_ (_31673_, _31672_, _06220_);
  or _81873_ (_31674_, _31658_, _06229_);
  and _81874_ (_31675_, _31674_, _06153_);
  and _81875_ (_31676_, _31675_, _31673_);
  and _81876_ (_31679_, _29992_, _07847_);
  or _81877_ (_31680_, _31679_, _31665_);
  and _81878_ (_31681_, _31680_, _06152_);
  or _81879_ (_31682_, _31681_, _06145_);
  or _81880_ (_31683_, _31682_, _31676_);
  or _81881_ (_31684_, _31665_, _29999_);
  and _81882_ (_31685_, _31684_, _31667_);
  or _81883_ (_31686_, _31685_, _06146_);
  and _81884_ (_31687_, _31686_, _06140_);
  and _81885_ (_31688_, _31687_, _31683_);
  and _81886_ (_31689_, _30005_, _07847_);
  or _81887_ (_31690_, _31689_, _31665_);
  and _81888_ (_31691_, _31690_, _06139_);
  or _81889_ (_31692_, _31691_, _09842_);
  or _81890_ (_31693_, _31692_, _31688_);
  and _81891_ (_31694_, _31693_, _31651_);
  or _81892_ (_31695_, _31694_, _06116_);
  and _81893_ (_31696_, _12789_, _09211_);
  or _81894_ (_31697_, _31648_, _06117_);
  or _81895_ (_31698_, _31697_, _31696_);
  and _81896_ (_31701_, _31698_, _06114_);
  and _81897_ (_31702_, _31701_, _31695_);
  and _81898_ (_31703_, _30029_, _12789_);
  or _81899_ (_31704_, _31648_, _31703_);
  and _81900_ (_31705_, _31704_, _05787_);
  or _81901_ (_31706_, _31705_, _31702_);
  or _81902_ (_31707_, _31706_, _11136_);
  and _81903_ (_31708_, _29948_, _29945_);
  and _81904_ (_31709_, _31708_, _12789_);
  or _81905_ (_31710_, _31648_, _07127_);
  or _81906_ (_31711_, _31710_, _31709_);
  and _81907_ (_31712_, _12789_, _08768_);
  or _81908_ (_31713_, _31712_, _31648_);
  or _81909_ (_31714_, _31713_, _06111_);
  and _81910_ (_31715_, _31714_, _07125_);
  and _81911_ (_31716_, _31715_, _31711_);
  and _81912_ (_31717_, _31716_, _31707_);
  and _81913_ (_31718_, _30043_, _12789_);
  and _81914_ (_31719_, _31718_, _30046_);
  or _81915_ (_31720_, _31719_, _31648_);
  and _81916_ (_31723_, _31720_, _06402_);
  or _81917_ (_31724_, _31723_, _31717_);
  and _81918_ (_31725_, _31724_, _07132_);
  or _81919_ (_31726_, _31648_, _12842_);
  and _81920_ (_31727_, _31713_, _06306_);
  and _81921_ (_31728_, _31727_, _31726_);
  or _81922_ (_31729_, _31728_, _31725_);
  and _81923_ (_31730_, _31729_, _07130_);
  and _81924_ (_31731_, _31658_, _06411_);
  and _81925_ (_31732_, _31731_, _31726_);
  or _81926_ (_31733_, _31732_, _06303_);
  or _81927_ (_31734_, _31733_, _31730_);
  and _81928_ (_31735_, _29945_, _12789_);
  or _81929_ (_31736_, _31648_, _08819_);
  or _81930_ (_31737_, _31736_, _31735_);
  and _81931_ (_31738_, _31737_, _08824_);
  and _81932_ (_31739_, _31738_, _31734_);
  or _81933_ (_31740_, _31718_, _31648_);
  and _81934_ (_31741_, _31740_, _06396_);
  or _81935_ (_31742_, _31741_, _06433_);
  or _81936_ (_31745_, _31742_, _31739_);
  or _81937_ (_31746_, _31653_, _06829_);
  and _81938_ (_31747_, _31746_, _05749_);
  and _81939_ (_31748_, _31747_, _31745_);
  and _81940_ (_31749_, _31680_, _05748_);
  or _81941_ (_31750_, _31749_, _06440_);
  or _81942_ (_31751_, _31750_, _31748_);
  and _81943_ (_31752_, _30077_, _12789_);
  or _81944_ (_31753_, _31648_, _06444_);
  or _81945_ (_31754_, _31753_, _31752_);
  and _81946_ (_31755_, _31754_, _01317_);
  and _81947_ (_31756_, _31755_, _31751_);
  or _81948_ (_43724_, _31756_, _31647_);
  and _81949_ (_31757_, _13096_, \oc8051_golden_model_1.P0 [3]);
  and _81950_ (_31758_, _12789_, _07544_);
  or _81951_ (_31759_, _31758_, _31757_);
  or _81952_ (_31760_, _31759_, _06132_);
  and _81953_ (_31761_, _13101_, \oc8051_golden_model_1.P0 [3]);
  and _81954_ (_31762_, _30100_, _07847_);
  or _81955_ (_31763_, _31762_, _31761_);
  and _81956_ (_31766_, _31763_, _06152_);
  and _81957_ (_31767_, _30106_, _12789_);
  or _81958_ (_31768_, _31767_, _31757_);
  or _81959_ (_31769_, _31768_, _06161_);
  and _81960_ (_31770_, _12789_, \oc8051_golden_model_1.ACC [3]);
  or _81961_ (_31771_, _31770_, _31757_);
  and _81962_ (_31772_, _31771_, _07056_);
  and _81963_ (_31773_, _07057_, \oc8051_golden_model_1.P0 [3]);
  or _81964_ (_31774_, _31773_, _06160_);
  or _81965_ (_31775_, _31774_, _31772_);
  and _81966_ (_31776_, _31775_, _06157_);
  and _81967_ (_31777_, _31776_, _31769_);
  and _81968_ (_31778_, _30119_, _07847_);
  or _81969_ (_31779_, _31778_, _31761_);
  and _81970_ (_31780_, _31779_, _06156_);
  or _81971_ (_31781_, _31780_, _06217_);
  or _81972_ (_31782_, _31781_, _31777_);
  or _81973_ (_31783_, _31759_, _07075_);
  and _81974_ (_31784_, _31783_, _31782_);
  or _81975_ (_31785_, _31784_, _06220_);
  or _81976_ (_31788_, _31771_, _06229_);
  and _81977_ (_31789_, _31788_, _06153_);
  and _81978_ (_31790_, _31789_, _31785_);
  or _81979_ (_31791_, _31790_, _31766_);
  and _81980_ (_31792_, _31791_, _06146_);
  or _81981_ (_31793_, _31761_, _30134_);
  and _81982_ (_31794_, _31779_, _06145_);
  and _81983_ (_31795_, _31794_, _31793_);
  or _81984_ (_31796_, _31795_, _31792_);
  and _81985_ (_31797_, _31796_, _06140_);
  and _81986_ (_31798_, _30141_, _07847_);
  or _81987_ (_31799_, _31798_, _31761_);
  and _81988_ (_31800_, _31799_, _06139_);
  or _81989_ (_31801_, _31800_, _09842_);
  or _81990_ (_31802_, _31801_, _31797_);
  and _81991_ (_31803_, _31802_, _31760_);
  or _81992_ (_31804_, _31803_, _06116_);
  and _81993_ (_31805_, _12789_, _09210_);
  or _81994_ (_31806_, _31757_, _06117_);
  or _81995_ (_31807_, _31806_, _31805_);
  and _81996_ (_31810_, _31807_, _06114_);
  and _81997_ (_31811_, _31810_, _31804_);
  and _81998_ (_31812_, _30163_, _12789_);
  or _81999_ (_31813_, _31812_, _31757_);
  and _82000_ (_31814_, _31813_, _05787_);
  or _82001_ (_31815_, _31814_, _11136_);
  or _82002_ (_31816_, _31815_, _31811_);
  and _82003_ (_31817_, _31042_, _12789_);
  or _82004_ (_31818_, _31757_, _07127_);
  or _82005_ (_31819_, _31818_, _31817_);
  and _82006_ (_31820_, _12789_, _08712_);
  or _82007_ (_31821_, _31820_, _31757_);
  or _82008_ (_31822_, _31821_, _06111_);
  and _82009_ (_31823_, _31822_, _07125_);
  and _82010_ (_31824_, _31823_, _31819_);
  and _82011_ (_31825_, _31824_, _31816_);
  and _82012_ (_31826_, _31053_, _12789_);
  or _82013_ (_31827_, _31826_, _31757_);
  and _82014_ (_31828_, _31827_, _06402_);
  or _82015_ (_31829_, _31828_, _31825_);
  and _82016_ (_31832_, _31829_, _07132_);
  or _82017_ (_31833_, _31757_, _12834_);
  and _82018_ (_31834_, _31821_, _06306_);
  and _82019_ (_31835_, _31834_, _31833_);
  or _82020_ (_31836_, _31835_, _31832_);
  and _82021_ (_31837_, _31836_, _07130_);
  and _82022_ (_31838_, _31771_, _06411_);
  and _82023_ (_31839_, _31838_, _31833_);
  or _82024_ (_31840_, _31839_, _06303_);
  or _82025_ (_31841_, _31840_, _31837_);
  and _82026_ (_31842_, _30175_, _12789_);
  or _82027_ (_31843_, _31757_, _08819_);
  or _82028_ (_31844_, _31843_, _31842_);
  and _82029_ (_31845_, _31844_, _08824_);
  and _82030_ (_31846_, _31845_, _31841_);
  and _82031_ (_31847_, _30185_, _12789_);
  or _82032_ (_31848_, _31847_, _31757_);
  and _82033_ (_31849_, _31848_, _06396_);
  or _82034_ (_31850_, _31849_, _06433_);
  or _82035_ (_31851_, _31850_, _31846_);
  or _82036_ (_31854_, _31768_, _06829_);
  and _82037_ (_31855_, _31854_, _05749_);
  and _82038_ (_31856_, _31855_, _31851_);
  and _82039_ (_31857_, _31763_, _05748_);
  or _82040_ (_31858_, _31857_, _06440_);
  or _82041_ (_31859_, _31858_, _31856_);
  and _82042_ (_31860_, _30219_, _12789_);
  or _82043_ (_31861_, _31757_, _06444_);
  or _82044_ (_31862_, _31861_, _31860_);
  and _82045_ (_31863_, _31862_, _01317_);
  and _82046_ (_31865_, _31863_, _31859_);
  nor _82047_ (_31866_, \oc8051_golden_model_1.P0 [3], rst);
  nor _82048_ (_31867_, _31866_, _00000_);
  or _82049_ (_43725_, _31867_, _31865_);
  and _82050_ (_31868_, _13096_, \oc8051_golden_model_1.P0 [4]);
  and _82051_ (_31869_, _12789_, _08336_);
  or _82052_ (_31870_, _31869_, _31868_);
  or _82053_ (_31871_, _31870_, _06132_);
  and _82054_ (_31872_, _13101_, \oc8051_golden_model_1.P0 [4]);
  and _82055_ (_31873_, _30242_, _07847_);
  or _82056_ (_31875_, _31873_, _31872_);
  and _82057_ (_31876_, _31875_, _06152_);
  and _82058_ (_31877_, _30248_, _12789_);
  or _82059_ (_31878_, _31877_, _31868_);
  or _82060_ (_31879_, _31878_, _06161_);
  and _82061_ (_31880_, _12789_, \oc8051_golden_model_1.ACC [4]);
  or _82062_ (_31881_, _31880_, _31868_);
  and _82063_ (_31882_, _31881_, _07056_);
  and _82064_ (_31883_, _07057_, \oc8051_golden_model_1.P0 [4]);
  or _82065_ (_31884_, _31883_, _06160_);
  or _82066_ (_31886_, _31884_, _31882_);
  and _82067_ (_31887_, _31886_, _06157_);
  and _82068_ (_31888_, _31887_, _31879_);
  and _82069_ (_31889_, _30261_, _07847_);
  or _82070_ (_31890_, _31889_, _31872_);
  and _82071_ (_31891_, _31890_, _06156_);
  or _82072_ (_31892_, _31891_, _06217_);
  or _82073_ (_31893_, _31892_, _31888_);
  or _82074_ (_31894_, _31870_, _07075_);
  and _82075_ (_31895_, _31894_, _31893_);
  or _82076_ (_31897_, _31895_, _06220_);
  or _82077_ (_31898_, _31881_, _06229_);
  and _82078_ (_31899_, _31898_, _06153_);
  and _82079_ (_31900_, _31899_, _31897_);
  or _82080_ (_31901_, _31900_, _31876_);
  and _82081_ (_31902_, _31901_, _06146_);
  or _82082_ (_31903_, _31872_, _30276_);
  and _82083_ (_31904_, _31890_, _06145_);
  and _82084_ (_31905_, _31904_, _31903_);
  or _82085_ (_31906_, _31905_, _31902_);
  and _82086_ (_31908_, _31906_, _06140_);
  and _82087_ (_31909_, _30283_, _07847_);
  or _82088_ (_31910_, _31909_, _31872_);
  and _82089_ (_31911_, _31910_, _06139_);
  or _82090_ (_31912_, _31911_, _09842_);
  or _82091_ (_31913_, _31912_, _31908_);
  and _82092_ (_31914_, _31913_, _31871_);
  or _82093_ (_31915_, _31914_, _06116_);
  and _82094_ (_31916_, _12789_, _09209_);
  or _82095_ (_31917_, _31868_, _06117_);
  or _82096_ (_31919_, _31917_, _31916_);
  and _82097_ (_31920_, _31919_, _06114_);
  and _82098_ (_31921_, _31920_, _31915_);
  and _82099_ (_31922_, _30305_, _12789_);
  or _82100_ (_31923_, _31922_, _31868_);
  and _82101_ (_31924_, _31923_, _05787_);
  or _82102_ (_31925_, _31924_, _11136_);
  or _82103_ (_31926_, _31925_, _31921_);
  and _82104_ (_31927_, _30317_, _12789_);
  and _82105_ (_31928_, _31927_, _30320_);
  or _82106_ (_31930_, _31868_, _07127_);
  or _82107_ (_31931_, _31930_, _31928_);
  and _82108_ (_31932_, _12789_, _08715_);
  or _82109_ (_31933_, _31932_, _31868_);
  or _82110_ (_31934_, _31933_, _06111_);
  and _82111_ (_31935_, _31934_, _07125_);
  and _82112_ (_31936_, _31935_, _31931_);
  and _82113_ (_31937_, _31936_, _31926_);
  and _82114_ (_31938_, _31172_, _12789_);
  or _82115_ (_31939_, _31938_, _31868_);
  and _82116_ (_31941_, _31939_, _06402_);
  or _82117_ (_31942_, _31941_, _31937_);
  and _82118_ (_31943_, _31942_, _07132_);
  or _82119_ (_31944_, _31868_, _12826_);
  and _82120_ (_31945_, _31933_, _06306_);
  and _82121_ (_31946_, _31945_, _31944_);
  or _82122_ (_31947_, _31946_, _31943_);
  and _82123_ (_31948_, _31947_, _07130_);
  and _82124_ (_31949_, _31881_, _06411_);
  and _82125_ (_31950_, _31949_, _31944_);
  or _82126_ (_31951_, _31950_, _06303_);
  or _82127_ (_31952_, _31951_, _31948_);
  or _82128_ (_31953_, _31868_, _08819_);
  or _82129_ (_31954_, _31953_, _31927_);
  and _82130_ (_31955_, _31954_, _08824_);
  and _82131_ (_31956_, _31955_, _31952_);
  and _82132_ (_31957_, _30327_, _12789_);
  or _82133_ (_31958_, _31957_, _31868_);
  and _82134_ (_31959_, _31958_, _06396_);
  or _82135_ (_31960_, _31959_, _06433_);
  or _82136_ (_31962_, _31960_, _31956_);
  or _82137_ (_31963_, _31878_, _06829_);
  and _82138_ (_31964_, _31963_, _05749_);
  and _82139_ (_31965_, _31964_, _31962_);
  and _82140_ (_31966_, _31875_, _05748_);
  or _82141_ (_31967_, _31966_, _06440_);
  or _82142_ (_31968_, _31967_, _31965_);
  and _82143_ (_31969_, _30361_, _12789_);
  or _82144_ (_31970_, _31868_, _06444_);
  or _82145_ (_31971_, _31970_, _31969_);
  and _82146_ (_31973_, _31971_, _01317_);
  and _82147_ (_31974_, _31973_, _31968_);
  nor _82148_ (_31975_, \oc8051_golden_model_1.P0 [4], rst);
  nor _82149_ (_31976_, _31975_, _00000_);
  or _82150_ (_43726_, _31976_, _31974_);
  and _82151_ (_31977_, _13096_, \oc8051_golden_model_1.P0 [5]);
  and _82152_ (_31978_, _12789_, _08101_);
  or _82153_ (_31979_, _31978_, _31977_);
  or _82154_ (_31980_, _31979_, _06132_);
  and _82155_ (_31981_, _30378_, _12789_);
  or _82156_ (_31983_, _31981_, _31977_);
  or _82157_ (_31984_, _31983_, _06161_);
  and _82158_ (_31985_, _12789_, \oc8051_golden_model_1.ACC [5]);
  or _82159_ (_31986_, _31985_, _31977_);
  and _82160_ (_31987_, _31986_, _07056_);
  and _82161_ (_31988_, _07057_, \oc8051_golden_model_1.P0 [5]);
  or _82162_ (_31989_, _31988_, _06160_);
  or _82163_ (_31990_, _31989_, _31987_);
  and _82164_ (_31991_, _31990_, _06157_);
  and _82165_ (_31992_, _31991_, _31984_);
  and _82166_ (_31994_, _13101_, \oc8051_golden_model_1.P0 [5]);
  and _82167_ (_31995_, _30400_, _07847_);
  or _82168_ (_31996_, _31995_, _31994_);
  and _82169_ (_31997_, _31996_, _06156_);
  or _82170_ (_31998_, _31997_, _06217_);
  or _82171_ (_31999_, _31998_, _31992_);
  or _82172_ (_32000_, _31979_, _07075_);
  and _82173_ (_32001_, _32000_, _31999_);
  or _82174_ (_32002_, _32001_, _06220_);
  or _82175_ (_32003_, _31986_, _06229_);
  and _82176_ (_32005_, _32003_, _06153_);
  and _82177_ (_32006_, _32005_, _32002_);
  and _82178_ (_32007_, _30414_, _07847_);
  or _82179_ (_32008_, _32007_, _31994_);
  and _82180_ (_32009_, _32008_, _06152_);
  or _82181_ (_32010_, _32009_, _06145_);
  or _82182_ (_32011_, _32010_, _32006_);
  or _82183_ (_32012_, _31994_, _30420_);
  and _82184_ (_32013_, _32012_, _31996_);
  or _82185_ (_32014_, _32013_, _06146_);
  and _82186_ (_32016_, _32014_, _06140_);
  and _82187_ (_32017_, _32016_, _32011_);
  and _82188_ (_32018_, _30426_, _07847_);
  or _82189_ (_32019_, _32018_, _31994_);
  and _82190_ (_32020_, _32019_, _06139_);
  or _82191_ (_32021_, _32020_, _09842_);
  or _82192_ (_32022_, _32021_, _32017_);
  and _82193_ (_32023_, _32022_, _31980_);
  or _82194_ (_32024_, _32023_, _06116_);
  and _82195_ (_32025_, _12789_, _09208_);
  or _82196_ (_32027_, _31977_, _06117_);
  or _82197_ (_32028_, _32027_, _32025_);
  and _82198_ (_32029_, _32028_, _06114_);
  and _82199_ (_32030_, _32029_, _32024_);
  and _82200_ (_32031_, _30449_, _12789_);
  or _82201_ (_32032_, _32031_, _31977_);
  and _82202_ (_32033_, _32032_, _05787_);
  or _82203_ (_32034_, _32033_, _11136_);
  or _82204_ (_32035_, _32034_, _32030_);
  and _82205_ (_32036_, _30464_, _30461_);
  and _82206_ (_32038_, _32036_, _12789_);
  or _82207_ (_32039_, _31977_, _07127_);
  or _82208_ (_32040_, _32039_, _32038_);
  and _82209_ (_32041_, _12789_, _08736_);
  or _82210_ (_32042_, _32041_, _31977_);
  or _82211_ (_32043_, _32042_, _06111_);
  and _82212_ (_32044_, _32043_, _07125_);
  and _82213_ (_32045_, _32044_, _32040_);
  and _82214_ (_32046_, _32045_, _32035_);
  and _82215_ (_32047_, _30474_, _30471_);
  and _82216_ (_32049_, _32047_, _12789_);
  or _82217_ (_32050_, _32049_, _31977_);
  and _82218_ (_32051_, _32050_, _06402_);
  or _82219_ (_32052_, _32051_, _32046_);
  and _82220_ (_32053_, _32052_, _07132_);
  or _82221_ (_32054_, _31977_, _12818_);
  and _82222_ (_32055_, _32042_, _06306_);
  and _82223_ (_32056_, _32055_, _32054_);
  or _82224_ (_32057_, _32056_, _32053_);
  and _82225_ (_32058_, _32057_, _07130_);
  and _82226_ (_32060_, _31986_, _06411_);
  and _82227_ (_32061_, _32060_, _32054_);
  or _82228_ (_32062_, _32061_, _06303_);
  or _82229_ (_32063_, _32062_, _32058_);
  and _82230_ (_32064_, _30461_, _12789_);
  or _82231_ (_32065_, _31977_, _08819_);
  or _82232_ (_32066_, _32065_, _32064_);
  and _82233_ (_32067_, _32066_, _08824_);
  and _82234_ (_32068_, _32067_, _32063_);
  and _82235_ (_32069_, _30471_, _12789_);
  or _82236_ (_32071_, _32069_, _31977_);
  and _82237_ (_32072_, _32071_, _06396_);
  or _82238_ (_32073_, _32072_, _06433_);
  or _82239_ (_32074_, _32073_, _32068_);
  or _82240_ (_32075_, _31983_, _06829_);
  and _82241_ (_32076_, _32075_, _05749_);
  and _82242_ (_32077_, _32076_, _32074_);
  and _82243_ (_32078_, _32008_, _05748_);
  or _82244_ (_32079_, _32078_, _06440_);
  or _82245_ (_32080_, _32079_, _32077_);
  and _82246_ (_32082_, _30505_, _12789_);
  or _82247_ (_32083_, _31977_, _06444_);
  or _82248_ (_32084_, _32083_, _32082_);
  and _82249_ (_32085_, _32084_, _01317_);
  and _82250_ (_32086_, _32085_, _32080_);
  nor _82251_ (_32087_, \oc8051_golden_model_1.P0 [5], rst);
  nor _82252_ (_32088_, _32087_, _00000_);
  or _82253_ (_43727_, _32088_, _32086_);
  nor _82254_ (_32089_, \oc8051_golden_model_1.P0 [6], rst);
  nor _82255_ (_32090_, _32089_, _00000_);
  and _82256_ (_32092_, _13096_, \oc8051_golden_model_1.P0 [6]);
  and _82257_ (_32093_, _12789_, _08012_);
  or _82258_ (_32094_, _32093_, _32092_);
  or _82259_ (_32095_, _32094_, _06132_);
  and _82260_ (_32096_, _13101_, \oc8051_golden_model_1.P0 [6]);
  and _82261_ (_32097_, _30526_, _07847_);
  or _82262_ (_32098_, _32097_, _32096_);
  and _82263_ (_32099_, _32098_, _06152_);
  and _82264_ (_32100_, _30532_, _12789_);
  or _82265_ (_32101_, _32100_, _32092_);
  or _82266_ (_32103_, _32101_, _06161_);
  and _82267_ (_32104_, _12789_, \oc8051_golden_model_1.ACC [6]);
  or _82268_ (_32105_, _32104_, _32092_);
  and _82269_ (_32106_, _32105_, _07056_);
  and _82270_ (_32107_, _07057_, \oc8051_golden_model_1.P0 [6]);
  or _82271_ (_32108_, _32107_, _06160_);
  or _82272_ (_32109_, _32108_, _32106_);
  and _82273_ (_32110_, _32109_, _06157_);
  and _82274_ (_32111_, _32110_, _32103_);
  and _82275_ (_32112_, _30545_, _07847_);
  or _82276_ (_32114_, _32112_, _32096_);
  and _82277_ (_32115_, _32114_, _06156_);
  or _82278_ (_32116_, _32115_, _06217_);
  or _82279_ (_32117_, _32116_, _32111_);
  or _82280_ (_32118_, _32094_, _07075_);
  and _82281_ (_32119_, _32118_, _32117_);
  or _82282_ (_32120_, _32119_, _06220_);
  or _82283_ (_32121_, _32105_, _06229_);
  and _82284_ (_32122_, _32121_, _06153_);
  and _82285_ (_32123_, _32122_, _32120_);
  or _82286_ (_32125_, _32123_, _32099_);
  and _82287_ (_32126_, _32125_, _06146_);
  or _82288_ (_32127_, _32096_, _30560_);
  and _82289_ (_32128_, _32114_, _06145_);
  and _82290_ (_32129_, _32128_, _32127_);
  or _82291_ (_32130_, _32129_, _32126_);
  and _82292_ (_32131_, _32130_, _06140_);
  and _82293_ (_32132_, _30567_, _07847_);
  or _82294_ (_32133_, _32132_, _32096_);
  and _82295_ (_32134_, _32133_, _06139_);
  or _82296_ (_32136_, _32134_, _09842_);
  or _82297_ (_32137_, _32136_, _32131_);
  and _82298_ (_32138_, _32137_, _32095_);
  or _82299_ (_32139_, _32138_, _06116_);
  and _82300_ (_32140_, _12789_, _09207_);
  or _82301_ (_32141_, _32092_, _06117_);
  or _82302_ (_32142_, _32141_, _32140_);
  and _82303_ (_32143_, _32142_, _06114_);
  and _82304_ (_32144_, _32143_, _32139_);
  and _82305_ (_32145_, _30589_, _12789_);
  or _82306_ (_32147_, _32145_, _32092_);
  and _82307_ (_32148_, _32147_, _05787_);
  or _82308_ (_32149_, _32148_, _11136_);
  or _82309_ (_32150_, _32149_, _32144_);
  and _82310_ (_32151_, _30604_, _30601_);
  and _82311_ (_32152_, _32151_, _12789_);
  or _82312_ (_32153_, _32092_, _07127_);
  or _82313_ (_32154_, _32153_, _32152_);
  and _82314_ (_32155_, _12789_, _15402_);
  or _82315_ (_32156_, _32155_, _32092_);
  or _82316_ (_32158_, _32156_, _06111_);
  and _82317_ (_32159_, _32158_, _07125_);
  and _82318_ (_32160_, _32159_, _32154_);
  and _82319_ (_32161_, _32160_, _32150_);
  and _82320_ (_32162_, _30613_, _12789_);
  or _82321_ (_32163_, _32162_, _32092_);
  and _82322_ (_32164_, _32163_, _06402_);
  or _82323_ (_32165_, _32164_, _32161_);
  and _82324_ (_32166_, _32165_, _07132_);
  or _82325_ (_32167_, _32092_, _12810_);
  and _82326_ (_32169_, _32156_, _06306_);
  and _82327_ (_32170_, _32169_, _32167_);
  or _82328_ (_32171_, _32170_, _32166_);
  and _82329_ (_32172_, _32171_, _07130_);
  and _82330_ (_32173_, _32105_, _06411_);
  and _82331_ (_32174_, _32173_, _32167_);
  or _82332_ (_32175_, _32174_, _06303_);
  or _82333_ (_32176_, _32175_, _32172_);
  and _82334_ (_32177_, _30601_, _12789_);
  or _82335_ (_32178_, _32092_, _08819_);
  or _82336_ (_32180_, _32178_, _32177_);
  and _82337_ (_32181_, _32180_, _08824_);
  and _82338_ (_32182_, _32181_, _32176_);
  and _82339_ (_32183_, _30611_, _12789_);
  or _82340_ (_32184_, _32183_, _32092_);
  and _82341_ (_32185_, _32184_, _06396_);
  or _82342_ (_32186_, _32185_, _06433_);
  or _82343_ (_32187_, _32186_, _32182_);
  or _82344_ (_32188_, _32101_, _06829_);
  and _82345_ (_32189_, _32188_, _05749_);
  and _82346_ (_32191_, _32189_, _32187_);
  and _82347_ (_32192_, _32098_, _05748_);
  or _82348_ (_32193_, _32192_, _06440_);
  or _82349_ (_32194_, _32193_, _32191_);
  and _82350_ (_32195_, _30646_, _12789_);
  or _82351_ (_32196_, _32092_, _06444_);
  or _82352_ (_32197_, _32196_, _32195_);
  and _82353_ (_32198_, _32197_, _01317_);
  and _82354_ (_32199_, _32198_, _32194_);
  or _82355_ (_43728_, _32199_, _32090_);
  nor _82356_ (_32201_, \oc8051_golden_model_1.P1 [0], rst);
  nor _82357_ (_32202_, _32201_, _00000_);
  and _82358_ (_32203_, _13196_, \oc8051_golden_model_1.P1 [0]);
  and _82359_ (_32204_, _29675_, _12792_);
  or _82360_ (_32205_, _32204_, _32203_);
  and _82361_ (_32206_, _32205_, _06402_);
  and _82362_ (_32207_, _12792_, _07049_);
  or _82363_ (_32208_, _32207_, _32203_);
  or _82364_ (_32209_, _32208_, _06132_);
  and _82365_ (_32210_, _13201_, \oc8051_golden_model_1.P1 [0]);
  and _82366_ (_32212_, _29705_, _12778_);
  or _82367_ (_32213_, _32212_, _32210_);
  or _82368_ (_32214_, _32213_, _06157_);
  nor _82369_ (_32215_, _12858_, _13196_);
  or _82370_ (_32216_, _32215_, _32203_);
  and _82371_ (_32217_, _32216_, _06160_);
  and _82372_ (_32218_, _07057_, \oc8051_golden_model_1.P1 [0]);
  and _82373_ (_32219_, _12792_, \oc8051_golden_model_1.ACC [0]);
  or _82374_ (_32220_, _32219_, _32203_);
  and _82375_ (_32221_, _32220_, _07056_);
  or _82376_ (_32223_, _32221_, _32218_);
  and _82377_ (_32224_, _32223_, _06161_);
  or _82378_ (_32225_, _32224_, _06156_);
  or _82379_ (_32226_, _32225_, _32217_);
  and _82380_ (_32227_, _32226_, _32214_);
  and _82381_ (_32228_, _32227_, _07075_);
  and _82382_ (_32229_, _32208_, _06217_);
  or _82383_ (_32230_, _32229_, _06220_);
  or _82384_ (_32231_, _32230_, _32228_);
  or _82385_ (_32232_, _32220_, _06229_);
  and _82386_ (_32234_, _32232_, _06153_);
  and _82387_ (_32235_, _32234_, _32231_);
  and _82388_ (_32236_, _32203_, _06152_);
  or _82389_ (_32237_, _32236_, _06145_);
  or _82390_ (_32238_, _32237_, _32235_);
  or _82391_ (_32239_, _32216_, _06146_);
  and _82392_ (_32240_, _32239_, _06140_);
  and _82393_ (_32241_, _32240_, _32238_);
  or _82394_ (_32242_, _32210_, _14170_);
  and _82395_ (_32243_, _32242_, _06139_);
  and _82396_ (_32245_, _32243_, _32213_);
  or _82397_ (_32246_, _32245_, _09842_);
  or _82398_ (_32247_, _32246_, _32241_);
  and _82399_ (_32248_, _32247_, _32209_);
  or _82400_ (_32249_, _32248_, _06116_);
  and _82401_ (_32250_, _12792_, _09160_);
  or _82402_ (_32251_, _32203_, _06117_);
  or _82403_ (_32252_, _32251_, _32250_);
  and _82404_ (_32253_, _32252_, _06114_);
  and _82405_ (_32254_, _32253_, _32249_);
  and _82406_ (_32256_, _29746_, _12792_);
  or _82407_ (_32257_, _32256_, _32203_);
  and _82408_ (_32258_, _32257_, _05787_);
  or _82409_ (_32259_, _32258_, _32254_);
  or _82410_ (_32260_, _32259_, _11136_);
  and _82411_ (_32261_, _29756_, _12792_);
  or _82412_ (_32262_, _32203_, _07127_);
  or _82413_ (_32263_, _32262_, _32261_);
  and _82414_ (_32264_, _12792_, _08708_);
  or _82415_ (_32265_, _32264_, _32203_);
  or _82416_ (_32267_, _32265_, _06111_);
  and _82417_ (_32268_, _32267_, _07125_);
  and _82418_ (_32269_, _32268_, _32263_);
  and _82419_ (_32270_, _32269_, _32260_);
  or _82420_ (_32271_, _32270_, _32206_);
  and _82421_ (_32272_, _32271_, _07132_);
  nand _82422_ (_32273_, _32265_, _06306_);
  nor _82423_ (_32274_, _32273_, _32215_);
  or _82424_ (_32275_, _32274_, _32272_);
  and _82425_ (_32276_, _32275_, _07130_);
  or _82426_ (_32278_, _32203_, _12858_);
  and _82427_ (_32279_, _32220_, _06411_);
  and _82428_ (_32280_, _32279_, _32278_);
  or _82429_ (_32281_, _32280_, _06303_);
  or _82430_ (_32282_, _32281_, _32276_);
  and _82431_ (_32283_, _29752_, _12792_);
  or _82432_ (_32284_, _32203_, _08819_);
  or _82433_ (_32285_, _32284_, _32283_);
  and _82434_ (_32286_, _32285_, _08824_);
  and _82435_ (_32287_, _32286_, _32282_);
  and _82436_ (_32289_, _29673_, _12792_);
  or _82437_ (_32290_, _32289_, _32203_);
  and _82438_ (_32291_, _32290_, _06396_);
  or _82439_ (_32292_, _32291_, _06433_);
  or _82440_ (_32293_, _32292_, _32287_);
  or _82441_ (_32294_, _32216_, _06829_);
  and _82442_ (_32295_, _32294_, _05749_);
  and _82443_ (_32296_, _32295_, _32293_);
  and _82444_ (_32297_, _32203_, _05748_);
  or _82445_ (_32298_, _32297_, _06440_);
  or _82446_ (_32300_, _32298_, _32296_);
  or _82447_ (_32301_, _32216_, _06444_);
  and _82448_ (_32302_, _32301_, _01317_);
  and _82449_ (_32303_, _32302_, _32300_);
  or _82450_ (_43730_, _32303_, _32202_);
  and _82451_ (_32304_, _29814_, _12778_);
  and _82452_ (_32305_, _32304_, _29813_);
  and _82453_ (_32306_, _13201_, \oc8051_golden_model_1.P1 [1]);
  or _82454_ (_32307_, _32306_, _06146_);
  or _82455_ (_32308_, _32307_, _32305_);
  or _82456_ (_32310_, _12792_, \oc8051_golden_model_1.P1 [1]);
  and _82457_ (_32311_, _29823_, _12792_);
  not _82458_ (_32312_, _32311_);
  and _82459_ (_32313_, _32312_, _32310_);
  or _82460_ (_32314_, _32313_, _06161_);
  nand _82461_ (_32315_, _12792_, _05887_);
  and _82462_ (_32316_, _32315_, _32310_);
  and _82463_ (_32317_, _32316_, _07056_);
  and _82464_ (_32318_, _07057_, \oc8051_golden_model_1.P1 [1]);
  or _82465_ (_32319_, _32318_, _06160_);
  or _82466_ (_32321_, _32319_, _32317_);
  and _82467_ (_32322_, _32321_, _06157_);
  and _82468_ (_32323_, _32322_, _32314_);
  or _82469_ (_32324_, _32306_, _06217_);
  or _82470_ (_32325_, _32324_, _32304_);
  and _82471_ (_32326_, _32325_, _13860_);
  or _82472_ (_32327_, _32326_, _32323_);
  and _82473_ (_32328_, _13196_, \oc8051_golden_model_1.P1 [1]);
  and _82474_ (_32329_, _12792_, _07306_);
  or _82475_ (_32330_, _32329_, _32328_);
  or _82476_ (_32332_, _32330_, _07075_);
  and _82477_ (_32333_, _32332_, _32327_);
  or _82478_ (_32334_, _32333_, _06220_);
  or _82479_ (_32335_, _32316_, _06229_);
  and _82480_ (_32336_, _32335_, _06153_);
  and _82481_ (_32337_, _32336_, _32334_);
  and _82482_ (_32338_, _29851_, _12778_);
  or _82483_ (_32339_, _32338_, _32306_);
  and _82484_ (_32340_, _32339_, _06152_);
  or _82485_ (_32341_, _32340_, _06145_);
  or _82486_ (_32343_, _32341_, _32337_);
  and _82487_ (_32344_, _32343_, _32308_);
  and _82488_ (_32345_, _32344_, _06140_);
  and _82489_ (_32346_, _29860_, _12778_);
  or _82490_ (_32347_, _32306_, _32346_);
  and _82491_ (_32348_, _32347_, _06139_);
  or _82492_ (_32349_, _32348_, _09842_);
  or _82493_ (_32350_, _32349_, _32345_);
  or _82494_ (_32351_, _32330_, _06132_);
  and _82495_ (_32352_, _32351_, _32350_);
  or _82496_ (_32354_, _32352_, _06116_);
  and _82497_ (_32355_, _12792_, _09115_);
  or _82498_ (_32356_, _32328_, _06117_);
  or _82499_ (_32357_, _32356_, _32355_);
  and _82500_ (_32358_, _32357_, _06114_);
  and _82501_ (_32359_, _32358_, _32354_);
  and _82502_ (_32360_, _29883_, _12792_);
  or _82503_ (_32361_, _32360_, _32328_);
  and _82504_ (_32362_, _32361_, _05787_);
  or _82505_ (_32363_, _32362_, _32359_);
  and _82506_ (_32365_, _32363_, _06298_);
  or _82507_ (_32366_, _30823_, _13196_);
  and _82508_ (_32367_, _32366_, _06297_);
  nand _82509_ (_32368_, _12792_, _06945_);
  and _82510_ (_32369_, _32368_, _06110_);
  or _82511_ (_32370_, _32369_, _32367_);
  and _82512_ (_32371_, _32370_, _32310_);
  or _82513_ (_32372_, _32371_, _32365_);
  and _82514_ (_32373_, _32372_, _07125_);
  or _82515_ (_32374_, _30833_, _13196_);
  and _82516_ (_32376_, _32310_, _06402_);
  and _82517_ (_32377_, _32376_, _32374_);
  or _82518_ (_32378_, _32377_, _32373_);
  and _82519_ (_32379_, _32378_, _07132_);
  or _82520_ (_32380_, _29896_, _13196_);
  and _82521_ (_32381_, _32310_, _06306_);
  and _82522_ (_32382_, _32381_, _32380_);
  or _82523_ (_32383_, _32382_, _32379_);
  and _82524_ (_32384_, _32383_, _07130_);
  or _82525_ (_32385_, _32328_, _12850_);
  and _82526_ (_32387_, _32316_, _06411_);
  and _82527_ (_32388_, _32387_, _32385_);
  or _82528_ (_32389_, _32388_, _32384_);
  and _82529_ (_32390_, _32389_, _06397_);
  or _82530_ (_32391_, _32368_, _12850_);
  and _82531_ (_32392_, _32310_, _06303_);
  and _82532_ (_32393_, _32392_, _32391_);
  or _82533_ (_32394_, _32315_, _12850_);
  and _82534_ (_32395_, _32310_, _06396_);
  and _82535_ (_32396_, _32395_, _32394_);
  or _82536_ (_32398_, _32396_, _06433_);
  or _82537_ (_32399_, _32398_, _32393_);
  or _82538_ (_32400_, _32399_, _32390_);
  or _82539_ (_32401_, _32313_, _06829_);
  and _82540_ (_32402_, _32401_, _05749_);
  and _82541_ (_32403_, _32402_, _32400_);
  and _82542_ (_32404_, _32339_, _05748_);
  or _82543_ (_32405_, _32404_, _06440_);
  or _82544_ (_32406_, _32405_, _32403_);
  or _82545_ (_32407_, _32328_, _06444_);
  or _82546_ (_32409_, _32407_, _32311_);
  and _82547_ (_32410_, _32409_, _01317_);
  and _82548_ (_32411_, _32410_, _32406_);
  nor _82549_ (_32412_, \oc8051_golden_model_1.P1 [1], rst);
  nor _82550_ (_32413_, _32412_, _00000_);
  or _82551_ (_43731_, _32413_, _32411_);
  and _82552_ (_32414_, _13196_, \oc8051_golden_model_1.P1 [2]);
  and _82553_ (_32415_, _12792_, _07708_);
  or _82554_ (_32416_, _32415_, _32414_);
  or _82555_ (_32417_, _32416_, _06132_);
  and _82556_ (_32419_, _29954_, _12792_);
  or _82557_ (_32420_, _32419_, _32414_);
  or _82558_ (_32421_, _32420_, _06161_);
  and _82559_ (_32422_, _12792_, \oc8051_golden_model_1.ACC [2]);
  or _82560_ (_32423_, _32422_, _32414_);
  and _82561_ (_32424_, _32423_, _07056_);
  and _82562_ (_32425_, _07057_, \oc8051_golden_model_1.P1 [2]);
  or _82563_ (_32426_, _32425_, _06160_);
  or _82564_ (_32427_, _32426_, _32424_);
  and _82565_ (_32428_, _32427_, _06157_);
  and _82566_ (_32430_, _32428_, _32421_);
  and _82567_ (_32431_, _13201_, \oc8051_golden_model_1.P1 [2]);
  and _82568_ (_32432_, _29976_, _12778_);
  or _82569_ (_32433_, _32432_, _32431_);
  and _82570_ (_32434_, _32433_, _06156_);
  or _82571_ (_32435_, _32434_, _06217_);
  or _82572_ (_32436_, _32435_, _32430_);
  or _82573_ (_32437_, _32416_, _07075_);
  and _82574_ (_32438_, _32437_, _32436_);
  or _82575_ (_32439_, _32438_, _06220_);
  or _82576_ (_32441_, _32423_, _06229_);
  and _82577_ (_32442_, _32441_, _06153_);
  and _82578_ (_32443_, _32442_, _32439_);
  and _82579_ (_32444_, _29992_, _12778_);
  or _82580_ (_32445_, _32444_, _32431_);
  and _82581_ (_32446_, _32445_, _06152_);
  or _82582_ (_32447_, _32446_, _06145_);
  or _82583_ (_32448_, _32447_, _32443_);
  or _82584_ (_32449_, _32431_, _29999_);
  and _82585_ (_32450_, _32449_, _32433_);
  or _82586_ (_32452_, _32450_, _06146_);
  and _82587_ (_32453_, _32452_, _06140_);
  and _82588_ (_32454_, _32453_, _32448_);
  and _82589_ (_32455_, _30005_, _12778_);
  or _82590_ (_32456_, _32455_, _32431_);
  and _82591_ (_32457_, _32456_, _06139_);
  or _82592_ (_32458_, _32457_, _09842_);
  or _82593_ (_32459_, _32458_, _32454_);
  and _82594_ (_32460_, _32459_, _32417_);
  or _82595_ (_32461_, _32460_, _06116_);
  and _82596_ (_32463_, _12792_, _09211_);
  or _82597_ (_32464_, _32414_, _06117_);
  or _82598_ (_32465_, _32464_, _32463_);
  and _82599_ (_32466_, _32465_, _06114_);
  and _82600_ (_32467_, _32466_, _32461_);
  and _82601_ (_32468_, _30029_, _12792_);
  or _82602_ (_32469_, _32414_, _32468_);
  and _82603_ (_32470_, _32469_, _05787_);
  or _82604_ (_32471_, _32470_, _32467_);
  or _82605_ (_32472_, _32471_, _11136_);
  and _82606_ (_32474_, _31708_, _12792_);
  or _82607_ (_32475_, _32414_, _07127_);
  or _82608_ (_32476_, _32475_, _32474_);
  and _82609_ (_32477_, _12792_, _08768_);
  or _82610_ (_32478_, _32477_, _32414_);
  or _82611_ (_32479_, _32478_, _06111_);
  and _82612_ (_32480_, _32479_, _07125_);
  and _82613_ (_32481_, _32480_, _32476_);
  and _82614_ (_32482_, _32481_, _32472_);
  and _82615_ (_32483_, _30043_, _12792_);
  or _82616_ (_32485_, _32483_, _32414_);
  or _82617_ (_32486_, _32414_, _30046_);
  and _82618_ (_32487_, _32486_, _06402_);
  and _82619_ (_32488_, _32487_, _32485_);
  or _82620_ (_32489_, _32488_, _32482_);
  and _82621_ (_32490_, _32489_, _07132_);
  or _82622_ (_32491_, _32414_, _12842_);
  and _82623_ (_32492_, _32478_, _06306_);
  and _82624_ (_32493_, _32492_, _32491_);
  or _82625_ (_32494_, _32493_, _32490_);
  and _82626_ (_32496_, _32494_, _07130_);
  and _82627_ (_32497_, _32423_, _06411_);
  and _82628_ (_32498_, _32497_, _32491_);
  or _82629_ (_32499_, _32498_, _06303_);
  or _82630_ (_32500_, _32499_, _32496_);
  and _82631_ (_32501_, _29945_, _12792_);
  or _82632_ (_32502_, _32414_, _08819_);
  or _82633_ (_32503_, _32502_, _32501_);
  and _82634_ (_32504_, _32503_, _08824_);
  and _82635_ (_32505_, _32504_, _32500_);
  and _82636_ (_32507_, _32485_, _06396_);
  or _82637_ (_32508_, _32507_, _06433_);
  or _82638_ (_32509_, _32508_, _32505_);
  or _82639_ (_32510_, _32420_, _06829_);
  and _82640_ (_32511_, _32510_, _05749_);
  and _82641_ (_32512_, _32511_, _32509_);
  and _82642_ (_32513_, _32445_, _05748_);
  or _82643_ (_32514_, _32513_, _06440_);
  or _82644_ (_32515_, _32514_, _32512_);
  and _82645_ (_32516_, _30077_, _12792_);
  or _82646_ (_32518_, _32414_, _06444_);
  or _82647_ (_32519_, _32518_, _32516_);
  and _82648_ (_32520_, _32519_, _01317_);
  and _82649_ (_32521_, _32520_, _32515_);
  nor _82650_ (_32522_, \oc8051_golden_model_1.P1 [2], rst);
  nor _82651_ (_32523_, _32522_, _00000_);
  or _82652_ (_43732_, _32523_, _32521_);
  nor _82653_ (_32524_, \oc8051_golden_model_1.P1 [3], rst);
  nor _82654_ (_32525_, _32524_, _00000_);
  and _82655_ (_32526_, _13196_, \oc8051_golden_model_1.P1 [3]);
  and _82656_ (_32528_, _12792_, _07544_);
  or _82657_ (_32529_, _32528_, _32526_);
  or _82658_ (_32530_, _32529_, _06132_);
  and _82659_ (_32531_, _13201_, \oc8051_golden_model_1.P1 [3]);
  and _82660_ (_32532_, _30100_, _12778_);
  or _82661_ (_32533_, _32532_, _32531_);
  and _82662_ (_32534_, _32533_, _06152_);
  and _82663_ (_32535_, _30106_, _12792_);
  or _82664_ (_32536_, _32535_, _32526_);
  or _82665_ (_32537_, _32536_, _06161_);
  and _82666_ (_32539_, _12792_, \oc8051_golden_model_1.ACC [3]);
  or _82667_ (_32540_, _32539_, _32526_);
  and _82668_ (_32541_, _32540_, _07056_);
  and _82669_ (_32542_, _07057_, \oc8051_golden_model_1.P1 [3]);
  or _82670_ (_32543_, _32542_, _06160_);
  or _82671_ (_32544_, _32543_, _32541_);
  and _82672_ (_32545_, _32544_, _06157_);
  and _82673_ (_32546_, _32545_, _32537_);
  and _82674_ (_32547_, _30119_, _12778_);
  or _82675_ (_32548_, _32547_, _32531_);
  and _82676_ (_32550_, _32548_, _06156_);
  or _82677_ (_32551_, _32550_, _06217_);
  or _82678_ (_32552_, _32551_, _32546_);
  or _82679_ (_32553_, _32529_, _07075_);
  and _82680_ (_32554_, _32553_, _32552_);
  or _82681_ (_32555_, _32554_, _06220_);
  or _82682_ (_32556_, _32540_, _06229_);
  and _82683_ (_32557_, _32556_, _06153_);
  and _82684_ (_32558_, _32557_, _32555_);
  or _82685_ (_32559_, _32558_, _32534_);
  and _82686_ (_32561_, _32559_, _06146_);
  or _82687_ (_32562_, _32531_, _30134_);
  and _82688_ (_32563_, _32548_, _06145_);
  and _82689_ (_32564_, _32563_, _32562_);
  or _82690_ (_32565_, _32564_, _32561_);
  and _82691_ (_32566_, _32565_, _06140_);
  and _82692_ (_32567_, _30141_, _12778_);
  or _82693_ (_32568_, _32567_, _32531_);
  and _82694_ (_32569_, _32568_, _06139_);
  or _82695_ (_32570_, _32569_, _09842_);
  or _82696_ (_32572_, _32570_, _32566_);
  and _82697_ (_32573_, _32572_, _32530_);
  or _82698_ (_32574_, _32573_, _06116_);
  and _82699_ (_32575_, _12792_, _09210_);
  or _82700_ (_32576_, _32526_, _06117_);
  or _82701_ (_32577_, _32576_, _32575_);
  and _82702_ (_32578_, _32577_, _06114_);
  and _82703_ (_32579_, _32578_, _32574_);
  and _82704_ (_32580_, _30163_, _12792_);
  or _82705_ (_32581_, _32580_, _32526_);
  and _82706_ (_32583_, _32581_, _05787_);
  or _82707_ (_32584_, _32583_, _11136_);
  or _82708_ (_32585_, _32584_, _32579_);
  and _82709_ (_32586_, _31042_, _12792_);
  or _82710_ (_32587_, _32526_, _07127_);
  or _82711_ (_32588_, _32587_, _32586_);
  and _82712_ (_32589_, _12792_, _08712_);
  or _82713_ (_32590_, _32589_, _32526_);
  or _82714_ (_32591_, _32590_, _06111_);
  and _82715_ (_32592_, _32591_, _07125_);
  and _82716_ (_32594_, _32592_, _32588_);
  and _82717_ (_32595_, _32594_, _32585_);
  and _82718_ (_32596_, _31053_, _12792_);
  or _82719_ (_32597_, _32596_, _32526_);
  and _82720_ (_32598_, _32597_, _06402_);
  or _82721_ (_32599_, _32598_, _32595_);
  and _82722_ (_32600_, _32599_, _07132_);
  or _82723_ (_32601_, _32526_, _12834_);
  and _82724_ (_32602_, _32590_, _06306_);
  and _82725_ (_32603_, _32602_, _32601_);
  or _82726_ (_32605_, _32603_, _32600_);
  and _82727_ (_32606_, _32605_, _07130_);
  and _82728_ (_32607_, _32540_, _06411_);
  and _82729_ (_32608_, _32607_, _32601_);
  or _82730_ (_32609_, _32608_, _06303_);
  or _82731_ (_32610_, _32609_, _32606_);
  and _82732_ (_32611_, _30175_, _12792_);
  or _82733_ (_32612_, _32526_, _08819_);
  or _82734_ (_32613_, _32612_, _32611_);
  and _82735_ (_32614_, _32613_, _08824_);
  and _82736_ (_32616_, _32614_, _32610_);
  and _82737_ (_32617_, _30185_, _12792_);
  or _82738_ (_32618_, _32617_, _32526_);
  and _82739_ (_32619_, _32618_, _06396_);
  or _82740_ (_32620_, _32619_, _06433_);
  or _82741_ (_32621_, _32620_, _32616_);
  or _82742_ (_32622_, _32536_, _06829_);
  and _82743_ (_32623_, _32622_, _05749_);
  and _82744_ (_32624_, _32623_, _32621_);
  and _82745_ (_32625_, _32533_, _05748_);
  or _82746_ (_32627_, _32625_, _06440_);
  or _82747_ (_32628_, _32627_, _32624_);
  and _82748_ (_32629_, _30219_, _12792_);
  or _82749_ (_32630_, _32526_, _06444_);
  or _82750_ (_32631_, _32630_, _32629_);
  and _82751_ (_32632_, _32631_, _01317_);
  and _82752_ (_32633_, _32632_, _32628_);
  or _82753_ (_43733_, _32633_, _32525_);
  and _82754_ (_32634_, _13196_, \oc8051_golden_model_1.P1 [4]);
  and _82755_ (_32635_, _12792_, _08336_);
  or _82756_ (_32637_, _32635_, _32634_);
  or _82757_ (_32638_, _32637_, _06132_);
  and _82758_ (_32639_, _13201_, \oc8051_golden_model_1.P1 [4]);
  and _82759_ (_32640_, _30242_, _12778_);
  or _82760_ (_32641_, _32640_, _32639_);
  and _82761_ (_32642_, _32641_, _06152_);
  and _82762_ (_32643_, _30248_, _12792_);
  or _82763_ (_32644_, _32643_, _32634_);
  or _82764_ (_32645_, _32644_, _06161_);
  and _82765_ (_32646_, _12792_, \oc8051_golden_model_1.ACC [4]);
  or _82766_ (_32648_, _32646_, _32634_);
  and _82767_ (_32649_, _32648_, _07056_);
  and _82768_ (_32650_, _07057_, \oc8051_golden_model_1.P1 [4]);
  or _82769_ (_32651_, _32650_, _06160_);
  or _82770_ (_32652_, _32651_, _32649_);
  and _82771_ (_32653_, _32652_, _06157_);
  and _82772_ (_32654_, _32653_, _32645_);
  and _82773_ (_32655_, _30261_, _12778_);
  or _82774_ (_32656_, _32655_, _32639_);
  and _82775_ (_32657_, _32656_, _06156_);
  or _82776_ (_32659_, _32657_, _06217_);
  or _82777_ (_32660_, _32659_, _32654_);
  or _82778_ (_32661_, _32637_, _07075_);
  and _82779_ (_32662_, _32661_, _32660_);
  or _82780_ (_32663_, _32662_, _06220_);
  or _82781_ (_32664_, _32648_, _06229_);
  and _82782_ (_32665_, _32664_, _06153_);
  and _82783_ (_32666_, _32665_, _32663_);
  or _82784_ (_32667_, _32666_, _32642_);
  and _82785_ (_32668_, _32667_, _06146_);
  or _82786_ (_32670_, _32639_, _30276_);
  and _82787_ (_32671_, _32656_, _06145_);
  and _82788_ (_32672_, _32671_, _32670_);
  or _82789_ (_32673_, _32672_, _32668_);
  and _82790_ (_32674_, _32673_, _06140_);
  and _82791_ (_32675_, _30283_, _12778_);
  or _82792_ (_32676_, _32675_, _32639_);
  and _82793_ (_32677_, _32676_, _06139_);
  or _82794_ (_32678_, _32677_, _09842_);
  or _82795_ (_32679_, _32678_, _32674_);
  and _82796_ (_32681_, _32679_, _32638_);
  or _82797_ (_32682_, _32681_, _06116_);
  and _82798_ (_32683_, _12792_, _09209_);
  or _82799_ (_32684_, _32634_, _06117_);
  or _82800_ (_32685_, _32684_, _32683_);
  and _82801_ (_32686_, _32685_, _06114_);
  and _82802_ (_32687_, _32686_, _32682_);
  and _82803_ (_32688_, _30305_, _12792_);
  or _82804_ (_32689_, _32688_, _32634_);
  and _82805_ (_32690_, _32689_, _05787_);
  or _82806_ (_32691_, _32690_, _06110_);
  or _82807_ (_32692_, _32691_, _32687_);
  and _82808_ (_32693_, _12792_, _08715_);
  or _82809_ (_32694_, _32693_, _32634_);
  or _82810_ (_32695_, _32694_, _06111_);
  and _82811_ (_32696_, _32695_, _07127_);
  and _82812_ (_32697_, _32696_, _32692_);
  and _82813_ (_32698_, _30317_, _12792_);
  or _82814_ (_32699_, _32698_, _32634_);
  or _82815_ (_32700_, _32634_, _30320_);
  and _82816_ (_32702_, _32700_, _06297_);
  and _82817_ (_32703_, _32702_, _32699_);
  or _82818_ (_32704_, _32703_, _06402_);
  or _82819_ (_32705_, _32704_, _32697_);
  and _82820_ (_32706_, _31172_, _12792_);
  or _82821_ (_32707_, _32634_, _07125_);
  or _82822_ (_32708_, _32707_, _32706_);
  and _82823_ (_32709_, _32708_, _07132_);
  and _82824_ (_32710_, _32709_, _32705_);
  or _82825_ (_32711_, _32634_, _12826_);
  and _82826_ (_32713_, _32694_, _06306_);
  and _82827_ (_32714_, _32713_, _32711_);
  or _82828_ (_32715_, _32714_, _32710_);
  and _82829_ (_32716_, _32715_, _07130_);
  and _82830_ (_32717_, _32648_, _06411_);
  and _82831_ (_32718_, _32717_, _32711_);
  or _82832_ (_32719_, _32718_, _06303_);
  or _82833_ (_32720_, _32719_, _32716_);
  or _82834_ (_32721_, _32699_, _08819_);
  and _82835_ (_32722_, _32721_, _08824_);
  and _82836_ (_32724_, _32722_, _32720_);
  and _82837_ (_32725_, _30327_, _12792_);
  or _82838_ (_32726_, _32725_, _32634_);
  and _82839_ (_32727_, _32726_, _06396_);
  or _82840_ (_32728_, _32727_, _06433_);
  or _82841_ (_32729_, _32728_, _32724_);
  or _82842_ (_32730_, _32644_, _06829_);
  and _82843_ (_32731_, _32730_, _05749_);
  and _82844_ (_32732_, _32731_, _32729_);
  and _82845_ (_32733_, _32641_, _05748_);
  or _82846_ (_32735_, _32733_, _06440_);
  or _82847_ (_32736_, _32735_, _32732_);
  and _82848_ (_32737_, _30361_, _12792_);
  or _82849_ (_32738_, _32634_, _06444_);
  or _82850_ (_32739_, _32738_, _32737_);
  and _82851_ (_32740_, _32739_, _01317_);
  and _82852_ (_32741_, _32740_, _32736_);
  nor _82853_ (_32742_, \oc8051_golden_model_1.P1 [4], rst);
  nor _82854_ (_32743_, _32742_, _00000_);
  or _82855_ (_43734_, _32743_, _32741_);
  and _82856_ (_32745_, _13196_, \oc8051_golden_model_1.P1 [5]);
  and _82857_ (_32746_, _12792_, _08101_);
  or _82858_ (_32747_, _32746_, _32745_);
  or _82859_ (_32748_, _32747_, _06132_);
  and _82860_ (_32749_, _30378_, _12792_);
  or _82861_ (_32750_, _32749_, _32745_);
  or _82862_ (_32751_, _32750_, _06161_);
  and _82863_ (_32752_, _12792_, \oc8051_golden_model_1.ACC [5]);
  or _82864_ (_32753_, _32752_, _32745_);
  and _82865_ (_32754_, _32753_, _07056_);
  and _82866_ (_32756_, _07057_, \oc8051_golden_model_1.P1 [5]);
  or _82867_ (_32757_, _32756_, _06160_);
  or _82868_ (_32758_, _32757_, _32754_);
  and _82869_ (_32759_, _32758_, _06157_);
  and _82870_ (_32760_, _32759_, _32751_);
  and _82871_ (_32761_, _13201_, \oc8051_golden_model_1.P1 [5]);
  and _82872_ (_32762_, _30400_, _12778_);
  or _82873_ (_32763_, _32762_, _32761_);
  and _82874_ (_32764_, _32763_, _06156_);
  or _82875_ (_32765_, _32764_, _06217_);
  or _82876_ (_32767_, _32765_, _32760_);
  or _82877_ (_32768_, _32747_, _07075_);
  and _82878_ (_32769_, _32768_, _32767_);
  or _82879_ (_32770_, _32769_, _06220_);
  or _82880_ (_32771_, _32753_, _06229_);
  and _82881_ (_32772_, _32771_, _06153_);
  and _82882_ (_32773_, _32772_, _32770_);
  and _82883_ (_32774_, _30414_, _12778_);
  or _82884_ (_32775_, _32774_, _32761_);
  and _82885_ (_32776_, _32775_, _06152_);
  or _82886_ (_32778_, _32776_, _06145_);
  or _82887_ (_32779_, _32778_, _32773_);
  or _82888_ (_32780_, _32761_, _30420_);
  and _82889_ (_32781_, _32780_, _32763_);
  or _82890_ (_32782_, _32781_, _06146_);
  and _82891_ (_32783_, _32782_, _06140_);
  and _82892_ (_32784_, _32783_, _32779_);
  and _82893_ (_32785_, _30426_, _12778_);
  or _82894_ (_32786_, _32785_, _32761_);
  and _82895_ (_32787_, _32786_, _06139_);
  or _82896_ (_32789_, _32787_, _09842_);
  or _82897_ (_32790_, _32789_, _32784_);
  and _82898_ (_32791_, _32790_, _32748_);
  or _82899_ (_32792_, _32791_, _06116_);
  and _82900_ (_32793_, _12792_, _09208_);
  or _82901_ (_32794_, _32745_, _06117_);
  or _82902_ (_32795_, _32794_, _32793_);
  and _82903_ (_32796_, _32795_, _06114_);
  and _82904_ (_32797_, _32796_, _32792_);
  and _82905_ (_32798_, _30449_, _12792_);
  or _82906_ (_32800_, _32798_, _32745_);
  and _82907_ (_32801_, _32800_, _05787_);
  or _82908_ (_32802_, _32801_, _11136_);
  or _82909_ (_32803_, _32802_, _32797_);
  and _82910_ (_32804_, _32036_, _12792_);
  or _82911_ (_32805_, _32745_, _07127_);
  or _82912_ (_32806_, _32805_, _32804_);
  and _82913_ (_32807_, _12792_, _08736_);
  or _82914_ (_32808_, _32807_, _32745_);
  or _82915_ (_32809_, _32808_, _06111_);
  and _82916_ (_32811_, _32809_, _07125_);
  and _82917_ (_32812_, _32811_, _32806_);
  and _82918_ (_32813_, _32812_, _32803_);
  and _82919_ (_32814_, _32047_, _12792_);
  or _82920_ (_32815_, _32814_, _32745_);
  and _82921_ (_32816_, _32815_, _06402_);
  or _82922_ (_32817_, _32816_, _32813_);
  and _82923_ (_32818_, _32817_, _07132_);
  or _82924_ (_32819_, _32745_, _12818_);
  and _82925_ (_32820_, _32808_, _06306_);
  and _82926_ (_32822_, _32820_, _32819_);
  or _82927_ (_32823_, _32822_, _32818_);
  and _82928_ (_32824_, _32823_, _07130_);
  and _82929_ (_32825_, _32753_, _06411_);
  and _82930_ (_32826_, _32825_, _32819_);
  or _82931_ (_32827_, _32826_, _06303_);
  or _82932_ (_32828_, _32827_, _32824_);
  and _82933_ (_32829_, _30461_, _12792_);
  or _82934_ (_32830_, _32745_, _08819_);
  or _82935_ (_32831_, _32830_, _32829_);
  and _82936_ (_32833_, _32831_, _08824_);
  and _82937_ (_32834_, _32833_, _32828_);
  and _82938_ (_32835_, _30471_, _12792_);
  or _82939_ (_32836_, _32835_, _32745_);
  and _82940_ (_32837_, _32836_, _06396_);
  or _82941_ (_32838_, _32837_, _06433_);
  or _82942_ (_32839_, _32838_, _32834_);
  or _82943_ (_32840_, _32750_, _06829_);
  and _82944_ (_32841_, _32840_, _05749_);
  and _82945_ (_32842_, _32841_, _32839_);
  and _82946_ (_32844_, _32775_, _05748_);
  or _82947_ (_32845_, _32844_, _06440_);
  or _82948_ (_32846_, _32845_, _32842_);
  and _82949_ (_32847_, _30505_, _12792_);
  or _82950_ (_32848_, _32745_, _06444_);
  or _82951_ (_32849_, _32848_, _32847_);
  and _82952_ (_32850_, _32849_, _01317_);
  and _82953_ (_32851_, _32850_, _32846_);
  nor _82954_ (_32852_, \oc8051_golden_model_1.P1 [5], rst);
  nor _82955_ (_32853_, _32852_, _00000_);
  or _82956_ (_43735_, _32853_, _32851_);
  and _82957_ (_32855_, _13196_, \oc8051_golden_model_1.P1 [6]);
  and _82958_ (_32856_, _12792_, _08012_);
  or _82959_ (_32857_, _32856_, _32855_);
  or _82960_ (_32858_, _32857_, _06132_);
  and _82961_ (_32859_, _13201_, \oc8051_golden_model_1.P1 [6]);
  and _82962_ (_32860_, _30526_, _12778_);
  or _82963_ (_32861_, _32860_, _32859_);
  and _82964_ (_32862_, _32861_, _06152_);
  and _82965_ (_32863_, _30532_, _12792_);
  or _82966_ (_32865_, _32863_, _32855_);
  or _82967_ (_32866_, _32865_, _06161_);
  and _82968_ (_32867_, _12792_, \oc8051_golden_model_1.ACC [6]);
  or _82969_ (_32868_, _32867_, _32855_);
  and _82970_ (_32869_, _32868_, _07056_);
  and _82971_ (_32870_, _07057_, \oc8051_golden_model_1.P1 [6]);
  or _82972_ (_32871_, _32870_, _06160_);
  or _82973_ (_32872_, _32871_, _32869_);
  and _82974_ (_32873_, _32872_, _06157_);
  and _82975_ (_32874_, _32873_, _32866_);
  and _82976_ (_32876_, _30545_, _12778_);
  or _82977_ (_32877_, _32876_, _32859_);
  and _82978_ (_32878_, _32877_, _06156_);
  or _82979_ (_32879_, _32878_, _06217_);
  or _82980_ (_32880_, _32879_, _32874_);
  or _82981_ (_32881_, _32857_, _07075_);
  and _82982_ (_32882_, _32881_, _32880_);
  or _82983_ (_32883_, _32882_, _06220_);
  or _82984_ (_32884_, _32868_, _06229_);
  and _82985_ (_32885_, _32884_, _06153_);
  and _82986_ (_32887_, _32885_, _32883_);
  or _82987_ (_32888_, _32887_, _32862_);
  and _82988_ (_32889_, _32888_, _06146_);
  or _82989_ (_32890_, _32859_, _30560_);
  and _82990_ (_32891_, _32877_, _06145_);
  and _82991_ (_32892_, _32891_, _32890_);
  or _82992_ (_32893_, _32892_, _32889_);
  and _82993_ (_32894_, _32893_, _06140_);
  and _82994_ (_32895_, _30567_, _12778_);
  or _82995_ (_32896_, _32895_, _32859_);
  and _82996_ (_32898_, _32896_, _06139_);
  or _82997_ (_32899_, _32898_, _09842_);
  or _82998_ (_32900_, _32899_, _32894_);
  and _82999_ (_32901_, _32900_, _32858_);
  or _83000_ (_32902_, _32901_, _06116_);
  and _83001_ (_32903_, _12792_, _09207_);
  or _83002_ (_32904_, _32855_, _06117_);
  or _83003_ (_32905_, _32904_, _32903_);
  and _83004_ (_32906_, _32905_, _06114_);
  and _83005_ (_32907_, _32906_, _32902_);
  and _83006_ (_32909_, _30589_, _12792_);
  or _83007_ (_32910_, _32909_, _32855_);
  and _83008_ (_32911_, _32910_, _05787_);
  or _83009_ (_32912_, _32911_, _11136_);
  or _83010_ (_32913_, _32912_, _32907_);
  and _83011_ (_32914_, _32151_, _12792_);
  or _83012_ (_32915_, _32855_, _07127_);
  or _83013_ (_32916_, _32915_, _32914_);
  and _83014_ (_32917_, _12792_, _15402_);
  or _83015_ (_32918_, _32917_, _32855_);
  or _83016_ (_32920_, _32918_, _06111_);
  and _83017_ (_32921_, _32920_, _07125_);
  and _83018_ (_32922_, _32921_, _32916_);
  and _83019_ (_32923_, _32922_, _32913_);
  and _83020_ (_32924_, _30613_, _12792_);
  or _83021_ (_32925_, _32924_, _32855_);
  and _83022_ (_32926_, _32925_, _06402_);
  or _83023_ (_32927_, _32926_, _32923_);
  and _83024_ (_32928_, _32927_, _07132_);
  or _83025_ (_32929_, _32855_, _12810_);
  and _83026_ (_32931_, _32918_, _06306_);
  and _83027_ (_32932_, _32931_, _32929_);
  or _83028_ (_32933_, _32932_, _32928_);
  and _83029_ (_32934_, _32933_, _07130_);
  and _83030_ (_32935_, _32868_, _06411_);
  and _83031_ (_32936_, _32935_, _32929_);
  or _83032_ (_32937_, _32936_, _06303_);
  or _83033_ (_32938_, _32937_, _32934_);
  and _83034_ (_32939_, _30601_, _12792_);
  or _83035_ (_32940_, _32855_, _08819_);
  or _83036_ (_32942_, _32940_, _32939_);
  and _83037_ (_32943_, _32942_, _08824_);
  and _83038_ (_32944_, _32943_, _32938_);
  and _83039_ (_32945_, _30611_, _12792_);
  or _83040_ (_32946_, _32945_, _32855_);
  and _83041_ (_32947_, _32946_, _06396_);
  or _83042_ (_32948_, _32947_, _06433_);
  or _83043_ (_32949_, _32948_, _32944_);
  or _83044_ (_32950_, _32865_, _06829_);
  and _83045_ (_32951_, _32950_, _05749_);
  and _83046_ (_32953_, _32951_, _32949_);
  and _83047_ (_32954_, _32861_, _05748_);
  or _83048_ (_32955_, _32954_, _06440_);
  or _83049_ (_32956_, _32955_, _32953_);
  and _83050_ (_32957_, _30646_, _12792_);
  or _83051_ (_32958_, _32855_, _06444_);
  or _83052_ (_32959_, _32958_, _32957_);
  and _83053_ (_32960_, _32959_, _01317_);
  and _83054_ (_32961_, _32960_, _32956_);
  nor _83055_ (_32962_, \oc8051_golden_model_1.P1 [6], rst);
  nor _83056_ (_32964_, _32962_, _00000_);
  or _83057_ (_43736_, _32964_, _32961_);
  not _83058_ (_32965_, \oc8051_golden_model_1.IP [0]);
  nor _83059_ (_32966_, _01317_, _32965_);
  nand _83060_ (_32967_, _10276_, _07830_);
  nor _83061_ (_32968_, _07830_, _32965_);
  nor _83062_ (_32969_, _32968_, _07130_);
  nand _83063_ (_32970_, _32969_, _32967_);
  and _83064_ (_32971_, _07830_, _07049_);
  or _83065_ (_32972_, _32971_, _32968_);
  or _83066_ (_32974_, _32972_, _06132_);
  nor _83067_ (_32975_, _08211_, _13300_);
  or _83068_ (_32976_, _32975_, _32968_);
  or _83069_ (_32977_, _32976_, _06161_);
  and _83070_ (_32978_, _07830_, \oc8051_golden_model_1.ACC [0]);
  or _83071_ (_32979_, _32978_, _32968_);
  and _83072_ (_32980_, _32979_, _07056_);
  nor _83073_ (_32981_, _07056_, _32965_);
  or _83074_ (_32982_, _32981_, _06160_);
  or _83075_ (_32983_, _32982_, _32980_);
  and _83076_ (_32985_, _32983_, _06157_);
  and _83077_ (_32986_, _32985_, _32977_);
  nor _83078_ (_32987_, _08415_, _32965_);
  and _83079_ (_32988_, _14169_, _08415_);
  or _83080_ (_32989_, _32988_, _32987_);
  and _83081_ (_32990_, _32989_, _06156_);
  or _83082_ (_32991_, _32990_, _32986_);
  and _83083_ (_32992_, _32991_, _07075_);
  and _83084_ (_32993_, _32972_, _06217_);
  or _83085_ (_32994_, _32993_, _06220_);
  or _83086_ (_32996_, _32994_, _32992_);
  or _83087_ (_32997_, _32979_, _06229_);
  and _83088_ (_32998_, _32997_, _06153_);
  and _83089_ (_32999_, _32998_, _32996_);
  and _83090_ (_33000_, _32968_, _06152_);
  or _83091_ (_33001_, _33000_, _06145_);
  or _83092_ (_33002_, _33001_, _32999_);
  or _83093_ (_33003_, _32976_, _06146_);
  and _83094_ (_33004_, _33003_, _06140_);
  and _83095_ (_33005_, _33004_, _33002_);
  or _83096_ (_33007_, _32987_, _14170_);
  and _83097_ (_33008_, _33007_, _06139_);
  and _83098_ (_33009_, _33008_, _32989_);
  or _83099_ (_33010_, _33009_, _09842_);
  or _83100_ (_33011_, _33010_, _33005_);
  and _83101_ (_33012_, _33011_, _32974_);
  or _83102_ (_33013_, _33012_, _06116_);
  and _83103_ (_33014_, _09160_, _07830_);
  or _83104_ (_33015_, _32968_, _06117_);
  or _83105_ (_33016_, _33015_, _33014_);
  and _83106_ (_33018_, _33016_, _06114_);
  and _83107_ (_33019_, _33018_, _33013_);
  and _83108_ (_33020_, _14260_, _07830_);
  or _83109_ (_33021_, _33020_, _32968_);
  and _83110_ (_33022_, _33021_, _05787_);
  or _83111_ (_33023_, _33022_, _33019_);
  or _83112_ (_33024_, _33023_, _11136_);
  and _83113_ (_33025_, _14275_, _07830_);
  or _83114_ (_33026_, _32968_, _07127_);
  or _83115_ (_33027_, _33026_, _33025_);
  and _83116_ (_33029_, _07830_, _08708_);
  or _83117_ (_33030_, _33029_, _32968_);
  or _83118_ (_33031_, _33030_, _06111_);
  and _83119_ (_33032_, _33031_, _07125_);
  and _83120_ (_33033_, _33032_, _33027_);
  and _83121_ (_33034_, _33033_, _33024_);
  nor _83122_ (_33035_, _12321_, _13300_);
  or _83123_ (_33036_, _33035_, _32968_);
  and _83124_ (_33037_, _32967_, _06402_);
  and _83125_ (_33038_, _33037_, _33036_);
  or _83126_ (_33040_, _33038_, _33034_);
  and _83127_ (_33041_, _33040_, _07132_);
  nand _83128_ (_33042_, _33030_, _06306_);
  nor _83129_ (_33043_, _33042_, _32975_);
  or _83130_ (_33044_, _33043_, _06411_);
  or _83131_ (_33045_, _33044_, _33041_);
  and _83132_ (_33046_, _33045_, _32970_);
  or _83133_ (_33047_, _33046_, _06303_);
  and _83134_ (_33048_, _14167_, _07830_);
  or _83135_ (_33049_, _32968_, _08819_);
  or _83136_ (_33051_, _33049_, _33048_);
  and _83137_ (_33052_, _33051_, _08824_);
  and _83138_ (_33053_, _33052_, _33047_);
  and _83139_ (_33054_, _33036_, _06396_);
  or _83140_ (_33055_, _33054_, _06433_);
  or _83141_ (_33056_, _33055_, _33053_);
  or _83142_ (_33057_, _32976_, _06829_);
  and _83143_ (_33058_, _33057_, _33056_);
  or _83144_ (_33059_, _33058_, _05748_);
  or _83145_ (_33060_, _32968_, _05749_);
  and _83146_ (_33062_, _33060_, _33059_);
  or _83147_ (_33063_, _33062_, _06440_);
  or _83148_ (_33064_, _32976_, _06444_);
  and _83149_ (_33065_, _33064_, _01317_);
  and _83150_ (_33066_, _33065_, _33063_);
  or _83151_ (_33067_, _33066_, _32966_);
  and _83152_ (_43738_, _33067_, _43100_);
  not _83153_ (_33068_, \oc8051_golden_model_1.IP [1]);
  nor _83154_ (_33069_, _01317_, _33068_);
  nor _83155_ (_33070_, _07830_, _33068_);
  nor _83156_ (_33072_, _10277_, _13300_);
  or _83157_ (_33073_, _33072_, _33070_);
  or _83158_ (_33074_, _33073_, _08824_);
  or _83159_ (_33075_, _14442_, _13300_);
  or _83160_ (_33076_, _07830_, \oc8051_golden_model_1.IP [1]);
  and _83161_ (_33077_, _33076_, _05787_);
  and _83162_ (_33078_, _33077_, _33075_);
  and _83163_ (_33079_, _07830_, _07306_);
  or _83164_ (_33080_, _33079_, _33070_);
  or _83165_ (_33081_, _33080_, _07075_);
  and _83166_ (_33083_, _14363_, _07830_);
  not _83167_ (_33084_, _33083_);
  and _83168_ (_33085_, _33084_, _33076_);
  or _83169_ (_33086_, _33085_, _06161_);
  and _83170_ (_33087_, _07830_, \oc8051_golden_model_1.ACC [1]);
  or _83171_ (_33088_, _33087_, _33070_);
  and _83172_ (_33089_, _33088_, _07056_);
  nor _83173_ (_33090_, _07056_, _33068_);
  or _83174_ (_33091_, _33090_, _06160_);
  or _83175_ (_33092_, _33091_, _33089_);
  and _83176_ (_33094_, _33092_, _06157_);
  and _83177_ (_33095_, _33094_, _33086_);
  nor _83178_ (_33096_, _08415_, _33068_);
  and _83179_ (_33097_, _14367_, _08415_);
  or _83180_ (_33098_, _33097_, _33096_);
  and _83181_ (_33099_, _33098_, _06156_);
  or _83182_ (_33100_, _33099_, _06217_);
  or _83183_ (_33101_, _33100_, _33095_);
  and _83184_ (_33102_, _33101_, _33081_);
  or _83185_ (_33103_, _33102_, _06220_);
  or _83186_ (_33105_, _33088_, _06229_);
  and _83187_ (_33106_, _33105_, _06153_);
  and _83188_ (_33107_, _33106_, _33103_);
  and _83189_ (_33108_, _14349_, _08415_);
  or _83190_ (_33109_, _33108_, _33096_);
  and _83191_ (_33110_, _33109_, _06152_);
  or _83192_ (_33111_, _33110_, _06145_);
  or _83193_ (_33112_, _33111_, _33107_);
  and _83194_ (_33113_, _33097_, _14382_);
  or _83195_ (_33114_, _33096_, _06146_);
  or _83196_ (_33116_, _33114_, _33113_);
  and _83197_ (_33117_, _33116_, _33112_);
  and _83198_ (_33118_, _33117_, _06140_);
  and _83199_ (_33119_, _14351_, _08415_);
  or _83200_ (_33120_, _33096_, _33119_);
  and _83201_ (_33121_, _33120_, _06139_);
  or _83202_ (_33122_, _33121_, _09842_);
  or _83203_ (_33123_, _33122_, _33118_);
  or _83204_ (_33124_, _33080_, _06132_);
  and _83205_ (_33125_, _33124_, _33123_);
  or _83206_ (_33127_, _33125_, _06116_);
  and _83207_ (_33128_, _09115_, _07830_);
  or _83208_ (_33129_, _33070_, _06117_);
  or _83209_ (_33130_, _33129_, _33128_);
  and _83210_ (_33131_, _33130_, _06114_);
  and _83211_ (_33132_, _33131_, _33127_);
  or _83212_ (_33133_, _33132_, _33078_);
  and _83213_ (_33134_, _33133_, _06298_);
  or _83214_ (_33135_, _14346_, _13300_);
  and _83215_ (_33136_, _33135_, _06297_);
  nand _83216_ (_33138_, _07830_, _06945_);
  and _83217_ (_33139_, _33138_, _06110_);
  or _83218_ (_33140_, _33139_, _33136_);
  and _83219_ (_33141_, _33140_, _33076_);
  or _83220_ (_33142_, _33141_, _06402_);
  or _83221_ (_33143_, _33142_, _33134_);
  nand _83222_ (_33144_, _10275_, _07830_);
  and _83223_ (_33145_, _33144_, _33073_);
  or _83224_ (_33146_, _33145_, _07125_);
  and _83225_ (_33147_, _33146_, _07132_);
  and _83226_ (_33149_, _33147_, _33143_);
  or _83227_ (_33150_, _14344_, _13300_);
  and _83228_ (_33151_, _33076_, _06306_);
  and _83229_ (_33152_, _33151_, _33150_);
  or _83230_ (_33153_, _33152_, _06411_);
  or _83231_ (_33154_, _33153_, _33149_);
  nor _83232_ (_33155_, _33070_, _07130_);
  nand _83233_ (_33156_, _33155_, _33144_);
  and _83234_ (_33157_, _33156_, _08819_);
  and _83235_ (_33158_, _33157_, _33154_);
  or _83236_ (_33160_, _33138_, _08176_);
  and _83237_ (_33161_, _33076_, _06303_);
  and _83238_ (_33162_, _33161_, _33160_);
  or _83239_ (_33163_, _33162_, _06396_);
  or _83240_ (_33164_, _33163_, _33158_);
  and _83241_ (_33165_, _33164_, _33074_);
  or _83242_ (_33166_, _33165_, _06433_);
  or _83243_ (_33167_, _33085_, _06829_);
  and _83244_ (_33168_, _33167_, _05749_);
  and _83245_ (_33169_, _33168_, _33166_);
  and _83246_ (_33171_, _33109_, _05748_);
  or _83247_ (_33172_, _33171_, _06440_);
  or _83248_ (_33173_, _33172_, _33169_);
  or _83249_ (_33174_, _33070_, _06444_);
  or _83250_ (_33175_, _33174_, _33083_);
  and _83251_ (_33176_, _33175_, _01317_);
  and _83252_ (_33177_, _33176_, _33173_);
  or _83253_ (_33178_, _33177_, _33069_);
  and _83254_ (_43739_, _33178_, _43100_);
  and _83255_ (_33179_, _01321_, \oc8051_golden_model_1.IP [2]);
  and _83256_ (_33181_, _13300_, \oc8051_golden_model_1.IP [2]);
  and _83257_ (_33182_, _07830_, _07708_);
  or _83258_ (_33183_, _33182_, _33181_);
  or _83259_ (_33184_, _33183_, _06132_);
  or _83260_ (_33185_, _33183_, _07075_);
  and _83261_ (_33186_, _14542_, _07830_);
  or _83262_ (_33187_, _33186_, _33181_);
  or _83263_ (_33188_, _33187_, _06161_);
  and _83264_ (_33189_, _07830_, \oc8051_golden_model_1.ACC [2]);
  or _83265_ (_33190_, _33189_, _33181_);
  and _83266_ (_33192_, _33190_, _07056_);
  and _83267_ (_33193_, _07057_, \oc8051_golden_model_1.IP [2]);
  or _83268_ (_33194_, _33193_, _06160_);
  or _83269_ (_33195_, _33194_, _33192_);
  and _83270_ (_33196_, _33195_, _06157_);
  and _83271_ (_33197_, _33196_, _33188_);
  and _83272_ (_33198_, _13305_, \oc8051_golden_model_1.IP [2]);
  and _83273_ (_33199_, _14538_, _08415_);
  or _83274_ (_33200_, _33199_, _33198_);
  and _83275_ (_33201_, _33200_, _06156_);
  or _83276_ (_33203_, _33201_, _06217_);
  or _83277_ (_33204_, _33203_, _33197_);
  and _83278_ (_33205_, _33204_, _33185_);
  or _83279_ (_33206_, _33205_, _06220_);
  or _83280_ (_33207_, _33190_, _06229_);
  and _83281_ (_33208_, _33207_, _06153_);
  and _83282_ (_33209_, _33208_, _33206_);
  and _83283_ (_33210_, _14536_, _08415_);
  or _83284_ (_33211_, _33210_, _33198_);
  and _83285_ (_33212_, _33211_, _06152_);
  or _83286_ (_33214_, _33212_, _06145_);
  or _83287_ (_33215_, _33214_, _33209_);
  and _83288_ (_33216_, _33199_, _14569_);
  or _83289_ (_33217_, _33198_, _06146_);
  or _83290_ (_33218_, _33217_, _33216_);
  and _83291_ (_33219_, _33218_, _06140_);
  and _83292_ (_33220_, _33219_, _33215_);
  and _83293_ (_33221_, _14583_, _08415_);
  or _83294_ (_33222_, _33221_, _33198_);
  and _83295_ (_33223_, _33222_, _06139_);
  or _83296_ (_33225_, _33223_, _09842_);
  or _83297_ (_33226_, _33225_, _33220_);
  and _83298_ (_33227_, _33226_, _33184_);
  or _83299_ (_33228_, _33227_, _06116_);
  and _83300_ (_33229_, _09211_, _07830_);
  or _83301_ (_33230_, _33181_, _06117_);
  or _83302_ (_33231_, _33230_, _33229_);
  and _83303_ (_33232_, _33231_, _06114_);
  and _83304_ (_33233_, _33232_, _33228_);
  and _83305_ (_33234_, _14630_, _07830_);
  or _83306_ (_33236_, _33181_, _33234_);
  and _83307_ (_33237_, _33236_, _05787_);
  or _83308_ (_33238_, _33237_, _33233_);
  or _83309_ (_33239_, _33238_, _11136_);
  and _83310_ (_33240_, _14646_, _07830_);
  or _83311_ (_33241_, _33181_, _07127_);
  or _83312_ (_33242_, _33241_, _33240_);
  and _83313_ (_33243_, _07830_, _08768_);
  or _83314_ (_33244_, _33243_, _33181_);
  or _83315_ (_33245_, _33244_, _06111_);
  and _83316_ (_33247_, _33245_, _07125_);
  and _83317_ (_33248_, _33247_, _33242_);
  and _83318_ (_33249_, _33248_, _33239_);
  and _83319_ (_33250_, _10282_, _07830_);
  or _83320_ (_33251_, _33250_, _33181_);
  and _83321_ (_33252_, _33251_, _06402_);
  or _83322_ (_33253_, _33252_, _33249_);
  and _83323_ (_33254_, _33253_, _07132_);
  or _83324_ (_33255_, _33181_, _08248_);
  and _83325_ (_33256_, _33244_, _06306_);
  and _83326_ (_33258_, _33256_, _33255_);
  or _83327_ (_33259_, _33258_, _33254_);
  and _83328_ (_33260_, _33259_, _07130_);
  and _83329_ (_33261_, _33190_, _06411_);
  and _83330_ (_33262_, _33261_, _33255_);
  or _83331_ (_33263_, _33262_, _06303_);
  or _83332_ (_33264_, _33263_, _33260_);
  and _83333_ (_33265_, _14643_, _07830_);
  or _83334_ (_33266_, _33181_, _08819_);
  or _83335_ (_33267_, _33266_, _33265_);
  and _83336_ (_33269_, _33267_, _08824_);
  and _83337_ (_33270_, _33269_, _33264_);
  nor _83338_ (_33271_, _10281_, _13300_);
  or _83339_ (_33272_, _33271_, _33181_);
  and _83340_ (_33273_, _33272_, _06396_);
  or _83341_ (_33274_, _33273_, _06433_);
  or _83342_ (_33275_, _33274_, _33270_);
  or _83343_ (_33276_, _33187_, _06829_);
  and _83344_ (_33277_, _33276_, _05749_);
  and _83345_ (_33278_, _33277_, _33275_);
  and _83346_ (_33280_, _33211_, _05748_);
  or _83347_ (_33281_, _33280_, _06440_);
  or _83348_ (_33282_, _33281_, _33278_);
  and _83349_ (_33283_, _14710_, _07830_);
  or _83350_ (_33284_, _33181_, _06444_);
  or _83351_ (_33285_, _33284_, _33283_);
  and _83352_ (_33286_, _33285_, _01317_);
  and _83353_ (_33287_, _33286_, _33282_);
  or _83354_ (_33288_, _33287_, _33179_);
  and _83355_ (_43740_, _33288_, _43100_);
  and _83356_ (_33290_, _01321_, \oc8051_golden_model_1.IP [3]);
  and _83357_ (_33291_, _13300_, \oc8051_golden_model_1.IP [3]);
  and _83358_ (_33292_, _07830_, _07544_);
  or _83359_ (_33293_, _33292_, _33291_);
  or _83360_ (_33294_, _33293_, _06132_);
  and _83361_ (_33295_, _14738_, _07830_);
  or _83362_ (_33296_, _33295_, _33291_);
  or _83363_ (_33297_, _33296_, _06161_);
  and _83364_ (_33298_, _07830_, \oc8051_golden_model_1.ACC [3]);
  or _83365_ (_33299_, _33298_, _33291_);
  and _83366_ (_33301_, _33299_, _07056_);
  and _83367_ (_33302_, _07057_, \oc8051_golden_model_1.IP [3]);
  or _83368_ (_33303_, _33302_, _06160_);
  or _83369_ (_33304_, _33303_, _33301_);
  and _83370_ (_33305_, _33304_, _06157_);
  and _83371_ (_33306_, _33305_, _33297_);
  and _83372_ (_33307_, _13305_, \oc8051_golden_model_1.IP [3]);
  and _83373_ (_33308_, _14735_, _08415_);
  or _83374_ (_33309_, _33308_, _33307_);
  and _83375_ (_33310_, _33309_, _06156_);
  or _83376_ (_33312_, _33310_, _06217_);
  or _83377_ (_33313_, _33312_, _33306_);
  or _83378_ (_33314_, _33293_, _07075_);
  and _83379_ (_33315_, _33314_, _33313_);
  or _83380_ (_33316_, _33315_, _06220_);
  or _83381_ (_33317_, _33299_, _06229_);
  and _83382_ (_33318_, _33317_, _06153_);
  and _83383_ (_33319_, _33318_, _33316_);
  and _83384_ (_33320_, _14731_, _08415_);
  or _83385_ (_33321_, _33320_, _33307_);
  and _83386_ (_33323_, _33321_, _06152_);
  or _83387_ (_33324_, _33323_, _06145_);
  or _83388_ (_33325_, _33324_, _33319_);
  or _83389_ (_33326_, _33307_, _14764_);
  and _83390_ (_33327_, _33326_, _33309_);
  or _83391_ (_33328_, _33327_, _06146_);
  and _83392_ (_33329_, _33328_, _06140_);
  and _83393_ (_33330_, _33329_, _33325_);
  and _83394_ (_33331_, _14732_, _08415_);
  or _83395_ (_33332_, _33331_, _33307_);
  and _83396_ (_33334_, _33332_, _06139_);
  or _83397_ (_33335_, _33334_, _09842_);
  or _83398_ (_33336_, _33335_, _33330_);
  and _83399_ (_33337_, _33336_, _33294_);
  or _83400_ (_33338_, _33337_, _06116_);
  and _83401_ (_33339_, _09210_, _07830_);
  or _83402_ (_33340_, _33291_, _06117_);
  or _83403_ (_33341_, _33340_, _33339_);
  and _83404_ (_33342_, _33341_, _06114_);
  and _83405_ (_33343_, _33342_, _33338_);
  and _83406_ (_33345_, _14825_, _07830_);
  or _83407_ (_33346_, _33291_, _33345_);
  and _83408_ (_33347_, _33346_, _05787_);
  or _83409_ (_33348_, _33347_, _33343_);
  or _83410_ (_33349_, _33348_, _11136_);
  and _83411_ (_33350_, _14727_, _07830_);
  or _83412_ (_33351_, _33291_, _07127_);
  or _83413_ (_33352_, _33351_, _33350_);
  and _83414_ (_33353_, _07830_, _08712_);
  or _83415_ (_33354_, _33353_, _33291_);
  or _83416_ (_33356_, _33354_, _06111_);
  and _83417_ (_33357_, _33356_, _07125_);
  and _83418_ (_33358_, _33357_, _33352_);
  and _83419_ (_33359_, _33358_, _33349_);
  and _83420_ (_33360_, _12318_, _07830_);
  or _83421_ (_33361_, _33360_, _33291_);
  and _83422_ (_33362_, _33361_, _06402_);
  or _83423_ (_33363_, _33362_, _33359_);
  and _83424_ (_33364_, _33363_, _07132_);
  or _83425_ (_33365_, _33291_, _08140_);
  and _83426_ (_33367_, _33354_, _06306_);
  and _83427_ (_33368_, _33367_, _33365_);
  or _83428_ (_33369_, _33368_, _33364_);
  and _83429_ (_33370_, _33369_, _07130_);
  and _83430_ (_33371_, _33299_, _06411_);
  and _83431_ (_33372_, _33371_, _33365_);
  or _83432_ (_33373_, _33372_, _06303_);
  or _83433_ (_33374_, _33373_, _33370_);
  and _83434_ (_33375_, _14724_, _07830_);
  or _83435_ (_33376_, _33291_, _08819_);
  or _83436_ (_33378_, _33376_, _33375_);
  and _83437_ (_33379_, _33378_, _08824_);
  and _83438_ (_33380_, _33379_, _33374_);
  nor _83439_ (_33381_, _10273_, _13300_);
  or _83440_ (_33382_, _33381_, _33291_);
  and _83441_ (_33383_, _33382_, _06396_);
  or _83442_ (_33384_, _33383_, _06433_);
  or _83443_ (_33385_, _33384_, _33380_);
  or _83444_ (_33386_, _33296_, _06829_);
  and _83445_ (_33387_, _33386_, _05749_);
  and _83446_ (_33389_, _33387_, _33385_);
  and _83447_ (_33390_, _33321_, _05748_);
  or _83448_ (_33391_, _33390_, _06440_);
  or _83449_ (_33392_, _33391_, _33389_);
  and _83450_ (_33393_, _14897_, _07830_);
  or _83451_ (_33394_, _33291_, _06444_);
  or _83452_ (_33395_, _33394_, _33393_);
  and _83453_ (_33396_, _33395_, _01317_);
  and _83454_ (_33397_, _33396_, _33392_);
  or _83455_ (_33398_, _33397_, _33290_);
  and _83456_ (_43742_, _33398_, _43100_);
  and _83457_ (_33400_, _01321_, \oc8051_golden_model_1.IP [4]);
  and _83458_ (_33401_, _13300_, \oc8051_golden_model_1.IP [4]);
  and _83459_ (_33402_, _08336_, _07830_);
  or _83460_ (_33403_, _33402_, _33401_);
  or _83461_ (_33404_, _33403_, _06132_);
  and _83462_ (_33405_, _13305_, \oc8051_golden_model_1.IP [4]);
  and _83463_ (_33406_, _14942_, _08415_);
  or _83464_ (_33407_, _33406_, _33405_);
  and _83465_ (_33408_, _33407_, _06152_);
  and _83466_ (_33410_, _14928_, _07830_);
  or _83467_ (_33411_, _33410_, _33401_);
  or _83468_ (_33412_, _33411_, _06161_);
  and _83469_ (_33413_, _07830_, \oc8051_golden_model_1.ACC [4]);
  or _83470_ (_33414_, _33413_, _33401_);
  and _83471_ (_33415_, _33414_, _07056_);
  and _83472_ (_33416_, _07057_, \oc8051_golden_model_1.IP [4]);
  or _83473_ (_33417_, _33416_, _06160_);
  or _83474_ (_33418_, _33417_, _33415_);
  and _83475_ (_33419_, _33418_, _06157_);
  and _83476_ (_33421_, _33419_, _33412_);
  and _83477_ (_33422_, _14932_, _08415_);
  or _83478_ (_33423_, _33422_, _33405_);
  and _83479_ (_33424_, _33423_, _06156_);
  or _83480_ (_33425_, _33424_, _06217_);
  or _83481_ (_33426_, _33425_, _33421_);
  or _83482_ (_33427_, _33403_, _07075_);
  and _83483_ (_33428_, _33427_, _33426_);
  or _83484_ (_33429_, _33428_, _06220_);
  or _83485_ (_33430_, _33414_, _06229_);
  and _83486_ (_33432_, _33430_, _06153_);
  and _83487_ (_33433_, _33432_, _33429_);
  or _83488_ (_33434_, _33433_, _33408_);
  and _83489_ (_33435_, _33434_, _06146_);
  and _83490_ (_33436_, _14950_, _08415_);
  or _83491_ (_33437_, _33436_, _33405_);
  and _83492_ (_33438_, _33437_, _06145_);
  or _83493_ (_33439_, _33438_, _33435_);
  and _83494_ (_33440_, _33439_, _06140_);
  and _83495_ (_33441_, _14966_, _08415_);
  or _83496_ (_33443_, _33441_, _33405_);
  and _83497_ (_33444_, _33443_, _06139_);
  or _83498_ (_33445_, _33444_, _09842_);
  or _83499_ (_33446_, _33445_, _33440_);
  and _83500_ (_33447_, _33446_, _33404_);
  or _83501_ (_33448_, _33447_, _06116_);
  and _83502_ (_33449_, _09209_, _07830_);
  or _83503_ (_33450_, _33401_, _06117_);
  or _83504_ (_33451_, _33450_, _33449_);
  and _83505_ (_33452_, _33451_, _06114_);
  and _83506_ (_33454_, _33452_, _33448_);
  and _83507_ (_33455_, _15013_, _07830_);
  or _83508_ (_33456_, _33455_, _33401_);
  and _83509_ (_33457_, _33456_, _05787_);
  or _83510_ (_33458_, _33457_, _11136_);
  or _83511_ (_33459_, _33458_, _33454_);
  and _83512_ (_33460_, _15029_, _07830_);
  or _83513_ (_33461_, _33401_, _07127_);
  or _83514_ (_33462_, _33461_, _33460_);
  and _83515_ (_33463_, _08715_, _07830_);
  or _83516_ (_33464_, _33463_, _33401_);
  or _83517_ (_33465_, _33464_, _06111_);
  and _83518_ (_33466_, _33465_, _07125_);
  and _83519_ (_33467_, _33466_, _33462_);
  and _83520_ (_33468_, _33467_, _33459_);
  and _83521_ (_33469_, _10289_, _07830_);
  or _83522_ (_33470_, _33469_, _33401_);
  and _83523_ (_33471_, _33470_, _06402_);
  or _83524_ (_33472_, _33471_, _33468_);
  and _83525_ (_33473_, _33472_, _07132_);
  or _83526_ (_33475_, _33401_, _08339_);
  and _83527_ (_33476_, _33464_, _06306_);
  and _83528_ (_33477_, _33476_, _33475_);
  or _83529_ (_33478_, _33477_, _33473_);
  and _83530_ (_33479_, _33478_, _07130_);
  and _83531_ (_33480_, _33414_, _06411_);
  and _83532_ (_33481_, _33480_, _33475_);
  or _83533_ (_33482_, _33481_, _06303_);
  or _83534_ (_33483_, _33482_, _33479_);
  and _83535_ (_33484_, _15026_, _07830_);
  or _83536_ (_33486_, _33401_, _08819_);
  or _83537_ (_33487_, _33486_, _33484_);
  and _83538_ (_33488_, _33487_, _08824_);
  and _83539_ (_33489_, _33488_, _33483_);
  nor _83540_ (_33490_, _10288_, _13300_);
  or _83541_ (_33491_, _33490_, _33401_);
  and _83542_ (_33492_, _33491_, _06396_);
  or _83543_ (_33493_, _33492_, _06433_);
  or _83544_ (_33494_, _33493_, _33489_);
  or _83545_ (_33495_, _33411_, _06829_);
  and _83546_ (_33497_, _33495_, _05749_);
  and _83547_ (_33498_, _33497_, _33494_);
  and _83548_ (_33499_, _33407_, _05748_);
  or _83549_ (_33500_, _33499_, _06440_);
  or _83550_ (_33501_, _33500_, _33498_);
  and _83551_ (_33502_, _15087_, _07830_);
  or _83552_ (_33503_, _33401_, _06444_);
  or _83553_ (_33504_, _33503_, _33502_);
  and _83554_ (_33505_, _33504_, _01317_);
  and _83555_ (_33506_, _33505_, _33501_);
  or _83556_ (_33508_, _33506_, _33400_);
  and _83557_ (_43743_, _33508_, _43100_);
  and _83558_ (_33509_, _01321_, \oc8051_golden_model_1.IP [5]);
  and _83559_ (_33510_, _13300_, \oc8051_golden_model_1.IP [5]);
  and _83560_ (_33511_, _15119_, _07830_);
  or _83561_ (_33512_, _33511_, _33510_);
  or _83562_ (_33513_, _33512_, _06161_);
  and _83563_ (_33514_, _07830_, \oc8051_golden_model_1.ACC [5]);
  or _83564_ (_33515_, _33514_, _33510_);
  and _83565_ (_33516_, _33515_, _07056_);
  and _83566_ (_33518_, _07057_, \oc8051_golden_model_1.IP [5]);
  or _83567_ (_33519_, _33518_, _06160_);
  or _83568_ (_33520_, _33519_, _33516_);
  and _83569_ (_33521_, _33520_, _06157_);
  and _83570_ (_33522_, _33521_, _33513_);
  and _83571_ (_33523_, _13305_, \oc8051_golden_model_1.IP [5]);
  and _83572_ (_33524_, _15123_, _08415_);
  or _83573_ (_33525_, _33524_, _33523_);
  and _83574_ (_33526_, _33525_, _06156_);
  or _83575_ (_33527_, _33526_, _06217_);
  or _83576_ (_33529_, _33527_, _33522_);
  and _83577_ (_33530_, _08101_, _07830_);
  or _83578_ (_33531_, _33530_, _33510_);
  or _83579_ (_33532_, _33531_, _07075_);
  and _83580_ (_33533_, _33532_, _33529_);
  or _83581_ (_33534_, _33533_, _06220_);
  or _83582_ (_33535_, _33515_, _06229_);
  and _83583_ (_33536_, _33535_, _06153_);
  and _83584_ (_33537_, _33536_, _33534_);
  and _83585_ (_33538_, _15104_, _08415_);
  or _83586_ (_33540_, _33538_, _33523_);
  and _83587_ (_33541_, _33540_, _06152_);
  or _83588_ (_33542_, _33541_, _06145_);
  or _83589_ (_33543_, _33542_, _33537_);
  or _83590_ (_33544_, _33523_, _15138_);
  and _83591_ (_33545_, _33544_, _33525_);
  or _83592_ (_33546_, _33545_, _06146_);
  and _83593_ (_33547_, _33546_, _06140_);
  and _83594_ (_33548_, _33547_, _33543_);
  and _83595_ (_33549_, _15155_, _08415_);
  or _83596_ (_33551_, _33549_, _33523_);
  and _83597_ (_33552_, _33551_, _06139_);
  or _83598_ (_33553_, _33552_, _09842_);
  or _83599_ (_33554_, _33553_, _33548_);
  or _83600_ (_33555_, _33531_, _06132_);
  and _83601_ (_33556_, _33555_, _33554_);
  or _83602_ (_33557_, _33556_, _06116_);
  and _83603_ (_33558_, _09208_, _07830_);
  or _83604_ (_33559_, _33510_, _06117_);
  or _83605_ (_33560_, _33559_, _33558_);
  and _83606_ (_33562_, _33560_, _06114_);
  and _83607_ (_33563_, _33562_, _33557_);
  and _83608_ (_33564_, _15203_, _07830_);
  or _83609_ (_33565_, _33564_, _33510_);
  and _83610_ (_33566_, _33565_, _05787_);
  or _83611_ (_33567_, _33566_, _11136_);
  or _83612_ (_33568_, _33567_, _33563_);
  and _83613_ (_33569_, _15219_, _07830_);
  or _83614_ (_33570_, _33510_, _07127_);
  or _83615_ (_33571_, _33570_, _33569_);
  and _83616_ (_33573_, _08736_, _07830_);
  or _83617_ (_33574_, _33573_, _33510_);
  or _83618_ (_33575_, _33574_, _06111_);
  and _83619_ (_33576_, _33575_, _07125_);
  and _83620_ (_33577_, _33576_, _33571_);
  and _83621_ (_33578_, _33577_, _33568_);
  and _83622_ (_33579_, _12325_, _07830_);
  or _83623_ (_33580_, _33579_, _33510_);
  and _83624_ (_33581_, _33580_, _06402_);
  or _83625_ (_33582_, _33581_, _33578_);
  and _83626_ (_33584_, _33582_, _07132_);
  or _83627_ (_33585_, _33510_, _08104_);
  and _83628_ (_33586_, _33574_, _06306_);
  and _83629_ (_33587_, _33586_, _33585_);
  or _83630_ (_33588_, _33587_, _33584_);
  and _83631_ (_33589_, _33588_, _07130_);
  and _83632_ (_33590_, _33515_, _06411_);
  and _83633_ (_33591_, _33590_, _33585_);
  or _83634_ (_33592_, _33591_, _06303_);
  or _83635_ (_33593_, _33592_, _33589_);
  and _83636_ (_33595_, _15216_, _07830_);
  or _83637_ (_33596_, _33510_, _08819_);
  or _83638_ (_33597_, _33596_, _33595_);
  and _83639_ (_33598_, _33597_, _08824_);
  and _83640_ (_33599_, _33598_, _33593_);
  nor _83641_ (_33600_, _10269_, _13300_);
  or _83642_ (_33601_, _33600_, _33510_);
  and _83643_ (_33602_, _33601_, _06396_);
  or _83644_ (_33603_, _33602_, _06433_);
  or _83645_ (_33604_, _33603_, _33599_);
  or _83646_ (_33606_, _33512_, _06829_);
  and _83647_ (_33607_, _33606_, _05749_);
  and _83648_ (_33608_, _33607_, _33604_);
  and _83649_ (_33609_, _33540_, _05748_);
  or _83650_ (_33610_, _33609_, _06440_);
  or _83651_ (_33611_, _33610_, _33608_);
  and _83652_ (_33612_, _15275_, _07830_);
  or _83653_ (_33613_, _33510_, _06444_);
  or _83654_ (_33614_, _33613_, _33612_);
  and _83655_ (_33615_, _33614_, _01317_);
  and _83656_ (_33617_, _33615_, _33611_);
  or _83657_ (_33618_, _33617_, _33509_);
  and _83658_ (_43744_, _33618_, _43100_);
  and _83659_ (_33619_, _01321_, \oc8051_golden_model_1.IP [6]);
  and _83660_ (_33620_, _13300_, \oc8051_golden_model_1.IP [6]);
  and _83661_ (_33621_, _15300_, _07830_);
  or _83662_ (_33622_, _33621_, _33620_);
  or _83663_ (_33623_, _33622_, _06161_);
  and _83664_ (_33624_, _07830_, \oc8051_golden_model_1.ACC [6]);
  or _83665_ (_33625_, _33624_, _33620_);
  and _83666_ (_33627_, _33625_, _07056_);
  and _83667_ (_33628_, _07057_, \oc8051_golden_model_1.IP [6]);
  or _83668_ (_33629_, _33628_, _06160_);
  or _83669_ (_33630_, _33629_, _33627_);
  and _83670_ (_33631_, _33630_, _06157_);
  and _83671_ (_33632_, _33631_, _33623_);
  and _83672_ (_33633_, _13305_, \oc8051_golden_model_1.IP [6]);
  and _83673_ (_33634_, _15316_, _08415_);
  or _83674_ (_33635_, _33634_, _33633_);
  and _83675_ (_33636_, _33635_, _06156_);
  or _83676_ (_33638_, _33636_, _06217_);
  or _83677_ (_33639_, _33638_, _33632_);
  and _83678_ (_33640_, _08012_, _07830_);
  or _83679_ (_33641_, _33640_, _33620_);
  or _83680_ (_33642_, _33641_, _07075_);
  and _83681_ (_33643_, _33642_, _33639_);
  or _83682_ (_33644_, _33643_, _06220_);
  or _83683_ (_33645_, _33625_, _06229_);
  and _83684_ (_33646_, _33645_, _06153_);
  and _83685_ (_33647_, _33646_, _33644_);
  and _83686_ (_33649_, _15297_, _08415_);
  or _83687_ (_33650_, _33649_, _33633_);
  and _83688_ (_33651_, _33650_, _06152_);
  or _83689_ (_33652_, _33651_, _06145_);
  or _83690_ (_33653_, _33652_, _33647_);
  or _83691_ (_33654_, _33633_, _15331_);
  and _83692_ (_33655_, _33654_, _33635_);
  or _83693_ (_33656_, _33655_, _06146_);
  and _83694_ (_33657_, _33656_, _06140_);
  and _83695_ (_33658_, _33657_, _33653_);
  and _83696_ (_33660_, _15348_, _08415_);
  or _83697_ (_33661_, _33660_, _33633_);
  and _83698_ (_33662_, _33661_, _06139_);
  or _83699_ (_33663_, _33662_, _09842_);
  or _83700_ (_33664_, _33663_, _33658_);
  or _83701_ (_33665_, _33641_, _06132_);
  and _83702_ (_33666_, _33665_, _33664_);
  or _83703_ (_33667_, _33666_, _06116_);
  and _83704_ (_33668_, _09207_, _07830_);
  or _83705_ (_33669_, _33620_, _06117_);
  or _83706_ (_33671_, _33669_, _33668_);
  and _83707_ (_33672_, _33671_, _06114_);
  and _83708_ (_33673_, _33672_, _33667_);
  and _83709_ (_33674_, _15395_, _07830_);
  or _83710_ (_33675_, _33674_, _33620_);
  and _83711_ (_33676_, _33675_, _05787_);
  or _83712_ (_33677_, _33676_, _11136_);
  or _83713_ (_33678_, _33677_, _33673_);
  and _83714_ (_33679_, _15413_, _07830_);
  or _83715_ (_33680_, _33620_, _07127_);
  or _83716_ (_33682_, _33680_, _33679_);
  and _83717_ (_33683_, _15402_, _07830_);
  or _83718_ (_33684_, _33683_, _33620_);
  or _83719_ (_33685_, _33684_, _06111_);
  and _83720_ (_33686_, _33685_, _07125_);
  and _83721_ (_33687_, _33686_, _33682_);
  and _83722_ (_33688_, _33687_, _33678_);
  and _83723_ (_33689_, _10295_, _07830_);
  or _83724_ (_33690_, _33689_, _33620_);
  and _83725_ (_33691_, _33690_, _06402_);
  or _83726_ (_33693_, _33691_, _33688_);
  and _83727_ (_33694_, _33693_, _07132_);
  or _83728_ (_33695_, _33620_, _08015_);
  and _83729_ (_33696_, _33684_, _06306_);
  and _83730_ (_33697_, _33696_, _33695_);
  or _83731_ (_33698_, _33697_, _33694_);
  and _83732_ (_33699_, _33698_, _07130_);
  and _83733_ (_33700_, _33625_, _06411_);
  and _83734_ (_33701_, _33700_, _33695_);
  or _83735_ (_33702_, _33701_, _06303_);
  or _83736_ (_33704_, _33702_, _33699_);
  and _83737_ (_33705_, _15410_, _07830_);
  or _83738_ (_33706_, _33620_, _08819_);
  or _83739_ (_33707_, _33706_, _33705_);
  and _83740_ (_33708_, _33707_, _08824_);
  and _83741_ (_33709_, _33708_, _33704_);
  nor _83742_ (_33710_, _10294_, _13300_);
  or _83743_ (_33711_, _33710_, _33620_);
  and _83744_ (_33712_, _33711_, _06396_);
  or _83745_ (_33713_, _33712_, _06433_);
  or _83746_ (_33715_, _33713_, _33709_);
  or _83747_ (_33716_, _33622_, _06829_);
  and _83748_ (_33717_, _33716_, _05749_);
  and _83749_ (_33718_, _33717_, _33715_);
  and _83750_ (_33719_, _33650_, _05748_);
  or _83751_ (_33720_, _33719_, _06440_);
  or _83752_ (_33721_, _33720_, _33718_);
  and _83753_ (_33722_, _15478_, _07830_);
  or _83754_ (_33723_, _33620_, _06444_);
  or _83755_ (_33724_, _33723_, _33722_);
  and _83756_ (_33726_, _33724_, _01317_);
  and _83757_ (_33727_, _33726_, _33721_);
  or _83758_ (_33728_, _33727_, _33619_);
  and _83759_ (_43745_, _33728_, _43100_);
  not _83760_ (_33729_, \oc8051_golden_model_1.IE [0]);
  nor _83761_ (_33730_, _01317_, _33729_);
  nand _83762_ (_33731_, _10276_, _07826_);
  nor _83763_ (_33732_, _07826_, _33729_);
  nor _83764_ (_33733_, _33732_, _07130_);
  nand _83765_ (_33734_, _33733_, _33731_);
  and _83766_ (_33736_, _07826_, _07049_);
  or _83767_ (_33737_, _33736_, _33732_);
  or _83768_ (_33738_, _33737_, _06132_);
  nor _83769_ (_33739_, _08211_, _13402_);
  or _83770_ (_33740_, _33739_, _33732_);
  or _83771_ (_33741_, _33740_, _06161_);
  and _83772_ (_33742_, _07826_, \oc8051_golden_model_1.ACC [0]);
  or _83773_ (_33743_, _33742_, _33732_);
  and _83774_ (_33744_, _33743_, _07056_);
  nor _83775_ (_33745_, _07056_, _33729_);
  or _83776_ (_33747_, _33745_, _06160_);
  or _83777_ (_33748_, _33747_, _33744_);
  and _83778_ (_33749_, _33748_, _06157_);
  and _83779_ (_33750_, _33749_, _33741_);
  nor _83780_ (_33751_, _08418_, _33729_);
  and _83781_ (_33752_, _14169_, _08418_);
  or _83782_ (_33753_, _33752_, _33751_);
  and _83783_ (_33754_, _33753_, _06156_);
  or _83784_ (_33755_, _33754_, _33750_);
  and _83785_ (_33756_, _33755_, _07075_);
  and _83786_ (_33758_, _33737_, _06217_);
  or _83787_ (_33759_, _33758_, _06220_);
  or _83788_ (_33760_, _33759_, _33756_);
  or _83789_ (_33761_, _33743_, _06229_);
  and _83790_ (_33762_, _33761_, _06153_);
  and _83791_ (_33763_, _33762_, _33760_);
  and _83792_ (_33764_, _33732_, _06152_);
  or _83793_ (_33765_, _33764_, _06145_);
  or _83794_ (_33766_, _33765_, _33763_);
  or _83795_ (_33767_, _33740_, _06146_);
  and _83796_ (_33769_, _33767_, _06140_);
  and _83797_ (_33770_, _33769_, _33766_);
  or _83798_ (_33771_, _33751_, _14170_);
  and _83799_ (_33772_, _33771_, _06139_);
  and _83800_ (_33773_, _33772_, _33753_);
  or _83801_ (_33774_, _33773_, _09842_);
  or _83802_ (_33775_, _33774_, _33770_);
  and _83803_ (_33776_, _33775_, _33738_);
  or _83804_ (_33777_, _33776_, _06116_);
  and _83805_ (_33778_, _09160_, _07826_);
  or _83806_ (_33780_, _33732_, _06117_);
  or _83807_ (_33781_, _33780_, _33778_);
  and _83808_ (_33782_, _33781_, _06114_);
  and _83809_ (_33783_, _33782_, _33777_);
  and _83810_ (_33784_, _14260_, _07826_);
  or _83811_ (_33785_, _33784_, _33732_);
  and _83812_ (_33786_, _33785_, _05787_);
  or _83813_ (_33787_, _33786_, _33783_);
  or _83814_ (_33788_, _33787_, _11136_);
  and _83815_ (_33789_, _14275_, _07826_);
  or _83816_ (_33791_, _33732_, _07127_);
  or _83817_ (_33792_, _33791_, _33789_);
  and _83818_ (_33793_, _07826_, _08708_);
  or _83819_ (_33794_, _33793_, _33732_);
  or _83820_ (_33795_, _33794_, _06111_);
  and _83821_ (_33796_, _33795_, _07125_);
  and _83822_ (_33797_, _33796_, _33792_);
  and _83823_ (_33798_, _33797_, _33788_);
  nor _83824_ (_33799_, _12321_, _13402_);
  or _83825_ (_33800_, _33799_, _33732_);
  and _83826_ (_33802_, _33731_, _06402_);
  and _83827_ (_33803_, _33802_, _33800_);
  or _83828_ (_33804_, _33803_, _33798_);
  and _83829_ (_33805_, _33804_, _07132_);
  nand _83830_ (_33806_, _33794_, _06306_);
  nor _83831_ (_33807_, _33806_, _33739_);
  or _83832_ (_33808_, _33807_, _06411_);
  or _83833_ (_33809_, _33808_, _33805_);
  and _83834_ (_33810_, _33809_, _33734_);
  or _83835_ (_33811_, _33810_, _06303_);
  and _83836_ (_33813_, _14167_, _07826_);
  or _83837_ (_33814_, _33732_, _08819_);
  or _83838_ (_33815_, _33814_, _33813_);
  and _83839_ (_33816_, _33815_, _08824_);
  and _83840_ (_33817_, _33816_, _33811_);
  and _83841_ (_33818_, _33800_, _06396_);
  or _83842_ (_33819_, _33818_, _06433_);
  or _83843_ (_33820_, _33819_, _33817_);
  or _83844_ (_33821_, _33740_, _06829_);
  and _83845_ (_33822_, _33821_, _33820_);
  or _83846_ (_33824_, _33822_, _05748_);
  or _83847_ (_33825_, _33732_, _05749_);
  and _83848_ (_33826_, _33825_, _33824_);
  or _83849_ (_33827_, _33826_, _06440_);
  or _83850_ (_33828_, _33740_, _06444_);
  and _83851_ (_33829_, _33828_, _01317_);
  and _83852_ (_33830_, _33829_, _33827_);
  or _83853_ (_33831_, _33830_, _33730_);
  and _83854_ (_43747_, _33831_, _43100_);
  not _83855_ (_33832_, \oc8051_golden_model_1.IE [1]);
  nor _83856_ (_33834_, _01317_, _33832_);
  nor _83857_ (_33835_, _07826_, _33832_);
  nor _83858_ (_33836_, _10277_, _13402_);
  or _83859_ (_33837_, _33836_, _33835_);
  or _83860_ (_33838_, _33837_, _08824_);
  and _83861_ (_33839_, _07826_, _07306_);
  or _83862_ (_33840_, _33839_, _33835_);
  or _83863_ (_33841_, _33840_, _07075_);
  or _83864_ (_33842_, _07826_, \oc8051_golden_model_1.IE [1]);
  and _83865_ (_33843_, _14363_, _07826_);
  not _83866_ (_33845_, _33843_);
  and _83867_ (_33846_, _33845_, _33842_);
  or _83868_ (_33847_, _33846_, _06161_);
  and _83869_ (_33848_, _07826_, \oc8051_golden_model_1.ACC [1]);
  or _83870_ (_33849_, _33848_, _33835_);
  and _83871_ (_33850_, _33849_, _07056_);
  nor _83872_ (_33851_, _07056_, _33832_);
  or _83873_ (_33852_, _33851_, _06160_);
  or _83874_ (_33853_, _33852_, _33850_);
  and _83875_ (_33854_, _33853_, _06157_);
  and _83876_ (_33856_, _33854_, _33847_);
  nor _83877_ (_33857_, _08418_, _33832_);
  and _83878_ (_33858_, _14367_, _08418_);
  or _83879_ (_33859_, _33858_, _33857_);
  and _83880_ (_33860_, _33859_, _06156_);
  or _83881_ (_33861_, _33860_, _06217_);
  or _83882_ (_33862_, _33861_, _33856_);
  and _83883_ (_33863_, _33862_, _33841_);
  or _83884_ (_33864_, _33863_, _06220_);
  or _83885_ (_33865_, _33849_, _06229_);
  and _83886_ (_33867_, _33865_, _06153_);
  and _83887_ (_33868_, _33867_, _33864_);
  and _83888_ (_33869_, _14349_, _08418_);
  or _83889_ (_33870_, _33869_, _33857_);
  and _83890_ (_33871_, _33870_, _06152_);
  or _83891_ (_33872_, _33871_, _06145_);
  or _83892_ (_33873_, _33872_, _33868_);
  and _83893_ (_33874_, _33858_, _14382_);
  or _83894_ (_33875_, _33857_, _06146_);
  or _83895_ (_33876_, _33875_, _33874_);
  and _83896_ (_33878_, _33876_, _33873_);
  and _83897_ (_33879_, _33878_, _06140_);
  and _83898_ (_33880_, _14351_, _08418_);
  or _83899_ (_33881_, _33857_, _33880_);
  and _83900_ (_33882_, _33881_, _06139_);
  or _83901_ (_33883_, _33882_, _09842_);
  or _83902_ (_33884_, _33883_, _33879_);
  or _83903_ (_33885_, _33840_, _06132_);
  and _83904_ (_33886_, _33885_, _33884_);
  or _83905_ (_33887_, _33886_, _06116_);
  and _83906_ (_33889_, _09115_, _07826_);
  or _83907_ (_33890_, _33835_, _06117_);
  or _83908_ (_33891_, _33890_, _33889_);
  and _83909_ (_33892_, _33891_, _06114_);
  and _83910_ (_33893_, _33892_, _33887_);
  and _83911_ (_33894_, _14442_, _07826_);
  or _83912_ (_33895_, _33894_, _33835_);
  and _83913_ (_33896_, _33895_, _05787_);
  or _83914_ (_33897_, _33896_, _33893_);
  and _83915_ (_33898_, _33897_, _06298_);
  or _83916_ (_33900_, _14346_, _13402_);
  and _83917_ (_33901_, _33900_, _06297_);
  nand _83918_ (_33902_, _07826_, _06945_);
  and _83919_ (_33903_, _33902_, _06110_);
  or _83920_ (_33904_, _33903_, _33901_);
  and _83921_ (_33905_, _33904_, _33842_);
  or _83922_ (_33906_, _33905_, _06402_);
  or _83923_ (_33907_, _33906_, _33898_);
  nand _83924_ (_33908_, _10275_, _07826_);
  and _83925_ (_33909_, _33908_, _33837_);
  or _83926_ (_33911_, _33909_, _07125_);
  and _83927_ (_33912_, _33911_, _07132_);
  and _83928_ (_33913_, _33912_, _33907_);
  or _83929_ (_33914_, _14344_, _13402_);
  and _83930_ (_33915_, _33842_, _06306_);
  and _83931_ (_33916_, _33915_, _33914_);
  or _83932_ (_33917_, _33916_, _06411_);
  or _83933_ (_33918_, _33917_, _33913_);
  nor _83934_ (_33919_, _33835_, _07130_);
  nand _83935_ (_33920_, _33919_, _33908_);
  and _83936_ (_33922_, _33920_, _08819_);
  and _83937_ (_33923_, _33922_, _33918_);
  or _83938_ (_33924_, _33902_, _08176_);
  and _83939_ (_33925_, _33842_, _06303_);
  and _83940_ (_33926_, _33925_, _33924_);
  or _83941_ (_33927_, _33926_, _06396_);
  or _83942_ (_33928_, _33927_, _33923_);
  and _83943_ (_33929_, _33928_, _33838_);
  or _83944_ (_33930_, _33929_, _06433_);
  or _83945_ (_33931_, _33846_, _06829_);
  and _83946_ (_33933_, _33931_, _05749_);
  and _83947_ (_33934_, _33933_, _33930_);
  and _83948_ (_33935_, _33870_, _05748_);
  or _83949_ (_33936_, _33935_, _06440_);
  or _83950_ (_33937_, _33936_, _33934_);
  or _83951_ (_33938_, _33835_, _06444_);
  or _83952_ (_33939_, _33938_, _33843_);
  and _83953_ (_33940_, _33939_, _01317_);
  and _83954_ (_33941_, _33940_, _33937_);
  or _83955_ (_33942_, _33941_, _33834_);
  and _83956_ (_43748_, _33942_, _43100_);
  and _83957_ (_33944_, _01321_, \oc8051_golden_model_1.IE [2]);
  and _83958_ (_33945_, _13402_, \oc8051_golden_model_1.IE [2]);
  and _83959_ (_33946_, _07826_, _07708_);
  or _83960_ (_33947_, _33946_, _33945_);
  or _83961_ (_33948_, _33947_, _06132_);
  or _83962_ (_33949_, _33947_, _07075_);
  and _83963_ (_33950_, _14542_, _07826_);
  or _83964_ (_33951_, _33950_, _33945_);
  or _83965_ (_33952_, _33951_, _06161_);
  and _83966_ (_33954_, _07826_, \oc8051_golden_model_1.ACC [2]);
  or _83967_ (_33955_, _33954_, _33945_);
  and _83968_ (_33956_, _33955_, _07056_);
  and _83969_ (_33957_, _07057_, \oc8051_golden_model_1.IE [2]);
  or _83970_ (_33958_, _33957_, _06160_);
  or _83971_ (_33959_, _33958_, _33956_);
  and _83972_ (_33960_, _33959_, _06157_);
  and _83973_ (_33961_, _33960_, _33952_);
  and _83974_ (_33962_, _13407_, \oc8051_golden_model_1.IE [2]);
  and _83975_ (_33963_, _14538_, _08418_);
  or _83976_ (_33965_, _33963_, _33962_);
  and _83977_ (_33966_, _33965_, _06156_);
  or _83978_ (_33967_, _33966_, _06217_);
  or _83979_ (_33968_, _33967_, _33961_);
  and _83980_ (_33969_, _33968_, _33949_);
  or _83981_ (_33970_, _33969_, _06220_);
  or _83982_ (_33971_, _33955_, _06229_);
  and _83983_ (_33972_, _33971_, _06153_);
  and _83984_ (_33973_, _33972_, _33970_);
  and _83985_ (_33974_, _14536_, _08418_);
  or _83986_ (_33976_, _33974_, _33962_);
  and _83987_ (_33977_, _33976_, _06152_);
  or _83988_ (_33978_, _33977_, _06145_);
  or _83989_ (_33979_, _33978_, _33973_);
  and _83990_ (_33980_, _33963_, _14569_);
  or _83991_ (_33981_, _33962_, _06146_);
  or _83992_ (_33982_, _33981_, _33980_);
  and _83993_ (_33983_, _33982_, _06140_);
  and _83994_ (_33984_, _33983_, _33979_);
  and _83995_ (_33985_, _14583_, _08418_);
  or _83996_ (_33987_, _33985_, _33962_);
  and _83997_ (_33988_, _33987_, _06139_);
  or _83998_ (_33989_, _33988_, _09842_);
  or _83999_ (_33990_, _33989_, _33984_);
  and _84000_ (_33991_, _33990_, _33948_);
  or _84001_ (_33992_, _33991_, _06116_);
  and _84002_ (_33993_, _09211_, _07826_);
  or _84003_ (_33994_, _33945_, _06117_);
  or _84004_ (_33995_, _33994_, _33993_);
  and _84005_ (_33996_, _33995_, _06114_);
  and _84006_ (_33998_, _33996_, _33992_);
  and _84007_ (_33999_, _14630_, _07826_);
  or _84008_ (_34000_, _33945_, _33999_);
  and _84009_ (_34001_, _34000_, _05787_);
  or _84010_ (_34002_, _34001_, _33998_);
  or _84011_ (_34003_, _34002_, _11136_);
  and _84012_ (_34004_, _14646_, _07826_);
  or _84013_ (_34005_, _33945_, _07127_);
  or _84014_ (_34006_, _34005_, _34004_);
  and _84015_ (_34007_, _07826_, _08768_);
  or _84016_ (_34009_, _34007_, _33945_);
  or _84017_ (_34010_, _34009_, _06111_);
  and _84018_ (_34011_, _34010_, _07125_);
  and _84019_ (_34012_, _34011_, _34006_);
  and _84020_ (_34013_, _34012_, _34003_);
  and _84021_ (_34014_, _10282_, _07826_);
  or _84022_ (_34015_, _34014_, _33945_);
  and _84023_ (_34016_, _34015_, _06402_);
  or _84024_ (_34017_, _34016_, _34013_);
  and _84025_ (_34018_, _34017_, _07132_);
  or _84026_ (_34020_, _33945_, _08248_);
  and _84027_ (_34021_, _34009_, _06306_);
  and _84028_ (_34022_, _34021_, _34020_);
  or _84029_ (_34023_, _34022_, _34018_);
  and _84030_ (_34024_, _34023_, _07130_);
  and _84031_ (_34025_, _33955_, _06411_);
  and _84032_ (_34026_, _34025_, _34020_);
  or _84033_ (_34027_, _34026_, _06303_);
  or _84034_ (_34028_, _34027_, _34024_);
  and _84035_ (_34029_, _14643_, _07826_);
  or _84036_ (_34031_, _33945_, _08819_);
  or _84037_ (_34032_, _34031_, _34029_);
  and _84038_ (_34033_, _34032_, _08824_);
  and _84039_ (_34034_, _34033_, _34028_);
  nor _84040_ (_34035_, _10281_, _13402_);
  or _84041_ (_34036_, _34035_, _33945_);
  and _84042_ (_34037_, _34036_, _06396_);
  or _84043_ (_34038_, _34037_, _06433_);
  or _84044_ (_34039_, _34038_, _34034_);
  or _84045_ (_34040_, _33951_, _06829_);
  and _84046_ (_34042_, _34040_, _05749_);
  and _84047_ (_34043_, _34042_, _34039_);
  and _84048_ (_34044_, _33976_, _05748_);
  or _84049_ (_34045_, _34044_, _06440_);
  or _84050_ (_34046_, _34045_, _34043_);
  and _84051_ (_34047_, _14710_, _07826_);
  or _84052_ (_34048_, _33945_, _06444_);
  or _84053_ (_34049_, _34048_, _34047_);
  and _84054_ (_34050_, _34049_, _01317_);
  and _84055_ (_34051_, _34050_, _34046_);
  or _84056_ (_34053_, _34051_, _33944_);
  and _84057_ (_43749_, _34053_, _43100_);
  and _84058_ (_34054_, _01321_, \oc8051_golden_model_1.IE [3]);
  and _84059_ (_34055_, _13402_, \oc8051_golden_model_1.IE [3]);
  and _84060_ (_34056_, _07826_, _07544_);
  or _84061_ (_34057_, _34056_, _34055_);
  or _84062_ (_34058_, _34057_, _06132_);
  and _84063_ (_34059_, _14738_, _07826_);
  or _84064_ (_34060_, _34059_, _34055_);
  or _84065_ (_34061_, _34060_, _06161_);
  and _84066_ (_34063_, _07826_, \oc8051_golden_model_1.ACC [3]);
  or _84067_ (_34064_, _34063_, _34055_);
  and _84068_ (_34065_, _34064_, _07056_);
  and _84069_ (_34066_, _07057_, \oc8051_golden_model_1.IE [3]);
  or _84070_ (_34067_, _34066_, _06160_);
  or _84071_ (_34068_, _34067_, _34065_);
  and _84072_ (_34069_, _34068_, _06157_);
  and _84073_ (_34070_, _34069_, _34061_);
  and _84074_ (_34071_, _13407_, \oc8051_golden_model_1.IE [3]);
  and _84075_ (_34072_, _14735_, _08418_);
  or _84076_ (_34074_, _34072_, _34071_);
  and _84077_ (_34075_, _34074_, _06156_);
  or _84078_ (_34076_, _34075_, _06217_);
  or _84079_ (_34077_, _34076_, _34070_);
  or _84080_ (_34078_, _34057_, _07075_);
  and _84081_ (_34079_, _34078_, _34077_);
  or _84082_ (_34080_, _34079_, _06220_);
  or _84083_ (_34081_, _34064_, _06229_);
  and _84084_ (_34082_, _34081_, _06153_);
  and _84085_ (_34083_, _34082_, _34080_);
  and _84086_ (_34085_, _14731_, _08418_);
  or _84087_ (_34086_, _34085_, _34071_);
  and _84088_ (_34087_, _34086_, _06152_);
  or _84089_ (_34088_, _34087_, _06145_);
  or _84090_ (_34089_, _34088_, _34083_);
  or _84091_ (_34090_, _34071_, _14764_);
  and _84092_ (_34091_, _34090_, _34074_);
  or _84093_ (_34092_, _34091_, _06146_);
  and _84094_ (_34093_, _34092_, _06140_);
  and _84095_ (_34094_, _34093_, _34089_);
  and _84096_ (_34096_, _14732_, _08418_);
  or _84097_ (_34097_, _34096_, _34071_);
  and _84098_ (_34098_, _34097_, _06139_);
  or _84099_ (_34099_, _34098_, _09842_);
  or _84100_ (_34100_, _34099_, _34094_);
  and _84101_ (_34101_, _34100_, _34058_);
  or _84102_ (_34102_, _34101_, _06116_);
  and _84103_ (_34103_, _09210_, _07826_);
  or _84104_ (_34104_, _34055_, _06117_);
  or _84105_ (_34105_, _34104_, _34103_);
  and _84106_ (_34107_, _34105_, _06114_);
  and _84107_ (_34108_, _34107_, _34102_);
  and _84108_ (_34109_, _14825_, _07826_);
  or _84109_ (_34110_, _34055_, _34109_);
  and _84110_ (_34111_, _34110_, _05787_);
  or _84111_ (_34112_, _34111_, _34108_);
  or _84112_ (_34113_, _34112_, _11136_);
  and _84113_ (_34114_, _14727_, _07826_);
  or _84114_ (_34115_, _34055_, _07127_);
  or _84115_ (_34116_, _34115_, _34114_);
  and _84116_ (_34118_, _07826_, _08712_);
  or _84117_ (_34119_, _34118_, _34055_);
  or _84118_ (_34120_, _34119_, _06111_);
  and _84119_ (_34121_, _34120_, _07125_);
  and _84120_ (_34122_, _34121_, _34116_);
  and _84121_ (_34123_, _34122_, _34113_);
  and _84122_ (_34124_, _12318_, _07826_);
  or _84123_ (_34125_, _34124_, _34055_);
  and _84124_ (_34126_, _34125_, _06402_);
  or _84125_ (_34127_, _34126_, _34123_);
  and _84126_ (_34129_, _34127_, _07132_);
  or _84127_ (_34130_, _34055_, _08140_);
  and _84128_ (_34131_, _34119_, _06306_);
  and _84129_ (_34132_, _34131_, _34130_);
  or _84130_ (_34133_, _34132_, _34129_);
  and _84131_ (_34134_, _34133_, _07130_);
  and _84132_ (_34135_, _34064_, _06411_);
  and _84133_ (_34136_, _34135_, _34130_);
  or _84134_ (_34137_, _34136_, _06303_);
  or _84135_ (_34138_, _34137_, _34134_);
  and _84136_ (_34140_, _14724_, _07826_);
  or _84137_ (_34141_, _34055_, _08819_);
  or _84138_ (_34142_, _34141_, _34140_);
  and _84139_ (_34143_, _34142_, _08824_);
  and _84140_ (_34144_, _34143_, _34138_);
  nor _84141_ (_34145_, _10273_, _13402_);
  or _84142_ (_34146_, _34145_, _34055_);
  and _84143_ (_34147_, _34146_, _06396_);
  or _84144_ (_34148_, _34147_, _06433_);
  or _84145_ (_34149_, _34148_, _34144_);
  or _84146_ (_34151_, _34060_, _06829_);
  and _84147_ (_34152_, _34151_, _05749_);
  and _84148_ (_34153_, _34152_, _34149_);
  and _84149_ (_34154_, _34086_, _05748_);
  or _84150_ (_34155_, _34154_, _06440_);
  or _84151_ (_34156_, _34155_, _34153_);
  and _84152_ (_34157_, _14897_, _07826_);
  or _84153_ (_34158_, _34055_, _06444_);
  or _84154_ (_34159_, _34158_, _34157_);
  and _84155_ (_34160_, _34159_, _01317_);
  and _84156_ (_34161_, _34160_, _34156_);
  or _84157_ (_34162_, _34161_, _34054_);
  and _84158_ (_43750_, _34162_, _43100_);
  and _84159_ (_34163_, _01321_, \oc8051_golden_model_1.IE [4]);
  and _84160_ (_34164_, _13402_, \oc8051_golden_model_1.IE [4]);
  and _84161_ (_34165_, _08336_, _07826_);
  or _84162_ (_34166_, _34165_, _34164_);
  or _84163_ (_34167_, _34166_, _06132_);
  and _84164_ (_34168_, _13407_, \oc8051_golden_model_1.IE [4]);
  and _84165_ (_34169_, _14942_, _08418_);
  or _84166_ (_34171_, _34169_, _34168_);
  and _84167_ (_34172_, _34171_, _06152_);
  and _84168_ (_34173_, _14928_, _07826_);
  or _84169_ (_34174_, _34173_, _34164_);
  or _84170_ (_34175_, _34174_, _06161_);
  and _84171_ (_34176_, _07826_, \oc8051_golden_model_1.ACC [4]);
  or _84172_ (_34177_, _34176_, _34164_);
  and _84173_ (_34178_, _34177_, _07056_);
  and _84174_ (_34179_, _07057_, \oc8051_golden_model_1.IE [4]);
  or _84175_ (_34180_, _34179_, _06160_);
  or _84176_ (_34182_, _34180_, _34178_);
  and _84177_ (_34183_, _34182_, _06157_);
  and _84178_ (_34184_, _34183_, _34175_);
  and _84179_ (_34185_, _14932_, _08418_);
  or _84180_ (_34186_, _34185_, _34168_);
  and _84181_ (_34187_, _34186_, _06156_);
  or _84182_ (_34188_, _34187_, _06217_);
  or _84183_ (_34189_, _34188_, _34184_);
  or _84184_ (_34190_, _34166_, _07075_);
  and _84185_ (_34191_, _34190_, _34189_);
  or _84186_ (_34193_, _34191_, _06220_);
  or _84187_ (_34194_, _34177_, _06229_);
  and _84188_ (_34195_, _34194_, _06153_);
  and _84189_ (_34196_, _34195_, _34193_);
  or _84190_ (_34197_, _34196_, _34172_);
  and _84191_ (_34198_, _34197_, _06146_);
  and _84192_ (_34199_, _14950_, _08418_);
  or _84193_ (_34200_, _34199_, _34168_);
  and _84194_ (_34201_, _34200_, _06145_);
  or _84195_ (_34202_, _34201_, _34198_);
  and _84196_ (_34204_, _34202_, _06140_);
  and _84197_ (_34205_, _14966_, _08418_);
  or _84198_ (_34206_, _34205_, _34168_);
  and _84199_ (_34207_, _34206_, _06139_);
  or _84200_ (_34208_, _34207_, _09842_);
  or _84201_ (_34209_, _34208_, _34204_);
  and _84202_ (_34210_, _34209_, _34167_);
  or _84203_ (_34211_, _34210_, _06116_);
  and _84204_ (_34212_, _09209_, _07826_);
  or _84205_ (_34213_, _34164_, _06117_);
  or _84206_ (_34215_, _34213_, _34212_);
  and _84207_ (_34216_, _34215_, _06114_);
  and _84208_ (_34217_, _34216_, _34211_);
  and _84209_ (_34218_, _15013_, _07826_);
  or _84210_ (_34219_, _34218_, _34164_);
  and _84211_ (_34220_, _34219_, _05787_);
  or _84212_ (_34221_, _34220_, _11136_);
  or _84213_ (_34222_, _34221_, _34217_);
  and _84214_ (_34223_, _15029_, _07826_);
  or _84215_ (_34224_, _34164_, _07127_);
  or _84216_ (_34226_, _34224_, _34223_);
  and _84217_ (_34227_, _08715_, _07826_);
  or _84218_ (_34228_, _34227_, _34164_);
  or _84219_ (_34229_, _34228_, _06111_);
  and _84220_ (_34230_, _34229_, _07125_);
  and _84221_ (_34231_, _34230_, _34226_);
  and _84222_ (_34232_, _34231_, _34222_);
  and _84223_ (_34233_, _10289_, _07826_);
  or _84224_ (_34234_, _34233_, _34164_);
  and _84225_ (_34235_, _34234_, _06402_);
  or _84226_ (_34237_, _34235_, _34232_);
  and _84227_ (_34238_, _34237_, _07132_);
  or _84228_ (_34239_, _34164_, _08339_);
  and _84229_ (_34240_, _34228_, _06306_);
  and _84230_ (_34241_, _34240_, _34239_);
  or _84231_ (_34242_, _34241_, _34238_);
  and _84232_ (_34243_, _34242_, _07130_);
  and _84233_ (_34244_, _34177_, _06411_);
  and _84234_ (_34245_, _34244_, _34239_);
  or _84235_ (_34246_, _34245_, _06303_);
  or _84236_ (_34248_, _34246_, _34243_);
  and _84237_ (_34249_, _15026_, _07826_);
  or _84238_ (_34250_, _34164_, _08819_);
  or _84239_ (_34251_, _34250_, _34249_);
  and _84240_ (_34252_, _34251_, _08824_);
  and _84241_ (_34253_, _34252_, _34248_);
  nor _84242_ (_34254_, _10288_, _13402_);
  or _84243_ (_34255_, _34254_, _34164_);
  and _84244_ (_34256_, _34255_, _06396_);
  or _84245_ (_34257_, _34256_, _06433_);
  or _84246_ (_34259_, _34257_, _34253_);
  or _84247_ (_34260_, _34174_, _06829_);
  and _84248_ (_34261_, _34260_, _05749_);
  and _84249_ (_34262_, _34261_, _34259_);
  and _84250_ (_34263_, _34171_, _05748_);
  or _84251_ (_34264_, _34263_, _06440_);
  or _84252_ (_34265_, _34264_, _34262_);
  and _84253_ (_34266_, _15087_, _07826_);
  or _84254_ (_34267_, _34164_, _06444_);
  or _84255_ (_34268_, _34267_, _34266_);
  and _84256_ (_34270_, _34268_, _01317_);
  and _84257_ (_34271_, _34270_, _34265_);
  or _84258_ (_34272_, _34271_, _34163_);
  and _84259_ (_43751_, _34272_, _43100_);
  and _84260_ (_34273_, _01321_, \oc8051_golden_model_1.IE [5]);
  and _84261_ (_34274_, _13402_, \oc8051_golden_model_1.IE [5]);
  and _84262_ (_34275_, _15119_, _07826_);
  or _84263_ (_34276_, _34275_, _34274_);
  or _84264_ (_34278_, _34276_, _06161_);
  and _84265_ (_34280_, _07826_, \oc8051_golden_model_1.ACC [5]);
  or _84266_ (_34283_, _34280_, _34274_);
  and _84267_ (_34285_, _34283_, _07056_);
  and _84268_ (_34287_, _07057_, \oc8051_golden_model_1.IE [5]);
  or _84269_ (_34289_, _34287_, _06160_);
  or _84270_ (_34291_, _34289_, _34285_);
  and _84271_ (_34293_, _34291_, _06157_);
  and _84272_ (_34295_, _34293_, _34278_);
  and _84273_ (_34297_, _13407_, \oc8051_golden_model_1.IE [5]);
  and _84274_ (_34298_, _15123_, _08418_);
  or _84275_ (_34299_, _34298_, _34297_);
  and _84276_ (_34301_, _34299_, _06156_);
  or _84277_ (_34302_, _34301_, _06217_);
  or _84278_ (_34303_, _34302_, _34295_);
  and _84279_ (_34304_, _08101_, _07826_);
  or _84280_ (_34305_, _34304_, _34274_);
  or _84281_ (_34306_, _34305_, _07075_);
  and _84282_ (_34307_, _34306_, _34303_);
  or _84283_ (_34308_, _34307_, _06220_);
  or _84284_ (_34309_, _34283_, _06229_);
  and _84285_ (_34310_, _34309_, _06153_);
  and _84286_ (_34312_, _34310_, _34308_);
  and _84287_ (_34313_, _15104_, _08418_);
  or _84288_ (_34314_, _34313_, _34297_);
  and _84289_ (_34315_, _34314_, _06152_);
  or _84290_ (_34316_, _34315_, _06145_);
  or _84291_ (_34317_, _34316_, _34312_);
  or _84292_ (_34318_, _34297_, _15138_);
  and _84293_ (_34319_, _34318_, _34299_);
  or _84294_ (_34320_, _34319_, _06146_);
  and _84295_ (_34321_, _34320_, _06140_);
  and _84296_ (_34323_, _34321_, _34317_);
  and _84297_ (_34324_, _15155_, _08418_);
  or _84298_ (_34325_, _34324_, _34297_);
  and _84299_ (_34326_, _34325_, _06139_);
  or _84300_ (_34327_, _34326_, _09842_);
  or _84301_ (_34328_, _34327_, _34323_);
  or _84302_ (_34329_, _34305_, _06132_);
  and _84303_ (_34330_, _34329_, _34328_);
  or _84304_ (_34331_, _34330_, _06116_);
  and _84305_ (_34332_, _09208_, _07826_);
  or _84306_ (_34334_, _34274_, _06117_);
  or _84307_ (_34335_, _34334_, _34332_);
  and _84308_ (_34336_, _34335_, _06114_);
  and _84309_ (_34337_, _34336_, _34331_);
  and _84310_ (_34338_, _15203_, _07826_);
  or _84311_ (_34339_, _34338_, _34274_);
  and _84312_ (_34340_, _34339_, _05787_);
  or _84313_ (_34341_, _34340_, _11136_);
  or _84314_ (_34342_, _34341_, _34337_);
  and _84315_ (_34343_, _15219_, _07826_);
  or _84316_ (_34345_, _34274_, _07127_);
  or _84317_ (_34346_, _34345_, _34343_);
  and _84318_ (_34347_, _08736_, _07826_);
  or _84319_ (_34348_, _34347_, _34274_);
  or _84320_ (_34349_, _34348_, _06111_);
  and _84321_ (_34350_, _34349_, _07125_);
  and _84322_ (_34351_, _34350_, _34346_);
  and _84323_ (_34352_, _34351_, _34342_);
  and _84324_ (_34353_, _12325_, _07826_);
  or _84325_ (_34354_, _34353_, _34274_);
  and _84326_ (_34356_, _34354_, _06402_);
  or _84327_ (_34357_, _34356_, _34352_);
  and _84328_ (_34358_, _34357_, _07132_);
  or _84329_ (_34359_, _34274_, _08104_);
  and _84330_ (_34360_, _34348_, _06306_);
  and _84331_ (_34361_, _34360_, _34359_);
  or _84332_ (_34362_, _34361_, _34358_);
  and _84333_ (_34363_, _34362_, _07130_);
  and _84334_ (_34364_, _34283_, _06411_);
  and _84335_ (_34365_, _34364_, _34359_);
  or _84336_ (_34367_, _34365_, _06303_);
  or _84337_ (_34368_, _34367_, _34363_);
  and _84338_ (_34369_, _15216_, _07826_);
  or _84339_ (_34370_, _34274_, _08819_);
  or _84340_ (_34371_, _34370_, _34369_);
  and _84341_ (_34372_, _34371_, _08824_);
  and _84342_ (_34373_, _34372_, _34368_);
  nor _84343_ (_34374_, _10269_, _13402_);
  or _84344_ (_34375_, _34374_, _34274_);
  and _84345_ (_34376_, _34375_, _06396_);
  or _84346_ (_34378_, _34376_, _06433_);
  or _84347_ (_34379_, _34378_, _34373_);
  or _84348_ (_34380_, _34276_, _06829_);
  and _84349_ (_34381_, _34380_, _05749_);
  and _84350_ (_34382_, _34381_, _34379_);
  and _84351_ (_34383_, _34314_, _05748_);
  or _84352_ (_34384_, _34383_, _06440_);
  or _84353_ (_34385_, _34384_, _34382_);
  and _84354_ (_34386_, _15275_, _07826_);
  or _84355_ (_34387_, _34274_, _06444_);
  or _84356_ (_34389_, _34387_, _34386_);
  and _84357_ (_34390_, _34389_, _01317_);
  and _84358_ (_34391_, _34390_, _34385_);
  or _84359_ (_34392_, _34391_, _34273_);
  and _84360_ (_43752_, _34392_, _43100_);
  and _84361_ (_34393_, _01321_, \oc8051_golden_model_1.IE [6]);
  and _84362_ (_34394_, _13402_, \oc8051_golden_model_1.IE [6]);
  and _84363_ (_34395_, _15300_, _07826_);
  or _84364_ (_34396_, _34395_, _34394_);
  or _84365_ (_34397_, _34396_, _06161_);
  and _84366_ (_34399_, _07826_, \oc8051_golden_model_1.ACC [6]);
  or _84367_ (_34400_, _34399_, _34394_);
  and _84368_ (_34401_, _34400_, _07056_);
  and _84369_ (_34402_, _07057_, \oc8051_golden_model_1.IE [6]);
  or _84370_ (_34403_, _34402_, _06160_);
  or _84371_ (_34404_, _34403_, _34401_);
  and _84372_ (_34405_, _34404_, _06157_);
  and _84373_ (_34406_, _34405_, _34397_);
  and _84374_ (_34407_, _13407_, \oc8051_golden_model_1.IE [6]);
  and _84375_ (_34408_, _15316_, _08418_);
  or _84376_ (_34410_, _34408_, _34407_);
  and _84377_ (_34411_, _34410_, _06156_);
  or _84378_ (_34412_, _34411_, _06217_);
  or _84379_ (_34413_, _34412_, _34406_);
  and _84380_ (_34414_, _08012_, _07826_);
  or _84381_ (_34415_, _34414_, _34394_);
  or _84382_ (_34416_, _34415_, _07075_);
  and _84383_ (_34417_, _34416_, _34413_);
  or _84384_ (_34418_, _34417_, _06220_);
  or _84385_ (_34419_, _34400_, _06229_);
  and _84386_ (_34421_, _34419_, _06153_);
  and _84387_ (_34422_, _34421_, _34418_);
  and _84388_ (_34423_, _15297_, _08418_);
  or _84389_ (_34424_, _34423_, _34407_);
  and _84390_ (_34425_, _34424_, _06152_);
  or _84391_ (_34426_, _34425_, _06145_);
  or _84392_ (_34427_, _34426_, _34422_);
  or _84393_ (_34428_, _34407_, _15331_);
  and _84394_ (_34429_, _34428_, _34410_);
  or _84395_ (_34430_, _34429_, _06146_);
  and _84396_ (_34432_, _34430_, _06140_);
  and _84397_ (_34433_, _34432_, _34427_);
  and _84398_ (_34434_, _15348_, _08418_);
  or _84399_ (_34435_, _34434_, _34407_);
  and _84400_ (_34436_, _34435_, _06139_);
  or _84401_ (_34437_, _34436_, _09842_);
  or _84402_ (_34438_, _34437_, _34433_);
  or _84403_ (_34439_, _34415_, _06132_);
  and _84404_ (_34440_, _34439_, _34438_);
  or _84405_ (_34441_, _34440_, _06116_);
  and _84406_ (_34443_, _09207_, _07826_);
  or _84407_ (_34444_, _34394_, _06117_);
  or _84408_ (_34445_, _34444_, _34443_);
  and _84409_ (_34446_, _34445_, _06114_);
  and _84410_ (_34447_, _34446_, _34441_);
  and _84411_ (_34448_, _15395_, _07826_);
  or _84412_ (_34449_, _34448_, _34394_);
  and _84413_ (_34450_, _34449_, _05787_);
  or _84414_ (_34451_, _34450_, _11136_);
  or _84415_ (_34452_, _34451_, _34447_);
  and _84416_ (_34454_, _15413_, _07826_);
  or _84417_ (_34455_, _34394_, _07127_);
  or _84418_ (_34456_, _34455_, _34454_);
  and _84419_ (_34457_, _15402_, _07826_);
  or _84420_ (_34458_, _34457_, _34394_);
  or _84421_ (_34459_, _34458_, _06111_);
  and _84422_ (_34460_, _34459_, _07125_);
  and _84423_ (_34461_, _34460_, _34456_);
  and _84424_ (_34462_, _34461_, _34452_);
  and _84425_ (_34463_, _10295_, _07826_);
  or _84426_ (_34465_, _34463_, _34394_);
  and _84427_ (_34466_, _34465_, _06402_);
  or _84428_ (_34467_, _34466_, _34462_);
  and _84429_ (_34468_, _34467_, _07132_);
  or _84430_ (_34469_, _34394_, _08015_);
  and _84431_ (_34470_, _34458_, _06306_);
  and _84432_ (_34471_, _34470_, _34469_);
  or _84433_ (_34472_, _34471_, _34468_);
  and _84434_ (_34473_, _34472_, _07130_);
  and _84435_ (_34474_, _34400_, _06411_);
  and _84436_ (_34476_, _34474_, _34469_);
  or _84437_ (_34477_, _34476_, _06303_);
  or _84438_ (_34478_, _34477_, _34473_);
  and _84439_ (_34479_, _15410_, _07826_);
  or _84440_ (_34480_, _34394_, _08819_);
  or _84441_ (_34481_, _34480_, _34479_);
  and _84442_ (_34482_, _34481_, _08824_);
  and _84443_ (_34483_, _34482_, _34478_);
  nor _84444_ (_34484_, _10294_, _13402_);
  or _84445_ (_34485_, _34484_, _34394_);
  and _84446_ (_34487_, _34485_, _06396_);
  or _84447_ (_34488_, _34487_, _06433_);
  or _84448_ (_34489_, _34488_, _34483_);
  or _84449_ (_34490_, _34396_, _06829_);
  and _84450_ (_34491_, _34490_, _05749_);
  and _84451_ (_34492_, _34491_, _34489_);
  and _84452_ (_34493_, _34424_, _05748_);
  or _84453_ (_34494_, _34493_, _06440_);
  or _84454_ (_34495_, _34494_, _34492_);
  and _84455_ (_34496_, _15478_, _07826_);
  or _84456_ (_34498_, _34394_, _06444_);
  or _84457_ (_34499_, _34498_, _34496_);
  and _84458_ (_34500_, _34499_, _01317_);
  and _84459_ (_34501_, _34500_, _34495_);
  or _84460_ (_34502_, _34501_, _34393_);
  and _84461_ (_43753_, _34502_, _43100_);
  not _84462_ (_34503_, \oc8051_golden_model_1.SCON [0]);
  nor _84463_ (_34504_, _01317_, _34503_);
  nor _84464_ (_34505_, _07778_, _34503_);
  and _84465_ (_34506_, _07778_, _07049_);
  or _84466_ (_34508_, _34506_, _34505_);
  or _84467_ (_34509_, _34508_, _06132_);
  nor _84468_ (_34510_, _08211_, _13504_);
  or _84469_ (_34511_, _34510_, _34505_);
  or _84470_ (_34512_, _34511_, _06161_);
  and _84471_ (_34513_, _07778_, \oc8051_golden_model_1.ACC [0]);
  or _84472_ (_34514_, _34513_, _34505_);
  and _84473_ (_34515_, _34514_, _07056_);
  nor _84474_ (_34516_, _07056_, _34503_);
  or _84475_ (_34517_, _34516_, _06160_);
  or _84476_ (_34519_, _34517_, _34515_);
  and _84477_ (_34520_, _34519_, _06157_);
  and _84478_ (_34521_, _34520_, _34512_);
  nor _84479_ (_34522_, _08413_, _34503_);
  and _84480_ (_34523_, _14169_, _08413_);
  or _84481_ (_34524_, _34523_, _34522_);
  and _84482_ (_34525_, _34524_, _06156_);
  or _84483_ (_34526_, _34525_, _34521_);
  and _84484_ (_34527_, _34526_, _07075_);
  and _84485_ (_34528_, _34508_, _06217_);
  or _84486_ (_34530_, _34528_, _06220_);
  or _84487_ (_34531_, _34530_, _34527_);
  or _84488_ (_34532_, _34514_, _06229_);
  and _84489_ (_34533_, _34532_, _06153_);
  and _84490_ (_34534_, _34533_, _34531_);
  and _84491_ (_34535_, _34505_, _06152_);
  or _84492_ (_34536_, _34535_, _06145_);
  or _84493_ (_34537_, _34536_, _34534_);
  or _84494_ (_34538_, _34511_, _06146_);
  and _84495_ (_34539_, _34538_, _06140_);
  and _84496_ (_34541_, _34539_, _34537_);
  or _84497_ (_34542_, _34522_, _14170_);
  and _84498_ (_34543_, _34542_, _06139_);
  and _84499_ (_34544_, _34543_, _34524_);
  or _84500_ (_34545_, _34544_, _09842_);
  or _84501_ (_34546_, _34545_, _34541_);
  and _84502_ (_34547_, _34546_, _34509_);
  or _84503_ (_34548_, _34547_, _06116_);
  and _84504_ (_34549_, _09160_, _07778_);
  or _84505_ (_34550_, _34505_, _06117_);
  or _84506_ (_34552_, _34550_, _34549_);
  and _84507_ (_34553_, _34552_, _06114_);
  and _84508_ (_34554_, _34553_, _34548_);
  and _84509_ (_34555_, _14260_, _07778_);
  or _84510_ (_34556_, _34555_, _34505_);
  and _84511_ (_34557_, _34556_, _05787_);
  or _84512_ (_34558_, _34557_, _34554_);
  or _84513_ (_34559_, _34558_, _11136_);
  and _84514_ (_34560_, _14275_, _07778_);
  or _84515_ (_34561_, _34505_, _07127_);
  or _84516_ (_34563_, _34561_, _34560_);
  and _84517_ (_34564_, _07778_, _08708_);
  or _84518_ (_34565_, _34564_, _34505_);
  or _84519_ (_34566_, _34565_, _06111_);
  and _84520_ (_34567_, _34566_, _07125_);
  and _84521_ (_34568_, _34567_, _34563_);
  and _84522_ (_34569_, _34568_, _34559_);
  nor _84523_ (_34570_, _12321_, _13504_);
  or _84524_ (_34571_, _34570_, _34505_);
  nand _84525_ (_34572_, _10276_, _07778_);
  and _84526_ (_34574_, _34572_, _06402_);
  and _84527_ (_34575_, _34574_, _34571_);
  or _84528_ (_34576_, _34575_, _34569_);
  and _84529_ (_34577_, _34576_, _07132_);
  nand _84530_ (_34578_, _34565_, _06306_);
  nor _84531_ (_34579_, _34578_, _34510_);
  or _84532_ (_34580_, _34579_, _06411_);
  or _84533_ (_34581_, _34580_, _34577_);
  nor _84534_ (_34582_, _34505_, _07130_);
  nand _84535_ (_34583_, _34582_, _34572_);
  and _84536_ (_34585_, _34583_, _34581_);
  or _84537_ (_34586_, _34585_, _06303_);
  and _84538_ (_34587_, _14167_, _07778_);
  or _84539_ (_34588_, _34505_, _08819_);
  or _84540_ (_34589_, _34588_, _34587_);
  and _84541_ (_34590_, _34589_, _08824_);
  and _84542_ (_34591_, _34590_, _34586_);
  and _84543_ (_34592_, _34571_, _06396_);
  or _84544_ (_34593_, _34592_, _06433_);
  or _84545_ (_34594_, _34593_, _34591_);
  or _84546_ (_34596_, _34511_, _06829_);
  and _84547_ (_34597_, _34596_, _34594_);
  or _84548_ (_34598_, _34597_, _05748_);
  or _84549_ (_34599_, _34505_, _05749_);
  and _84550_ (_34600_, _34599_, _34598_);
  or _84551_ (_34601_, _34600_, _06440_);
  or _84552_ (_34602_, _34511_, _06444_);
  and _84553_ (_34603_, _34602_, _01317_);
  and _84554_ (_34604_, _34603_, _34601_);
  or _84555_ (_34605_, _34604_, _34504_);
  and _84556_ (_43755_, _34605_, _43100_);
  not _84557_ (_34607_, \oc8051_golden_model_1.SCON [1]);
  nor _84558_ (_34608_, _01317_, _34607_);
  nor _84559_ (_34609_, _07778_, _34607_);
  and _84560_ (_34610_, _07778_, _07306_);
  or _84561_ (_34611_, _34610_, _34609_);
  or _84562_ (_34612_, _34611_, _07075_);
  or _84563_ (_34613_, _07778_, \oc8051_golden_model_1.SCON [1]);
  and _84564_ (_34614_, _14363_, _07778_);
  not _84565_ (_34615_, _34614_);
  and _84566_ (_34617_, _34615_, _34613_);
  or _84567_ (_34618_, _34617_, _06161_);
  and _84568_ (_34619_, _07778_, \oc8051_golden_model_1.ACC [1]);
  or _84569_ (_34620_, _34619_, _34609_);
  and _84570_ (_34621_, _34620_, _07056_);
  nor _84571_ (_34622_, _07056_, _34607_);
  or _84572_ (_34623_, _34622_, _06160_);
  or _84573_ (_34624_, _34623_, _34621_);
  and _84574_ (_34625_, _34624_, _06157_);
  and _84575_ (_34626_, _34625_, _34618_);
  nor _84576_ (_34628_, _08413_, _34607_);
  and _84577_ (_34629_, _14367_, _08413_);
  or _84578_ (_34630_, _34629_, _34628_);
  and _84579_ (_34631_, _34630_, _06156_);
  or _84580_ (_34632_, _34631_, _06217_);
  or _84581_ (_34633_, _34632_, _34626_);
  and _84582_ (_34634_, _34633_, _34612_);
  or _84583_ (_34635_, _34634_, _06220_);
  or _84584_ (_34636_, _34620_, _06229_);
  and _84585_ (_34637_, _34636_, _06153_);
  and _84586_ (_34639_, _34637_, _34635_);
  and _84587_ (_34640_, _14349_, _08413_);
  or _84588_ (_34641_, _34640_, _34628_);
  and _84589_ (_34642_, _34641_, _06152_);
  or _84590_ (_34643_, _34642_, _06145_);
  or _84591_ (_34644_, _34643_, _34639_);
  and _84592_ (_34645_, _34629_, _14382_);
  or _84593_ (_34646_, _34628_, _06146_);
  or _84594_ (_34647_, _34646_, _34645_);
  and _84595_ (_34648_, _34647_, _34644_);
  and _84596_ (_34650_, _34648_, _06140_);
  and _84597_ (_34651_, _14351_, _08413_);
  or _84598_ (_34652_, _34628_, _34651_);
  and _84599_ (_34653_, _34652_, _06139_);
  or _84600_ (_34654_, _34653_, _09842_);
  or _84601_ (_34655_, _34654_, _34650_);
  or _84602_ (_34656_, _34611_, _06132_);
  and _84603_ (_34657_, _34656_, _34655_);
  or _84604_ (_34658_, _34657_, _06116_);
  and _84605_ (_34659_, _09115_, _07778_);
  or _84606_ (_34661_, _34609_, _06117_);
  or _84607_ (_34662_, _34661_, _34659_);
  and _84608_ (_34663_, _34662_, _06114_);
  and _84609_ (_34664_, _34663_, _34658_);
  and _84610_ (_34665_, _14442_, _07778_);
  or _84611_ (_34666_, _34665_, _34609_);
  and _84612_ (_34667_, _34666_, _05787_);
  or _84613_ (_34668_, _34667_, _34664_);
  and _84614_ (_34669_, _34668_, _06298_);
  or _84615_ (_34670_, _14346_, _13504_);
  and _84616_ (_34672_, _34613_, _06297_);
  and _84617_ (_34673_, _34672_, _34670_);
  nand _84618_ (_34674_, _07778_, _06945_);
  and _84619_ (_34675_, _34674_, _06110_);
  and _84620_ (_34676_, _34675_, _34613_);
  or _84621_ (_34677_, _34676_, _06402_);
  or _84622_ (_34678_, _34677_, _34673_);
  or _84623_ (_34679_, _34678_, _34669_);
  nor _84624_ (_34680_, _10277_, _13504_);
  or _84625_ (_34681_, _34680_, _34609_);
  nand _84626_ (_34683_, _10275_, _07778_);
  and _84627_ (_34684_, _34683_, _34681_);
  or _84628_ (_34685_, _34684_, _07125_);
  and _84629_ (_34686_, _34685_, _07132_);
  and _84630_ (_34687_, _34686_, _34679_);
  or _84631_ (_34688_, _14344_, _13504_);
  and _84632_ (_34689_, _34613_, _06306_);
  and _84633_ (_34690_, _34689_, _34688_);
  or _84634_ (_34691_, _34690_, _06411_);
  or _84635_ (_34692_, _34691_, _34687_);
  nor _84636_ (_34694_, _34609_, _07130_);
  nand _84637_ (_34695_, _34694_, _34683_);
  and _84638_ (_34696_, _34695_, _08819_);
  and _84639_ (_34697_, _34696_, _34692_);
  or _84640_ (_34698_, _34674_, _08176_);
  and _84641_ (_34699_, _34613_, _06303_);
  and _84642_ (_34700_, _34699_, _34698_);
  or _84643_ (_34701_, _34700_, _06396_);
  or _84644_ (_34702_, _34701_, _34697_);
  or _84645_ (_34703_, _34681_, _08824_);
  and _84646_ (_34705_, _34703_, _34702_);
  or _84647_ (_34706_, _34705_, _06433_);
  or _84648_ (_34707_, _34617_, _06829_);
  and _84649_ (_34708_, _34707_, _05749_);
  and _84650_ (_34709_, _34708_, _34706_);
  and _84651_ (_34710_, _34641_, _05748_);
  or _84652_ (_34711_, _34710_, _06440_);
  or _84653_ (_34712_, _34711_, _34709_);
  or _84654_ (_34713_, _34609_, _06444_);
  or _84655_ (_34714_, _34713_, _34614_);
  and _84656_ (_34716_, _34714_, _01317_);
  and _84657_ (_34717_, _34716_, _34712_);
  or _84658_ (_34718_, _34717_, _34608_);
  and _84659_ (_43756_, _34718_, _43100_);
  and _84660_ (_34719_, _01321_, \oc8051_golden_model_1.SCON [2]);
  and _84661_ (_34720_, _13504_, \oc8051_golden_model_1.SCON [2]);
  and _84662_ (_34721_, _07778_, _07708_);
  or _84663_ (_34722_, _34721_, _34720_);
  or _84664_ (_34723_, _34722_, _06132_);
  or _84665_ (_34724_, _34722_, _07075_);
  and _84666_ (_34726_, _14542_, _07778_);
  or _84667_ (_34727_, _34726_, _34720_);
  or _84668_ (_34728_, _34727_, _06161_);
  and _84669_ (_34729_, _07778_, \oc8051_golden_model_1.ACC [2]);
  or _84670_ (_34730_, _34729_, _34720_);
  and _84671_ (_34731_, _34730_, _07056_);
  and _84672_ (_34732_, _07057_, \oc8051_golden_model_1.SCON [2]);
  or _84673_ (_34733_, _34732_, _06160_);
  or _84674_ (_34734_, _34733_, _34731_);
  and _84675_ (_34735_, _34734_, _06157_);
  and _84676_ (_34737_, _34735_, _34728_);
  and _84677_ (_34738_, _13509_, \oc8051_golden_model_1.SCON [2]);
  and _84678_ (_34739_, _14538_, _08413_);
  or _84679_ (_34740_, _34739_, _34738_);
  and _84680_ (_34741_, _34740_, _06156_);
  or _84681_ (_34742_, _34741_, _06217_);
  or _84682_ (_34743_, _34742_, _34737_);
  and _84683_ (_34744_, _34743_, _34724_);
  or _84684_ (_34745_, _34744_, _06220_);
  or _84685_ (_34746_, _34730_, _06229_);
  and _84686_ (_34748_, _34746_, _06153_);
  and _84687_ (_34749_, _34748_, _34745_);
  and _84688_ (_34750_, _14536_, _08413_);
  or _84689_ (_34751_, _34750_, _34738_);
  and _84690_ (_34752_, _34751_, _06152_);
  or _84691_ (_34753_, _34752_, _06145_);
  or _84692_ (_34754_, _34753_, _34749_);
  and _84693_ (_34755_, _34739_, _14569_);
  or _84694_ (_34756_, _34738_, _06146_);
  or _84695_ (_34757_, _34756_, _34755_);
  and _84696_ (_34759_, _34757_, _06140_);
  and _84697_ (_34760_, _34759_, _34754_);
  and _84698_ (_34761_, _14583_, _08413_);
  or _84699_ (_34762_, _34761_, _34738_);
  and _84700_ (_34763_, _34762_, _06139_);
  or _84701_ (_34764_, _34763_, _09842_);
  or _84702_ (_34765_, _34764_, _34760_);
  and _84703_ (_34766_, _34765_, _34723_);
  or _84704_ (_34767_, _34766_, _06116_);
  and _84705_ (_34768_, _09211_, _07778_);
  or _84706_ (_34770_, _34720_, _06117_);
  or _84707_ (_34771_, _34770_, _34768_);
  and _84708_ (_34772_, _34771_, _06114_);
  and _84709_ (_34773_, _34772_, _34767_);
  and _84710_ (_34774_, _14630_, _07778_);
  or _84711_ (_34775_, _34720_, _34774_);
  and _84712_ (_34776_, _34775_, _05787_);
  or _84713_ (_34777_, _34776_, _34773_);
  or _84714_ (_34778_, _34777_, _11136_);
  and _84715_ (_34779_, _14646_, _07778_);
  or _84716_ (_34781_, _34720_, _07127_);
  or _84717_ (_34782_, _34781_, _34779_);
  and _84718_ (_34783_, _07778_, _08768_);
  or _84719_ (_34784_, _34783_, _34720_);
  or _84720_ (_34785_, _34784_, _06111_);
  and _84721_ (_34786_, _34785_, _07125_);
  and _84722_ (_34787_, _34786_, _34782_);
  and _84723_ (_34788_, _34787_, _34778_);
  and _84724_ (_34789_, _10282_, _07778_);
  or _84725_ (_34790_, _34789_, _34720_);
  and _84726_ (_34792_, _34790_, _06402_);
  or _84727_ (_34793_, _34792_, _34788_);
  and _84728_ (_34794_, _34793_, _07132_);
  or _84729_ (_34795_, _34720_, _08248_);
  and _84730_ (_34796_, _34784_, _06306_);
  and _84731_ (_34797_, _34796_, _34795_);
  or _84732_ (_34798_, _34797_, _34794_);
  and _84733_ (_34799_, _34798_, _07130_);
  and _84734_ (_34800_, _34730_, _06411_);
  and _84735_ (_34801_, _34800_, _34795_);
  or _84736_ (_34803_, _34801_, _06303_);
  or _84737_ (_34804_, _34803_, _34799_);
  and _84738_ (_34805_, _14643_, _07778_);
  or _84739_ (_34806_, _34720_, _08819_);
  or _84740_ (_34807_, _34806_, _34805_);
  and _84741_ (_34808_, _34807_, _08824_);
  and _84742_ (_34809_, _34808_, _34804_);
  nor _84743_ (_34810_, _10281_, _13504_);
  or _84744_ (_34811_, _34810_, _34720_);
  and _84745_ (_34812_, _34811_, _06396_);
  or _84746_ (_34814_, _34812_, _06433_);
  or _84747_ (_34815_, _34814_, _34809_);
  or _84748_ (_34816_, _34727_, _06829_);
  and _84749_ (_34817_, _34816_, _05749_);
  and _84750_ (_34818_, _34817_, _34815_);
  and _84751_ (_34819_, _34751_, _05748_);
  or _84752_ (_34820_, _34819_, _06440_);
  or _84753_ (_34821_, _34820_, _34818_);
  and _84754_ (_34822_, _14710_, _07778_);
  or _84755_ (_34823_, _34720_, _06444_);
  or _84756_ (_34825_, _34823_, _34822_);
  and _84757_ (_34826_, _34825_, _01317_);
  and _84758_ (_34827_, _34826_, _34821_);
  or _84759_ (_34828_, _34827_, _34719_);
  and _84760_ (_43757_, _34828_, _43100_);
  and _84761_ (_34829_, _01321_, \oc8051_golden_model_1.SCON [3]);
  and _84762_ (_34830_, _13504_, \oc8051_golden_model_1.SCON [3]);
  and _84763_ (_34831_, _07778_, _07544_);
  or _84764_ (_34832_, _34831_, _34830_);
  or _84765_ (_34833_, _34832_, _06132_);
  and _84766_ (_34835_, _14738_, _07778_);
  or _84767_ (_34836_, _34835_, _34830_);
  or _84768_ (_34837_, _34836_, _06161_);
  and _84769_ (_34838_, _07778_, \oc8051_golden_model_1.ACC [3]);
  or _84770_ (_34839_, _34838_, _34830_);
  and _84771_ (_34840_, _34839_, _07056_);
  and _84772_ (_34841_, _07057_, \oc8051_golden_model_1.SCON [3]);
  or _84773_ (_34842_, _34841_, _06160_);
  or _84774_ (_34843_, _34842_, _34840_);
  and _84775_ (_34844_, _34843_, _06157_);
  and _84776_ (_34846_, _34844_, _34837_);
  and _84777_ (_34847_, _13509_, \oc8051_golden_model_1.SCON [3]);
  and _84778_ (_34848_, _14735_, _08413_);
  or _84779_ (_34849_, _34848_, _34847_);
  and _84780_ (_34850_, _34849_, _06156_);
  or _84781_ (_34851_, _34850_, _06217_);
  or _84782_ (_34852_, _34851_, _34846_);
  or _84783_ (_34853_, _34832_, _07075_);
  and _84784_ (_34854_, _34853_, _34852_);
  or _84785_ (_34855_, _34854_, _06220_);
  or _84786_ (_34857_, _34839_, _06229_);
  and _84787_ (_34858_, _34857_, _06153_);
  and _84788_ (_34859_, _34858_, _34855_);
  and _84789_ (_34860_, _14731_, _08413_);
  or _84790_ (_34861_, _34860_, _34847_);
  and _84791_ (_34862_, _34861_, _06152_);
  or _84792_ (_34863_, _34862_, _06145_);
  or _84793_ (_34864_, _34863_, _34859_);
  or _84794_ (_34865_, _34847_, _14764_);
  and _84795_ (_34866_, _34865_, _34849_);
  or _84796_ (_34868_, _34866_, _06146_);
  and _84797_ (_34869_, _34868_, _06140_);
  and _84798_ (_34870_, _34869_, _34864_);
  and _84799_ (_34871_, _14732_, _08413_);
  or _84800_ (_34872_, _34871_, _34847_);
  and _84801_ (_34873_, _34872_, _06139_);
  or _84802_ (_34874_, _34873_, _09842_);
  or _84803_ (_34875_, _34874_, _34870_);
  and _84804_ (_34876_, _34875_, _34833_);
  or _84805_ (_34877_, _34876_, _06116_);
  and _84806_ (_34879_, _09210_, _07778_);
  or _84807_ (_34880_, _34830_, _06117_);
  or _84808_ (_34881_, _34880_, _34879_);
  and _84809_ (_34882_, _34881_, _06114_);
  and _84810_ (_34883_, _34882_, _34877_);
  and _84811_ (_34884_, _14825_, _07778_);
  or _84812_ (_34885_, _34830_, _34884_);
  and _84813_ (_34886_, _34885_, _05787_);
  or _84814_ (_34887_, _34886_, _34883_);
  or _84815_ (_34888_, _34887_, _11136_);
  and _84816_ (_34890_, _14727_, _07778_);
  or _84817_ (_34891_, _34830_, _07127_);
  or _84818_ (_34892_, _34891_, _34890_);
  and _84819_ (_34893_, _07778_, _08712_);
  or _84820_ (_34894_, _34893_, _34830_);
  or _84821_ (_34895_, _34894_, _06111_);
  and _84822_ (_34896_, _34895_, _07125_);
  and _84823_ (_34897_, _34896_, _34892_);
  and _84824_ (_34898_, _34897_, _34888_);
  and _84825_ (_34899_, _12318_, _07778_);
  or _84826_ (_34901_, _34899_, _34830_);
  and _84827_ (_34902_, _34901_, _06402_);
  or _84828_ (_34903_, _34902_, _34898_);
  and _84829_ (_34904_, _34903_, _07132_);
  or _84830_ (_34905_, _34830_, _08140_);
  and _84831_ (_34906_, _34894_, _06306_);
  and _84832_ (_34907_, _34906_, _34905_);
  or _84833_ (_34908_, _34907_, _34904_);
  and _84834_ (_34909_, _34908_, _07130_);
  and _84835_ (_34910_, _34839_, _06411_);
  and _84836_ (_34912_, _34910_, _34905_);
  or _84837_ (_34913_, _34912_, _06303_);
  or _84838_ (_34914_, _34913_, _34909_);
  and _84839_ (_34915_, _14724_, _07778_);
  or _84840_ (_34916_, _34830_, _08819_);
  or _84841_ (_34917_, _34916_, _34915_);
  and _84842_ (_34918_, _34917_, _08824_);
  and _84843_ (_34919_, _34918_, _34914_);
  nor _84844_ (_34920_, _10273_, _13504_);
  or _84845_ (_34921_, _34920_, _34830_);
  and _84846_ (_34923_, _34921_, _06396_);
  or _84847_ (_34924_, _34923_, _06433_);
  or _84848_ (_34925_, _34924_, _34919_);
  or _84849_ (_34926_, _34836_, _06829_);
  and _84850_ (_34927_, _34926_, _05749_);
  and _84851_ (_34928_, _34927_, _34925_);
  and _84852_ (_34929_, _34861_, _05748_);
  or _84853_ (_34930_, _34929_, _06440_);
  or _84854_ (_34931_, _34930_, _34928_);
  and _84855_ (_34932_, _14897_, _07778_);
  or _84856_ (_34933_, _34830_, _06444_);
  or _84857_ (_34934_, _34933_, _34932_);
  and _84858_ (_34935_, _34934_, _01317_);
  and _84859_ (_34936_, _34935_, _34931_);
  or _84860_ (_34937_, _34936_, _34829_);
  and _84861_ (_43758_, _34937_, _43100_);
  and _84862_ (_34938_, _01321_, \oc8051_golden_model_1.SCON [4]);
  and _84863_ (_34939_, _13504_, \oc8051_golden_model_1.SCON [4]);
  and _84864_ (_34940_, _08336_, _07778_);
  or _84865_ (_34941_, _34940_, _34939_);
  or _84866_ (_34943_, _34941_, _06132_);
  and _84867_ (_34944_, _13509_, \oc8051_golden_model_1.SCON [4]);
  and _84868_ (_34945_, _14942_, _08413_);
  or _84869_ (_34946_, _34945_, _34944_);
  and _84870_ (_34947_, _34946_, _06152_);
  and _84871_ (_34948_, _14928_, _07778_);
  or _84872_ (_34949_, _34948_, _34939_);
  or _84873_ (_34950_, _34949_, _06161_);
  and _84874_ (_34951_, _07778_, \oc8051_golden_model_1.ACC [4]);
  or _84875_ (_34952_, _34951_, _34939_);
  and _84876_ (_34954_, _34952_, _07056_);
  and _84877_ (_34955_, _07057_, \oc8051_golden_model_1.SCON [4]);
  or _84878_ (_34956_, _34955_, _06160_);
  or _84879_ (_34957_, _34956_, _34954_);
  and _84880_ (_34958_, _34957_, _06157_);
  and _84881_ (_34959_, _34958_, _34950_);
  and _84882_ (_34960_, _14932_, _08413_);
  or _84883_ (_34961_, _34960_, _34944_);
  and _84884_ (_34962_, _34961_, _06156_);
  or _84885_ (_34963_, _34962_, _06217_);
  or _84886_ (_34965_, _34963_, _34959_);
  or _84887_ (_34966_, _34941_, _07075_);
  and _84888_ (_34967_, _34966_, _34965_);
  or _84889_ (_34968_, _34967_, _06220_);
  or _84890_ (_34969_, _34952_, _06229_);
  and _84891_ (_34970_, _34969_, _06153_);
  and _84892_ (_34971_, _34970_, _34968_);
  or _84893_ (_34972_, _34971_, _34947_);
  and _84894_ (_34973_, _34972_, _06146_);
  and _84895_ (_34974_, _14950_, _08413_);
  or _84896_ (_34976_, _34974_, _34944_);
  and _84897_ (_34977_, _34976_, _06145_);
  or _84898_ (_34978_, _34977_, _34973_);
  and _84899_ (_34979_, _34978_, _06140_);
  and _84900_ (_34980_, _14966_, _08413_);
  or _84901_ (_34981_, _34980_, _34944_);
  and _84902_ (_34982_, _34981_, _06139_);
  or _84903_ (_34983_, _34982_, _09842_);
  or _84904_ (_34984_, _34983_, _34979_);
  and _84905_ (_34985_, _34984_, _34943_);
  or _84906_ (_34987_, _34985_, _06116_);
  and _84907_ (_34988_, _09209_, _07778_);
  or _84908_ (_34989_, _34939_, _06117_);
  or _84909_ (_34990_, _34989_, _34988_);
  and _84910_ (_34991_, _34990_, _06114_);
  and _84911_ (_34992_, _34991_, _34987_);
  and _84912_ (_34993_, _15013_, _07778_);
  or _84913_ (_34994_, _34993_, _34939_);
  and _84914_ (_34995_, _34994_, _05787_);
  or _84915_ (_34996_, _34995_, _11136_);
  or _84916_ (_34998_, _34996_, _34992_);
  and _84917_ (_34999_, _15029_, _07778_);
  or _84918_ (_35000_, _34939_, _07127_);
  or _84919_ (_35001_, _35000_, _34999_);
  and _84920_ (_35002_, _08715_, _07778_);
  or _84921_ (_35003_, _35002_, _34939_);
  or _84922_ (_35004_, _35003_, _06111_);
  and _84923_ (_35005_, _35004_, _07125_);
  and _84924_ (_35006_, _35005_, _35001_);
  and _84925_ (_35007_, _35006_, _34998_);
  and _84926_ (_35009_, _10289_, _07778_);
  or _84927_ (_35010_, _35009_, _34939_);
  and _84928_ (_35011_, _35010_, _06402_);
  or _84929_ (_35012_, _35011_, _35007_);
  and _84930_ (_35013_, _35012_, _07132_);
  or _84931_ (_35014_, _34939_, _08339_);
  and _84932_ (_35015_, _35003_, _06306_);
  and _84933_ (_35016_, _35015_, _35014_);
  or _84934_ (_35017_, _35016_, _35013_);
  and _84935_ (_35018_, _35017_, _07130_);
  and _84936_ (_35020_, _34952_, _06411_);
  and _84937_ (_35021_, _35020_, _35014_);
  or _84938_ (_35022_, _35021_, _06303_);
  or _84939_ (_35023_, _35022_, _35018_);
  and _84940_ (_35024_, _15026_, _07778_);
  or _84941_ (_35025_, _34939_, _08819_);
  or _84942_ (_35026_, _35025_, _35024_);
  and _84943_ (_35027_, _35026_, _08824_);
  and _84944_ (_35028_, _35027_, _35023_);
  nor _84945_ (_35029_, _10288_, _13504_);
  or _84946_ (_35031_, _35029_, _34939_);
  and _84947_ (_35032_, _35031_, _06396_);
  or _84948_ (_35033_, _35032_, _06433_);
  or _84949_ (_35034_, _35033_, _35028_);
  or _84950_ (_35035_, _34949_, _06829_);
  and _84951_ (_35036_, _35035_, _05749_);
  and _84952_ (_35037_, _35036_, _35034_);
  and _84953_ (_35038_, _34946_, _05748_);
  or _84954_ (_35039_, _35038_, _06440_);
  or _84955_ (_35040_, _35039_, _35037_);
  and _84956_ (_35042_, _15087_, _07778_);
  or _84957_ (_35043_, _34939_, _06444_);
  or _84958_ (_35044_, _35043_, _35042_);
  and _84959_ (_35045_, _35044_, _01317_);
  and _84960_ (_35046_, _35045_, _35040_);
  or _84961_ (_35047_, _35046_, _34938_);
  and _84962_ (_43759_, _35047_, _43100_);
  and _84963_ (_35048_, _01321_, \oc8051_golden_model_1.SCON [5]);
  and _84964_ (_35049_, _13504_, \oc8051_golden_model_1.SCON [5]);
  and _84965_ (_35050_, _15119_, _07778_);
  or _84966_ (_35052_, _35050_, _35049_);
  or _84967_ (_35053_, _35052_, _06161_);
  and _84968_ (_35054_, _07778_, \oc8051_golden_model_1.ACC [5]);
  or _84969_ (_35055_, _35054_, _35049_);
  and _84970_ (_35056_, _35055_, _07056_);
  and _84971_ (_35057_, _07057_, \oc8051_golden_model_1.SCON [5]);
  or _84972_ (_35058_, _35057_, _06160_);
  or _84973_ (_35059_, _35058_, _35056_);
  and _84974_ (_35060_, _35059_, _06157_);
  and _84975_ (_35061_, _35060_, _35053_);
  and _84976_ (_35063_, _13509_, \oc8051_golden_model_1.SCON [5]);
  and _84977_ (_35064_, _15123_, _08413_);
  or _84978_ (_35065_, _35064_, _35063_);
  and _84979_ (_35066_, _35065_, _06156_);
  or _84980_ (_35067_, _35066_, _06217_);
  or _84981_ (_35068_, _35067_, _35061_);
  and _84982_ (_35069_, _08101_, _07778_);
  or _84983_ (_35070_, _35069_, _35049_);
  or _84984_ (_35071_, _35070_, _07075_);
  and _84985_ (_35072_, _35071_, _35068_);
  or _84986_ (_35074_, _35072_, _06220_);
  or _84987_ (_35075_, _35055_, _06229_);
  and _84988_ (_35076_, _35075_, _06153_);
  and _84989_ (_35077_, _35076_, _35074_);
  and _84990_ (_35078_, _15104_, _08413_);
  or _84991_ (_35079_, _35078_, _35063_);
  and _84992_ (_35080_, _35079_, _06152_);
  or _84993_ (_35081_, _35080_, _06145_);
  or _84994_ (_35082_, _35081_, _35077_);
  or _84995_ (_35083_, _35063_, _15138_);
  and _84996_ (_35085_, _35083_, _35065_);
  or _84997_ (_35086_, _35085_, _06146_);
  and _84998_ (_35087_, _35086_, _06140_);
  and _84999_ (_35088_, _35087_, _35082_);
  and _85000_ (_35089_, _15155_, _08413_);
  or _85001_ (_35090_, _35089_, _35063_);
  and _85002_ (_35091_, _35090_, _06139_);
  or _85003_ (_35092_, _35091_, _09842_);
  or _85004_ (_35093_, _35092_, _35088_);
  or _85005_ (_35094_, _35070_, _06132_);
  and _85006_ (_35096_, _35094_, _35093_);
  or _85007_ (_35097_, _35096_, _06116_);
  and _85008_ (_35098_, _09208_, _07778_);
  or _85009_ (_35099_, _35049_, _06117_);
  or _85010_ (_35100_, _35099_, _35098_);
  and _85011_ (_35101_, _35100_, _06114_);
  and _85012_ (_35102_, _35101_, _35097_);
  and _85013_ (_35103_, _15203_, _07778_);
  or _85014_ (_35104_, _35103_, _35049_);
  and _85015_ (_35105_, _35104_, _05787_);
  or _85016_ (_35107_, _35105_, _11136_);
  or _85017_ (_35108_, _35107_, _35102_);
  and _85018_ (_35109_, _15219_, _07778_);
  or _85019_ (_35110_, _35049_, _07127_);
  or _85020_ (_35111_, _35110_, _35109_);
  and _85021_ (_35112_, _08736_, _07778_);
  or _85022_ (_35113_, _35112_, _35049_);
  or _85023_ (_35114_, _35113_, _06111_);
  and _85024_ (_35115_, _35114_, _07125_);
  and _85025_ (_35116_, _35115_, _35111_);
  and _85026_ (_35118_, _35116_, _35108_);
  and _85027_ (_35119_, _12325_, _07778_);
  or _85028_ (_35120_, _35119_, _35049_);
  and _85029_ (_35121_, _35120_, _06402_);
  or _85030_ (_35122_, _35121_, _35118_);
  and _85031_ (_35123_, _35122_, _07132_);
  or _85032_ (_35124_, _35049_, _08104_);
  and _85033_ (_35125_, _35113_, _06306_);
  and _85034_ (_35126_, _35125_, _35124_);
  or _85035_ (_35127_, _35126_, _35123_);
  and _85036_ (_35129_, _35127_, _07130_);
  and _85037_ (_35130_, _35055_, _06411_);
  and _85038_ (_35131_, _35130_, _35124_);
  or _85039_ (_35132_, _35131_, _06303_);
  or _85040_ (_35133_, _35132_, _35129_);
  and _85041_ (_35134_, _15216_, _07778_);
  or _85042_ (_35135_, _35049_, _08819_);
  or _85043_ (_35136_, _35135_, _35134_);
  and _85044_ (_35137_, _35136_, _08824_);
  and _85045_ (_35138_, _35137_, _35133_);
  nor _85046_ (_35140_, _10269_, _13504_);
  or _85047_ (_35141_, _35140_, _35049_);
  and _85048_ (_35142_, _35141_, _06396_);
  or _85049_ (_35143_, _35142_, _06433_);
  or _85050_ (_35144_, _35143_, _35138_);
  or _85051_ (_35145_, _35052_, _06829_);
  and _85052_ (_35146_, _35145_, _05749_);
  and _85053_ (_35147_, _35146_, _35144_);
  and _85054_ (_35148_, _35079_, _05748_);
  or _85055_ (_35149_, _35148_, _06440_);
  or _85056_ (_35151_, _35149_, _35147_);
  and _85057_ (_35152_, _15275_, _07778_);
  or _85058_ (_35153_, _35049_, _06444_);
  or _85059_ (_35154_, _35153_, _35152_);
  and _85060_ (_35155_, _35154_, _01317_);
  and _85061_ (_35156_, _35155_, _35151_);
  or _85062_ (_35157_, _35156_, _35048_);
  and _85063_ (_43761_, _35157_, _43100_);
  and _85064_ (_35158_, _01321_, \oc8051_golden_model_1.SCON [6]);
  and _85065_ (_35159_, _13504_, \oc8051_golden_model_1.SCON [6]);
  and _85066_ (_35161_, _15300_, _07778_);
  or _85067_ (_35162_, _35161_, _35159_);
  or _85068_ (_35163_, _35162_, _06161_);
  and _85069_ (_35164_, _07778_, \oc8051_golden_model_1.ACC [6]);
  or _85070_ (_35165_, _35164_, _35159_);
  and _85071_ (_35166_, _35165_, _07056_);
  and _85072_ (_35167_, _07057_, \oc8051_golden_model_1.SCON [6]);
  or _85073_ (_35168_, _35167_, _06160_);
  or _85074_ (_35169_, _35168_, _35166_);
  and _85075_ (_35170_, _35169_, _06157_);
  and _85076_ (_35172_, _35170_, _35163_);
  and _85077_ (_35173_, _13509_, \oc8051_golden_model_1.SCON [6]);
  and _85078_ (_35174_, _15316_, _08413_);
  or _85079_ (_35175_, _35174_, _35173_);
  and _85080_ (_35176_, _35175_, _06156_);
  or _85081_ (_35177_, _35176_, _06217_);
  or _85082_ (_35178_, _35177_, _35172_);
  and _85083_ (_35179_, _08012_, _07778_);
  or _85084_ (_35180_, _35179_, _35159_);
  or _85085_ (_35181_, _35180_, _07075_);
  and _85086_ (_35183_, _35181_, _35178_);
  or _85087_ (_35184_, _35183_, _06220_);
  or _85088_ (_35185_, _35165_, _06229_);
  and _85089_ (_35186_, _35185_, _06153_);
  and _85090_ (_35187_, _35186_, _35184_);
  and _85091_ (_35188_, _15297_, _08413_);
  or _85092_ (_35189_, _35188_, _35173_);
  and _85093_ (_35190_, _35189_, _06152_);
  or _85094_ (_35191_, _35190_, _06145_);
  or _85095_ (_35192_, _35191_, _35187_);
  or _85096_ (_35194_, _35173_, _15331_);
  and _85097_ (_35195_, _35194_, _35175_);
  or _85098_ (_35196_, _35195_, _06146_);
  and _85099_ (_35197_, _35196_, _06140_);
  and _85100_ (_35198_, _35197_, _35192_);
  and _85101_ (_35199_, _15348_, _08413_);
  or _85102_ (_35200_, _35199_, _35173_);
  and _85103_ (_35201_, _35200_, _06139_);
  or _85104_ (_35202_, _35201_, _09842_);
  or _85105_ (_35203_, _35202_, _35198_);
  or _85106_ (_35205_, _35180_, _06132_);
  and _85107_ (_35206_, _35205_, _35203_);
  or _85108_ (_35207_, _35206_, _06116_);
  and _85109_ (_35208_, _09207_, _07778_);
  or _85110_ (_35209_, _35159_, _06117_);
  or _85111_ (_35210_, _35209_, _35208_);
  and _85112_ (_35211_, _35210_, _06114_);
  and _85113_ (_35212_, _35211_, _35207_);
  and _85114_ (_35213_, _15395_, _07778_);
  or _85115_ (_35214_, _35213_, _35159_);
  and _85116_ (_35216_, _35214_, _05787_);
  or _85117_ (_35217_, _35216_, _11136_);
  or _85118_ (_35218_, _35217_, _35212_);
  and _85119_ (_35219_, _15413_, _07778_);
  or _85120_ (_35220_, _35159_, _07127_);
  or _85121_ (_35221_, _35220_, _35219_);
  and _85122_ (_35222_, _15402_, _07778_);
  or _85123_ (_35223_, _35222_, _35159_);
  or _85124_ (_35224_, _35223_, _06111_);
  and _85125_ (_35225_, _35224_, _07125_);
  and _85126_ (_35227_, _35225_, _35221_);
  and _85127_ (_35228_, _35227_, _35218_);
  and _85128_ (_35229_, _10295_, _07778_);
  or _85129_ (_35230_, _35229_, _35159_);
  and _85130_ (_35231_, _35230_, _06402_);
  or _85131_ (_35232_, _35231_, _35228_);
  and _85132_ (_35233_, _35232_, _07132_);
  or _85133_ (_35234_, _35159_, _08015_);
  and _85134_ (_35235_, _35223_, _06306_);
  and _85135_ (_35236_, _35235_, _35234_);
  or _85136_ (_35238_, _35236_, _35233_);
  and _85137_ (_35239_, _35238_, _07130_);
  and _85138_ (_35240_, _35165_, _06411_);
  and _85139_ (_35241_, _35240_, _35234_);
  or _85140_ (_35242_, _35241_, _06303_);
  or _85141_ (_35243_, _35242_, _35239_);
  and _85142_ (_35244_, _15410_, _07778_);
  or _85143_ (_35245_, _35159_, _08819_);
  or _85144_ (_35246_, _35245_, _35244_);
  and _85145_ (_35247_, _35246_, _08824_);
  and _85146_ (_35249_, _35247_, _35243_);
  nor _85147_ (_35250_, _10294_, _13504_);
  or _85148_ (_35251_, _35250_, _35159_);
  and _85149_ (_35252_, _35251_, _06396_);
  or _85150_ (_35253_, _35252_, _06433_);
  or _85151_ (_35254_, _35253_, _35249_);
  or _85152_ (_35255_, _35162_, _06829_);
  and _85153_ (_35256_, _35255_, _05749_);
  and _85154_ (_35257_, _35256_, _35254_);
  and _85155_ (_35258_, _35189_, _05748_);
  or _85156_ (_35260_, _35258_, _06440_);
  or _85157_ (_35261_, _35260_, _35257_);
  and _85158_ (_35262_, _15478_, _07778_);
  or _85159_ (_35263_, _35159_, _06444_);
  or _85160_ (_35264_, _35263_, _35262_);
  and _85161_ (_35265_, _35264_, _01317_);
  and _85162_ (_35266_, _35265_, _35261_);
  or _85163_ (_35267_, _35266_, _35158_);
  and _85164_ (_43762_, _35267_, _43100_);
  nor _85165_ (_35268_, _01317_, _06142_);
  nor _85166_ (_35270_, _13615_, _06142_);
  and _85167_ (_35271_, _13615_, \oc8051_golden_model_1.ACC [0]);
  and _85168_ (_35272_, _35271_, _08211_);
  or _85169_ (_35273_, _35272_, _35270_);
  or _85170_ (_35274_, _35273_, _07130_);
  nor _85171_ (_35275_, _08211_, _13718_);
  or _85172_ (_35276_, _35275_, _35270_);
  or _85173_ (_35277_, _35276_, _06161_);
  or _85174_ (_35278_, _35271_, _35270_);
  and _85175_ (_35279_, _35278_, _07056_);
  nor _85176_ (_35281_, _07056_, _06142_);
  or _85177_ (_35282_, _35281_, _06160_);
  or _85178_ (_35283_, _35282_, _35279_);
  and _85179_ (_35284_, _35283_, _07075_);
  and _85180_ (_35285_, _35284_, _35277_);
  or _85181_ (_35286_, _35285_, _06671_);
  or _85182_ (_35287_, _35278_, _06229_);
  and _85183_ (_35288_, _35287_, _07191_);
  and _85184_ (_35289_, _35288_, _35286_);
  nand _85185_ (_35290_, _06132_, _07093_);
  or _85186_ (_35292_, _35290_, _35289_);
  and _85187_ (_35293_, _07858_, _07049_);
  or _85188_ (_35294_, _35270_, _06132_);
  or _85189_ (_35295_, _35294_, _35293_);
  and _85190_ (_35296_, _35295_, _35292_);
  or _85191_ (_35297_, _35296_, _06116_);
  or _85192_ (_35298_, _35270_, _06117_);
  and _85193_ (_35299_, _09160_, _13615_);
  or _85194_ (_35300_, _35299_, _35298_);
  and _85195_ (_35301_, _35300_, _35297_);
  or _85196_ (_35303_, _35301_, _05787_);
  and _85197_ (_35304_, _14260_, _07858_);
  or _85198_ (_35305_, _35270_, _06114_);
  or _85199_ (_35306_, _35305_, _35304_);
  and _85200_ (_35307_, _35306_, _06111_);
  and _85201_ (_35308_, _35307_, _35303_);
  and _85202_ (_35309_, _13615_, _08708_);
  or _85203_ (_35310_, _35309_, _35270_);
  and _85204_ (_35311_, _35310_, _06110_);
  or _85205_ (_35312_, _35311_, _06297_);
  or _85206_ (_35314_, _35312_, _35308_);
  and _85207_ (_35315_, _14275_, _13615_);
  or _85208_ (_35316_, _35315_, _35270_);
  or _85209_ (_35317_, _35316_, _07127_);
  and _85210_ (_35318_, _35317_, _07125_);
  and _85211_ (_35319_, _35318_, _35314_);
  nor _85212_ (_35320_, _12321_, _13718_);
  or _85213_ (_35321_, _35320_, _35270_);
  nor _85214_ (_35322_, _35272_, _07125_);
  and _85215_ (_35323_, _35322_, _35321_);
  or _85216_ (_35325_, _35323_, _35319_);
  and _85217_ (_35326_, _35325_, _07132_);
  nand _85218_ (_35327_, _35310_, _06306_);
  nor _85219_ (_35328_, _35327_, _35275_);
  or _85220_ (_35329_, _35328_, _06411_);
  or _85221_ (_35330_, _35329_, _35326_);
  and _85222_ (_35331_, _35330_, _35274_);
  or _85223_ (_35332_, _35331_, _06303_);
  and _85224_ (_35333_, _14167_, _07858_);
  or _85225_ (_35334_, _35270_, _08819_);
  or _85226_ (_35336_, _35334_, _35333_);
  and _85227_ (_35337_, _35336_, _08824_);
  and _85228_ (_35338_, _35337_, _35332_);
  and _85229_ (_35339_, _35321_, _06396_);
  or _85230_ (_35340_, _35339_, _19287_);
  or _85231_ (_35341_, _35340_, _35338_);
  or _85232_ (_35342_, _35276_, _06630_);
  and _85233_ (_35343_, _35342_, _01317_);
  and _85234_ (_35344_, _35343_, _35341_);
  or _85235_ (_35345_, _35344_, _35268_);
  and _85236_ (_43763_, _35345_, _43100_);
  nand _85237_ (_35347_, _06417_, \oc8051_golden_model_1.SP [1]);
  nand _85238_ (_35348_, _07858_, _06945_);
  or _85239_ (_35349_, _35348_, _08176_);
  or _85240_ (_35350_, _13615_, \oc8051_golden_model_1.SP [1]);
  and _85241_ (_35351_, _35350_, _06303_);
  and _85242_ (_35352_, _35351_, _35349_);
  and _85243_ (_35353_, _35350_, _05787_);
  or _85244_ (_35354_, _14442_, _13718_);
  and _85245_ (_35355_, _35354_, _35353_);
  and _85246_ (_35357_, _14363_, _07858_);
  not _85247_ (_35358_, _35357_);
  and _85248_ (_35359_, _35358_, _35350_);
  or _85249_ (_35360_, _35359_, _06161_);
  nor _85250_ (_35361_, _13615_, _06979_);
  and _85251_ (_35362_, _13615_, \oc8051_golden_model_1.ACC [1]);
  or _85252_ (_35363_, _35362_, _35361_);
  or _85253_ (_35364_, _35363_, _07057_);
  or _85254_ (_35365_, _07056_, \oc8051_golden_model_1.SP [1]);
  and _85255_ (_35366_, _35365_, _06582_);
  and _85256_ (_35368_, _35366_, _35364_);
  and _85257_ (_35369_, _06581_, _06979_);
  or _85258_ (_35370_, _35369_, _06160_);
  or _85259_ (_35371_, _35370_, _35368_);
  and _85260_ (_35372_, _35371_, _05764_);
  and _85261_ (_35373_, _35372_, _35360_);
  nor _85262_ (_35374_, _05764_, \oc8051_golden_model_1.SP [1]);
  or _85263_ (_35375_, _35374_, _06217_);
  or _85264_ (_35376_, _35375_, _35373_);
  nand _85265_ (_35377_, _07189_, _06217_);
  and _85266_ (_35379_, _35377_, _35376_);
  or _85267_ (_35380_, _35379_, _06220_);
  or _85268_ (_35381_, _35363_, _06229_);
  and _85269_ (_35382_, _35381_, _07191_);
  and _85270_ (_35383_, _35382_, _35380_);
  not _85271_ (_35384_, _07389_);
  or _85272_ (_35385_, _35384_, _07190_);
  or _85273_ (_35386_, _35385_, _35383_);
  or _85274_ (_35387_, _07389_, _06979_);
  and _85275_ (_35388_, _35387_, _06132_);
  and _85276_ (_35390_, _35388_, _35386_);
  or _85277_ (_35391_, _13718_, _07306_);
  and _85278_ (_35392_, _35350_, _09842_);
  and _85279_ (_35393_, _35392_, _35391_);
  or _85280_ (_35394_, _35393_, _06116_);
  or _85281_ (_35395_, _35394_, _35390_);
  or _85282_ (_35396_, _35361_, _06117_);
  and _85283_ (_35397_, _09115_, _13615_);
  or _85284_ (_35398_, _35397_, _35396_);
  and _85285_ (_35399_, _35398_, _06114_);
  and _85286_ (_35401_, _35399_, _35395_);
  or _85287_ (_35402_, _35401_, _35355_);
  and _85288_ (_35403_, _35402_, _06111_);
  and _85289_ (_35404_, _35350_, _06110_);
  and _85290_ (_35405_, _35404_, _35348_);
  or _85291_ (_35406_, _35405_, _06076_);
  or _85292_ (_35407_, _35406_, _35403_);
  or _85293_ (_35408_, _05836_, _06979_);
  and _85294_ (_35409_, _35408_, _07127_);
  and _85295_ (_35410_, _35409_, _35407_);
  or _85296_ (_35412_, _14346_, _13718_);
  and _85297_ (_35413_, _35350_, _06297_);
  and _85298_ (_35414_, _35413_, _35412_);
  or _85299_ (_35415_, _35414_, _06402_);
  or _85300_ (_35416_, _35415_, _35410_);
  and _85301_ (_35417_, _10278_, _13615_);
  or _85302_ (_35418_, _35417_, _35361_);
  or _85303_ (_35419_, _35418_, _07125_);
  and _85304_ (_35420_, _35419_, _07132_);
  and _85305_ (_35421_, _35420_, _35416_);
  or _85306_ (_35423_, _14344_, _13718_);
  and _85307_ (_35424_, _35350_, _06306_);
  and _85308_ (_35425_, _35424_, _35423_);
  or _85309_ (_35426_, _35425_, _06411_);
  or _85310_ (_35427_, _35426_, _35421_);
  and _85311_ (_35428_, _35362_, _08176_);
  or _85312_ (_35429_, _35428_, _35361_);
  or _85313_ (_35430_, _35429_, _07130_);
  and _85314_ (_35431_, _35430_, _35427_);
  or _85315_ (_35432_, _35431_, _07124_);
  nor _85316_ (_35434_, _05848_, _06979_);
  nor _85317_ (_35435_, _35434_, _06303_);
  and _85318_ (_35436_, _35435_, _35432_);
  or _85319_ (_35437_, _35436_, _35352_);
  and _85320_ (_35438_, _35437_, _08824_);
  nor _85321_ (_35439_, _10277_, _13718_);
  or _85322_ (_35440_, _35439_, _35361_);
  and _85323_ (_35441_, _35440_, _06396_);
  or _85324_ (_35442_, _35441_, _06417_);
  or _85325_ (_35443_, _35442_, _35438_);
  nand _85326_ (_35445_, _35443_, _35347_);
  nor _85327_ (_35446_, _06167_, _07142_);
  nand _85328_ (_35447_, _35446_, _35445_);
  or _85329_ (_35448_, _35446_, _06979_);
  and _85330_ (_35449_, _35448_, _06829_);
  and _85331_ (_35450_, _35449_, _35447_);
  and _85332_ (_35451_, _35359_, _06433_);
  or _85333_ (_35452_, _35451_, _07577_);
  or _85334_ (_35453_, _35452_, _35450_);
  or _85335_ (_35454_, _07160_, _06979_);
  and _85336_ (_35456_, _35454_, _06444_);
  and _85337_ (_35457_, _35456_, _35453_);
  or _85338_ (_35458_, _35357_, _35361_);
  and _85339_ (_35459_, _35458_, _06440_);
  or _85340_ (_35460_, _35459_, _01321_);
  or _85341_ (_35461_, _35460_, _35457_);
  or _85342_ (_35462_, _01317_, \oc8051_golden_model_1.SP [1]);
  and _85343_ (_35463_, _35462_, _43100_);
  and _85344_ (_43765_, _35463_, _35461_);
  nor _85345_ (_35464_, _01317_, _06566_);
  or _85346_ (_35466_, _07755_, _05836_);
  and _85347_ (_35467_, _07858_, _07708_);
  nor _85348_ (_35468_, _13615_, _06566_);
  or _85349_ (_35469_, _35468_, _06132_);
  or _85350_ (_35470_, _35469_, _35467_);
  and _85351_ (_35471_, _14542_, _07858_);
  or _85352_ (_35472_, _35471_, _35468_);
  or _85353_ (_35473_, _35472_, _06161_);
  and _85354_ (_35474_, _13615_, \oc8051_golden_model_1.ACC [2]);
  or _85355_ (_35475_, _35474_, _35468_);
  or _85356_ (_35477_, _35475_, _07057_);
  or _85357_ (_35478_, _07056_, \oc8051_golden_model_1.SP [2]);
  and _85358_ (_35479_, _35478_, _06582_);
  and _85359_ (_35480_, _35479_, _35477_);
  and _85360_ (_35481_, _07755_, _06581_);
  or _85361_ (_35482_, _35481_, _06160_);
  or _85362_ (_35483_, _35482_, _35480_);
  and _85363_ (_35484_, _35483_, _05764_);
  and _85364_ (_35485_, _35484_, _35473_);
  nor _85365_ (_35486_, _15819_, _05764_);
  or _85366_ (_35488_, _35486_, _06217_);
  or _85367_ (_35489_, _35488_, _35485_);
  nand _85368_ (_35490_, _08465_, _06217_);
  and _85369_ (_35491_, _35490_, _35489_);
  or _85370_ (_35492_, _35491_, _06220_);
  or _85371_ (_35493_, _35475_, _06229_);
  and _85372_ (_35494_, _35493_, _07191_);
  and _85373_ (_35495_, _35494_, _35492_);
  or _85374_ (_35496_, _07601_, _07388_);
  or _85375_ (_35497_, _35496_, _35495_);
  nor _85376_ (_35499_, _07755_, _05760_);
  nor _85377_ (_35500_, _35499_, _05791_);
  and _85378_ (_35501_, _35500_, _35497_);
  nand _85379_ (_35502_, _07755_, _05791_);
  nand _85380_ (_35503_, _35502_, _06132_);
  or _85381_ (_35504_, _35503_, _35501_);
  and _85382_ (_35505_, _35504_, _35470_);
  or _85383_ (_35506_, _35505_, _06116_);
  or _85384_ (_35507_, _35468_, _06117_);
  and _85385_ (_35508_, _09211_, _13615_);
  or _85386_ (_35510_, _35508_, _35507_);
  and _85387_ (_35511_, _35510_, _06114_);
  and _85388_ (_35512_, _35511_, _35506_);
  and _85389_ (_35513_, _14630_, _13615_);
  or _85390_ (_35514_, _35513_, _35468_);
  and _85391_ (_35515_, _35514_, _05787_);
  or _85392_ (_35516_, _35515_, _06110_);
  or _85393_ (_35517_, _35516_, _35512_);
  and _85394_ (_35518_, _13615_, _08768_);
  or _85395_ (_35519_, _35518_, _35468_);
  or _85396_ (_35521_, _35519_, _06111_);
  and _85397_ (_35522_, _35521_, _35517_);
  or _85398_ (_35523_, _35522_, _06076_);
  and _85399_ (_35524_, _35523_, _35466_);
  or _85400_ (_35525_, _35524_, _06297_);
  and _85401_ (_35526_, _14646_, _13615_);
  or _85402_ (_35527_, _35526_, _35468_);
  or _85403_ (_35528_, _35527_, _07127_);
  and _85404_ (_35529_, _35528_, _07125_);
  and _85405_ (_35530_, _35529_, _35525_);
  and _85406_ (_35532_, _10282_, _13615_);
  or _85407_ (_35533_, _35532_, _35468_);
  and _85408_ (_35534_, _35533_, _06402_);
  or _85409_ (_35535_, _35534_, _35530_);
  and _85410_ (_35536_, _35535_, _07132_);
  or _85411_ (_35537_, _35468_, _08248_);
  and _85412_ (_35538_, _35519_, _06306_);
  and _85413_ (_35539_, _35538_, _35537_);
  or _85414_ (_35540_, _35539_, _35536_);
  and _85415_ (_35541_, _35540_, _12514_);
  and _85416_ (_35543_, _35475_, _06411_);
  and _85417_ (_35544_, _35543_, _35537_);
  nor _85418_ (_35545_, _15819_, _05848_);
  or _85419_ (_35546_, _35545_, _06303_);
  or _85420_ (_35547_, _35546_, _35544_);
  or _85421_ (_35548_, _35547_, _35541_);
  and _85422_ (_35549_, _14643_, _07858_);
  or _85423_ (_35550_, _35468_, _08819_);
  or _85424_ (_35551_, _35550_, _35549_);
  and _85425_ (_35552_, _35551_, _35548_);
  or _85426_ (_35554_, _35552_, _06396_);
  nor _85427_ (_35555_, _10281_, _13718_);
  or _85428_ (_35556_, _35555_, _35468_);
  or _85429_ (_35557_, _35556_, _08824_);
  and _85430_ (_35558_, _35557_, _12558_);
  and _85431_ (_35559_, _35558_, _35554_);
  and _85432_ (_35560_, _15819_, _06417_);
  or _85433_ (_35561_, _35560_, _07142_);
  or _85434_ (_35562_, _35561_, _35559_);
  or _85435_ (_35563_, _07755_, _05846_);
  and _85436_ (_35565_, _35563_, _06168_);
  and _85437_ (_35566_, _35565_, _35562_);
  and _85438_ (_35567_, _15819_, _06167_);
  or _85439_ (_35568_, _35567_, _06433_);
  or _85440_ (_35569_, _35568_, _35566_);
  or _85441_ (_35570_, _35472_, _06829_);
  and _85442_ (_35571_, _35570_, _07160_);
  and _85443_ (_35572_, _35571_, _35569_);
  nor _85444_ (_35573_, _15819_, _07160_);
  or _85445_ (_35574_, _35573_, _06440_);
  or _85446_ (_35576_, _35574_, _35572_);
  and _85447_ (_35577_, _14710_, _07858_);
  or _85448_ (_35578_, _35468_, _06444_);
  or _85449_ (_35579_, _35578_, _35577_);
  and _85450_ (_35580_, _35579_, _01317_);
  and _85451_ (_35581_, _35580_, _35576_);
  or _85452_ (_35582_, _35581_, _35464_);
  and _85453_ (_43766_, _35582_, _43100_);
  nor _85454_ (_35583_, _01317_, _06216_);
  or _85455_ (_35584_, _07759_, _07160_);
  or _85456_ (_35586_, _07759_, _05836_);
  and _85457_ (_35587_, _07858_, _07544_);
  nor _85458_ (_35588_, _13615_, _06216_);
  or _85459_ (_35589_, _35588_, _06116_);
  or _85460_ (_35590_, _35589_, _35587_);
  and _85461_ (_35591_, _35590_, _13620_);
  and _85462_ (_35592_, _14738_, _07858_);
  or _85463_ (_35593_, _35592_, _35588_);
  or _85464_ (_35594_, _35593_, _06161_);
  and _85465_ (_35595_, _13615_, \oc8051_golden_model_1.ACC [3]);
  or _85466_ (_35597_, _35595_, _35588_);
  or _85467_ (_35598_, _35597_, _07057_);
  or _85468_ (_35599_, _07056_, \oc8051_golden_model_1.SP [3]);
  and _85469_ (_35600_, _35599_, _06582_);
  and _85470_ (_35601_, _35600_, _35598_);
  and _85471_ (_35602_, _07759_, _06581_);
  or _85472_ (_35603_, _35602_, _06160_);
  or _85473_ (_35604_, _35603_, _35601_);
  and _85474_ (_35605_, _35604_, _05764_);
  and _85475_ (_35606_, _35605_, _35594_);
  nor _85476_ (_35608_, _15639_, _05764_);
  or _85477_ (_35609_, _35608_, _06217_);
  or _85478_ (_35610_, _35609_, _35606_);
  nand _85479_ (_35611_, _08455_, _06217_);
  and _85480_ (_35612_, _35611_, _35610_);
  or _85481_ (_35613_, _35612_, _06220_);
  or _85482_ (_35614_, _35597_, _06229_);
  and _85483_ (_35615_, _35614_, _07191_);
  and _85484_ (_35616_, _35615_, _35613_);
  or _85485_ (_35617_, _07525_, _35384_);
  or _85486_ (_35619_, _35617_, _35616_);
  or _85487_ (_35620_, _07759_, _07389_);
  and _85488_ (_35621_, _35620_, _06132_);
  and _85489_ (_35622_, _35621_, _35619_);
  or _85490_ (_35623_, _35622_, _35591_);
  or _85491_ (_35624_, _35588_, _06117_);
  and _85492_ (_35625_, _09210_, _13615_);
  or _85493_ (_35626_, _35625_, _35624_);
  and _85494_ (_35627_, _35626_, _06114_);
  and _85495_ (_35628_, _35627_, _35623_);
  and _85496_ (_35630_, _14825_, _13615_);
  or _85497_ (_35631_, _35630_, _35588_);
  and _85498_ (_35632_, _35631_, _05787_);
  or _85499_ (_35633_, _35632_, _06110_);
  or _85500_ (_35634_, _35633_, _35628_);
  and _85501_ (_35635_, _13615_, _08712_);
  or _85502_ (_35636_, _35635_, _35588_);
  or _85503_ (_35637_, _35636_, _06111_);
  and _85504_ (_35638_, _35637_, _35634_);
  or _85505_ (_35639_, _35638_, _06076_);
  and _85506_ (_35641_, _35639_, _35586_);
  or _85507_ (_35642_, _35641_, _06297_);
  and _85508_ (_35643_, _14727_, _13615_);
  or _85509_ (_35644_, _35643_, _35588_);
  or _85510_ (_35645_, _35644_, _07127_);
  and _85511_ (_35646_, _35645_, _07125_);
  and _85512_ (_35647_, _35646_, _35642_);
  and _85513_ (_35648_, _12318_, _13615_);
  or _85514_ (_35649_, _35648_, _35588_);
  and _85515_ (_35650_, _35649_, _06402_);
  or _85516_ (_35652_, _35650_, _35647_);
  and _85517_ (_35653_, _35652_, _07132_);
  or _85518_ (_35654_, _35588_, _08140_);
  and _85519_ (_35655_, _35636_, _06306_);
  and _85520_ (_35656_, _35655_, _35654_);
  or _85521_ (_35657_, _35656_, _35653_);
  and _85522_ (_35658_, _35657_, _12514_);
  and _85523_ (_35659_, _35597_, _06411_);
  and _85524_ (_35660_, _35659_, _35654_);
  nor _85525_ (_35661_, _15639_, _05848_);
  or _85526_ (_35663_, _35661_, _06303_);
  or _85527_ (_35664_, _35663_, _35660_);
  or _85528_ (_35665_, _35664_, _35658_);
  and _85529_ (_35666_, _14724_, _07858_);
  or _85530_ (_35667_, _35588_, _08819_);
  or _85531_ (_35668_, _35667_, _35666_);
  and _85532_ (_35669_, _35668_, _35665_);
  or _85533_ (_35670_, _35669_, _06396_);
  nor _85534_ (_35671_, _10273_, _13718_);
  or _85535_ (_35672_, _35671_, _35588_);
  or _85536_ (_35674_, _35672_, _08824_);
  and _85537_ (_35675_, _35674_, _12558_);
  and _85538_ (_35676_, _35675_, _35670_);
  nor _85539_ (_35677_, _08452_, _06216_);
  or _85540_ (_35678_, _35677_, _08453_);
  and _85541_ (_35679_, _35678_, _06417_);
  or _85542_ (_35680_, _35679_, _07142_);
  or _85543_ (_35681_, _35680_, _35676_);
  or _85544_ (_35682_, _07759_, _05846_);
  and _85545_ (_35683_, _35682_, _35681_);
  or _85546_ (_35685_, _35683_, _06167_);
  or _85547_ (_35686_, _35678_, _06168_);
  and _85548_ (_35687_, _35686_, _06829_);
  and _85549_ (_35688_, _35687_, _35685_);
  and _85550_ (_35689_, _35593_, _06433_);
  or _85551_ (_35690_, _35689_, _07577_);
  or _85552_ (_35691_, _35690_, _35688_);
  and _85553_ (_35692_, _35691_, _35584_);
  or _85554_ (_35693_, _35692_, _06440_);
  and _85555_ (_35694_, _14897_, _07858_);
  or _85556_ (_35695_, _35588_, _06444_);
  or _85557_ (_35696_, _35695_, _35694_);
  and _85558_ (_35697_, _35696_, _01317_);
  and _85559_ (_35698_, _35697_, _35693_);
  or _85560_ (_35699_, _35698_, _35583_);
  and _85561_ (_43767_, _35699_, _43100_);
  nor _85562_ (_35700_, _01317_, _13644_);
  nor _85563_ (_35701_, _07756_, \oc8051_golden_model_1.SP [4]);
  nor _85564_ (_35702_, _35701_, _13607_);
  or _85565_ (_35703_, _35702_, _07160_);
  or _85566_ (_35705_, _35702_, _05846_);
  and _85567_ (_35706_, _08336_, _07858_);
  nor _85568_ (_35707_, _13615_, _13644_);
  or _85569_ (_35708_, _35707_, _06116_);
  or _85570_ (_35709_, _35708_, _35706_);
  and _85571_ (_35710_, _35709_, _13620_);
  and _85572_ (_35711_, _14928_, _07858_);
  or _85573_ (_35712_, _35711_, _35707_);
  or _85574_ (_35713_, _35712_, _06161_);
  and _85575_ (_35714_, _13615_, \oc8051_golden_model_1.ACC [4]);
  or _85576_ (_35716_, _35714_, _35707_);
  or _85577_ (_35717_, _35716_, _07057_);
  or _85578_ (_35718_, _07056_, \oc8051_golden_model_1.SP [4]);
  and _85579_ (_35719_, _35718_, _06582_);
  and _85580_ (_35720_, _35719_, _35717_);
  and _85581_ (_35721_, _35702_, _06581_);
  or _85582_ (_35722_, _35721_, _06160_);
  or _85583_ (_35723_, _35722_, _35720_);
  and _85584_ (_35724_, _35723_, _05764_);
  and _85585_ (_35725_, _35724_, _35713_);
  and _85586_ (_35727_, _35702_, _07485_);
  or _85587_ (_35728_, _35727_, _06217_);
  or _85588_ (_35729_, _35728_, _35725_);
  and _85589_ (_35730_, _13645_, _06142_);
  nor _85590_ (_35731_, _08454_, _13644_);
  nor _85591_ (_35732_, _35731_, _35730_);
  nand _85592_ (_35733_, _35732_, _06217_);
  and _85593_ (_35734_, _35733_, _35729_);
  or _85594_ (_35735_, _35734_, _06220_);
  or _85595_ (_35736_, _35716_, _06229_);
  and _85596_ (_35738_, _35736_, _07191_);
  and _85597_ (_35739_, _35738_, _35735_);
  and _85598_ (_35740_, _07479_, \oc8051_golden_model_1.SP [4]);
  nor _85599_ (_35741_, _07479_, \oc8051_golden_model_1.SP [4]);
  nor _85600_ (_35742_, _35741_, _35740_);
  nand _85601_ (_35743_, _35742_, _06151_);
  nand _85602_ (_35744_, _35743_, _07389_);
  or _85603_ (_35745_, _35744_, _35739_);
  or _85604_ (_35746_, _35702_, _07389_);
  and _85605_ (_35747_, _35746_, _06132_);
  and _85606_ (_35749_, _35747_, _35745_);
  or _85607_ (_35750_, _35749_, _35710_);
  or _85608_ (_35751_, _35707_, _06117_);
  and _85609_ (_35752_, _09209_, _13615_);
  or _85610_ (_35753_, _35752_, _35751_);
  and _85611_ (_35754_, _35753_, _06114_);
  and _85612_ (_35755_, _35754_, _35750_);
  and _85613_ (_35756_, _15013_, _13615_);
  or _85614_ (_35757_, _35756_, _35707_);
  and _85615_ (_35758_, _35757_, _05787_);
  or _85616_ (_35760_, _35758_, _06110_);
  or _85617_ (_35761_, _35760_, _35755_);
  and _85618_ (_35762_, _08715_, _13615_);
  or _85619_ (_35763_, _35762_, _35707_);
  or _85620_ (_35764_, _35763_, _06111_);
  and _85621_ (_35765_, _35764_, _35761_);
  or _85622_ (_35766_, _35765_, _06076_);
  or _85623_ (_35767_, _35702_, _05836_);
  and _85624_ (_35768_, _35767_, _35766_);
  or _85625_ (_35769_, _35768_, _06297_);
  and _85626_ (_35771_, _15029_, _07858_);
  or _85627_ (_35772_, _35707_, _07127_);
  or _85628_ (_35773_, _35772_, _35771_);
  and _85629_ (_35774_, _35773_, _07125_);
  and _85630_ (_35775_, _35774_, _35769_);
  and _85631_ (_35776_, _10289_, _13615_);
  or _85632_ (_35777_, _35776_, _35707_);
  and _85633_ (_35778_, _35777_, _06402_);
  or _85634_ (_35779_, _35778_, _35775_);
  and _85635_ (_35780_, _35779_, _07132_);
  or _85636_ (_35782_, _35707_, _08339_);
  and _85637_ (_35783_, _35763_, _06306_);
  and _85638_ (_35784_, _35783_, _35782_);
  or _85639_ (_35785_, _35784_, _35780_);
  and _85640_ (_35786_, _35785_, _12514_);
  and _85641_ (_35787_, _35716_, _06411_);
  and _85642_ (_35788_, _35787_, _35782_);
  and _85643_ (_35789_, _35702_, _07124_);
  or _85644_ (_35790_, _35789_, _06303_);
  or _85645_ (_35791_, _35790_, _35788_);
  or _85646_ (_35793_, _35791_, _35786_);
  and _85647_ (_35794_, _15026_, _07858_);
  or _85648_ (_35795_, _35707_, _08819_);
  or _85649_ (_35796_, _35795_, _35794_);
  and _85650_ (_35797_, _35796_, _35793_);
  or _85651_ (_35798_, _35797_, _06396_);
  nor _85652_ (_35799_, _10288_, _13718_);
  or _85653_ (_35800_, _35799_, _35707_);
  or _85654_ (_35801_, _35800_, _08824_);
  and _85655_ (_35802_, _35801_, _12558_);
  and _85656_ (_35804_, _35802_, _35798_);
  nor _85657_ (_35805_, _08453_, _13644_);
  or _85658_ (_35806_, _35805_, _13645_);
  and _85659_ (_35807_, _35806_, _06417_);
  or _85660_ (_35808_, _35807_, _07142_);
  or _85661_ (_35809_, _35808_, _35804_);
  and _85662_ (_35810_, _35809_, _35705_);
  or _85663_ (_35811_, _35810_, _06167_);
  or _85664_ (_35812_, _35806_, _06168_);
  and _85665_ (_35813_, _35812_, _06829_);
  and _85666_ (_35815_, _35813_, _35811_);
  and _85667_ (_35816_, _35712_, _06433_);
  or _85668_ (_35817_, _35816_, _07577_);
  or _85669_ (_35818_, _35817_, _35815_);
  and _85670_ (_35819_, _35818_, _35703_);
  or _85671_ (_35820_, _35819_, _06440_);
  and _85672_ (_35821_, _15087_, _07858_);
  or _85673_ (_35822_, _35707_, _06444_);
  or _85674_ (_35823_, _35822_, _35821_);
  and _85675_ (_35824_, _35823_, _01317_);
  and _85676_ (_35826_, _35824_, _35820_);
  or _85677_ (_35827_, _35826_, _35700_);
  and _85678_ (_43768_, _35827_, _43100_);
  nor _85679_ (_35828_, _01317_, _13643_);
  nor _85680_ (_35829_, _13607_, \oc8051_golden_model_1.SP [5]);
  nor _85681_ (_35830_, _35829_, _13608_);
  or _85682_ (_35831_, _35830_, _07160_);
  and _85683_ (_35832_, _08101_, _07858_);
  nor _85684_ (_35833_, _13615_, _13643_);
  or _85685_ (_35834_, _35833_, _06116_);
  or _85686_ (_35836_, _35834_, _35832_);
  and _85687_ (_35837_, _35836_, _13620_);
  and _85688_ (_35838_, _15119_, _07858_);
  or _85689_ (_35839_, _35838_, _35833_);
  or _85690_ (_35840_, _35839_, _06161_);
  and _85691_ (_35841_, _13615_, \oc8051_golden_model_1.ACC [5]);
  or _85692_ (_35842_, _35841_, _35833_);
  or _85693_ (_35843_, _35842_, _07057_);
  or _85694_ (_35844_, _07056_, \oc8051_golden_model_1.SP [5]);
  and _85695_ (_35845_, _35844_, _06582_);
  and _85696_ (_35847_, _35845_, _35843_);
  and _85697_ (_35848_, _35830_, _06581_);
  or _85698_ (_35849_, _35848_, _06160_);
  or _85699_ (_35850_, _35849_, _35847_);
  and _85700_ (_35851_, _35850_, _05764_);
  and _85701_ (_35852_, _35851_, _35840_);
  and _85702_ (_35853_, _35830_, _07485_);
  or _85703_ (_35854_, _35853_, _06217_);
  or _85704_ (_35855_, _35854_, _35852_);
  and _85705_ (_35856_, _13646_, _06142_);
  nor _85706_ (_35858_, _35730_, _13643_);
  nor _85707_ (_35859_, _35858_, _35856_);
  nand _85708_ (_35860_, _35859_, _06217_);
  and _85709_ (_35861_, _35860_, _35855_);
  or _85710_ (_35862_, _35861_, _06220_);
  or _85711_ (_35863_, _35842_, _06229_);
  and _85712_ (_35864_, _35863_, _07191_);
  and _85713_ (_35865_, _35864_, _35862_);
  nor _85714_ (_35866_, _35740_, \oc8051_golden_model_1.SP [5]);
  nor _85715_ (_35867_, _35866_, _13659_);
  nand _85716_ (_35869_, _35867_, _06151_);
  nand _85717_ (_35870_, _35869_, _07389_);
  or _85718_ (_35871_, _35870_, _35865_);
  or _85719_ (_35872_, _35830_, _07389_);
  and _85720_ (_35873_, _35872_, _06132_);
  and _85721_ (_35874_, _35873_, _35871_);
  or _85722_ (_35875_, _35874_, _35837_);
  or _85723_ (_35876_, _35833_, _06117_);
  and _85724_ (_35877_, _09208_, _13615_);
  or _85725_ (_35878_, _35877_, _35876_);
  and _85726_ (_35880_, _35878_, _06114_);
  and _85727_ (_35881_, _35880_, _35875_);
  and _85728_ (_35882_, _15203_, _13615_);
  or _85729_ (_35883_, _35882_, _35833_);
  and _85730_ (_35884_, _35883_, _05787_);
  or _85731_ (_35885_, _35884_, _06110_);
  or _85732_ (_35886_, _35885_, _35881_);
  and _85733_ (_35887_, _08736_, _13615_);
  or _85734_ (_35888_, _35887_, _35833_);
  or _85735_ (_35889_, _35888_, _06111_);
  and _85736_ (_35891_, _35889_, _35886_);
  or _85737_ (_35892_, _35891_, _06076_);
  or _85738_ (_35893_, _35830_, _05836_);
  and _85739_ (_35894_, _35893_, _35892_);
  or _85740_ (_35895_, _35894_, _06297_);
  and _85741_ (_35896_, _15219_, _07858_);
  or _85742_ (_35897_, _35833_, _07127_);
  or _85743_ (_35898_, _35897_, _35896_);
  and _85744_ (_35899_, _35898_, _07125_);
  and _85745_ (_35900_, _35899_, _35895_);
  and _85746_ (_35902_, _12325_, _13615_);
  or _85747_ (_35903_, _35902_, _35833_);
  and _85748_ (_35904_, _35903_, _06402_);
  or _85749_ (_35905_, _35904_, _35900_);
  and _85750_ (_35906_, _35905_, _07132_);
  or _85751_ (_35907_, _35833_, _08104_);
  and _85752_ (_35908_, _35888_, _06306_);
  and _85753_ (_35909_, _35908_, _35907_);
  or _85754_ (_35910_, _35909_, _35906_);
  and _85755_ (_35911_, _35910_, _12514_);
  and _85756_ (_35913_, _35842_, _06411_);
  and _85757_ (_35914_, _35913_, _35907_);
  and _85758_ (_35915_, _35830_, _07124_);
  or _85759_ (_35916_, _35915_, _06303_);
  or _85760_ (_35917_, _35916_, _35914_);
  or _85761_ (_35918_, _35917_, _35911_);
  and _85762_ (_35919_, _15216_, _07858_);
  or _85763_ (_35920_, _35833_, _08819_);
  or _85764_ (_35921_, _35920_, _35919_);
  and _85765_ (_35922_, _35921_, _35918_);
  or _85766_ (_35924_, _35922_, _06396_);
  nor _85767_ (_35925_, _10269_, _13718_);
  or _85768_ (_35926_, _35925_, _35833_);
  or _85769_ (_35927_, _35926_, _08824_);
  and _85770_ (_35928_, _35927_, _12558_);
  and _85771_ (_35929_, _35928_, _35924_);
  nor _85772_ (_35930_, _13645_, _13643_);
  or _85773_ (_35931_, _35930_, _13646_);
  and _85774_ (_35932_, _35931_, _06417_);
  or _85775_ (_35933_, _35932_, _07142_);
  or _85776_ (_35935_, _35933_, _35929_);
  or _85777_ (_35936_, _35830_, _05846_);
  and _85778_ (_35937_, _35936_, _35935_);
  or _85779_ (_35938_, _35937_, _06167_);
  or _85780_ (_35939_, _35931_, _06168_);
  and _85781_ (_35940_, _35939_, _06829_);
  and _85782_ (_35941_, _35940_, _35938_);
  and _85783_ (_35942_, _35839_, _06433_);
  or _85784_ (_35943_, _35942_, _07577_);
  or _85785_ (_35944_, _35943_, _35941_);
  and _85786_ (_35946_, _35944_, _35831_);
  or _85787_ (_35947_, _35946_, _06440_);
  and _85788_ (_35948_, _15275_, _07858_);
  or _85789_ (_35949_, _35833_, _06444_);
  or _85790_ (_35950_, _35949_, _35948_);
  and _85791_ (_35951_, _35950_, _01317_);
  and _85792_ (_35952_, _35951_, _35947_);
  or _85793_ (_35953_, _35952_, _35828_);
  and _85794_ (_43769_, _35953_, _43100_);
  nor _85795_ (_35954_, _01317_, _13642_);
  nor _85796_ (_35956_, _13615_, _13642_);
  and _85797_ (_35957_, _15300_, _07858_);
  or _85798_ (_35958_, _35957_, _35956_);
  or _85799_ (_35959_, _35958_, _06161_);
  and _85800_ (_35960_, _13615_, \oc8051_golden_model_1.ACC [6]);
  or _85801_ (_35961_, _35960_, _35956_);
  or _85802_ (_35962_, _35961_, _07057_);
  or _85803_ (_35963_, _07056_, \oc8051_golden_model_1.SP [6]);
  and _85804_ (_35964_, _35963_, _06582_);
  and _85805_ (_35965_, _35964_, _35962_);
  nor _85806_ (_35967_, _13608_, \oc8051_golden_model_1.SP [6]);
  nor _85807_ (_35968_, _35967_, _13609_);
  and _85808_ (_35969_, _35968_, _06581_);
  or _85809_ (_35970_, _35969_, _06160_);
  or _85810_ (_35971_, _35970_, _35965_);
  and _85811_ (_35972_, _35971_, _05764_);
  and _85812_ (_35973_, _35972_, _35959_);
  and _85813_ (_35974_, _35968_, _07485_);
  or _85814_ (_35975_, _35974_, _06217_);
  or _85815_ (_35976_, _35975_, _35973_);
  nor _85816_ (_35978_, _35856_, _13642_);
  nor _85817_ (_35979_, _35978_, _13648_);
  nand _85818_ (_35980_, _35979_, _06217_);
  and _85819_ (_35981_, _35980_, _35976_);
  or _85820_ (_35982_, _35981_, _06220_);
  or _85821_ (_35983_, _35961_, _06229_);
  and _85822_ (_35984_, _35983_, _07191_);
  and _85823_ (_35985_, _35984_, _35982_);
  nor _85824_ (_35986_, _13659_, \oc8051_golden_model_1.SP [6]);
  nor _85825_ (_35987_, _35986_, _13661_);
  and _85826_ (_35989_, _35987_, _06151_);
  or _85827_ (_35990_, _35989_, _35985_);
  and _85828_ (_35991_, _35990_, _07389_);
  nand _85829_ (_35992_, _35968_, _35384_);
  nand _85830_ (_35993_, _35992_, _06132_);
  or _85831_ (_35994_, _35993_, _35991_);
  and _85832_ (_35995_, _08012_, _07858_);
  or _85833_ (_35996_, _35956_, _06132_);
  or _85834_ (_35997_, _35996_, _35995_);
  and _85835_ (_35998_, _35997_, _35994_);
  or _85836_ (_36000_, _35998_, _06116_);
  and _85837_ (_36001_, _09207_, _13615_);
  or _85838_ (_36002_, _35956_, _06117_);
  or _85839_ (_36003_, _36002_, _36001_);
  and _85840_ (_36004_, _36003_, _06114_);
  and _85841_ (_36005_, _36004_, _36000_);
  and _85842_ (_36006_, _15395_, _07858_);
  or _85843_ (_36007_, _36006_, _35956_);
  and _85844_ (_36008_, _36007_, _05787_);
  or _85845_ (_36009_, _36008_, _06110_);
  or _85846_ (_36011_, _36009_, _36005_);
  and _85847_ (_36012_, _15402_, _13615_);
  or _85848_ (_36013_, _36012_, _35956_);
  or _85849_ (_36014_, _36013_, _06111_);
  and _85850_ (_36015_, _36014_, _36011_);
  or _85851_ (_36016_, _36015_, _06076_);
  or _85852_ (_36017_, _35968_, _05836_);
  and _85853_ (_36018_, _36017_, _36016_);
  or _85854_ (_36019_, _36018_, _06297_);
  and _85855_ (_36020_, _15413_, _07858_);
  or _85856_ (_36022_, _35956_, _07127_);
  or _85857_ (_36023_, _36022_, _36020_);
  and _85858_ (_36024_, _36023_, _07125_);
  and _85859_ (_36025_, _36024_, _36019_);
  and _85860_ (_36026_, _10295_, _13615_);
  or _85861_ (_36027_, _36026_, _35956_);
  and _85862_ (_36028_, _36027_, _06402_);
  or _85863_ (_36029_, _36028_, _36025_);
  and _85864_ (_36030_, _36029_, _07132_);
  or _85865_ (_36031_, _35956_, _08015_);
  and _85866_ (_36033_, _36013_, _06306_);
  and _85867_ (_36034_, _36033_, _36031_);
  or _85868_ (_36035_, _36034_, _36030_);
  and _85869_ (_36036_, _36035_, _12514_);
  and _85870_ (_36037_, _35961_, _06411_);
  and _85871_ (_36038_, _36037_, _36031_);
  and _85872_ (_36039_, _35968_, _07124_);
  or _85873_ (_36040_, _36039_, _06303_);
  or _85874_ (_36041_, _36040_, _36038_);
  or _85875_ (_36042_, _36041_, _36036_);
  and _85876_ (_36044_, _15410_, _07858_);
  or _85877_ (_36045_, _35956_, _08819_);
  or _85878_ (_36046_, _36045_, _36044_);
  and _85879_ (_36047_, _36046_, _36042_);
  or _85880_ (_36048_, _36047_, _06396_);
  nor _85881_ (_36049_, _10294_, _13718_);
  or _85882_ (_36050_, _36049_, _35956_);
  or _85883_ (_36051_, _36050_, _08824_);
  and _85884_ (_36052_, _36051_, _12558_);
  and _85885_ (_36053_, _36052_, _36048_);
  nor _85886_ (_36055_, _13646_, _13642_);
  or _85887_ (_36056_, _36055_, _13647_);
  and _85888_ (_36057_, _36056_, _06417_);
  or _85889_ (_36058_, _36057_, _07142_);
  or _85890_ (_36059_, _36058_, _36053_);
  or _85891_ (_36060_, _35968_, _05846_);
  and _85892_ (_36061_, _36060_, _06168_);
  and _85893_ (_36062_, _36061_, _36059_);
  and _85894_ (_36063_, _36056_, _06167_);
  or _85895_ (_36064_, _36063_, _06433_);
  or _85896_ (_36066_, _36064_, _36062_);
  or _85897_ (_36067_, _35958_, _06829_);
  and _85898_ (_36068_, _36067_, _07160_);
  and _85899_ (_36069_, _36068_, _36066_);
  and _85900_ (_36070_, _35968_, _07577_);
  or _85901_ (_36071_, _36070_, _06440_);
  or _85902_ (_36072_, _36071_, _36069_);
  and _85903_ (_36073_, _15478_, _07858_);
  or _85904_ (_36074_, _35956_, _06444_);
  or _85905_ (_36075_, _36074_, _36073_);
  and _85906_ (_36077_, _36075_, _01317_);
  and _85907_ (_36078_, _36077_, _36072_);
  or _85908_ (_36079_, _36078_, _35954_);
  and _85909_ (_43770_, _36079_, _43100_);
  not _85910_ (_36080_, \oc8051_golden_model_1.SBUF [0]);
  nor _85911_ (_36081_, _01317_, _36080_);
  nor _85912_ (_36082_, _07783_, _36080_);
  nor _85913_ (_36083_, _08211_, _13750_);
  or _85914_ (_36084_, _36083_, _36082_);
  or _85915_ (_36085_, _36084_, _06161_);
  and _85916_ (_36087_, _07783_, \oc8051_golden_model_1.ACC [0]);
  or _85917_ (_36088_, _36087_, _36082_);
  and _85918_ (_36089_, _36088_, _07056_);
  nor _85919_ (_36090_, _07056_, _36080_);
  or _85920_ (_36091_, _36090_, _06160_);
  or _85921_ (_36092_, _36091_, _36089_);
  and _85922_ (_36093_, _36092_, _07075_);
  and _85923_ (_36094_, _36093_, _36085_);
  and _85924_ (_36095_, _07783_, _07049_);
  or _85925_ (_36096_, _36095_, _36082_);
  and _85926_ (_36098_, _36096_, _06217_);
  or _85927_ (_36099_, _36098_, _36094_);
  and _85928_ (_36100_, _36099_, _06229_);
  and _85929_ (_36101_, _36088_, _06220_);
  or _85930_ (_36102_, _36101_, _09842_);
  or _85931_ (_36103_, _36102_, _36100_);
  or _85932_ (_36104_, _36096_, _06132_);
  and _85933_ (_36105_, _36104_, _36103_);
  or _85934_ (_36106_, _36105_, _06116_);
  and _85935_ (_36107_, _09160_, _07783_);
  or _85936_ (_36109_, _36082_, _06117_);
  or _85937_ (_36110_, _36109_, _36107_);
  and _85938_ (_36111_, _36110_, _36106_);
  or _85939_ (_36112_, _36111_, _05787_);
  and _85940_ (_36113_, _14260_, _07783_);
  or _85941_ (_36114_, _36082_, _06114_);
  or _85942_ (_36115_, _36114_, _36113_);
  and _85943_ (_36116_, _36115_, _06111_);
  and _85944_ (_36117_, _36116_, _36112_);
  and _85945_ (_36118_, _07783_, _08708_);
  or _85946_ (_36120_, _36118_, _36082_);
  and _85947_ (_36121_, _36120_, _06110_);
  or _85948_ (_36122_, _36121_, _06297_);
  or _85949_ (_36123_, _36122_, _36117_);
  and _85950_ (_36124_, _14275_, _07783_);
  or _85951_ (_36125_, _36082_, _07127_);
  or _85952_ (_36126_, _36125_, _36124_);
  and _85953_ (_36127_, _36126_, _07125_);
  and _85954_ (_36128_, _36127_, _36123_);
  nor _85955_ (_36129_, _12321_, _13750_);
  or _85956_ (_36131_, _36129_, _36082_);
  nand _85957_ (_36132_, _10276_, _07783_);
  and _85958_ (_36133_, _36132_, _06402_);
  and _85959_ (_36134_, _36133_, _36131_);
  or _85960_ (_36135_, _36134_, _36128_);
  and _85961_ (_36136_, _36135_, _07132_);
  nand _85962_ (_36137_, _36120_, _06306_);
  nor _85963_ (_36138_, _36137_, _36083_);
  or _85964_ (_36139_, _36138_, _06411_);
  or _85965_ (_36140_, _36139_, _36136_);
  nor _85966_ (_36142_, _36082_, _07130_);
  nand _85967_ (_36143_, _36142_, _36132_);
  and _85968_ (_36144_, _36143_, _36140_);
  or _85969_ (_36145_, _36144_, _06303_);
  and _85970_ (_36146_, _14167_, _07783_);
  or _85971_ (_36147_, _36082_, _08819_);
  or _85972_ (_36148_, _36147_, _36146_);
  and _85973_ (_36149_, _36148_, _08824_);
  and _85974_ (_36150_, _36149_, _36145_);
  and _85975_ (_36151_, _36131_, _06396_);
  or _85976_ (_36153_, _36151_, _19287_);
  or _85977_ (_36154_, _36153_, _36150_);
  or _85978_ (_36155_, _36084_, _06630_);
  and _85979_ (_36156_, _36155_, _01317_);
  and _85980_ (_36157_, _36156_, _36154_);
  or _85981_ (_36158_, _36157_, _36081_);
  and _85982_ (_43772_, _36158_, _43100_);
  not _85983_ (_36159_, \oc8051_golden_model_1.SBUF [1]);
  nor _85984_ (_36160_, _01317_, _36159_);
  or _85985_ (_36161_, _14442_, _13750_);
  or _85986_ (_36163_, _07783_, \oc8051_golden_model_1.SBUF [1]);
  and _85987_ (_36164_, _36163_, _05787_);
  and _85988_ (_36165_, _36164_, _36161_);
  and _85989_ (_36166_, _09115_, _07783_);
  nor _85990_ (_36167_, _07783_, _36159_);
  or _85991_ (_36168_, _36167_, _06117_);
  or _85992_ (_36169_, _36168_, _36166_);
  and _85993_ (_36170_, _14363_, _07783_);
  not _85994_ (_36171_, _36170_);
  and _85995_ (_36172_, _36171_, _36163_);
  or _85996_ (_36174_, _36172_, _06161_);
  and _85997_ (_36175_, _07783_, \oc8051_golden_model_1.ACC [1]);
  or _85998_ (_36176_, _36175_, _36167_);
  and _85999_ (_36177_, _36176_, _07056_);
  nor _86000_ (_36178_, _07056_, _36159_);
  or _86001_ (_36179_, _36178_, _06160_);
  or _86002_ (_36180_, _36179_, _36177_);
  and _86003_ (_36181_, _36180_, _07075_);
  and _86004_ (_36182_, _36181_, _36174_);
  and _86005_ (_36183_, _07783_, _07306_);
  or _86006_ (_36185_, _36183_, _36167_);
  and _86007_ (_36186_, _36185_, _06217_);
  or _86008_ (_36187_, _36186_, _36182_);
  and _86009_ (_36188_, _36187_, _06229_);
  and _86010_ (_36189_, _36176_, _06220_);
  or _86011_ (_36190_, _36189_, _09842_);
  or _86012_ (_36191_, _36190_, _36188_);
  or _86013_ (_36192_, _36185_, _06132_);
  and _86014_ (_36193_, _36192_, _36191_);
  or _86015_ (_36194_, _36193_, _06116_);
  and _86016_ (_36196_, _36194_, _06114_);
  and _86017_ (_36197_, _36196_, _36169_);
  or _86018_ (_36198_, _36197_, _36165_);
  and _86019_ (_36199_, _36198_, _06298_);
  or _86020_ (_36200_, _14346_, _13750_);
  and _86021_ (_36201_, _36163_, _06297_);
  and _86022_ (_36202_, _36201_, _36200_);
  nand _86023_ (_36203_, _07783_, _06945_);
  and _86024_ (_36204_, _36163_, _06110_);
  and _86025_ (_36205_, _36204_, _36203_);
  or _86026_ (_36207_, _36205_, _06402_);
  or _86027_ (_36208_, _36207_, _36202_);
  or _86028_ (_36209_, _36208_, _36199_);
  nor _86029_ (_36210_, _10277_, _13750_);
  or _86030_ (_36211_, _36210_, _36167_);
  nand _86031_ (_36212_, _10275_, _07783_);
  and _86032_ (_36213_, _36212_, _36211_);
  or _86033_ (_36214_, _36213_, _07125_);
  and _86034_ (_36215_, _36214_, _07132_);
  and _86035_ (_36216_, _36215_, _36209_);
  or _86036_ (_36218_, _14344_, _13750_);
  and _86037_ (_36219_, _36163_, _06306_);
  and _86038_ (_36220_, _36219_, _36218_);
  or _86039_ (_36221_, _36220_, _06411_);
  or _86040_ (_36222_, _36221_, _36216_);
  nor _86041_ (_36223_, _36167_, _07130_);
  nand _86042_ (_36224_, _36223_, _36212_);
  and _86043_ (_36225_, _36224_, _08819_);
  and _86044_ (_36226_, _36225_, _36222_);
  or _86045_ (_36227_, _36203_, _08176_);
  and _86046_ (_36229_, _36163_, _06303_);
  and _86047_ (_36230_, _36229_, _36227_);
  or _86048_ (_36231_, _36230_, _06396_);
  or _86049_ (_36232_, _36231_, _36226_);
  or _86050_ (_36233_, _36211_, _08824_);
  and _86051_ (_36234_, _36233_, _36232_);
  and _86052_ (_36235_, _36234_, _06829_);
  and _86053_ (_36236_, _36172_, _06433_);
  or _86054_ (_36237_, _36236_, _06440_);
  or _86055_ (_36238_, _36237_, _36235_);
  or _86056_ (_36240_, _36167_, _06444_);
  or _86057_ (_36241_, _36240_, _36170_);
  and _86058_ (_36242_, _36241_, _01317_);
  and _86059_ (_36243_, _36242_, _36238_);
  or _86060_ (_36244_, _36243_, _36160_);
  and _86061_ (_43773_, _36244_, _43100_);
  and _86062_ (_36245_, _01321_, \oc8051_golden_model_1.SBUF [2]);
  and _86063_ (_36246_, _13750_, \oc8051_golden_model_1.SBUF [2]);
  or _86064_ (_36247_, _36246_, _08248_);
  and _86065_ (_36248_, _07783_, _08768_);
  or _86066_ (_36250_, _36248_, _36246_);
  and _86067_ (_36251_, _36250_, _06306_);
  and _86068_ (_36252_, _36251_, _36247_);
  and _86069_ (_36253_, _09211_, _07783_);
  or _86070_ (_36254_, _36253_, _36246_);
  and _86071_ (_36255_, _36254_, _06116_);
  and _86072_ (_36256_, _14542_, _07783_);
  or _86073_ (_36257_, _36256_, _36246_);
  or _86074_ (_36258_, _36257_, _06161_);
  and _86075_ (_36259_, _07783_, \oc8051_golden_model_1.ACC [2]);
  or _86076_ (_36261_, _36259_, _36246_);
  and _86077_ (_36262_, _36261_, _07056_);
  and _86078_ (_36263_, _07057_, \oc8051_golden_model_1.SBUF [2]);
  or _86079_ (_36264_, _36263_, _06160_);
  or _86080_ (_36265_, _36264_, _36262_);
  and _86081_ (_36266_, _36265_, _07075_);
  and _86082_ (_36267_, _36266_, _36258_);
  and _86083_ (_36268_, _07783_, _07708_);
  or _86084_ (_36269_, _36268_, _36246_);
  and _86085_ (_36270_, _36269_, _06217_);
  or _86086_ (_36272_, _36270_, _36267_);
  and _86087_ (_36273_, _36272_, _06229_);
  and _86088_ (_36274_, _36261_, _06220_);
  or _86089_ (_36275_, _36274_, _09842_);
  or _86090_ (_36276_, _36275_, _36273_);
  or _86091_ (_36277_, _36269_, _06132_);
  and _86092_ (_36278_, _36277_, _06117_);
  and _86093_ (_36279_, _36278_, _36276_);
  or _86094_ (_36280_, _36279_, _05787_);
  or _86095_ (_36281_, _36280_, _36255_);
  and _86096_ (_36283_, _14630_, _07783_);
  or _86097_ (_36284_, _36283_, _36246_);
  or _86098_ (_36285_, _36284_, _06114_);
  and _86099_ (_36286_, _36285_, _06111_);
  and _86100_ (_36287_, _36286_, _36281_);
  and _86101_ (_36288_, _36250_, _06110_);
  or _86102_ (_36289_, _36288_, _06297_);
  or _86103_ (_36290_, _36289_, _36287_);
  and _86104_ (_36291_, _14646_, _07783_);
  or _86105_ (_36292_, _36246_, _07127_);
  or _86106_ (_36294_, _36292_, _36291_);
  and _86107_ (_36295_, _36294_, _07125_);
  and _86108_ (_36296_, _36295_, _36290_);
  and _86109_ (_36297_, _10282_, _07783_);
  or _86110_ (_36298_, _36297_, _36246_);
  and _86111_ (_36299_, _36298_, _06402_);
  or _86112_ (_36300_, _36299_, _36296_);
  and _86113_ (_36301_, _36300_, _07132_);
  or _86114_ (_36302_, _36301_, _36252_);
  and _86115_ (_36303_, _36302_, _07130_);
  and _86116_ (_36305_, _36261_, _06411_);
  and _86117_ (_36306_, _36305_, _36247_);
  or _86118_ (_36307_, _36306_, _06303_);
  or _86119_ (_36308_, _36307_, _36303_);
  and _86120_ (_36309_, _14643_, _07783_);
  or _86121_ (_36310_, _36246_, _08819_);
  or _86122_ (_36311_, _36310_, _36309_);
  and _86123_ (_36312_, _36311_, _08824_);
  and _86124_ (_36313_, _36312_, _36308_);
  nor _86125_ (_36314_, _10281_, _13750_);
  or _86126_ (_36316_, _36314_, _36246_);
  and _86127_ (_36317_, _36316_, _06396_);
  or _86128_ (_36318_, _36317_, _36313_);
  and _86129_ (_36319_, _36318_, _06829_);
  and _86130_ (_36320_, _36257_, _06433_);
  or _86131_ (_36321_, _36320_, _06440_);
  or _86132_ (_36322_, _36321_, _36319_);
  and _86133_ (_36323_, _14710_, _07783_);
  or _86134_ (_36324_, _36246_, _06444_);
  or _86135_ (_36325_, _36324_, _36323_);
  and _86136_ (_36327_, _36325_, _01317_);
  and _86137_ (_36328_, _36327_, _36322_);
  or _86138_ (_36329_, _36328_, _36245_);
  and _86139_ (_43774_, _36329_, _43100_);
  and _86140_ (_36330_, _13750_, \oc8051_golden_model_1.SBUF [3]);
  or _86141_ (_36331_, _36330_, _08140_);
  and _86142_ (_36332_, _07783_, _08712_);
  or _86143_ (_36333_, _36332_, _36330_);
  and _86144_ (_36334_, _36333_, _06306_);
  and _86145_ (_36335_, _36334_, _36331_);
  and _86146_ (_36337_, _14738_, _07783_);
  or _86147_ (_36338_, _36337_, _36330_);
  or _86148_ (_36339_, _36338_, _06161_);
  and _86149_ (_36340_, _07783_, \oc8051_golden_model_1.ACC [3]);
  or _86150_ (_36341_, _36340_, _36330_);
  and _86151_ (_36342_, _36341_, _07056_);
  and _86152_ (_36343_, _07057_, \oc8051_golden_model_1.SBUF [3]);
  or _86153_ (_36344_, _36343_, _06160_);
  or _86154_ (_36345_, _36344_, _36342_);
  and _86155_ (_36346_, _36345_, _07075_);
  and _86156_ (_36348_, _36346_, _36339_);
  and _86157_ (_36349_, _07783_, _07544_);
  or _86158_ (_36350_, _36349_, _36330_);
  and _86159_ (_36351_, _36350_, _06217_);
  or _86160_ (_36352_, _36351_, _36348_);
  and _86161_ (_36353_, _36352_, _06229_);
  and _86162_ (_36354_, _36341_, _06220_);
  or _86163_ (_36355_, _36354_, _09842_);
  or _86164_ (_36356_, _36355_, _36353_);
  and _86165_ (_36357_, _36350_, _06117_);
  or _86166_ (_36359_, _36357_, _06133_);
  and _86167_ (_36360_, _36359_, _36356_);
  and _86168_ (_36361_, _09210_, _07783_);
  or _86169_ (_36362_, _36361_, _36330_);
  and _86170_ (_36363_, _36362_, _06116_);
  or _86171_ (_36364_, _36363_, _05787_);
  or _86172_ (_36365_, _36364_, _36360_);
  and _86173_ (_36366_, _14825_, _07783_);
  or _86174_ (_36367_, _36330_, _06114_);
  or _86175_ (_36368_, _36367_, _36366_);
  and _86176_ (_36370_, _36368_, _06111_);
  and _86177_ (_36371_, _36370_, _36365_);
  and _86178_ (_36372_, _36333_, _06110_);
  or _86179_ (_36373_, _36372_, _06297_);
  or _86180_ (_36374_, _36373_, _36371_);
  and _86181_ (_36375_, _14727_, _07783_);
  or _86182_ (_36376_, _36330_, _07127_);
  or _86183_ (_36377_, _36376_, _36375_);
  and _86184_ (_36378_, _36377_, _07125_);
  and _86185_ (_36379_, _36378_, _36374_);
  and _86186_ (_36381_, _12318_, _07783_);
  or _86187_ (_36382_, _36381_, _36330_);
  and _86188_ (_36383_, _36382_, _06402_);
  or _86189_ (_36384_, _36383_, _36379_);
  and _86190_ (_36385_, _36384_, _07132_);
  or _86191_ (_36386_, _36385_, _36335_);
  and _86192_ (_36387_, _36386_, _07130_);
  and _86193_ (_36388_, _36341_, _06411_);
  and _86194_ (_36389_, _36388_, _36331_);
  or _86195_ (_36390_, _36389_, _06303_);
  or _86196_ (_36392_, _36390_, _36387_);
  and _86197_ (_36393_, _14724_, _07783_);
  or _86198_ (_36394_, _36330_, _08819_);
  or _86199_ (_36395_, _36394_, _36393_);
  and _86200_ (_36396_, _36395_, _08824_);
  and _86201_ (_36397_, _36396_, _36392_);
  nor _86202_ (_36398_, _10273_, _13750_);
  or _86203_ (_36399_, _36398_, _36330_);
  and _86204_ (_36400_, _36399_, _06396_);
  or _86205_ (_36401_, _36400_, _06433_);
  or _86206_ (_36403_, _36401_, _36397_);
  or _86207_ (_36404_, _36338_, _06829_);
  and _86208_ (_36405_, _36404_, _06444_);
  and _86209_ (_36406_, _36405_, _36403_);
  and _86210_ (_36407_, _14897_, _07783_);
  or _86211_ (_36408_, _36407_, _36330_);
  and _86212_ (_36409_, _36408_, _06440_);
  or _86213_ (_36410_, _36409_, _01321_);
  or _86214_ (_36411_, _36410_, _36406_);
  or _86215_ (_36412_, _01317_, \oc8051_golden_model_1.SBUF [3]);
  and _86216_ (_36414_, _36412_, _43100_);
  and _86217_ (_43775_, _36414_, _36411_);
  and _86218_ (_36415_, _13750_, \oc8051_golden_model_1.SBUF [4]);
  and _86219_ (_36416_, _14928_, _07783_);
  or _86220_ (_36417_, _36416_, _36415_);
  or _86221_ (_36418_, _36417_, _06161_);
  and _86222_ (_36419_, _07783_, \oc8051_golden_model_1.ACC [4]);
  or _86223_ (_36420_, _36419_, _36415_);
  and _86224_ (_36421_, _36420_, _07056_);
  and _86225_ (_36422_, _07057_, \oc8051_golden_model_1.SBUF [4]);
  or _86226_ (_36423_, _36422_, _06160_);
  or _86227_ (_36424_, _36423_, _36421_);
  and _86228_ (_36425_, _36424_, _07075_);
  and _86229_ (_36426_, _36425_, _36418_);
  and _86230_ (_36427_, _08336_, _07783_);
  or _86231_ (_36428_, _36427_, _36415_);
  and _86232_ (_36429_, _36428_, _06217_);
  or _86233_ (_36430_, _36429_, _36426_);
  and _86234_ (_36431_, _36430_, _06229_);
  and _86235_ (_36432_, _36420_, _06220_);
  or _86236_ (_36434_, _36432_, _09842_);
  or _86237_ (_36435_, _36434_, _36431_);
  or _86238_ (_36436_, _36428_, _06132_);
  and _86239_ (_36437_, _36436_, _36435_);
  or _86240_ (_36438_, _36437_, _06116_);
  and _86241_ (_36439_, _09209_, _07783_);
  or _86242_ (_36440_, _36415_, _06117_);
  or _86243_ (_36441_, _36440_, _36439_);
  and _86244_ (_36442_, _36441_, _06114_);
  and _86245_ (_36443_, _36442_, _36438_);
  and _86246_ (_36445_, _15013_, _07783_);
  or _86247_ (_36446_, _36445_, _36415_);
  and _86248_ (_36447_, _36446_, _05787_);
  or _86249_ (_36448_, _36447_, _36443_);
  or _86250_ (_36449_, _36448_, _11136_);
  and _86251_ (_36450_, _15029_, _07783_);
  or _86252_ (_36451_, _36415_, _07127_);
  or _86253_ (_36452_, _36451_, _36450_);
  and _86254_ (_36453_, _08715_, _07783_);
  or _86255_ (_36454_, _36453_, _36415_);
  or _86256_ (_36456_, _36454_, _06111_);
  and _86257_ (_36457_, _36456_, _07125_);
  and _86258_ (_36458_, _36457_, _36452_);
  and _86259_ (_36459_, _36458_, _36449_);
  and _86260_ (_36460_, _10289_, _07783_);
  or _86261_ (_36461_, _36460_, _36415_);
  and _86262_ (_36462_, _36461_, _06402_);
  or _86263_ (_36463_, _36462_, _36459_);
  and _86264_ (_36464_, _36463_, _07132_);
  or _86265_ (_36465_, _36415_, _08339_);
  and _86266_ (_36467_, _36454_, _06306_);
  and _86267_ (_36468_, _36467_, _36465_);
  or _86268_ (_36469_, _36468_, _36464_);
  and _86269_ (_36470_, _36469_, _07130_);
  and _86270_ (_36471_, _36420_, _06411_);
  and _86271_ (_36472_, _36471_, _36465_);
  or _86272_ (_36473_, _36472_, _06303_);
  or _86273_ (_36474_, _36473_, _36470_);
  and _86274_ (_36475_, _15026_, _07783_);
  or _86275_ (_36476_, _36415_, _08819_);
  or _86276_ (_36478_, _36476_, _36475_);
  and _86277_ (_36479_, _36478_, _08824_);
  and _86278_ (_36480_, _36479_, _36474_);
  nor _86279_ (_36481_, _10288_, _13750_);
  or _86280_ (_36482_, _36481_, _36415_);
  and _86281_ (_36483_, _36482_, _06396_);
  or _86282_ (_36484_, _36483_, _06433_);
  or _86283_ (_36485_, _36484_, _36480_);
  or _86284_ (_36486_, _36417_, _06829_);
  and _86285_ (_36487_, _36486_, _06444_);
  and _86286_ (_36489_, _36487_, _36485_);
  and _86287_ (_36490_, _15087_, _07783_);
  or _86288_ (_36491_, _36490_, _36415_);
  and _86289_ (_36492_, _36491_, _06440_);
  or _86290_ (_36493_, _36492_, _01321_);
  or _86291_ (_36494_, _36493_, _36489_);
  or _86292_ (_36495_, _01317_, \oc8051_golden_model_1.SBUF [4]);
  and _86293_ (_36496_, _36495_, _43100_);
  and _86294_ (_43776_, _36496_, _36494_);
  and _86295_ (_36497_, _13750_, \oc8051_golden_model_1.SBUF [5]);
  or _86296_ (_36499_, _36497_, _08104_);
  and _86297_ (_36500_, _08736_, _07783_);
  or _86298_ (_36501_, _36500_, _36497_);
  and _86299_ (_36502_, _36501_, _06306_);
  and _86300_ (_36503_, _36502_, _36499_);
  and _86301_ (_36504_, _15119_, _07783_);
  or _86302_ (_36505_, _36504_, _36497_);
  or _86303_ (_36506_, _36505_, _06161_);
  and _86304_ (_36507_, _07783_, \oc8051_golden_model_1.ACC [5]);
  or _86305_ (_36508_, _36507_, _36497_);
  and _86306_ (_36510_, _36508_, _07056_);
  and _86307_ (_36511_, _07057_, \oc8051_golden_model_1.SBUF [5]);
  or _86308_ (_36512_, _36511_, _06160_);
  or _86309_ (_36513_, _36512_, _36510_);
  and _86310_ (_36514_, _36513_, _07075_);
  and _86311_ (_36515_, _36514_, _36506_);
  and _86312_ (_36516_, _08101_, _07783_);
  or _86313_ (_36517_, _36516_, _36497_);
  and _86314_ (_36518_, _36517_, _06217_);
  or _86315_ (_36519_, _36518_, _36515_);
  and _86316_ (_36521_, _36519_, _06229_);
  and _86317_ (_36522_, _36508_, _06220_);
  or _86318_ (_36523_, _36522_, _09842_);
  or _86319_ (_36524_, _36523_, _36521_);
  or _86320_ (_36525_, _36517_, _06132_);
  and _86321_ (_36526_, _36525_, _36524_);
  or _86322_ (_36527_, _36526_, _06116_);
  and _86323_ (_36528_, _09208_, _07783_);
  or _86324_ (_36529_, _36497_, _06117_);
  or _86325_ (_36530_, _36529_, _36528_);
  and _86326_ (_36532_, _36530_, _06114_);
  and _86327_ (_36533_, _36532_, _36527_);
  and _86328_ (_36534_, _15203_, _07783_);
  or _86329_ (_36535_, _36534_, _36497_);
  and _86330_ (_36536_, _36535_, _05787_);
  or _86331_ (_36537_, _36536_, _11136_);
  or _86332_ (_36538_, _36537_, _36533_);
  and _86333_ (_36539_, _15219_, _07783_);
  or _86334_ (_36540_, _36497_, _07127_);
  or _86335_ (_36541_, _36540_, _36539_);
  or _86336_ (_36543_, _36501_, _06111_);
  and _86337_ (_36544_, _36543_, _07125_);
  and _86338_ (_36545_, _36544_, _36541_);
  and _86339_ (_36546_, _36545_, _36538_);
  and _86340_ (_36547_, _12325_, _07783_);
  or _86341_ (_36548_, _36547_, _36497_);
  and _86342_ (_36549_, _36548_, _06402_);
  or _86343_ (_36550_, _36549_, _36546_);
  and _86344_ (_36551_, _36550_, _07132_);
  or _86345_ (_36552_, _36551_, _36503_);
  and _86346_ (_36554_, _36552_, _07130_);
  and _86347_ (_36555_, _36508_, _06411_);
  and _86348_ (_36556_, _36555_, _36499_);
  or _86349_ (_36557_, _36556_, _06303_);
  or _86350_ (_36558_, _36557_, _36554_);
  and _86351_ (_36559_, _15216_, _07783_);
  or _86352_ (_36560_, _36497_, _08819_);
  or _86353_ (_36561_, _36560_, _36559_);
  and _86354_ (_36562_, _36561_, _08824_);
  and _86355_ (_36563_, _36562_, _36558_);
  nor _86356_ (_36565_, _10269_, _13750_);
  or _86357_ (_36566_, _36565_, _36497_);
  and _86358_ (_36567_, _36566_, _06396_);
  or _86359_ (_36568_, _36567_, _06433_);
  or _86360_ (_36569_, _36568_, _36563_);
  or _86361_ (_36570_, _36505_, _06829_);
  and _86362_ (_36571_, _36570_, _06444_);
  and _86363_ (_36572_, _36571_, _36569_);
  and _86364_ (_36573_, _15275_, _07783_);
  or _86365_ (_36574_, _36573_, _36497_);
  and _86366_ (_36576_, _36574_, _06440_);
  or _86367_ (_36577_, _36576_, _01321_);
  or _86368_ (_36578_, _36577_, _36572_);
  or _86369_ (_36579_, _01317_, \oc8051_golden_model_1.SBUF [5]);
  and _86370_ (_36580_, _36579_, _43100_);
  and _86371_ (_43777_, _36580_, _36578_);
  and _86372_ (_36581_, _13750_, \oc8051_golden_model_1.SBUF [6]);
  and _86373_ (_36582_, _15300_, _07783_);
  or _86374_ (_36583_, _36582_, _36581_);
  or _86375_ (_36584_, _36583_, _06161_);
  and _86376_ (_36586_, _07783_, \oc8051_golden_model_1.ACC [6]);
  or _86377_ (_36587_, _36586_, _36581_);
  and _86378_ (_36588_, _36587_, _07056_);
  and _86379_ (_36589_, _07057_, \oc8051_golden_model_1.SBUF [6]);
  or _86380_ (_36590_, _36589_, _06160_);
  or _86381_ (_36591_, _36590_, _36588_);
  and _86382_ (_36592_, _36591_, _07075_);
  and _86383_ (_36593_, _36592_, _36584_);
  and _86384_ (_36594_, _08012_, _07783_);
  or _86385_ (_36595_, _36594_, _36581_);
  and _86386_ (_36597_, _36595_, _06217_);
  or _86387_ (_36598_, _36597_, _36593_);
  and _86388_ (_36599_, _36598_, _06229_);
  and _86389_ (_36600_, _36587_, _06220_);
  or _86390_ (_36601_, _36600_, _09842_);
  or _86391_ (_36602_, _36601_, _36599_);
  or _86392_ (_36603_, _36595_, _06132_);
  and _86393_ (_36604_, _36603_, _36602_);
  or _86394_ (_36605_, _36604_, _06116_);
  and _86395_ (_36606_, _09207_, _07783_);
  or _86396_ (_36608_, _36581_, _06117_);
  or _86397_ (_36609_, _36608_, _36606_);
  and _86398_ (_36610_, _36609_, _06114_);
  and _86399_ (_36611_, _36610_, _36605_);
  and _86400_ (_36612_, _15395_, _07783_);
  or _86401_ (_36613_, _36612_, _36581_);
  and _86402_ (_36614_, _36613_, _05787_);
  or _86403_ (_36615_, _36614_, _11136_);
  or _86404_ (_36616_, _36615_, _36611_);
  and _86405_ (_36617_, _15413_, _07783_);
  or _86406_ (_36619_, _36581_, _07127_);
  or _86407_ (_36620_, _36619_, _36617_);
  and _86408_ (_36621_, _15402_, _07783_);
  or _86409_ (_36622_, _36621_, _36581_);
  or _86410_ (_36623_, _36622_, _06111_);
  and _86411_ (_36624_, _36623_, _07125_);
  and _86412_ (_36625_, _36624_, _36620_);
  and _86413_ (_36626_, _36625_, _36616_);
  and _86414_ (_36627_, _10295_, _07783_);
  or _86415_ (_36628_, _36627_, _36581_);
  and _86416_ (_36630_, _36628_, _06402_);
  or _86417_ (_36631_, _36630_, _36626_);
  and _86418_ (_36632_, _36631_, _07132_);
  or _86419_ (_36633_, _36581_, _08015_);
  and _86420_ (_36634_, _36622_, _06306_);
  and _86421_ (_36635_, _36634_, _36633_);
  or _86422_ (_36636_, _36635_, _36632_);
  and _86423_ (_36637_, _36636_, _07130_);
  and _86424_ (_36638_, _36587_, _06411_);
  and _86425_ (_36639_, _36638_, _36633_);
  or _86426_ (_36641_, _36639_, _06303_);
  or _86427_ (_36642_, _36641_, _36637_);
  and _86428_ (_36643_, _15410_, _07783_);
  or _86429_ (_36644_, _36581_, _08819_);
  or _86430_ (_36645_, _36644_, _36643_);
  and _86431_ (_36646_, _36645_, _08824_);
  and _86432_ (_36647_, _36646_, _36642_);
  nor _86433_ (_36648_, _10294_, _13750_);
  or _86434_ (_36649_, _36648_, _36581_);
  and _86435_ (_36650_, _36649_, _06396_);
  or _86436_ (_36652_, _36650_, _06433_);
  or _86437_ (_36653_, _36652_, _36647_);
  or _86438_ (_36654_, _36583_, _06829_);
  and _86439_ (_36655_, _36654_, _06444_);
  and _86440_ (_36656_, _36655_, _36653_);
  and _86441_ (_36657_, _15478_, _07783_);
  or _86442_ (_36658_, _36657_, _36581_);
  and _86443_ (_36659_, _36658_, _06440_);
  or _86444_ (_36660_, _36659_, _01321_);
  or _86445_ (_36661_, _36660_, _36656_);
  or _86446_ (_36663_, _01317_, \oc8051_golden_model_1.SBUF [6]);
  and _86447_ (_36664_, _36663_, _43100_);
  and _86448_ (_43778_, _36664_, _36661_);
  not _86449_ (_36665_, \oc8051_golden_model_1.PSW [0]);
  nor _86450_ (_36666_, _01317_, _36665_);
  nand _86451_ (_36667_, _10276_, _07794_);
  nor _86452_ (_36668_, _07794_, _36665_);
  nor _86453_ (_36669_, _36668_, _07130_);
  nand _86454_ (_36670_, _36669_, _36667_);
  nor _86455_ (_36671_, _08404_, _36665_);
  and _86456_ (_36673_, _14169_, _08404_);
  or _86457_ (_36674_, _36673_, _36671_);
  or _86458_ (_36675_, _36674_, _06157_);
  nor _86459_ (_36676_, _08211_, _14076_);
  or _86460_ (_36677_, _36676_, _36668_);
  and _86461_ (_36678_, _36677_, _06160_);
  nor _86462_ (_36679_, _07056_, _36665_);
  and _86463_ (_36680_, _07794_, \oc8051_golden_model_1.ACC [0]);
  or _86464_ (_36681_, _36680_, _36668_);
  and _86465_ (_36682_, _36681_, _07056_);
  or _86466_ (_36684_, _36682_, _36679_);
  and _86467_ (_36685_, _36684_, _06161_);
  or _86468_ (_36686_, _36685_, _06156_);
  or _86469_ (_36687_, _36686_, _36678_);
  and _86470_ (_36688_, _36687_, _36675_);
  and _86471_ (_36689_, _36688_, _07075_);
  and _86472_ (_36690_, _07794_, _07049_);
  or _86473_ (_36691_, _36690_, _36668_);
  and _86474_ (_36692_, _36691_, _06217_);
  or _86475_ (_36693_, _36692_, _06220_);
  or _86476_ (_36695_, _36693_, _36689_);
  or _86477_ (_36696_, _36681_, _06229_);
  and _86478_ (_36697_, _36696_, _06153_);
  and _86479_ (_36698_, _36697_, _36695_);
  and _86480_ (_36699_, _36668_, _06152_);
  or _86481_ (_36700_, _36699_, _06145_);
  or _86482_ (_36701_, _36700_, _36698_);
  or _86483_ (_36702_, _36677_, _06146_);
  and _86484_ (_36703_, _36702_, _06140_);
  and _86485_ (_36704_, _36703_, _36701_);
  or _86486_ (_36706_, _36671_, _14170_);
  and _86487_ (_36707_, _36706_, _06139_);
  and _86488_ (_36708_, _36707_, _36674_);
  or _86489_ (_36709_, _36708_, _09842_);
  or _86490_ (_36710_, _36709_, _36704_);
  or _86491_ (_36711_, _36691_, _06132_);
  and _86492_ (_36712_, _36711_, _36710_);
  or _86493_ (_36713_, _36712_, _06116_);
  and _86494_ (_36714_, _09160_, _07794_);
  or _86495_ (_36715_, _36668_, _06117_);
  or _86496_ (_36717_, _36715_, _36714_);
  and _86497_ (_36718_, _36717_, _06114_);
  and _86498_ (_36719_, _36718_, _36713_);
  and _86499_ (_36720_, _14260_, _07794_);
  or _86500_ (_36721_, _36720_, _36668_);
  and _86501_ (_36722_, _36721_, _05787_);
  or _86502_ (_36723_, _36722_, _36719_);
  or _86503_ (_36724_, _36723_, _11136_);
  and _86504_ (_36725_, _14275_, _07794_);
  or _86505_ (_36726_, _36668_, _07127_);
  or _86506_ (_36728_, _36726_, _36725_);
  and _86507_ (_36729_, _07794_, _08708_);
  or _86508_ (_36730_, _36729_, _36668_);
  or _86509_ (_36731_, _36730_, _06111_);
  and _86510_ (_36732_, _36731_, _07125_);
  and _86511_ (_36733_, _36732_, _36728_);
  and _86512_ (_36734_, _36733_, _36724_);
  nor _86513_ (_36735_, _12321_, _14076_);
  or _86514_ (_36736_, _36735_, _36668_);
  and _86515_ (_36737_, _36667_, _06402_);
  and _86516_ (_36739_, _36737_, _36736_);
  or _86517_ (_36740_, _36739_, _36734_);
  and _86518_ (_36741_, _36740_, _07132_);
  nand _86519_ (_36742_, _36730_, _06306_);
  nor _86520_ (_36743_, _36742_, _36676_);
  or _86521_ (_36744_, _36743_, _06411_);
  or _86522_ (_36745_, _36744_, _36741_);
  and _86523_ (_36746_, _36745_, _36670_);
  or _86524_ (_36747_, _36746_, _06303_);
  and _86525_ (_36748_, _14167_, _07794_);
  or _86526_ (_36750_, _36668_, _08819_);
  or _86527_ (_36751_, _36750_, _36748_);
  and _86528_ (_36752_, _36751_, _08824_);
  and _86529_ (_36753_, _36752_, _36747_);
  and _86530_ (_36754_, _36736_, _06396_);
  or _86531_ (_36755_, _36754_, _06433_);
  or _86532_ (_36756_, _36755_, _36753_);
  or _86533_ (_36757_, _36677_, _06829_);
  and _86534_ (_36758_, _36757_, _36756_);
  or _86535_ (_36759_, _36758_, _05748_);
  or _86536_ (_36761_, _36668_, _05749_);
  and _86537_ (_36762_, _36761_, _36759_);
  or _86538_ (_36763_, _36762_, _06440_);
  or _86539_ (_36764_, _36677_, _06444_);
  and _86540_ (_36765_, _36764_, _01317_);
  and _86541_ (_36766_, _36765_, _36763_);
  or _86542_ (_36767_, _36766_, _36666_);
  and _86543_ (_43779_, _36767_, _43100_);
  not _86544_ (_36768_, \oc8051_golden_model_1.PSW [1]);
  nor _86545_ (_36769_, _01317_, _36768_);
  or _86546_ (_36771_, _14442_, _14076_);
  or _86547_ (_36772_, _07794_, \oc8051_golden_model_1.PSW [1]);
  and _86548_ (_36773_, _36772_, _05787_);
  and _86549_ (_36774_, _36773_, _36771_);
  nor _86550_ (_36775_, _07794_, _36768_);
  and _86551_ (_36776_, _07794_, _07306_);
  or _86552_ (_36777_, _36776_, _36775_);
  or _86553_ (_36778_, _36777_, _07075_);
  and _86554_ (_36779_, _14363_, _07794_);
  not _86555_ (_36780_, _36779_);
  and _86556_ (_36782_, _36780_, _36772_);
  or _86557_ (_36783_, _36782_, _06161_);
  and _86558_ (_36784_, _07794_, \oc8051_golden_model_1.ACC [1]);
  or _86559_ (_36785_, _36784_, _36775_);
  and _86560_ (_36786_, _36785_, _07056_);
  nor _86561_ (_36787_, _07056_, _36768_);
  or _86562_ (_36788_, _36787_, _06160_);
  or _86563_ (_36789_, _36788_, _36786_);
  and _86564_ (_36790_, _36789_, _06157_);
  and _86565_ (_36791_, _36790_, _36783_);
  nor _86566_ (_36793_, _08404_, _36768_);
  and _86567_ (_36794_, _14367_, _08404_);
  or _86568_ (_36795_, _36794_, _36793_);
  and _86569_ (_36796_, _36795_, _06156_);
  or _86570_ (_36797_, _36796_, _06217_);
  or _86571_ (_36798_, _36797_, _36791_);
  and _86572_ (_36799_, _36798_, _36778_);
  or _86573_ (_36800_, _36799_, _06220_);
  or _86574_ (_36801_, _36785_, _06229_);
  and _86575_ (_36802_, _36801_, _06153_);
  and _86576_ (_36804_, _36802_, _36800_);
  and _86577_ (_36805_, _14349_, _08404_);
  or _86578_ (_36806_, _36805_, _36793_);
  and _86579_ (_36807_, _36806_, _06152_);
  or _86580_ (_36808_, _36807_, _06145_);
  or _86581_ (_36809_, _36808_, _36804_);
  and _86582_ (_36810_, _36794_, _14382_);
  or _86583_ (_36811_, _36793_, _06146_);
  or _86584_ (_36812_, _36811_, _36810_);
  and _86585_ (_36813_, _36812_, _36809_);
  and _86586_ (_36815_, _36813_, _06140_);
  and _86587_ (_36816_, _14351_, _08404_);
  or _86588_ (_36817_, _36793_, _36816_);
  and _86589_ (_36818_, _36817_, _06139_);
  or _86590_ (_36819_, _36818_, _09842_);
  or _86591_ (_36820_, _36819_, _36815_);
  or _86592_ (_36821_, _36777_, _06132_);
  and _86593_ (_36822_, _36821_, _36820_);
  or _86594_ (_36823_, _36822_, _06116_);
  and _86595_ (_36824_, _09115_, _07794_);
  or _86596_ (_36826_, _36775_, _06117_);
  or _86597_ (_36827_, _36826_, _36824_);
  and _86598_ (_36828_, _36827_, _06114_);
  and _86599_ (_36829_, _36828_, _36823_);
  or _86600_ (_36830_, _36829_, _36774_);
  and _86601_ (_36831_, _36830_, _06298_);
  or _86602_ (_36832_, _14346_, _14076_);
  and _86603_ (_36833_, _36772_, _06297_);
  and _86604_ (_36834_, _36833_, _36832_);
  nand _86605_ (_36835_, _07794_, _06945_);
  and _86606_ (_36837_, _36835_, _06110_);
  and _86607_ (_36838_, _36837_, _36772_);
  or _86608_ (_36839_, _36838_, _06402_);
  or _86609_ (_36840_, _36839_, _36834_);
  or _86610_ (_36841_, _36840_, _36831_);
  nor _86611_ (_36842_, _10277_, _14076_);
  or _86612_ (_36843_, _36842_, _36775_);
  nand _86613_ (_36844_, _10275_, _07794_);
  and _86614_ (_36845_, _36844_, _36843_);
  or _86615_ (_36846_, _36845_, _07125_);
  and _86616_ (_36848_, _36846_, _07132_);
  and _86617_ (_36849_, _36848_, _36841_);
  or _86618_ (_36850_, _14344_, _14076_);
  and _86619_ (_36851_, _36772_, _06306_);
  and _86620_ (_36852_, _36851_, _36850_);
  or _86621_ (_36853_, _36852_, _06411_);
  or _86622_ (_36854_, _36853_, _36849_);
  nor _86623_ (_36855_, _36775_, _07130_);
  nand _86624_ (_36856_, _36855_, _36844_);
  and _86625_ (_36857_, _36856_, _08819_);
  and _86626_ (_36859_, _36857_, _36854_);
  or _86627_ (_36860_, _36835_, _08176_);
  and _86628_ (_36861_, _36772_, _06303_);
  and _86629_ (_36862_, _36861_, _36860_);
  or _86630_ (_36863_, _36862_, _06396_);
  or _86631_ (_36864_, _36863_, _36859_);
  or _86632_ (_36865_, _36843_, _08824_);
  and _86633_ (_36866_, _36865_, _36864_);
  or _86634_ (_36867_, _36866_, _06433_);
  or _86635_ (_36868_, _36782_, _06829_);
  and _86636_ (_36870_, _36868_, _05749_);
  and _86637_ (_36871_, _36870_, _36867_);
  and _86638_ (_36872_, _36806_, _05748_);
  or _86639_ (_36873_, _36872_, _06440_);
  or _86640_ (_36874_, _36873_, _36871_);
  or _86641_ (_36875_, _36775_, _06444_);
  or _86642_ (_36876_, _36875_, _36779_);
  and _86643_ (_36877_, _36876_, _01317_);
  and _86644_ (_36878_, _36877_, _36874_);
  or _86645_ (_36879_, _36878_, _36769_);
  and _86646_ (_43780_, _36879_, _43100_);
  and _86647_ (_36881_, _01321_, \oc8051_golden_model_1.PSW [2]);
  or _86648_ (_36882_, _14118_, _11038_);
  or _86649_ (_36883_, _11039_, _10781_);
  and _86650_ (_36884_, _36883_, _36882_);
  and _86651_ (_36885_, _36884_, _17199_);
  nor _86652_ (_36886_, _10657_, _06172_);
  or _86653_ (_36887_, _36886_, \oc8051_golden_model_1.ACC [7]);
  nor _86654_ (_36888_, _10657_, _14131_);
  not _86655_ (_36889_, _36888_);
  and _86656_ (_36891_, _36889_, _36887_);
  not _86657_ (_36892_, _36891_);
  or _86658_ (_36893_, _36892_, _14100_);
  and _86659_ (_36894_, _36889_, _10951_);
  and _86660_ (_36895_, _36894_, _36893_);
  and _86661_ (_36896_, _36888_, _10948_);
  or _86662_ (_36897_, _36896_, _36895_);
  and _86663_ (_36898_, _36897_, _10895_);
  and _86664_ (_36899_, _06122_, _06300_);
  not _86665_ (_36900_, _36899_);
  not _86666_ (_36902_, _10765_);
  nor _86667_ (_36903_, _36902_, _10302_);
  nor _86668_ (_36904_, _10303_, \oc8051_golden_model_1.ACC [7]);
  nor _86669_ (_36905_, _36903_, _36904_);
  not _86670_ (_36906_, _36905_);
  nor _86671_ (_36907_, _36906_, _14087_);
  nor _86672_ (_36908_, _36907_, _36903_);
  and _86673_ (_36909_, _36908_, _10370_);
  and _86674_ (_36910_, _36903_, _10367_);
  or _86675_ (_36911_, _36910_, _36909_);
  or _86676_ (_36913_, _36911_, _36900_);
  and _86677_ (_36914_, _14076_, \oc8051_golden_model_1.PSW [2]);
  and _86678_ (_36915_, _14630_, _07794_);
  or _86679_ (_36916_, _36915_, _36914_);
  and _86680_ (_36917_, _36916_, _05787_);
  and _86681_ (_36918_, _07794_, _07708_);
  or _86682_ (_36919_, _36918_, _36914_);
  or _86683_ (_36920_, _36919_, _06132_);
  and _86684_ (_36921_, _10584_, \oc8051_golden_model_1.ACC [7]);
  nor _86685_ (_36922_, _10584_, \oc8051_golden_model_1.ACC [7]);
  or _86686_ (_36924_, _36922_, _36921_);
  and _86687_ (_36925_, _36924_, _14007_);
  nor _86688_ (_36926_, _36924_, _14007_);
  nor _86689_ (_36927_, _36926_, _36925_);
  not _86690_ (_36928_, _36927_);
  nor _86691_ (_36929_, _36928_, _10646_);
  and _86692_ (_36930_, _36928_, _10646_);
  or _86693_ (_36931_, _36930_, _12380_);
  or _86694_ (_36932_, _36931_, _36929_);
  or _86695_ (_36933_, _36906_, _13995_);
  nand _86696_ (_36935_, _36906_, _13995_);
  and _86697_ (_36936_, _36935_, _36933_);
  and _86698_ (_36937_, _36936_, _10577_);
  nor _86699_ (_36938_, _36936_, _10577_);
  or _86700_ (_36939_, _36938_, _36937_);
  and _86701_ (_36940_, _36939_, _10557_);
  not _86702_ (_36941_, _08404_);
  and _86703_ (_36942_, _36941_, \oc8051_golden_model_1.PSW [2]);
  and _86704_ (_36943_, _14536_, _08404_);
  or _86705_ (_36944_, _36943_, _36942_);
  and _86706_ (_36946_, _36944_, _06152_);
  or _86707_ (_36947_, _36919_, _07075_);
  and _86708_ (_36948_, _14542_, _07794_);
  or _86709_ (_36949_, _36948_, _36914_);
  or _86710_ (_36950_, _36949_, _06161_);
  and _86711_ (_36951_, _07794_, \oc8051_golden_model_1.ACC [2]);
  or _86712_ (_36952_, _36951_, _36914_);
  and _86713_ (_36953_, _36952_, _07056_);
  and _86714_ (_36954_, _07057_, \oc8051_golden_model_1.PSW [2]);
  or _86715_ (_36955_, _36954_, _06160_);
  or _86716_ (_36957_, _36955_, _36953_);
  and _86717_ (_36958_, _36957_, _06157_);
  and _86718_ (_36959_, _36958_, _36950_);
  and _86719_ (_36960_, _14538_, _08404_);
  or _86720_ (_36961_, _36960_, _36942_);
  and _86721_ (_36962_, _36961_, _06156_);
  or _86722_ (_36963_, _36962_, _06217_);
  or _86723_ (_36964_, _36963_, _36959_);
  and _86724_ (_36965_, _36964_, _36947_);
  or _86725_ (_36966_, _36965_, _06220_);
  or _86726_ (_36968_, _36952_, _06229_);
  and _86727_ (_36969_, _36968_, _06153_);
  and _86728_ (_36970_, _36969_, _36966_);
  or _86729_ (_36971_, _36970_, _36946_);
  and _86730_ (_36972_, _36971_, _06146_);
  and _86731_ (_36973_, _36960_, _14569_);
  or _86732_ (_36974_, _36973_, _36942_);
  and _86733_ (_36975_, _36974_, _06145_);
  or _86734_ (_36976_, _36975_, _09295_);
  or _86735_ (_36977_, _36976_, _36972_);
  or _86736_ (_36979_, _16326_, _16210_);
  or _86737_ (_36980_, _36979_, _16438_);
  or _86738_ (_36981_, _36980_, _16556_);
  or _86739_ (_36982_, _36981_, _16673_);
  or _86740_ (_36983_, _36982_, _16790_);
  or _86741_ (_36984_, _36983_, _09838_);
  or _86742_ (_36985_, _36984_, _16908_);
  and _86743_ (_36986_, _36985_, _10554_);
  and _86744_ (_36987_, _36986_, _36977_);
  or _86745_ (_36988_, _36987_, _12379_);
  or _86746_ (_36990_, _36988_, _36940_);
  and _86747_ (_36991_, _36990_, _06265_);
  and _86748_ (_36992_, _36991_, _36932_);
  nor _86749_ (_36993_, _10396_, \oc8051_golden_model_1.ACC [7]);
  nor _86750_ (_36994_, _10395_, _14125_);
  nor _86751_ (_36995_, _36994_, _36993_);
  nor _86752_ (_36996_, _36995_, _10401_);
  nor _86753_ (_36997_, _14017_, _10397_);
  or _86754_ (_36998_, _36997_, _36996_);
  or _86755_ (_36999_, _36998_, _10450_);
  nand _86756_ (_37001_, _36998_, _10450_);
  and _86757_ (_37002_, _37001_, _06260_);
  and _86758_ (_37003_, _37002_, _36999_);
  or _86759_ (_37004_, _37003_, _10387_);
  or _86760_ (_37005_, _37004_, _36992_);
  and _86761_ (_37006_, _36891_, _14027_);
  nor _86762_ (_37007_, _36891_, _14027_);
  nor _86763_ (_37008_, _37007_, _37006_);
  and _86764_ (_37009_, _37008_, _10719_);
  nor _86765_ (_37010_, _37008_, _10719_);
  or _86766_ (_37012_, _37010_, _37009_);
  or _86767_ (_37013_, _37012_, _10388_);
  and _86768_ (_37014_, _37013_, _06140_);
  and _86769_ (_37015_, _37014_, _37005_);
  and _86770_ (_37016_, _14583_, _08404_);
  or _86771_ (_37017_, _37016_, _36942_);
  and _86772_ (_37018_, _37017_, _06139_);
  or _86773_ (_37019_, _37018_, _09842_);
  or _86774_ (_37020_, _37019_, _37015_);
  and _86775_ (_37021_, _37020_, _36920_);
  or _86776_ (_37023_, _37021_, _06116_);
  and _86777_ (_37024_, _09211_, _07794_);
  or _86778_ (_37025_, _36914_, _06117_);
  or _86779_ (_37026_, _37025_, _37024_);
  and _86780_ (_37027_, _37026_, _06114_);
  and _86781_ (_37028_, _37027_, _37023_);
  or _86782_ (_37029_, _37028_, _36917_);
  and _86783_ (_37030_, _37029_, _09861_);
  nor _86784_ (_37031_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and _86785_ (_37032_, _37031_, _09882_);
  nand _86786_ (_37034_, _37032_, _09855_);
  nand _86787_ (_37035_, _37034_, _06298_);
  or _86788_ (_37036_, _37035_, _37030_);
  and _86789_ (_37037_, _14646_, _07794_);
  or _86790_ (_37038_, _36914_, _07127_);
  or _86791_ (_37039_, _37038_, _37037_);
  and _86792_ (_37040_, _07794_, _08768_);
  or _86793_ (_37041_, _37040_, _36914_);
  or _86794_ (_37042_, _37041_, _06111_);
  and _86795_ (_37043_, _37042_, _07125_);
  and _86796_ (_37045_, _37043_, _37039_);
  and _86797_ (_37046_, _37045_, _37036_);
  and _86798_ (_37047_, _10282_, _07794_);
  or _86799_ (_37048_, _37047_, _36914_);
  and _86800_ (_37049_, _37048_, _06402_);
  or _86801_ (_37050_, _37049_, _37046_);
  and _86802_ (_37051_, _37050_, _07132_);
  or _86803_ (_37052_, _36914_, _08248_);
  and _86804_ (_37053_, _37041_, _06306_);
  and _86805_ (_37054_, _37053_, _37052_);
  or _86806_ (_37056_, _37054_, _37051_);
  and _86807_ (_37057_, _37056_, _07130_);
  and _86808_ (_37058_, _36952_, _06411_);
  and _86809_ (_37059_, _37058_, _37052_);
  or _86810_ (_37060_, _37059_, _06303_);
  or _86811_ (_37061_, _37060_, _37057_);
  and _86812_ (_37062_, _14643_, _07794_);
  or _86813_ (_37063_, _36914_, _08819_);
  or _86814_ (_37064_, _37063_, _37062_);
  and _86815_ (_37065_, _37064_, _08824_);
  and _86816_ (_37067_, _37065_, _37061_);
  nor _86817_ (_37068_, _10281_, _14076_);
  or _86818_ (_37069_, _37068_, _36914_);
  and _86819_ (_37070_, _37069_, _06396_);
  or _86820_ (_37071_, _37070_, _36899_);
  or _86821_ (_37072_, _37071_, _37067_);
  nand _86822_ (_37073_, _37072_, _36913_);
  and _86823_ (_37074_, _06288_, _06300_);
  nor _86824_ (_37075_, _37074_, _06976_);
  nand _86825_ (_37076_, _37075_, _37073_);
  or _86826_ (_37078_, _37075_, _36911_);
  and _86827_ (_37079_, _37078_, _06791_);
  and _86828_ (_37080_, _37079_, _37076_);
  and _86829_ (_37081_, _36911_, _06790_);
  or _86830_ (_37082_, _37081_, _10865_);
  or _86831_ (_37083_, _37082_, _37080_);
  nor _86832_ (_37084_, _36924_, _14083_);
  nor _86833_ (_37085_, _37084_, _36921_);
  and _86834_ (_37086_, _37085_, _10891_);
  and _86835_ (_37087_, _36921_, _10888_);
  or _86836_ (_37089_, _37087_, _10867_);
  or _86837_ (_37090_, _37089_, _37086_);
  and _86838_ (_37091_, _37090_, _37083_);
  or _86839_ (_37092_, _37091_, _06406_);
  nor _86840_ (_37093_, _36993_, _14094_);
  nor _86841_ (_37094_, _37093_, _36994_);
  and _86842_ (_37095_, _37094_, _10921_);
  and _86843_ (_37096_, _36994_, _10918_);
  or _86844_ (_37097_, _37096_, _06407_);
  or _86845_ (_37098_, _37097_, _37095_);
  and _86846_ (_37100_, _37098_, _10927_);
  and _86847_ (_37101_, _37100_, _37092_);
  or _86848_ (_37102_, _37101_, _36898_);
  and _86849_ (_37103_, _37102_, _10963_);
  nand _86850_ (_37104_, _10997_, _36902_);
  nand _86851_ (_37105_, _37104_, _18454_);
  nor _86852_ (_37106_, _37105_, _14108_);
  or _86853_ (_37107_, _37106_, _17195_);
  or _86854_ (_37108_, _37107_, _37103_);
  and _86855_ (_37109_, _36884_, _06276_);
  or _86856_ (_37111_, _37109_, _11041_);
  and _86857_ (_37112_, _37111_, _37108_);
  or _86858_ (_37113_, _37112_, _36885_);
  and _86859_ (_37114_, _37113_, _12690_);
  or _86860_ (_37115_, _10297_, _08809_);
  and _86861_ (_37116_, _14127_, _37115_);
  nand _86862_ (_37117_, _11080_, _14131_);
  and _86863_ (_37118_, _37117_, _14133_);
  or _86864_ (_37119_, _37118_, _06433_);
  or _86865_ (_37120_, _37119_, _37116_);
  or _86866_ (_37122_, _37120_, _37114_);
  or _86867_ (_37123_, _36949_, _06829_);
  and _86868_ (_37124_, _37123_, _05749_);
  and _86869_ (_37125_, _37124_, _37122_);
  and _86870_ (_37126_, _36944_, _05748_);
  or _86871_ (_37127_, _37126_, _06440_);
  or _86872_ (_37128_, _37127_, _37125_);
  and _86873_ (_37129_, _14710_, _07794_);
  or _86874_ (_37130_, _36914_, _06444_);
  or _86875_ (_37131_, _37130_, _37129_);
  and _86876_ (_37133_, _37131_, _01317_);
  and _86877_ (_37134_, _37133_, _37128_);
  or _86878_ (_37135_, _37134_, _36881_);
  and _86879_ (_43781_, _37135_, _43100_);
  and _86880_ (_37136_, _01321_, \oc8051_golden_model_1.PSW [3]);
  and _86881_ (_37137_, _14076_, \oc8051_golden_model_1.PSW [3]);
  and _86882_ (_37138_, _07794_, _07544_);
  or _86883_ (_37139_, _37138_, _37137_);
  or _86884_ (_37140_, _37139_, _06132_);
  and _86885_ (_37141_, _14738_, _07794_);
  or _86886_ (_37143_, _37141_, _37137_);
  or _86887_ (_37144_, _37143_, _06161_);
  and _86888_ (_37145_, _07794_, \oc8051_golden_model_1.ACC [3]);
  or _86889_ (_37146_, _37145_, _37137_);
  and _86890_ (_37147_, _37146_, _07056_);
  and _86891_ (_37148_, _07057_, \oc8051_golden_model_1.PSW [3]);
  or _86892_ (_37149_, _37148_, _06160_);
  or _86893_ (_37150_, _37149_, _37147_);
  and _86894_ (_37151_, _37150_, _06157_);
  and _86895_ (_37152_, _37151_, _37144_);
  and _86896_ (_37154_, _36941_, \oc8051_golden_model_1.PSW [3]);
  and _86897_ (_37155_, _14735_, _08404_);
  or _86898_ (_37156_, _37155_, _37154_);
  and _86899_ (_37157_, _37156_, _06156_);
  or _86900_ (_37158_, _37157_, _06217_);
  or _86901_ (_37159_, _37158_, _37152_);
  or _86902_ (_37160_, _37139_, _07075_);
  and _86903_ (_37161_, _37160_, _37159_);
  or _86904_ (_37162_, _37161_, _06220_);
  or _86905_ (_37163_, _37146_, _06229_);
  and _86906_ (_37165_, _37163_, _06153_);
  and _86907_ (_37166_, _37165_, _37162_);
  and _86908_ (_37167_, _14731_, _08404_);
  or _86909_ (_37168_, _37167_, _37154_);
  and _86910_ (_37169_, _37168_, _06152_);
  or _86911_ (_37170_, _37169_, _06145_);
  or _86912_ (_37171_, _37170_, _37166_);
  or _86913_ (_37172_, _37154_, _14764_);
  and _86914_ (_37173_, _37172_, _37156_);
  or _86915_ (_37174_, _37173_, _06146_);
  and _86916_ (_37176_, _37174_, _06140_);
  and _86917_ (_37177_, _37176_, _37171_);
  and _86918_ (_37178_, _14732_, _08404_);
  or _86919_ (_37179_, _37178_, _37154_);
  and _86920_ (_37180_, _37179_, _06139_);
  or _86921_ (_37181_, _37180_, _09842_);
  or _86922_ (_37182_, _37181_, _37177_);
  and _86923_ (_37183_, _37182_, _37140_);
  or _86924_ (_37184_, _37183_, _06116_);
  and _86925_ (_37185_, _09210_, _07794_);
  or _86926_ (_37187_, _37137_, _06117_);
  or _86927_ (_37188_, _37187_, _37185_);
  and _86928_ (_37189_, _37188_, _06114_);
  and _86929_ (_37190_, _37189_, _37184_);
  and _86930_ (_37191_, _14825_, _07794_);
  or _86931_ (_37192_, _37137_, _37191_);
  and _86932_ (_37193_, _37192_, _05787_);
  or _86933_ (_37194_, _37193_, _37190_);
  or _86934_ (_37195_, _37194_, _11136_);
  and _86935_ (_37196_, _14727_, _07794_);
  or _86936_ (_37198_, _37137_, _07127_);
  or _86937_ (_37199_, _37198_, _37196_);
  and _86938_ (_37200_, _07794_, _08712_);
  or _86939_ (_37201_, _37200_, _37137_);
  or _86940_ (_37202_, _37201_, _06111_);
  and _86941_ (_37203_, _37202_, _07125_);
  and _86942_ (_37204_, _37203_, _37199_);
  and _86943_ (_37205_, _37204_, _37195_);
  and _86944_ (_37206_, _12318_, _07794_);
  or _86945_ (_37207_, _37206_, _37137_);
  and _86946_ (_37209_, _37207_, _06402_);
  or _86947_ (_37210_, _37209_, _37205_);
  and _86948_ (_37211_, _37210_, _07132_);
  or _86949_ (_37212_, _37137_, _08140_);
  and _86950_ (_37213_, _37201_, _06306_);
  and _86951_ (_37214_, _37213_, _37212_);
  or _86952_ (_37215_, _37214_, _37211_);
  and _86953_ (_37216_, _37215_, _07130_);
  and _86954_ (_37217_, _37146_, _06411_);
  and _86955_ (_37218_, _37217_, _37212_);
  or _86956_ (_37220_, _37218_, _06303_);
  or _86957_ (_37221_, _37220_, _37216_);
  and _86958_ (_37222_, _14724_, _07794_);
  or _86959_ (_37223_, _37137_, _08819_);
  or _86960_ (_37224_, _37223_, _37222_);
  and _86961_ (_37225_, _37224_, _08824_);
  and _86962_ (_37226_, _37225_, _37221_);
  nor _86963_ (_37227_, _10273_, _14076_);
  or _86964_ (_37228_, _37227_, _37137_);
  and _86965_ (_37229_, _37228_, _06396_);
  or _86966_ (_37231_, _37229_, _06433_);
  or _86967_ (_37232_, _37231_, _37226_);
  or _86968_ (_37233_, _37143_, _06829_);
  and _86969_ (_37234_, _37233_, _05749_);
  and _86970_ (_37235_, _37234_, _37232_);
  and _86971_ (_37236_, _37168_, _05748_);
  or _86972_ (_37237_, _37236_, _06440_);
  or _86973_ (_37238_, _37237_, _37235_);
  and _86974_ (_37239_, _14897_, _07794_);
  or _86975_ (_37240_, _37137_, _06444_);
  or _86976_ (_37242_, _37240_, _37239_);
  and _86977_ (_37243_, _37242_, _01317_);
  and _86978_ (_37244_, _37243_, _37238_);
  or _86979_ (_37245_, _37244_, _37136_);
  and _86980_ (_43783_, _37245_, _43100_);
  and _86981_ (_37246_, _01321_, \oc8051_golden_model_1.PSW [4]);
  and _86982_ (_37247_, _06284_, _05781_);
  and _86983_ (_37248_, _14076_, \oc8051_golden_model_1.PSW [4]);
  and _86984_ (_37249_, _08336_, _07794_);
  or _86985_ (_37250_, _37249_, _37248_);
  or _86986_ (_37252_, _37250_, _06132_);
  and _86987_ (_37253_, _14928_, _07794_);
  or _86988_ (_37254_, _37253_, _37248_);
  or _86989_ (_37255_, _37254_, _06161_);
  and _86990_ (_37256_, _07794_, \oc8051_golden_model_1.ACC [4]);
  or _86991_ (_37257_, _37256_, _37248_);
  and _86992_ (_37258_, _37257_, _07056_);
  and _86993_ (_37259_, _07057_, \oc8051_golden_model_1.PSW [4]);
  or _86994_ (_37260_, _37259_, _06160_);
  or _86995_ (_37261_, _37260_, _37258_);
  and _86996_ (_37263_, _37261_, _06157_);
  and _86997_ (_37264_, _37263_, _37255_);
  and _86998_ (_37265_, _36941_, \oc8051_golden_model_1.PSW [4]);
  and _86999_ (_37266_, _14932_, _08404_);
  or _87000_ (_37267_, _37266_, _37265_);
  and _87001_ (_37268_, _37267_, _06156_);
  or _87002_ (_37269_, _37268_, _06217_);
  or _87003_ (_37270_, _37269_, _37264_);
  or _87004_ (_37271_, _37250_, _07075_);
  and _87005_ (_37272_, _37271_, _37270_);
  or _87006_ (_37274_, _37272_, _06220_);
  or _87007_ (_37275_, _37257_, _06229_);
  and _87008_ (_37276_, _37275_, _06153_);
  and _87009_ (_37277_, _37276_, _37274_);
  and _87010_ (_37278_, _14942_, _08404_);
  or _87011_ (_37279_, _37278_, _37265_);
  and _87012_ (_37280_, _37279_, _06152_);
  or _87013_ (_37281_, _37280_, _06145_);
  or _87014_ (_37282_, _37281_, _37277_);
  or _87015_ (_37283_, _37265_, _14949_);
  and _87016_ (_37285_, _37283_, _37267_);
  or _87017_ (_37286_, _37285_, _06146_);
  and _87018_ (_37287_, _37286_, _06140_);
  and _87019_ (_37288_, _37287_, _37282_);
  and _87020_ (_37289_, _14966_, _08404_);
  or _87021_ (_37290_, _37289_, _37265_);
  and _87022_ (_37291_, _37290_, _06139_);
  or _87023_ (_37292_, _37291_, _09842_);
  or _87024_ (_37293_, _37292_, _37288_);
  and _87025_ (_37294_, _37293_, _37252_);
  or _87026_ (_37296_, _37294_, _37247_);
  and _87027_ (_37297_, _09209_, _07794_);
  or _87028_ (_37298_, _37297_, _37248_);
  and _87029_ (_37299_, _37298_, _06276_);
  or _87030_ (_37300_, _37299_, _06117_);
  and _87031_ (_37301_, _37300_, _37296_);
  and _87032_ (_37302_, _06281_, _05781_);
  and _87033_ (_37303_, _37298_, _37302_);
  or _87034_ (_37304_, _37303_, _05787_);
  or _87035_ (_37305_, _37304_, _37301_);
  and _87036_ (_37307_, _15013_, _07794_);
  or _87037_ (_37308_, _37248_, _06114_);
  or _87038_ (_37309_, _37308_, _37307_);
  and _87039_ (_37310_, _37309_, _06111_);
  and _87040_ (_37311_, _37310_, _37305_);
  and _87041_ (_37312_, _08715_, _07794_);
  or _87042_ (_37313_, _37312_, _37248_);
  and _87043_ (_37314_, _37313_, _06110_);
  or _87044_ (_37315_, _37314_, _06297_);
  or _87045_ (_37316_, _37315_, _37311_);
  and _87046_ (_37318_, _15029_, _07794_);
  or _87047_ (_37319_, _37248_, _07127_);
  or _87048_ (_37320_, _37319_, _37318_);
  and _87049_ (_37321_, _37320_, _07125_);
  and _87050_ (_37322_, _37321_, _37316_);
  and _87051_ (_37323_, _10289_, _07794_);
  or _87052_ (_37324_, _37323_, _37248_);
  and _87053_ (_37325_, _37324_, _06402_);
  or _87054_ (_37326_, _37325_, _37322_);
  and _87055_ (_37327_, _37326_, _07132_);
  or _87056_ (_37329_, _37248_, _08339_);
  and _87057_ (_37330_, _37313_, _06306_);
  and _87058_ (_37331_, _37330_, _37329_);
  or _87059_ (_37332_, _37331_, _37327_);
  and _87060_ (_37333_, _37332_, _07130_);
  and _87061_ (_37334_, _37257_, _06411_);
  and _87062_ (_37335_, _37334_, _37329_);
  or _87063_ (_37336_, _37335_, _06303_);
  or _87064_ (_37337_, _37336_, _37333_);
  and _87065_ (_37338_, _15026_, _07794_);
  or _87066_ (_37340_, _37248_, _08819_);
  or _87067_ (_37341_, _37340_, _37338_);
  and _87068_ (_37342_, _37341_, _08824_);
  and _87069_ (_37343_, _37342_, _37337_);
  nor _87070_ (_37344_, _10288_, _14076_);
  or _87071_ (_37345_, _37344_, _37248_);
  and _87072_ (_37346_, _37345_, _06396_);
  or _87073_ (_37347_, _37346_, _06433_);
  or _87074_ (_37348_, _37347_, _37343_);
  or _87075_ (_37349_, _37254_, _06829_);
  and _87076_ (_37351_, _37349_, _05749_);
  and _87077_ (_37352_, _37351_, _37348_);
  and _87078_ (_37353_, _37279_, _05748_);
  or _87079_ (_37354_, _37353_, _06440_);
  or _87080_ (_37355_, _37354_, _37352_);
  and _87081_ (_37356_, _15087_, _07794_);
  or _87082_ (_37357_, _37248_, _06444_);
  or _87083_ (_37358_, _37357_, _37356_);
  and _87084_ (_37359_, _37358_, _01317_);
  and _87085_ (_37360_, _37359_, _37355_);
  or _87086_ (_37362_, _37360_, _37246_);
  and _87087_ (_43784_, _37362_, _43100_);
  and _87088_ (_37363_, _01321_, \oc8051_golden_model_1.PSW [5]);
  and _87089_ (_37364_, _14076_, \oc8051_golden_model_1.PSW [5]);
  and _87090_ (_37365_, _15119_, _07794_);
  or _87091_ (_37366_, _37365_, _37364_);
  or _87092_ (_37367_, _37366_, _06161_);
  and _87093_ (_37368_, _07794_, \oc8051_golden_model_1.ACC [5]);
  or _87094_ (_37369_, _37368_, _37364_);
  and _87095_ (_37370_, _37369_, _07056_);
  and _87096_ (_37372_, _07057_, \oc8051_golden_model_1.PSW [5]);
  or _87097_ (_37373_, _37372_, _06160_);
  or _87098_ (_37374_, _37373_, _37370_);
  and _87099_ (_37375_, _37374_, _06157_);
  and _87100_ (_37376_, _37375_, _37367_);
  and _87101_ (_37377_, _36941_, \oc8051_golden_model_1.PSW [5]);
  and _87102_ (_37378_, _15123_, _08404_);
  or _87103_ (_37379_, _37378_, _37377_);
  and _87104_ (_37380_, _37379_, _06156_);
  or _87105_ (_37381_, _37380_, _06217_);
  or _87106_ (_37383_, _37381_, _37376_);
  and _87107_ (_37384_, _08101_, _07794_);
  or _87108_ (_37385_, _37384_, _37364_);
  or _87109_ (_37386_, _37385_, _07075_);
  and _87110_ (_37387_, _37386_, _37383_);
  or _87111_ (_37388_, _37387_, _06220_);
  or _87112_ (_37389_, _37369_, _06229_);
  and _87113_ (_37390_, _37389_, _06153_);
  and _87114_ (_37391_, _37390_, _37388_);
  and _87115_ (_37392_, _15104_, _08404_);
  or _87116_ (_37394_, _37392_, _37377_);
  and _87117_ (_37395_, _37394_, _06152_);
  or _87118_ (_37396_, _37395_, _06145_);
  or _87119_ (_37397_, _37396_, _37391_);
  or _87120_ (_37398_, _37377_, _15138_);
  and _87121_ (_37399_, _37398_, _37379_);
  or _87122_ (_37400_, _37399_, _06146_);
  and _87123_ (_37401_, _37400_, _06140_);
  and _87124_ (_37402_, _37401_, _37397_);
  and _87125_ (_37403_, _15155_, _08404_);
  or _87126_ (_37405_, _37403_, _37377_);
  and _87127_ (_37406_, _37405_, _06139_);
  or _87128_ (_37407_, _37406_, _09842_);
  or _87129_ (_37408_, _37407_, _37402_);
  or _87130_ (_37409_, _37385_, _06132_);
  and _87131_ (_37410_, _37409_, _37408_);
  or _87132_ (_37411_, _37410_, _06116_);
  and _87133_ (_37412_, _09208_, _07794_);
  or _87134_ (_37413_, _37364_, _06117_);
  or _87135_ (_37414_, _37413_, _37412_);
  and _87136_ (_37416_, _37414_, _06114_);
  and _87137_ (_37417_, _37416_, _37411_);
  and _87138_ (_37418_, _15203_, _07794_);
  or _87139_ (_37419_, _37418_, _37364_);
  and _87140_ (_37420_, _37419_, _05787_);
  or _87141_ (_37421_, _37420_, _11136_);
  or _87142_ (_37422_, _37421_, _37417_);
  and _87143_ (_37423_, _15219_, _07794_);
  or _87144_ (_37424_, _37364_, _07127_);
  or _87145_ (_37425_, _37424_, _37423_);
  and _87146_ (_37427_, _08736_, _07794_);
  or _87147_ (_37428_, _37427_, _37364_);
  or _87148_ (_37429_, _37428_, _06111_);
  and _87149_ (_37430_, _37429_, _07125_);
  and _87150_ (_37431_, _37430_, _37425_);
  and _87151_ (_37432_, _37431_, _37422_);
  and _87152_ (_37433_, _12325_, _07794_);
  or _87153_ (_37434_, _37433_, _37364_);
  and _87154_ (_37435_, _37434_, _06402_);
  or _87155_ (_37436_, _37435_, _37432_);
  and _87156_ (_37438_, _37436_, _07132_);
  or _87157_ (_37439_, _37364_, _08104_);
  and _87158_ (_37440_, _37428_, _06306_);
  and _87159_ (_37441_, _37440_, _37439_);
  or _87160_ (_37442_, _37441_, _37438_);
  and _87161_ (_37443_, _37442_, _07130_);
  and _87162_ (_37444_, _37369_, _06411_);
  and _87163_ (_37445_, _37444_, _37439_);
  or _87164_ (_37446_, _37445_, _06303_);
  or _87165_ (_37447_, _37446_, _37443_);
  and _87166_ (_37449_, _15216_, _07794_);
  or _87167_ (_37450_, _37364_, _08819_);
  or _87168_ (_37451_, _37450_, _37449_);
  and _87169_ (_37452_, _37451_, _08824_);
  and _87170_ (_37453_, _37452_, _37447_);
  nor _87171_ (_37454_, _10269_, _14076_);
  or _87172_ (_37455_, _37454_, _37364_);
  and _87173_ (_37456_, _37455_, _06396_);
  or _87174_ (_37457_, _37456_, _06433_);
  or _87175_ (_37458_, _37457_, _37453_);
  or _87176_ (_37460_, _37366_, _06829_);
  and _87177_ (_37461_, _37460_, _05749_);
  and _87178_ (_37462_, _37461_, _37458_);
  and _87179_ (_37463_, _37394_, _05748_);
  or _87180_ (_37464_, _37463_, _06440_);
  or _87181_ (_37465_, _37464_, _37462_);
  and _87182_ (_37466_, _15275_, _07794_);
  or _87183_ (_37467_, _37364_, _06444_);
  or _87184_ (_37468_, _37467_, _37466_);
  and _87185_ (_37469_, _37468_, _01317_);
  and _87186_ (_37471_, _37469_, _37465_);
  or _87187_ (_37472_, _37471_, _37363_);
  and _87188_ (_43785_, _37472_, _43100_);
  nor _87189_ (_37473_, _01317_, _17884_);
  or _87190_ (_37474_, _10942_, _10654_);
  and _87191_ (_37475_, _37474_, _10895_);
  nor _87192_ (_37476_, _10882_, _10601_);
  nand _87193_ (_37477_, _37476_, _17240_);
  not _87194_ (_37478_, _10372_);
  or _87195_ (_37479_, _10361_, _10324_);
  and _87196_ (_37481_, _37479_, _37478_);
  and _87197_ (_37482_, _15410_, _07794_);
  nor _87198_ (_37483_, _07794_, _17884_);
  or _87199_ (_37484_, _37483_, _08819_);
  or _87200_ (_37485_, _37484_, _37482_);
  and _87201_ (_37486_, _08012_, _07794_);
  or _87202_ (_37487_, _37486_, _37483_);
  or _87203_ (_37488_, _37487_, _06132_);
  or _87204_ (_37489_, _10634_, _10601_);
  or _87205_ (_37490_, _37489_, _12380_);
  nor _87206_ (_37492_, _08404_, _17884_);
  and _87207_ (_37493_, _15297_, _08404_);
  or _87208_ (_37494_, _37493_, _37492_);
  and _87209_ (_37495_, _37494_, _06152_);
  and _87210_ (_37496_, _15300_, _07794_);
  or _87211_ (_37497_, _37496_, _37483_);
  or _87212_ (_37498_, _37497_, _06161_);
  and _87213_ (_37499_, _07794_, \oc8051_golden_model_1.ACC [6]);
  or _87214_ (_37500_, _37499_, _37483_);
  and _87215_ (_37501_, _37500_, _07056_);
  nor _87216_ (_37503_, _07056_, _17884_);
  or _87217_ (_37504_, _37503_, _06160_);
  or _87218_ (_37505_, _37504_, _37501_);
  and _87219_ (_37506_, _37505_, _06157_);
  and _87220_ (_37507_, _37506_, _37498_);
  and _87221_ (_37508_, _15316_, _08404_);
  or _87222_ (_37509_, _37508_, _37492_);
  and _87223_ (_37510_, _37509_, _06156_);
  or _87224_ (_37511_, _37510_, _06217_);
  or _87225_ (_37512_, _37511_, _37507_);
  or _87226_ (_37514_, _37487_, _07075_);
  and _87227_ (_37515_, _37514_, _37512_);
  or _87228_ (_37516_, _37515_, _06220_);
  or _87229_ (_37517_, _37500_, _06229_);
  and _87230_ (_37518_, _37517_, _06153_);
  and _87231_ (_37519_, _37518_, _37516_);
  or _87232_ (_37520_, _37519_, _37495_);
  and _87233_ (_37521_, _37520_, _06146_);
  or _87234_ (_37522_, _37492_, _15331_);
  and _87235_ (_37523_, _37522_, _06145_);
  and _87236_ (_37525_, _37523_, _37509_);
  or _87237_ (_37526_, _37525_, _10557_);
  or _87238_ (_37527_, _37526_, _37521_);
  or _87239_ (_37528_, _10554_, _10324_);
  or _87240_ (_37529_, _37528_, _10568_);
  and _87241_ (_37530_, _37529_, _37527_);
  or _87242_ (_37531_, _37530_, _12379_);
  and _87243_ (_37532_, _37531_, _37490_);
  and _87244_ (_37533_, _37532_, _06265_);
  or _87245_ (_37534_, _10441_, _10392_);
  and _87246_ (_37536_, _37534_, _06260_);
  or _87247_ (_37537_, _37536_, _10387_);
  or _87248_ (_37538_, _37537_, _37533_);
  or _87249_ (_37539_, _10654_, _10388_);
  or _87250_ (_37540_, _37539_, _10708_);
  and _87251_ (_37541_, _37540_, _06140_);
  and _87252_ (_37542_, _37541_, _37538_);
  and _87253_ (_37543_, _15348_, _08404_);
  or _87254_ (_37544_, _37543_, _37492_);
  and _87255_ (_37545_, _37544_, _06139_);
  or _87256_ (_37547_, _37545_, _09842_);
  or _87257_ (_37548_, _37547_, _37542_);
  and _87258_ (_37549_, _37548_, _37488_);
  or _87259_ (_37550_, _37549_, _06116_);
  and _87260_ (_37551_, _09207_, _07794_);
  or _87261_ (_37552_, _37483_, _06117_);
  or _87262_ (_37553_, _37552_, _37551_);
  and _87263_ (_37554_, _37553_, _06114_);
  and _87264_ (_37555_, _37554_, _37550_);
  and _87265_ (_37556_, _15395_, _07794_);
  or _87266_ (_37558_, _37556_, _37483_);
  and _87267_ (_37559_, _37558_, _05787_);
  or _87268_ (_37560_, _37559_, _11136_);
  or _87269_ (_37561_, _37560_, _37555_);
  and _87270_ (_37562_, _15413_, _07794_);
  or _87271_ (_37563_, _37483_, _07127_);
  or _87272_ (_37564_, _37563_, _37562_);
  and _87273_ (_37565_, _15402_, _07794_);
  or _87274_ (_37566_, _37565_, _37483_);
  or _87275_ (_37567_, _37566_, _06111_);
  and _87276_ (_37569_, _37567_, _07125_);
  and _87277_ (_37570_, _37569_, _37564_);
  and _87278_ (_37571_, _37570_, _37561_);
  and _87279_ (_37572_, _10295_, _07794_);
  or _87280_ (_37573_, _37572_, _37483_);
  and _87281_ (_37574_, _37573_, _06402_);
  or _87282_ (_37575_, _37574_, _37571_);
  and _87283_ (_37576_, _37575_, _07132_);
  or _87284_ (_37577_, _37483_, _08015_);
  and _87285_ (_37578_, _37566_, _06306_);
  and _87286_ (_37580_, _37578_, _37577_);
  or _87287_ (_37581_, _37580_, _37576_);
  and _87288_ (_37582_, _37581_, _07130_);
  and _87289_ (_37583_, _37500_, _06411_);
  and _87290_ (_37584_, _37583_, _37577_);
  or _87291_ (_37585_, _37584_, _06303_);
  or _87292_ (_37586_, _37585_, _37582_);
  and _87293_ (_37587_, _37586_, _37485_);
  or _87294_ (_37588_, _37587_, _06396_);
  nor _87295_ (_37589_, _10294_, _14076_);
  or _87296_ (_37591_, _37589_, _37483_);
  or _87297_ (_37592_, _37591_, _08824_);
  and _87298_ (_37593_, _37592_, _10372_);
  and _87299_ (_37594_, _37593_, _37588_);
  or _87300_ (_37595_, _37594_, _37481_);
  and _87301_ (_37596_, _37595_, _10375_);
  and _87302_ (_37597_, _37479_, _06794_);
  nor _87303_ (_37598_, _37597_, _37596_);
  nor _87304_ (_37599_, _37598_, _10376_);
  and _87305_ (_37600_, _37479_, _10376_);
  or _87306_ (_37602_, _37600_, _06795_);
  or _87307_ (_37603_, _37602_, _37599_);
  not _87308_ (_37604_, _06795_);
  or _87309_ (_37605_, _37479_, _37604_);
  and _87310_ (_37606_, _37605_, _10374_);
  and _87311_ (_37607_, _37606_, _37603_);
  and _87312_ (_37608_, _37479_, _10373_);
  or _87313_ (_37609_, _37608_, _37607_);
  or _87314_ (_37610_, _37609_, _17240_);
  and _87315_ (_37611_, _37610_, _37477_);
  or _87316_ (_37613_, _37611_, _06792_);
  nand _87317_ (_37614_, _37476_, _06792_);
  and _87318_ (_37615_, _37614_, _37613_);
  or _87319_ (_37616_, _37615_, _06406_);
  nor _87320_ (_37617_, _10901_, _10392_);
  nand _87321_ (_37618_, _37617_, _18090_);
  and _87322_ (_37619_, _37618_, _10927_);
  and _87323_ (_37620_, _37619_, _37616_);
  or _87324_ (_37621_, _37620_, _37475_);
  and _87325_ (_37622_, _37621_, _10963_);
  and _87326_ (_37624_, _10991_, _18454_);
  or _87327_ (_37625_, _37624_, _11003_);
  or _87328_ (_37626_, _37625_, _37622_);
  or _87329_ (_37627_, _11033_, _11041_);
  and _87330_ (_37628_, _37627_, _06171_);
  and _87331_ (_37629_, _37628_, _37626_);
  and _87332_ (_37630_, _10287_, _06169_);
  or _87333_ (_37631_, _37630_, _10264_);
  or _87334_ (_37632_, _37631_, _37629_);
  or _87335_ (_37633_, _11074_, _10265_);
  and _87336_ (_37635_, _37633_, _37632_);
  or _87337_ (_37636_, _37635_, _06433_);
  or _87338_ (_37637_, _37497_, _06829_);
  and _87339_ (_37638_, _37637_, _05749_);
  and _87340_ (_37639_, _37638_, _37636_);
  and _87341_ (_37640_, _37494_, _05748_);
  or _87342_ (_37641_, _37640_, _06440_);
  or _87343_ (_37642_, _37641_, _37639_);
  and _87344_ (_37643_, _15478_, _07794_);
  or _87345_ (_37644_, _37483_, _06444_);
  or _87346_ (_37646_, _37644_, _37643_);
  and _87347_ (_37647_, _37646_, _01317_);
  and _87348_ (_37648_, _37647_, _37642_);
  or _87349_ (_37649_, _37648_, _37473_);
  and _87350_ (_43786_, _37649_, _43100_);
  and _87351_ (_37650_, _05820_, op0_cnst);
  or _87352_ (_00001_, _37650_, rst);
  and _87353_ (_37651_, inst_finished_r, op0_cnst);
  not _87354_ (_37652_, word_in[1]);
  and _87355_ (_37653_, _37652_, word_in[0]);
  and _87356_ (_37655_, _37653_, \oc8051_golden_model_1.IRAM[1] [3]);
  nor _87357_ (_37656_, _37652_, word_in[0]);
  and _87358_ (_37657_, _37656_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor _87359_ (_37658_, _37657_, _37655_);
  nor _87360_ (_37659_, word_in[1], word_in[0]);
  and _87361_ (_37660_, _37659_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _87362_ (_37661_, word_in[1], word_in[0]);
  and _87363_ (_37662_, _37661_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor _87364_ (_37663_, _37662_, _37660_);
  and _87365_ (_37664_, _37663_, _37658_);
  nor _87366_ (_37666_, word_in[3], word_in[2]);
  not _87367_ (_37667_, _37666_);
  nor _87368_ (_37668_, _37667_, _37664_);
  and _87369_ (_37669_, _37653_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _87370_ (_37670_, _37656_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor _87371_ (_37671_, _37670_, _37669_);
  and _87372_ (_37672_, _37659_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _87373_ (_37673_, _37661_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor _87374_ (_37674_, _37673_, _37672_);
  and _87375_ (_37675_, _37674_, _37671_);
  and _87376_ (_37677_, word_in[3], word_in[2]);
  not _87377_ (_37678_, _37677_);
  nor _87378_ (_37679_, _37678_, _37675_);
  nor _87379_ (_37680_, _37679_, _37668_);
  and _87380_ (_37681_, _37653_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _87381_ (_37682_, _37656_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor _87382_ (_37683_, _37682_, _37681_);
  and _87383_ (_37684_, _37659_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _87384_ (_37685_, _37661_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor _87385_ (_37686_, _37685_, _37684_);
  and _87386_ (_37688_, _37686_, _37683_);
  not _87387_ (_37689_, word_in[3]);
  and _87388_ (_37690_, _37689_, word_in[2]);
  not _87389_ (_37691_, _37690_);
  nor _87390_ (_37692_, _37691_, _37688_);
  and _87391_ (_37693_, _37653_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _87392_ (_37694_, _37656_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor _87393_ (_37695_, _37694_, _37693_);
  and _87394_ (_37696_, _37659_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _87395_ (_37697_, _37661_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor _87396_ (_37699_, _37697_, _37696_);
  and _87397_ (_37700_, _37699_, _37695_);
  nor _87398_ (_37701_, _37689_, word_in[2]);
  not _87399_ (_37702_, _37701_);
  nor _87400_ (_37703_, _37702_, _37700_);
  nor _87401_ (_37704_, _37703_, _37692_);
  and _87402_ (_37705_, _37704_, _37680_);
  and _87403_ (_37706_, _37690_, _37661_);
  and _87404_ (_37707_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and _87405_ (_37708_, _37666_, _37661_);
  and _87406_ (_37710_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _87407_ (_37711_, _37710_, _37707_);
  and _87408_ (_37712_, _37677_, _37656_);
  and _87409_ (_37713_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and _87410_ (_37714_, _37677_, _37659_);
  and _87411_ (_37715_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _87412_ (_37716_, _37715_, _37713_);
  and _87413_ (_37717_, _37716_, _37711_);
  and _87414_ (_37718_, _37666_, _37656_);
  and _87415_ (_37719_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and _87416_ (_37721_, _37666_, _37653_);
  and _87417_ (_37722_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _87418_ (_37723_, _37722_, _37719_);
  and _87419_ (_37724_, _37690_, _37653_);
  and _87420_ (_37725_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and _87421_ (_37726_, _37690_, _37659_);
  and _87422_ (_37727_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _87423_ (_37728_, _37727_, _37725_);
  and _87424_ (_37729_, _37728_, _37723_);
  and _87425_ (_37730_, _37729_, _37717_);
  and _87426_ (_37732_, _37701_, _37656_);
  and _87427_ (_37733_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and _87428_ (_37734_, _37701_, _37659_);
  and _87429_ (_37735_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _87430_ (_37736_, _37735_, _37733_);
  and _87431_ (_37737_, _37677_, _37661_);
  and _87432_ (_37738_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _87433_ (_37739_, _37677_, _37653_);
  and _87434_ (_37740_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor _87435_ (_37741_, _37740_, _37738_);
  and _87436_ (_37743_, _37741_, _37736_);
  and _87437_ (_37744_, _37690_, _37656_);
  and _87438_ (_37745_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _87439_ (_37746_, _37666_, _37659_);
  and _87440_ (_37747_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _87441_ (_37748_, _37747_, _37745_);
  and _87442_ (_37749_, _37701_, _37661_);
  and _87443_ (_37750_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _87444_ (_37751_, _37701_, _37653_);
  and _87445_ (_37752_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor _87446_ (_37754_, _37752_, _37750_);
  and _87447_ (_37755_, _37754_, _37748_);
  and _87448_ (_37756_, _37755_, _37743_);
  and _87449_ (_37757_, _37756_, _37730_);
  nand _87450_ (_37758_, _37757_, _37705_);
  or _87451_ (_37759_, _37757_, _37705_);
  and _87452_ (_37760_, _37759_, _37758_);
  and _87453_ (_37761_, _37653_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _87454_ (_37762_, _37656_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor _87455_ (_37763_, _37762_, _37761_);
  and _87456_ (_37765_, _37659_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _87457_ (_37766_, _37661_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor _87458_ (_37767_, _37766_, _37765_);
  and _87459_ (_37768_, _37767_, _37763_);
  nor _87460_ (_37769_, _37768_, _37667_);
  and _87461_ (_37770_, _37653_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _87462_ (_37771_, _37656_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor _87463_ (_37772_, _37771_, _37770_);
  and _87464_ (_37773_, _37659_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _87465_ (_37774_, _37661_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor _87466_ (_37776_, _37774_, _37773_);
  and _87467_ (_37777_, _37776_, _37772_);
  nor _87468_ (_37778_, _37777_, _37678_);
  nor _87469_ (_37779_, _37778_, _37769_);
  and _87470_ (_37780_, _37653_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _87471_ (_37781_, _37656_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor _87472_ (_37782_, _37781_, _37780_);
  and _87473_ (_37783_, _37659_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _87474_ (_37784_, _37661_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor _87475_ (_37785_, _37784_, _37783_);
  and _87476_ (_37787_, _37785_, _37782_);
  nor _87477_ (_37788_, _37787_, _37691_);
  and _87478_ (_37789_, _37653_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _87479_ (_37790_, _37656_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor _87480_ (_37791_, _37790_, _37789_);
  and _87481_ (_37792_, _37659_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _87482_ (_37793_, _37661_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor _87483_ (_37794_, _37793_, _37792_);
  and _87484_ (_37795_, _37794_, _37791_);
  nor _87485_ (_37796_, _37795_, _37702_);
  nor _87486_ (_37798_, _37796_, _37788_);
  and _87487_ (_37799_, _37798_, _37779_);
  and _87488_ (_37800_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _87489_ (_37801_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor _87490_ (_37802_, _37801_, _37800_);
  and _87491_ (_37803_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and _87492_ (_37804_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor _87493_ (_37805_, _37804_, _37803_);
  and _87494_ (_37806_, _37805_, _37802_);
  and _87495_ (_37807_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _87496_ (_37809_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _87497_ (_37810_, _37809_, _37807_);
  and _87498_ (_37811_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _87499_ (_37812_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _87500_ (_37813_, _37812_, _37811_);
  and _87501_ (_37814_, _37813_, _37810_);
  and _87502_ (_37815_, _37814_, _37806_);
  and _87503_ (_37816_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and _87504_ (_37817_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _87505_ (_37818_, _37817_, _37816_);
  and _87506_ (_37820_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _87507_ (_37821_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _87508_ (_37822_, _37821_, _37820_);
  and _87509_ (_37823_, _37822_, _37818_);
  and _87510_ (_37824_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and _87511_ (_37825_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _87512_ (_37826_, _37825_, _37824_);
  and _87513_ (_37827_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _87514_ (_37828_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _87515_ (_37829_, _37828_, _37827_);
  and _87516_ (_37831_, _37829_, _37826_);
  and _87517_ (_37832_, _37831_, _37823_);
  and _87518_ (_37833_, _37832_, _37815_);
  nand _87519_ (_37834_, _37833_, _37799_);
  or _87520_ (_37835_, _37833_, _37799_);
  and _87521_ (_37836_, _37835_, _37834_);
  or _87522_ (_37837_, _37836_, _37760_);
  and _87523_ (_37838_, _37653_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _87524_ (_37839_, _37656_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor _87525_ (_37840_, _37839_, _37838_);
  and _87526_ (_37842_, _37659_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _87527_ (_37843_, _37661_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor _87528_ (_37844_, _37843_, _37842_);
  and _87529_ (_37845_, _37844_, _37840_);
  nor _87530_ (_37846_, _37845_, _37691_);
  and _87531_ (_37847_, _37653_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _87532_ (_37848_, _37656_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor _87533_ (_37849_, _37848_, _37847_);
  and _87534_ (_37850_, _37659_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _87535_ (_37851_, _37661_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor _87536_ (_37853_, _37851_, _37850_);
  and _87537_ (_37854_, _37853_, _37849_);
  nor _87538_ (_37855_, _37854_, _37678_);
  nor _87539_ (_37856_, _37855_, _37846_);
  and _87540_ (_37857_, _37653_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _87541_ (_37858_, _37656_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor _87542_ (_37859_, _37858_, _37857_);
  and _87543_ (_37860_, _37659_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _87544_ (_37861_, _37661_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor _87545_ (_37862_, _37861_, _37860_);
  and _87546_ (_37864_, _37862_, _37859_);
  nor _87547_ (_37865_, _37864_, _37667_);
  and _87548_ (_37866_, _37653_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _87549_ (_37867_, _37656_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor _87550_ (_37868_, _37867_, _37866_);
  and _87551_ (_37869_, _37659_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _87552_ (_37870_, _37661_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor _87553_ (_37871_, _37870_, _37869_);
  and _87554_ (_37872_, _37871_, _37868_);
  nor _87555_ (_37873_, _37872_, _37702_);
  nor _87556_ (_37875_, _37873_, _37865_);
  and _87557_ (_37876_, _37875_, _37856_);
  and _87558_ (_37877_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and _87559_ (_37878_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _87560_ (_37879_, _37878_, _37877_);
  and _87561_ (_37880_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _87562_ (_37881_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _87563_ (_37882_, _37881_, _37880_);
  and _87564_ (_37883_, _37882_, _37879_);
  and _87565_ (_37884_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and _87566_ (_37886_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _87567_ (_37887_, _37886_, _37884_);
  and _87568_ (_37888_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and _87569_ (_37889_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _87570_ (_37890_, _37889_, _37888_);
  and _87571_ (_37891_, _37890_, _37887_);
  and _87572_ (_37892_, _37891_, _37883_);
  and _87573_ (_37893_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _87574_ (_37894_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _87575_ (_37895_, _37894_, _37893_);
  and _87576_ (_37897_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and _87577_ (_37898_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor _87578_ (_37899_, _37898_, _37897_);
  and _87579_ (_37900_, _37899_, _37895_);
  and _87580_ (_37901_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _87581_ (_37902_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _87582_ (_37903_, _37902_, _37901_);
  and _87583_ (_37904_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and _87584_ (_37905_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _87585_ (_37906_, _37905_, _37904_);
  and _87586_ (_37908_, _37906_, _37903_);
  and _87587_ (_37909_, _37908_, _37900_);
  and _87588_ (_37910_, _37909_, _37892_);
  nand _87589_ (_37911_, _37910_, _37876_);
  or _87590_ (_37912_, _37910_, _37876_);
  and _87591_ (_37913_, _37912_, _37911_);
  and _87592_ (_37914_, _37653_, \oc8051_golden_model_1.IRAM[1] [0]);
  and _87593_ (_37915_, _37656_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor _87594_ (_37916_, _37915_, _37914_);
  and _87595_ (_37917_, _37659_, \oc8051_golden_model_1.IRAM[0] [0]);
  and _87596_ (_37919_, _37661_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor _87597_ (_37920_, _37919_, _37917_);
  and _87598_ (_37921_, _37920_, _37916_);
  nor _87599_ (_37922_, _37921_, _37667_);
  and _87600_ (_37923_, _37653_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _87601_ (_37924_, _37656_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor _87602_ (_37925_, _37924_, _37923_);
  and _87603_ (_37926_, _37659_, \oc8051_golden_model_1.IRAM[8] [0]);
  and _87604_ (_37927_, _37661_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor _87605_ (_37928_, _37927_, _37926_);
  and _87606_ (_37930_, _37928_, _37925_);
  nor _87607_ (_37931_, _37930_, _37702_);
  nor _87608_ (_37932_, _37931_, _37922_);
  and _87609_ (_37933_, _37653_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _87610_ (_37934_, _37656_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor _87611_ (_37935_, _37934_, _37933_);
  and _87612_ (_37936_, _37659_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _87613_ (_37937_, _37661_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor _87614_ (_37938_, _37937_, _37936_);
  and _87615_ (_37939_, _37938_, _37935_);
  nor _87616_ (_37941_, _37939_, _37691_);
  and _87617_ (_37942_, _37653_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _87618_ (_37943_, _37656_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor _87619_ (_37944_, _37943_, _37942_);
  and _87620_ (_37945_, _37659_, \oc8051_golden_model_1.IRAM[12] [0]);
  and _87621_ (_37946_, _37661_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor _87622_ (_37947_, _37946_, _37945_);
  and _87623_ (_37948_, _37947_, _37944_);
  nor _87624_ (_37949_, _37948_, _37678_);
  nor _87625_ (_37950_, _37949_, _37941_);
  and _87626_ (_37952_, _37950_, _37932_);
  and _87627_ (_37953_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _87628_ (_37954_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _87629_ (_37955_, _37954_, _37953_);
  and _87630_ (_37956_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _87631_ (_37957_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _87632_ (_37958_, _37957_, _37956_);
  and _87633_ (_37959_, _37958_, _37955_);
  and _87634_ (_37960_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and _87635_ (_37961_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _87636_ (_37963_, _37961_, _37960_);
  and _87637_ (_37964_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and _87638_ (_37965_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _87639_ (_37966_, _37965_, _37964_);
  and _87640_ (_37967_, _37966_, _37963_);
  and _87641_ (_37968_, _37967_, _37959_);
  and _87642_ (_37969_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and _87643_ (_37970_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _87644_ (_37971_, _37970_, _37969_);
  and _87645_ (_37972_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and _87646_ (_37974_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor _87647_ (_37975_, _37974_, _37972_);
  and _87648_ (_37976_, _37975_, _37971_);
  and _87649_ (_37977_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _87650_ (_37978_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _87651_ (_37979_, _37978_, _37977_);
  and _87652_ (_37980_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _87653_ (_37981_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _87654_ (_37982_, _37981_, _37980_);
  and _87655_ (_37983_, _37982_, _37979_);
  and _87656_ (_37985_, _37983_, _37976_);
  and _87657_ (_37986_, _37985_, _37968_);
  nand _87658_ (_37987_, _37986_, _37952_);
  or _87659_ (_37988_, _37986_, _37952_);
  and _87660_ (_37989_, _37988_, _37987_);
  or _87661_ (_37990_, _37989_, _37913_);
  or _87662_ (_37991_, _37990_, _37837_);
  and _87663_ (_37992_, _37653_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _87664_ (_37993_, _37656_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor _87665_ (_37994_, _37993_, _37992_);
  and _87666_ (_37996_, _37659_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _87667_ (_37997_, _37661_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor _87668_ (_37998_, _37997_, _37996_);
  and _87669_ (_37999_, _37998_, _37994_);
  nor _87670_ (_38000_, _37999_, _37691_);
  and _87671_ (_38001_, _37653_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _87672_ (_38002_, _37656_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor _87673_ (_38003_, _38002_, _38001_);
  and _87674_ (_38004_, _37659_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _87675_ (_38005_, _37661_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor _87676_ (_38007_, _38005_, _38004_);
  and _87677_ (_38008_, _38007_, _38003_);
  nor _87678_ (_38009_, _38008_, _37678_);
  nor _87679_ (_38010_, _38009_, _38000_);
  and _87680_ (_38011_, _37653_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _87681_ (_38012_, _37656_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor _87682_ (_38013_, _38012_, _38011_);
  and _87683_ (_38014_, _37659_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _87684_ (_38015_, _37661_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor _87685_ (_38016_, _38015_, _38014_);
  and _87686_ (_38018_, _38016_, _38013_);
  nor _87687_ (_38019_, _38018_, _37667_);
  and _87688_ (_38020_, _37653_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _87689_ (_38021_, _37656_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor _87690_ (_38022_, _38021_, _38020_);
  and _87691_ (_38023_, _37659_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _87692_ (_38024_, _37661_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor _87693_ (_38025_, _38024_, _38023_);
  and _87694_ (_38026_, _38025_, _38022_);
  nor _87695_ (_38027_, _38026_, _37702_);
  nor _87696_ (_38029_, _38027_, _38019_);
  and _87697_ (_38030_, _38029_, _38010_);
  and _87698_ (_38031_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _87699_ (_38032_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _87700_ (_38033_, _38032_, _38031_);
  and _87701_ (_38034_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _87702_ (_38035_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _87703_ (_38036_, _38035_, _38034_);
  and _87704_ (_38037_, _38036_, _38033_);
  and _87705_ (_38038_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and _87706_ (_38040_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _87707_ (_38041_, _38040_, _38038_);
  and _87708_ (_38042_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and _87709_ (_38043_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _87710_ (_38044_, _38043_, _38042_);
  and _87711_ (_38045_, _38044_, _38041_);
  and _87712_ (_38046_, _38045_, _38037_);
  and _87713_ (_38047_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and _87714_ (_38048_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _87715_ (_38049_, _38048_, _38047_);
  and _87716_ (_38051_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and _87717_ (_38052_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _87718_ (_38053_, _38052_, _38051_);
  and _87719_ (_38054_, _38053_, _38049_);
  and _87720_ (_38055_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and _87721_ (_38056_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _87722_ (_38057_, _38056_, _38055_);
  and _87723_ (_38058_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and _87724_ (_38059_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _87725_ (_38060_, _38059_, _38058_);
  and _87726_ (_38062_, _38060_, _38057_);
  and _87727_ (_38063_, _38062_, _38054_);
  and _87728_ (_38064_, _38063_, _38046_);
  nand _87729_ (_38065_, _38064_, _38030_);
  or _87730_ (_38066_, _38064_, _38030_);
  and _87731_ (_38067_, _38066_, _38065_);
  and _87732_ (_38068_, _37653_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _87733_ (_38069_, _37656_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor _87734_ (_38070_, _38069_, _38068_);
  and _87735_ (_38071_, _37659_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _87736_ (_38073_, _37661_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor _87737_ (_38074_, _38073_, _38071_);
  and _87738_ (_38075_, _38074_, _38070_);
  nor _87739_ (_38076_, _38075_, _37667_);
  and _87740_ (_38077_, _37653_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _87741_ (_38078_, _37656_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor _87742_ (_38079_, _38078_, _38077_);
  and _87743_ (_38080_, _37659_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _87744_ (_38081_, _37661_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor _87745_ (_38082_, _38081_, _38080_);
  and _87746_ (_38084_, _38082_, _38079_);
  nor _87747_ (_38085_, _38084_, _37678_);
  nor _87748_ (_38086_, _38085_, _38076_);
  and _87749_ (_38087_, _37653_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _87750_ (_38088_, _37656_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor _87751_ (_38089_, _38088_, _38087_);
  and _87752_ (_38090_, _37659_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _87753_ (_38091_, _37661_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor _87754_ (_38092_, _38091_, _38090_);
  and _87755_ (_38093_, _38092_, _38089_);
  nor _87756_ (_38095_, _38093_, _37691_);
  and _87757_ (_38096_, _37653_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _87758_ (_38097_, _37656_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor _87759_ (_38098_, _38097_, _38096_);
  and _87760_ (_38099_, _37659_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _87761_ (_38100_, _37661_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor _87762_ (_38101_, _38100_, _38099_);
  and _87763_ (_38102_, _38101_, _38098_);
  nor _87764_ (_38103_, _38102_, _37702_);
  nor _87765_ (_38104_, _38103_, _38095_);
  and _87766_ (_38106_, _38104_, _38086_);
  and _87767_ (_38107_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _87768_ (_38108_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _87769_ (_38109_, _38108_, _38107_);
  and _87770_ (_38110_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _87771_ (_38111_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _87772_ (_38112_, _38111_, _38110_);
  and _87773_ (_38113_, _38112_, _38109_);
  and _87774_ (_38114_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and _87775_ (_38115_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _87776_ (_38117_, _38115_, _38114_);
  and _87777_ (_38118_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and _87778_ (_38119_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor _87779_ (_38120_, _38119_, _38118_);
  and _87780_ (_38121_, _38120_, _38117_);
  and _87781_ (_38122_, _38121_, _38113_);
  and _87782_ (_38123_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and _87783_ (_38124_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _87784_ (_38125_, _38124_, _38123_);
  and _87785_ (_38126_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _87786_ (_38128_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _87787_ (_38129_, _38128_, _38126_);
  and _87788_ (_38130_, _38129_, _38125_);
  and _87789_ (_38131_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and _87790_ (_38132_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _87791_ (_38133_, _38132_, _38131_);
  and _87792_ (_38134_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _87793_ (_38135_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor _87794_ (_38136_, _38135_, _38134_);
  and _87795_ (_38137_, _38136_, _38133_);
  and _87796_ (_38139_, _38137_, _38130_);
  and _87797_ (_38140_, _38139_, _38122_);
  nand _87798_ (_38141_, _38140_, _38106_);
  or _87799_ (_38142_, _38140_, _38106_);
  and _87800_ (_38143_, _38142_, _38141_);
  or _87801_ (_38144_, _38143_, _38067_);
  and _87802_ (_38145_, _37653_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _87803_ (_38146_, _37656_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor _87804_ (_38147_, _38146_, _38145_);
  and _87805_ (_38148_, _37659_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _87806_ (_38150_, _37661_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor _87807_ (_38151_, _38150_, _38148_);
  and _87808_ (_38152_, _38151_, _38147_);
  nor _87809_ (_38153_, _38152_, _37691_);
  and _87810_ (_38154_, _37653_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _87811_ (_38155_, _37656_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor _87812_ (_38156_, _38155_, _38154_);
  and _87813_ (_38157_, _37659_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _87814_ (_38158_, _37661_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor _87815_ (_38159_, _38158_, _38157_);
  and _87816_ (_38161_, _38159_, _38156_);
  nor _87817_ (_38162_, _38161_, _37678_);
  nor _87818_ (_38163_, _38162_, _38153_);
  and _87819_ (_38164_, _37653_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _87820_ (_38165_, _37656_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor _87821_ (_38166_, _38165_, _38164_);
  and _87822_ (_38167_, _37659_, \oc8051_golden_model_1.IRAM[0] [7]);
  and _87823_ (_38168_, _37661_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor _87824_ (_38169_, _38168_, _38167_);
  and _87825_ (_38170_, _38169_, _38166_);
  nor _87826_ (_38172_, _38170_, _37667_);
  and _87827_ (_38173_, _37653_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _87828_ (_38174_, _37656_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor _87829_ (_38175_, _38174_, _38173_);
  and _87830_ (_38176_, _37659_, \oc8051_golden_model_1.IRAM[8] [7]);
  and _87831_ (_38177_, _37661_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor _87832_ (_38178_, _38177_, _38176_);
  and _87833_ (_38179_, _38178_, _38175_);
  nor _87834_ (_38180_, _38179_, _37702_);
  nor _87835_ (_38181_, _38180_, _38172_);
  and _87836_ (_38183_, _38181_, _38163_);
  and _87837_ (_38184_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and _87838_ (_38185_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _87839_ (_38186_, _38185_, _38184_);
  and _87840_ (_38187_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _87841_ (_38188_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor _87842_ (_38189_, _38188_, _38187_);
  and _87843_ (_38190_, _38189_, _38186_);
  and _87844_ (_38191_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _87845_ (_38192_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _87846_ (_38194_, _38192_, _38191_);
  and _87847_ (_38195_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and _87848_ (_38196_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _87849_ (_38197_, _38196_, _38195_);
  and _87850_ (_38198_, _38197_, _38194_);
  and _87851_ (_38199_, _38198_, _38190_);
  and _87852_ (_38200_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _87853_ (_38201_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor _87854_ (_38202_, _38201_, _38200_);
  and _87855_ (_38203_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _87856_ (_38205_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor _87857_ (_38206_, _38205_, _38203_);
  and _87858_ (_38207_, _38206_, _38202_);
  and _87859_ (_38208_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and _87860_ (_38209_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _87861_ (_38210_, _38209_, _38208_);
  and _87862_ (_38211_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and _87863_ (_38212_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _87864_ (_38213_, _38212_, _38211_);
  and _87865_ (_38214_, _38213_, _38210_);
  and _87866_ (_38216_, _38214_, _38207_);
  and _87867_ (_38217_, _38216_, _38199_);
  nand _87868_ (_38218_, _38217_, _38183_);
  or _87869_ (_38219_, _38217_, _38183_);
  and _87870_ (_38220_, _38219_, _38218_);
  and _87871_ (_38221_, _37653_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _87872_ (_38222_, _37656_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor _87873_ (_38223_, _38222_, _38221_);
  and _87874_ (_38224_, _37659_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _87875_ (_38225_, _37661_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor _87876_ (_38227_, _38225_, _38224_);
  and _87877_ (_38228_, _38227_, _38223_);
  nor _87878_ (_38229_, _38228_, _37667_);
  and _87879_ (_38230_, _37653_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _87880_ (_38231_, _37656_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor _87881_ (_38232_, _38231_, _38230_);
  and _87882_ (_38233_, _37659_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _87883_ (_38234_, _37661_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor _87884_ (_38235_, _38234_, _38233_);
  and _87885_ (_38236_, _38235_, _38232_);
  nor _87886_ (_38238_, _38236_, _37702_);
  nor _87887_ (_38239_, _38238_, _38229_);
  and _87888_ (_38240_, _37653_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _87889_ (_38241_, _37656_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor _87890_ (_38242_, _38241_, _38240_);
  and _87891_ (_38243_, _37659_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _87892_ (_38244_, _37661_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor _87893_ (_38245_, _38244_, _38243_);
  and _87894_ (_38246_, _38245_, _38242_);
  nor _87895_ (_38247_, _38246_, _37691_);
  and _87896_ (_38249_, _37653_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _87897_ (_38250_, _37656_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor _87898_ (_38251_, _38250_, _38249_);
  and _87899_ (_38252_, _37659_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _87900_ (_38253_, _37661_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor _87901_ (_38254_, _38253_, _38252_);
  and _87902_ (_38255_, _38254_, _38251_);
  nor _87903_ (_38256_, _38255_, _37678_);
  nor _87904_ (_38257_, _38256_, _38247_);
  and _87905_ (_38258_, _38257_, _38239_);
  and _87906_ (_38260_, _37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and _87907_ (_38261_, _37721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _87908_ (_38262_, _38261_, _38260_);
  and _87909_ (_38263_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _87910_ (_38264_, _37718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _87911_ (_38265_, _38264_, _38263_);
  and _87912_ (_38266_, _38265_, _38262_);
  and _87913_ (_38267_, _37739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _87914_ (_38268_, _37714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _87915_ (_38269_, _38268_, _38267_);
  and _87916_ (_38271_, _37724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _87917_ (_38272_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _87918_ (_38273_, _38272_, _38271_);
  and _87919_ (_38274_, _38273_, _38269_);
  and _87920_ (_38275_, _38274_, _38266_);
  and _87921_ (_38276_, _37712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and _87922_ (_38277_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _87923_ (_38278_, _38277_, _38276_);
  and _87924_ (_38279_, _37708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and _87925_ (_38280_, _37746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _87926_ (_38282_, _38280_, _38279_);
  and _87927_ (_38283_, _38282_, _38278_);
  and _87928_ (_38284_, _37737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _87929_ (_38285_, _37744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _87930_ (_38286_, _38285_, _38284_);
  and _87931_ (_38287_, _37732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and _87932_ (_38288_, _37734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _87933_ (_38289_, _38288_, _38287_);
  and _87934_ (_38290_, _38289_, _38286_);
  and _87935_ (_38291_, _38290_, _38283_);
  and _87936_ (_38293_, _38291_, _38275_);
  not _87937_ (_38294_, _38293_);
  nor _87938_ (_38295_, _38294_, _38258_);
  and _87939_ (_38296_, _38294_, _38258_);
  or _87940_ (_38297_, _38296_, _38295_);
  or _87941_ (_38298_, _38297_, _38220_);
  or _87942_ (_38299_, _38298_, _38144_);
  or _87943_ (_38300_, _38299_, _37991_);
  and _87944_ (property_invalid_iram, _38300_, _37651_);
  nor _87945_ (_38301_, _09981_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _87946_ (_38303_, _09981_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _87947_ (_38304_, _38303_, _38301_);
  nand _87948_ (_38305_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _87949_ (_38306_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _87950_ (_38307_, _38306_, _38305_);
  or _87951_ (_38308_, _38307_, _38304_);
  and _87952_ (_38309_, _05887_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _87953_ (_38310_, _05887_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _87954_ (_38311_, _38310_, _38309_);
  and _87955_ (_38312_, _05855_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _87956_ (_38314_, \oc8051_golden_model_1.ACC [0], _39264_);
  or _87957_ (_38315_, _38314_, _38312_);
  or _87958_ (_38316_, _38315_, _38311_);
  or _87959_ (_38317_, _38316_, _38308_);
  or _87960_ (_38318_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _87961_ (_38319_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _87962_ (_38320_, _38319_, _38318_);
  or _87963_ (_38321_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _87964_ (_38322_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _87965_ (_38323_, _38322_, _38321_);
  or _87966_ (_38325_, _38323_, _38320_);
  nand _87967_ (_38326_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _87968_ (_38327_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _87969_ (_38328_, _38327_, _38326_);
  and _87970_ (_38329_, _08430_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _87971_ (_38330_, _08430_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _87972_ (_38331_, _38330_, _38329_);
  or _87973_ (_38332_, _38331_, _38328_);
  or _87974_ (_38333_, _38332_, _38325_);
  or _87975_ (_38334_, _38333_, _38317_);
  and _87976_ (property_invalid_acc, _38334_, _37651_);
  nor _87977_ (_38336_, _25393_, _01950_);
  and _87978_ (_38337_, _26427_, _01962_);
  and _87979_ (_38338_, _25393_, _01950_);
  or _87980_ (_38339_, _38338_, _38337_);
  or _87981_ (_38340_, _38339_, _38336_);
  nor _87982_ (_38341_, _27478_, _01973_);
  and _87983_ (_38342_, _27478_, _01973_);
  nor _87984_ (_38343_, _26780_, _01966_);
  or _87985_ (_38344_, _38343_, _38342_);
  or _87986_ (_38346_, _38344_, _38341_);
  nor _87987_ (_38347_, _26427_, _01962_);
  and _87988_ (_38348_, _26780_, _01966_);
  nand _87989_ (_38349_, _27123_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _87990_ (_38350_, _27123_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _87991_ (_38351_, _38350_, _38349_);
  nor _87992_ (_38352_, _26084_, _01958_);
  and _87993_ (_38353_, _26084_, _01958_);
  nor _87994_ (_38354_, _28124_, _38782_);
  and _87995_ (_38355_, _28124_, _38782_);
  nor _87996_ (_38357_, _12760_, _38760_);
  nor _87997_ (_38358_, _28439_, _38787_);
  and _87998_ (_38359_, _12760_, _38760_);
  or _87999_ (_38360_, _38359_, _38358_);
  or _88000_ (_38361_, _38360_, _38357_);
  and _88001_ (_38362_, _28742_, _38772_);
  nor _88002_ (_38363_, _28742_, _38772_);
  or _88003_ (_38364_, _38363_, _38362_);
  and _88004_ (_38365_, _29365_, _38768_);
  and _88005_ (_38366_, _28439_, _38787_);
  or _88006_ (_38368_, _38366_, _38365_);
  or _88007_ (_38369_, _38368_, _38364_);
  nand _88008_ (_38370_, _27800_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _88009_ (_38371_, _27800_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _88010_ (_38372_, _38371_, _38370_);
  nor _88011_ (_38373_, _29365_, _38768_);
  nor _88012_ (_38374_, _29666_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _88013_ (_38375_, _29666_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _88014_ (_38376_, _25025_, _01946_);
  nor _88015_ (_38377_, _25025_, _01946_);
  or _88016_ (_38379_, _38377_, _38376_);
  or _88017_ (_38380_, _38379_, _38375_);
  or _88018_ (_38381_, _38380_, _38374_);
  nor _88019_ (_38382_, _29057_, _38793_);
  and _88020_ (_38383_, _29057_, _38793_);
  or _88021_ (_38384_, _38383_, _38382_);
  or _88022_ (_38385_, _38384_, _38381_);
  or _88023_ (_38386_, _38385_, _38373_);
  or _88024_ (_38387_, _38386_, _38372_);
  or _88025_ (_38388_, _38387_, _38369_);
  or _88026_ (_38390_, _38388_, _38361_);
  or _88027_ (_38391_, _38390_, _38355_);
  or _88028_ (_38392_, _38391_, _38354_);
  or _88029_ (_38393_, _38392_, _38353_);
  or _88030_ (_38394_, _38393_, _38352_);
  or _88031_ (_38395_, _38394_, _38351_);
  or _88032_ (_38396_, _38395_, _38348_);
  or _88033_ (_38397_, _38396_, _38347_);
  or _88034_ (_38398_, _38397_, _38346_);
  or _88035_ (_38399_, _38398_, _38340_);
  and _88036_ (_38401_, _25749_, _01954_);
  nor _88037_ (_38402_, _25749_, _01954_);
  or _88038_ (_38403_, _38402_, _38401_);
  or _88039_ (_38404_, _38403_, _38399_);
  and _88040_ (_38405_, _37650_, _01317_);
  and _88041_ (property_invalid_pc, _38405_, _38404_);
  buf _88042_ (_00544_, _43102_);
  buf _88043_ (_05108_, _43100_);
  buf _88044_ (_05159_, _43100_);
  buf _88045_ (_05211_, _43100_);
  buf _88046_ (_05262_, _43100_);
  buf _88047_ (_05314_, _43100_);
  buf _88048_ (_05365_, _43100_);
  buf _88049_ (_05417_, _43100_);
  buf _88050_ (_05470_, _43100_);
  buf _88051_ (_05523_, _43100_);
  buf _88052_ (_05576_, _43100_);
  buf _88053_ (_05629_, _43100_);
  buf _88054_ (_05682_, _43100_);
  buf _88055_ (_05735_, _43100_);
  buf _88056_ (_05788_, _43100_);
  buf _88057_ (_05841_, _43100_);
  buf _88058_ (_05894_, _43100_);
  buf _88059_ (_39277_, _39174_);
  buf _88060_ (_39279_, _39176_);
  buf _88061_ (_39292_, _39174_);
  buf _88062_ (_39293_, _39176_);
  buf _88063_ (_39605_, _39194_);
  buf _88064_ (_39606_, _39195_);
  buf _88065_ (_39607_, _39197_);
  buf _88066_ (_39608_, _39198_);
  buf _88067_ (_39609_, _39199_);
  buf _88068_ (_39610_, _39200_);
  buf _88069_ (_39611_, _39201_);
  buf _88070_ (_39612_, _39203_);
  buf _88071_ (_39613_, _39204_);
  buf _88072_ (_39615_, _39205_);
  buf _88073_ (_39616_, _39206_);
  buf _88074_ (_39617_, _39207_);
  buf _88075_ (_39618_, _39209_);
  buf _88076_ (_39619_, _39210_);
  buf _88077_ (_39670_, _39194_);
  buf _88078_ (_39671_, _39195_);
  buf _88079_ (_39672_, _39197_);
  buf _88080_ (_39673_, _39198_);
  buf _88081_ (_39674_, _39199_);
  buf _88082_ (_39675_, _39200_);
  buf _88083_ (_39676_, _39201_);
  buf _88084_ (_39677_, _39203_);
  buf _88085_ (_39678_, _39204_);
  buf _88086_ (_39680_, _39205_);
  buf _88087_ (_39681_, _39206_);
  buf _88088_ (_39682_, _39207_);
  buf _88089_ (_39683_, _39209_);
  buf _88090_ (_39684_, _39210_);
  buf _88091_ (_40076_, _39980_);
  buf _88092_ (_40240_, _39980_);
  dff _88093_ (op0_cnst, _00001_, clk);
  dff _88094_ (inst_finished_r, _00000_, clk);
  dff _88095_ (\oc8051_gm_cxrom_1.cell0.data [0], _05111_, clk);
  dff _88096_ (\oc8051_gm_cxrom_1.cell0.data [1], _05115_, clk);
  dff _88097_ (\oc8051_gm_cxrom_1.cell0.data [2], _05119_, clk);
  dff _88098_ (\oc8051_gm_cxrom_1.cell0.data [3], _05123_, clk);
  dff _88099_ (\oc8051_gm_cxrom_1.cell0.data [4], _05127_, clk);
  dff _88100_ (\oc8051_gm_cxrom_1.cell0.data [5], _05131_, clk);
  dff _88101_ (\oc8051_gm_cxrom_1.cell0.data [6], _05135_, clk);
  dff _88102_ (\oc8051_gm_cxrom_1.cell0.data [7], _05105_, clk);
  dff _88103_ (\oc8051_gm_cxrom_1.cell0.valid , _05108_, clk);
  dff _88104_ (\oc8051_gm_cxrom_1.cell1.data [0], _05163_, clk);
  dff _88105_ (\oc8051_gm_cxrom_1.cell1.data [1], _05167_, clk);
  dff _88106_ (\oc8051_gm_cxrom_1.cell1.data [2], _05171_, clk);
  dff _88107_ (\oc8051_gm_cxrom_1.cell1.data [3], _05175_, clk);
  dff _88108_ (\oc8051_gm_cxrom_1.cell1.data [4], _05179_, clk);
  dff _88109_ (\oc8051_gm_cxrom_1.cell1.data [5], _05183_, clk);
  dff _88110_ (\oc8051_gm_cxrom_1.cell1.data [6], _05186_, clk);
  dff _88111_ (\oc8051_gm_cxrom_1.cell1.data [7], _05156_, clk);
  dff _88112_ (\oc8051_gm_cxrom_1.cell1.valid , _05159_, clk);
  dff _88113_ (\oc8051_gm_cxrom_1.cell10.data [0], _05633_, clk);
  dff _88114_ (\oc8051_gm_cxrom_1.cell10.data [1], _05637_, clk);
  dff _88115_ (\oc8051_gm_cxrom_1.cell10.data [2], _05641_, clk);
  dff _88116_ (\oc8051_gm_cxrom_1.cell10.data [3], _05645_, clk);
  dff _88117_ (\oc8051_gm_cxrom_1.cell10.data [4], _05649_, clk);
  dff _88118_ (\oc8051_gm_cxrom_1.cell10.data [5], _05653_, clk);
  dff _88119_ (\oc8051_gm_cxrom_1.cell10.data [6], _05657_, clk);
  dff _88120_ (\oc8051_gm_cxrom_1.cell10.data [7], _05626_, clk);
  dff _88121_ (\oc8051_gm_cxrom_1.cell10.valid , _05629_, clk);
  dff _88122_ (\oc8051_gm_cxrom_1.cell11.data [0], _05686_, clk);
  dff _88123_ (\oc8051_gm_cxrom_1.cell11.data [1], _05690_, clk);
  dff _88124_ (\oc8051_gm_cxrom_1.cell11.data [2], _05694_, clk);
  dff _88125_ (\oc8051_gm_cxrom_1.cell11.data [3], _05698_, clk);
  dff _88126_ (\oc8051_gm_cxrom_1.cell11.data [4], _05702_, clk);
  dff _88127_ (\oc8051_gm_cxrom_1.cell11.data [5], _05706_, clk);
  dff _88128_ (\oc8051_gm_cxrom_1.cell11.data [6], _05710_, clk);
  dff _88129_ (\oc8051_gm_cxrom_1.cell11.data [7], _05679_, clk);
  dff _88130_ (\oc8051_gm_cxrom_1.cell11.valid , _05682_, clk);
  dff _88131_ (\oc8051_gm_cxrom_1.cell12.data [0], _05739_, clk);
  dff _88132_ (\oc8051_gm_cxrom_1.cell12.data [1], _05743_, clk);
  dff _88133_ (\oc8051_gm_cxrom_1.cell12.data [2], _05747_, clk);
  dff _88134_ (\oc8051_gm_cxrom_1.cell12.data [3], _05751_, clk);
  dff _88135_ (\oc8051_gm_cxrom_1.cell12.data [4], _05755_, clk);
  dff _88136_ (\oc8051_gm_cxrom_1.cell12.data [5], _05759_, clk);
  dff _88137_ (\oc8051_gm_cxrom_1.cell12.data [6], _05763_, clk);
  dff _88138_ (\oc8051_gm_cxrom_1.cell12.data [7], _05732_, clk);
  dff _88139_ (\oc8051_gm_cxrom_1.cell12.valid , _05735_, clk);
  dff _88140_ (\oc8051_gm_cxrom_1.cell13.data [0], _05792_, clk);
  dff _88141_ (\oc8051_gm_cxrom_1.cell13.data [1], _05796_, clk);
  dff _88142_ (\oc8051_gm_cxrom_1.cell13.data [2], _05800_, clk);
  dff _88143_ (\oc8051_gm_cxrom_1.cell13.data [3], _05804_, clk);
  dff _88144_ (\oc8051_gm_cxrom_1.cell13.data [4], _05808_, clk);
  dff _88145_ (\oc8051_gm_cxrom_1.cell13.data [5], _05812_, clk);
  dff _88146_ (\oc8051_gm_cxrom_1.cell13.data [6], _05816_, clk);
  dff _88147_ (\oc8051_gm_cxrom_1.cell13.data [7], _05785_, clk);
  dff _88148_ (\oc8051_gm_cxrom_1.cell13.valid , _05788_, clk);
  dff _88149_ (\oc8051_gm_cxrom_1.cell14.data [0], _05845_, clk);
  dff _88150_ (\oc8051_gm_cxrom_1.cell14.data [1], _05849_, clk);
  dff _88151_ (\oc8051_gm_cxrom_1.cell14.data [2], _05853_, clk);
  dff _88152_ (\oc8051_gm_cxrom_1.cell14.data [3], _05857_, clk);
  dff _88153_ (\oc8051_gm_cxrom_1.cell14.data [4], _05861_, clk);
  dff _88154_ (\oc8051_gm_cxrom_1.cell14.data [5], _05865_, clk);
  dff _88155_ (\oc8051_gm_cxrom_1.cell14.data [6], _05869_, clk);
  dff _88156_ (\oc8051_gm_cxrom_1.cell14.data [7], _05838_, clk);
  dff _88157_ (\oc8051_gm_cxrom_1.cell14.valid , _05841_, clk);
  dff _88158_ (\oc8051_gm_cxrom_1.cell15.data [0], _05898_, clk);
  dff _88159_ (\oc8051_gm_cxrom_1.cell15.data [1], _05902_, clk);
  dff _88160_ (\oc8051_gm_cxrom_1.cell15.data [2], _05906_, clk);
  dff _88161_ (\oc8051_gm_cxrom_1.cell15.data [3], _05910_, clk);
  dff _88162_ (\oc8051_gm_cxrom_1.cell15.data [4], _05914_, clk);
  dff _88163_ (\oc8051_gm_cxrom_1.cell15.data [5], _05918_, clk);
  dff _88164_ (\oc8051_gm_cxrom_1.cell15.data [6], _05922_, clk);
  dff _88165_ (\oc8051_gm_cxrom_1.cell15.data [7], _05891_, clk);
  dff _88166_ (\oc8051_gm_cxrom_1.cell15.valid , _05894_, clk);
  dff _88167_ (\oc8051_gm_cxrom_1.cell2.data [0], _05215_, clk);
  dff _88168_ (\oc8051_gm_cxrom_1.cell2.data [1], _05219_, clk);
  dff _88169_ (\oc8051_gm_cxrom_1.cell2.data [2], _05222_, clk);
  dff _88170_ (\oc8051_gm_cxrom_1.cell2.data [3], _05226_, clk);
  dff _88171_ (\oc8051_gm_cxrom_1.cell2.data [4], _05230_, clk);
  dff _88172_ (\oc8051_gm_cxrom_1.cell2.data [5], _05234_, clk);
  dff _88173_ (\oc8051_gm_cxrom_1.cell2.data [6], _05238_, clk);
  dff _88174_ (\oc8051_gm_cxrom_1.cell2.data [7], _05208_, clk);
  dff _88175_ (\oc8051_gm_cxrom_1.cell2.valid , _05211_, clk);
  dff _88176_ (\oc8051_gm_cxrom_1.cell3.data [0], _05266_, clk);
  dff _88177_ (\oc8051_gm_cxrom_1.cell3.data [1], _05270_, clk);
  dff _88178_ (\oc8051_gm_cxrom_1.cell3.data [2], _05274_, clk);
  dff _88179_ (\oc8051_gm_cxrom_1.cell3.data [3], _05278_, clk);
  dff _88180_ (\oc8051_gm_cxrom_1.cell3.data [4], _05282_, clk);
  dff _88181_ (\oc8051_gm_cxrom_1.cell3.data [5], _05286_, clk);
  dff _88182_ (\oc8051_gm_cxrom_1.cell3.data [6], _05290_, clk);
  dff _88183_ (\oc8051_gm_cxrom_1.cell3.data [7], _05259_, clk);
  dff _88184_ (\oc8051_gm_cxrom_1.cell3.valid , _05262_, clk);
  dff _88185_ (\oc8051_gm_cxrom_1.cell4.data [0], _05318_, clk);
  dff _88186_ (\oc8051_gm_cxrom_1.cell4.data [1], _05322_, clk);
  dff _88187_ (\oc8051_gm_cxrom_1.cell4.data [2], _05326_, clk);
  dff _88188_ (\oc8051_gm_cxrom_1.cell4.data [3], _05329_, clk);
  dff _88189_ (\oc8051_gm_cxrom_1.cell4.data [4], _05333_, clk);
  dff _88190_ (\oc8051_gm_cxrom_1.cell4.data [5], _05337_, clk);
  dff _88191_ (\oc8051_gm_cxrom_1.cell4.data [6], _05341_, clk);
  dff _88192_ (\oc8051_gm_cxrom_1.cell4.data [7], _05311_, clk);
  dff _88193_ (\oc8051_gm_cxrom_1.cell4.valid , _05314_, clk);
  dff _88194_ (\oc8051_gm_cxrom_1.cell5.data [0], _05369_, clk);
  dff _88195_ (\oc8051_gm_cxrom_1.cell5.data [1], _05373_, clk);
  dff _88196_ (\oc8051_gm_cxrom_1.cell5.data [2], _05377_, clk);
  dff _88197_ (\oc8051_gm_cxrom_1.cell5.data [3], _05381_, clk);
  dff _88198_ (\oc8051_gm_cxrom_1.cell5.data [4], _05385_, clk);
  dff _88199_ (\oc8051_gm_cxrom_1.cell5.data [5], _05389_, clk);
  dff _88200_ (\oc8051_gm_cxrom_1.cell5.data [6], _05393_, clk);
  dff _88201_ (\oc8051_gm_cxrom_1.cell5.data [7], _05363_, clk);
  dff _88202_ (\oc8051_gm_cxrom_1.cell5.valid , _05365_, clk);
  dff _88203_ (\oc8051_gm_cxrom_1.cell6.data [0], _05421_, clk);
  dff _88204_ (\oc8051_gm_cxrom_1.cell6.data [1], _05425_, clk);
  dff _88205_ (\oc8051_gm_cxrom_1.cell6.data [2], _05429_, clk);
  dff _88206_ (\oc8051_gm_cxrom_1.cell6.data [3], _05433_, clk);
  dff _88207_ (\oc8051_gm_cxrom_1.cell6.data [4], _05437_, clk);
  dff _88208_ (\oc8051_gm_cxrom_1.cell6.data [5], _05441_, clk);
  dff _88209_ (\oc8051_gm_cxrom_1.cell6.data [6], _05445_, clk);
  dff _88210_ (\oc8051_gm_cxrom_1.cell6.data [7], _05414_, clk);
  dff _88211_ (\oc8051_gm_cxrom_1.cell6.valid , _05417_, clk);
  dff _88212_ (\oc8051_gm_cxrom_1.cell7.data [0], _05474_, clk);
  dff _88213_ (\oc8051_gm_cxrom_1.cell7.data [1], _05478_, clk);
  dff _88214_ (\oc8051_gm_cxrom_1.cell7.data [2], _05482_, clk);
  dff _88215_ (\oc8051_gm_cxrom_1.cell7.data [3], _05486_, clk);
  dff _88216_ (\oc8051_gm_cxrom_1.cell7.data [4], _05490_, clk);
  dff _88217_ (\oc8051_gm_cxrom_1.cell7.data [5], _05494_, clk);
  dff _88218_ (\oc8051_gm_cxrom_1.cell7.data [6], _05498_, clk);
  dff _88219_ (\oc8051_gm_cxrom_1.cell7.data [7], _05467_, clk);
  dff _88220_ (\oc8051_gm_cxrom_1.cell7.valid , _05470_, clk);
  dff _88221_ (\oc8051_gm_cxrom_1.cell8.data [0], _05527_, clk);
  dff _88222_ (\oc8051_gm_cxrom_1.cell8.data [1], _05531_, clk);
  dff _88223_ (\oc8051_gm_cxrom_1.cell8.data [2], _05535_, clk);
  dff _88224_ (\oc8051_gm_cxrom_1.cell8.data [3], _05539_, clk);
  dff _88225_ (\oc8051_gm_cxrom_1.cell8.data [4], _05543_, clk);
  dff _88226_ (\oc8051_gm_cxrom_1.cell8.data [5], _05547_, clk);
  dff _88227_ (\oc8051_gm_cxrom_1.cell8.data [6], _05551_, clk);
  dff _88228_ (\oc8051_gm_cxrom_1.cell8.data [7], _05520_, clk);
  dff _88229_ (\oc8051_gm_cxrom_1.cell8.valid , _05523_, clk);
  dff _88230_ (\oc8051_gm_cxrom_1.cell9.data [0], _05580_, clk);
  dff _88231_ (\oc8051_gm_cxrom_1.cell9.data [1], _05584_, clk);
  dff _88232_ (\oc8051_gm_cxrom_1.cell9.data [2], _05588_, clk);
  dff _88233_ (\oc8051_gm_cxrom_1.cell9.data [3], _05592_, clk);
  dff _88234_ (\oc8051_gm_cxrom_1.cell9.data [4], _05596_, clk);
  dff _88235_ (\oc8051_gm_cxrom_1.cell9.data [5], _05600_, clk);
  dff _88236_ (\oc8051_gm_cxrom_1.cell9.data [6], _05604_, clk);
  dff _88237_ (\oc8051_gm_cxrom_1.cell9.data [7], _05573_, clk);
  dff _88238_ (\oc8051_gm_cxrom_1.cell9.valid , _05576_, clk);
  dff _88239_ (\oc8051_golden_model_1.IRAM[15] [0], _41193_, clk);
  dff _88240_ (\oc8051_golden_model_1.IRAM[15] [1], _41194_, clk);
  dff _88241_ (\oc8051_golden_model_1.IRAM[15] [2], _41196_, clk);
  dff _88242_ (\oc8051_golden_model_1.IRAM[15] [3], _41197_, clk);
  dff _88243_ (\oc8051_golden_model_1.IRAM[15] [4], _41198_, clk);
  dff _88244_ (\oc8051_golden_model_1.IRAM[15] [5], _41199_, clk);
  dff _88245_ (\oc8051_golden_model_1.IRAM[15] [6], _41200_, clk);
  dff _88246_ (\oc8051_golden_model_1.IRAM[15] [7], _40979_, clk);
  dff _88247_ (\oc8051_golden_model_1.IRAM[14] [0], _41181_, clk);
  dff _88248_ (\oc8051_golden_model_1.IRAM[14] [1], _41182_, clk);
  dff _88249_ (\oc8051_golden_model_1.IRAM[14] [2], _41184_, clk);
  dff _88250_ (\oc8051_golden_model_1.IRAM[14] [3], _41185_, clk);
  dff _88251_ (\oc8051_golden_model_1.IRAM[14] [4], _41186_, clk);
  dff _88252_ (\oc8051_golden_model_1.IRAM[14] [5], _41187_, clk);
  dff _88253_ (\oc8051_golden_model_1.IRAM[14] [6], _41188_, clk);
  dff _88254_ (\oc8051_golden_model_1.IRAM[14] [7], _41190_, clk);
  dff _88255_ (\oc8051_golden_model_1.IRAM[13] [0], _41169_, clk);
  dff _88256_ (\oc8051_golden_model_1.IRAM[13] [1], _41170_, clk);
  dff _88257_ (\oc8051_golden_model_1.IRAM[13] [2], _41171_, clk);
  dff _88258_ (\oc8051_golden_model_1.IRAM[13] [3], _41173_, clk);
  dff _88259_ (\oc8051_golden_model_1.IRAM[13] [4], _41174_, clk);
  dff _88260_ (\oc8051_golden_model_1.IRAM[13] [5], _41175_, clk);
  dff _88261_ (\oc8051_golden_model_1.IRAM[13] [6], _41176_, clk);
  dff _88262_ (\oc8051_golden_model_1.IRAM[13] [7], _41177_, clk);
  dff _88263_ (\oc8051_golden_model_1.IRAM[12] [0], _41158_, clk);
  dff _88264_ (\oc8051_golden_model_1.IRAM[12] [1], _41159_, clk);
  dff _88265_ (\oc8051_golden_model_1.IRAM[12] [2], _41160_, clk);
  dff _88266_ (\oc8051_golden_model_1.IRAM[12] [3], _41162_, clk);
  dff _88267_ (\oc8051_golden_model_1.IRAM[12] [4], _41163_, clk);
  dff _88268_ (\oc8051_golden_model_1.IRAM[12] [5], _41164_, clk);
  dff _88269_ (\oc8051_golden_model_1.IRAM[12] [6], _41165_, clk);
  dff _88270_ (\oc8051_golden_model_1.IRAM[12] [7], _41166_, clk);
  dff _88271_ (\oc8051_golden_model_1.IRAM[11] [0], _41148_, clk);
  dff _88272_ (\oc8051_golden_model_1.IRAM[11] [1], _41149_, clk);
  dff _88273_ (\oc8051_golden_model_1.IRAM[11] [2], _41150_, clk);
  dff _88274_ (\oc8051_golden_model_1.IRAM[11] [3], _41151_, clk);
  dff _88275_ (\oc8051_golden_model_1.IRAM[11] [4], _41152_, clk);
  dff _88276_ (\oc8051_golden_model_1.IRAM[11] [5], _41153_, clk);
  dff _88277_ (\oc8051_golden_model_1.IRAM[11] [6], _41154_, clk);
  dff _88278_ (\oc8051_golden_model_1.IRAM[11] [7], _41155_, clk);
  dff _88279_ (\oc8051_golden_model_1.IRAM[10] [0], _41136_, clk);
  dff _88280_ (\oc8051_golden_model_1.IRAM[10] [1], _41137_, clk);
  dff _88281_ (\oc8051_golden_model_1.IRAM[10] [2], _41138_, clk);
  dff _88282_ (\oc8051_golden_model_1.IRAM[10] [3], _41139_, clk);
  dff _88283_ (\oc8051_golden_model_1.IRAM[10] [4], _41140_, clk);
  dff _88284_ (\oc8051_golden_model_1.IRAM[10] [5], _41142_, clk);
  dff _88285_ (\oc8051_golden_model_1.IRAM[10] [6], _41143_, clk);
  dff _88286_ (\oc8051_golden_model_1.IRAM[10] [7], _41144_, clk);
  dff _88287_ (\oc8051_golden_model_1.IRAM[9] [0], _41123_, clk);
  dff _88288_ (\oc8051_golden_model_1.IRAM[9] [1], _41124_, clk);
  dff _88289_ (\oc8051_golden_model_1.IRAM[9] [2], _41125_, clk);
  dff _88290_ (\oc8051_golden_model_1.IRAM[9] [3], _41126_, clk);
  dff _88291_ (\oc8051_golden_model_1.IRAM[9] [4], _41127_, clk);
  dff _88292_ (\oc8051_golden_model_1.IRAM[9] [5], _41128_, clk);
  dff _88293_ (\oc8051_golden_model_1.IRAM[9] [6], _41131_, clk);
  dff _88294_ (\oc8051_golden_model_1.IRAM[9] [7], _41132_, clk);
  dff _88295_ (\oc8051_golden_model_1.IRAM[8] [0], _41112_, clk);
  dff _88296_ (\oc8051_golden_model_1.IRAM[8] [1], _41114_, clk);
  dff _88297_ (\oc8051_golden_model_1.IRAM[8] [2], _41115_, clk);
  dff _88298_ (\oc8051_golden_model_1.IRAM[8] [3], _41116_, clk);
  dff _88299_ (\oc8051_golden_model_1.IRAM[8] [4], _41117_, clk);
  dff _88300_ (\oc8051_golden_model_1.IRAM[8] [5], _41118_, clk);
  dff _88301_ (\oc8051_golden_model_1.IRAM[8] [6], _41120_, clk);
  dff _88302_ (\oc8051_golden_model_1.IRAM[8] [7], _41121_, clk);
  dff _88303_ (\oc8051_golden_model_1.IRAM[7] [0], _41100_, clk);
  dff _88304_ (\oc8051_golden_model_1.IRAM[7] [1], _41101_, clk);
  dff _88305_ (\oc8051_golden_model_1.IRAM[7] [2], _41102_, clk);
  dff _88306_ (\oc8051_golden_model_1.IRAM[7] [3], _41103_, clk);
  dff _88307_ (\oc8051_golden_model_1.IRAM[7] [4], _41104_, clk);
  dff _88308_ (\oc8051_golden_model_1.IRAM[7] [5], _41106_, clk);
  dff _88309_ (\oc8051_golden_model_1.IRAM[7] [6], _41107_, clk);
  dff _88310_ (\oc8051_golden_model_1.IRAM[7] [7], _41108_, clk);
  dff _88311_ (\oc8051_golden_model_1.IRAM[6] [0], _41088_, clk);
  dff _88312_ (\oc8051_golden_model_1.IRAM[6] [1], _41089_, clk);
  dff _88313_ (\oc8051_golden_model_1.IRAM[6] [2], _41090_, clk);
  dff _88314_ (\oc8051_golden_model_1.IRAM[6] [3], _41091_, clk);
  dff _88315_ (\oc8051_golden_model_1.IRAM[6] [4], _41092_, clk);
  dff _88316_ (\oc8051_golden_model_1.IRAM[6] [5], _41094_, clk);
  dff _88317_ (\oc8051_golden_model_1.IRAM[6] [6], _41095_, clk);
  dff _88318_ (\oc8051_golden_model_1.IRAM[6] [7], _41096_, clk);
  dff _88319_ (\oc8051_golden_model_1.IRAM[5] [0], _41075_, clk);
  dff _88320_ (\oc8051_golden_model_1.IRAM[5] [1], _41077_, clk);
  dff _88321_ (\oc8051_golden_model_1.IRAM[5] [2], _41078_, clk);
  dff _88322_ (\oc8051_golden_model_1.IRAM[5] [3], _41079_, clk);
  dff _88323_ (\oc8051_golden_model_1.IRAM[5] [4], _41080_, clk);
  dff _88324_ (\oc8051_golden_model_1.IRAM[5] [5], _41081_, clk);
  dff _88325_ (\oc8051_golden_model_1.IRAM[5] [6], _41083_, clk);
  dff _88326_ (\oc8051_golden_model_1.IRAM[5] [7], _41084_, clk);
  dff _88327_ (\oc8051_golden_model_1.IRAM[4] [0], _41063_, clk);
  dff _88328_ (\oc8051_golden_model_1.IRAM[4] [1], _41066_, clk);
  dff _88329_ (\oc8051_golden_model_1.IRAM[4] [2], _41067_, clk);
  dff _88330_ (\oc8051_golden_model_1.IRAM[4] [3], _41068_, clk);
  dff _88331_ (\oc8051_golden_model_1.IRAM[4] [4], _41069_, clk);
  dff _88332_ (\oc8051_golden_model_1.IRAM[4] [5], _41070_, clk);
  dff _88333_ (\oc8051_golden_model_1.IRAM[4] [6], _41071_, clk);
  dff _88334_ (\oc8051_golden_model_1.IRAM[4] [7], _41072_, clk);
  dff _88335_ (\oc8051_golden_model_1.IRAM[3] [0], _41052_, clk);
  dff _88336_ (\oc8051_golden_model_1.IRAM[3] [1], _41053_, clk);
  dff _88337_ (\oc8051_golden_model_1.IRAM[3] [2], _41054_, clk);
  dff _88338_ (\oc8051_golden_model_1.IRAM[3] [3], _41055_, clk);
  dff _88339_ (\oc8051_golden_model_1.IRAM[3] [4], _41056_, clk);
  dff _88340_ (\oc8051_golden_model_1.IRAM[3] [5], _41058_, clk);
  dff _88341_ (\oc8051_golden_model_1.IRAM[3] [6], _41059_, clk);
  dff _88342_ (\oc8051_golden_model_1.IRAM[3] [7], _41060_, clk);
  dff _88343_ (\oc8051_golden_model_1.IRAM[2] [0], _41038_, clk);
  dff _88344_ (\oc8051_golden_model_1.IRAM[2] [1], _41041_, clk);
  dff _88345_ (\oc8051_golden_model_1.IRAM[2] [2], _41042_, clk);
  dff _88346_ (\oc8051_golden_model_1.IRAM[2] [3], _41043_, clk);
  dff _88347_ (\oc8051_golden_model_1.IRAM[2] [4], _41044_, clk);
  dff _88348_ (\oc8051_golden_model_1.IRAM[2] [5], _41045_, clk);
  dff _88349_ (\oc8051_golden_model_1.IRAM[2] [6], _41047_, clk);
  dff _88350_ (\oc8051_golden_model_1.IRAM[2] [7], _41048_, clk);
  dff _88351_ (\oc8051_golden_model_1.IRAM[1] [0], _41027_, clk);
  dff _88352_ (\oc8051_golden_model_1.IRAM[1] [1], _41028_, clk);
  dff _88353_ (\oc8051_golden_model_1.IRAM[1] [2], _41029_, clk);
  dff _88354_ (\oc8051_golden_model_1.IRAM[1] [3], _41030_, clk);
  dff _88355_ (\oc8051_golden_model_1.IRAM[1] [4], _41031_, clk);
  dff _88356_ (\oc8051_golden_model_1.IRAM[1] [5], _41033_, clk);
  dff _88357_ (\oc8051_golden_model_1.IRAM[1] [6], _41034_, clk);
  dff _88358_ (\oc8051_golden_model_1.IRAM[1] [7], _41035_, clk);
  dff _88359_ (\oc8051_golden_model_1.IRAM[0] [0], _41013_, clk);
  dff _88360_ (\oc8051_golden_model_1.IRAM[0] [1], _41014_, clk);
  dff _88361_ (\oc8051_golden_model_1.IRAM[0] [2], _41016_, clk);
  dff _88362_ (\oc8051_golden_model_1.IRAM[0] [3], _41017_, clk);
  dff _88363_ (\oc8051_golden_model_1.IRAM[0] [4], _41018_, clk);
  dff _88364_ (\oc8051_golden_model_1.IRAM[0] [5], _41020_, clk);
  dff _88365_ (\oc8051_golden_model_1.IRAM[0] [6], _41021_, clk);
  dff _88366_ (\oc8051_golden_model_1.IRAM[0] [7], _41022_, clk);
  dff _88367_ (\oc8051_golden_model_1.B [0], _43594_, clk);
  dff _88368_ (\oc8051_golden_model_1.B [1], _43595_, clk);
  dff _88369_ (\oc8051_golden_model_1.B [2], _43596_, clk);
  dff _88370_ (\oc8051_golden_model_1.B [3], _43598_, clk);
  dff _88371_ (\oc8051_golden_model_1.B [4], _43599_, clk);
  dff _88372_ (\oc8051_golden_model_1.B [5], _43600_, clk);
  dff _88373_ (\oc8051_golden_model_1.B [6], _43601_, clk);
  dff _88374_ (\oc8051_golden_model_1.B [7], _40980_, clk);
  dff _88375_ (\oc8051_golden_model_1.ACC [0], _43603_, clk);
  dff _88376_ (\oc8051_golden_model_1.ACC [1], _43604_, clk);
  dff _88377_ (\oc8051_golden_model_1.ACC [2], _43605_, clk);
  dff _88378_ (\oc8051_golden_model_1.ACC [3], _43606_, clk);
  dff _88379_ (\oc8051_golden_model_1.ACC [4], _43607_, clk);
  dff _88380_ (\oc8051_golden_model_1.ACC [5], _43608_, clk);
  dff _88381_ (\oc8051_golden_model_1.ACC [6], _43609_, clk);
  dff _88382_ (\oc8051_golden_model_1.ACC [7], _40981_, clk);
  dff _88383_ (\oc8051_golden_model_1.PCON [0], _43611_, clk);
  dff _88384_ (\oc8051_golden_model_1.PCON [1], _43612_, clk);
  dff _88385_ (\oc8051_golden_model_1.PCON [2], _43613_, clk);
  dff _88386_ (\oc8051_golden_model_1.PCON [3], _43614_, clk);
  dff _88387_ (\oc8051_golden_model_1.PCON [4], _43615_, clk);
  dff _88388_ (\oc8051_golden_model_1.PCON [5], _43617_, clk);
  dff _88389_ (\oc8051_golden_model_1.PCON [6], _43618_, clk);
  dff _88390_ (\oc8051_golden_model_1.PCON [7], _40982_, clk);
  dff _88391_ (\oc8051_golden_model_1.TMOD [0], _43619_, clk);
  dff _88392_ (\oc8051_golden_model_1.TMOD [1], _43621_, clk);
  dff _88393_ (\oc8051_golden_model_1.TMOD [2], _43622_, clk);
  dff _88394_ (\oc8051_golden_model_1.TMOD [3], _43623_, clk);
  dff _88395_ (\oc8051_golden_model_1.TMOD [4], _43624_, clk);
  dff _88396_ (\oc8051_golden_model_1.TMOD [5], _43625_, clk);
  dff _88397_ (\oc8051_golden_model_1.TMOD [6], _43626_, clk);
  dff _88398_ (\oc8051_golden_model_1.TMOD [7], _40983_, clk);
  dff _88399_ (\oc8051_golden_model_1.DPL [0], _43628_, clk);
  dff _88400_ (\oc8051_golden_model_1.DPL [1], _43629_, clk);
  dff _88401_ (\oc8051_golden_model_1.DPL [2], _43630_, clk);
  dff _88402_ (\oc8051_golden_model_1.DPL [3], _43631_, clk);
  dff _88403_ (\oc8051_golden_model_1.DPL [4], _43632_, clk);
  dff _88404_ (\oc8051_golden_model_1.DPL [5], _43633_, clk);
  dff _88405_ (\oc8051_golden_model_1.DPL [6], _43634_, clk);
  dff _88406_ (\oc8051_golden_model_1.DPL [7], _40985_, clk);
  dff _88407_ (\oc8051_golden_model_1.DPH [0], _43636_, clk);
  dff _88408_ (\oc8051_golden_model_1.DPH [1], _43637_, clk);
  dff _88409_ (\oc8051_golden_model_1.DPH [2], _43638_, clk);
  dff _88410_ (\oc8051_golden_model_1.DPH [3], _43640_, clk);
  dff _88411_ (\oc8051_golden_model_1.DPH [4], _43641_, clk);
  dff _88412_ (\oc8051_golden_model_1.DPH [5], _43642_, clk);
  dff _88413_ (\oc8051_golden_model_1.DPH [6], _43643_, clk);
  dff _88414_ (\oc8051_golden_model_1.DPH [7], _40986_, clk);
  dff _88415_ (\oc8051_golden_model_1.TL1 [0], _43645_, clk);
  dff _88416_ (\oc8051_golden_model_1.TL1 [1], _43646_, clk);
  dff _88417_ (\oc8051_golden_model_1.TL1 [2], _43647_, clk);
  dff _88418_ (\oc8051_golden_model_1.TL1 [3], _43648_, clk);
  dff _88419_ (\oc8051_golden_model_1.TL1 [4], _43649_, clk);
  dff _88420_ (\oc8051_golden_model_1.TL1 [5], _43650_, clk);
  dff _88421_ (\oc8051_golden_model_1.TL1 [6], _43651_, clk);
  dff _88422_ (\oc8051_golden_model_1.TL1 [7], _40987_, clk);
  dff _88423_ (\oc8051_golden_model_1.TL0 [0], _43653_, clk);
  dff _88424_ (\oc8051_golden_model_1.TL0 [1], _43654_, clk);
  dff _88425_ (\oc8051_golden_model_1.TL0 [2], _43655_, clk);
  dff _88426_ (\oc8051_golden_model_1.TL0 [3], _43656_, clk);
  dff _88427_ (\oc8051_golden_model_1.TL0 [4], _43657_, clk);
  dff _88428_ (\oc8051_golden_model_1.TL0 [5], _43659_, clk);
  dff _88429_ (\oc8051_golden_model_1.TL0 [6], _43660_, clk);
  dff _88430_ (\oc8051_golden_model_1.TL0 [7], _40988_, clk);
  dff _88431_ (\oc8051_golden_model_1.TCON [0], _43661_, clk);
  dff _88432_ (\oc8051_golden_model_1.TCON [1], _43663_, clk);
  dff _88433_ (\oc8051_golden_model_1.TCON [2], _43664_, clk);
  dff _88434_ (\oc8051_golden_model_1.TCON [3], _43665_, clk);
  dff _88435_ (\oc8051_golden_model_1.TCON [4], _43666_, clk);
  dff _88436_ (\oc8051_golden_model_1.TCON [5], _43667_, clk);
  dff _88437_ (\oc8051_golden_model_1.TCON [6], _43668_, clk);
  dff _88438_ (\oc8051_golden_model_1.TCON [7], _40989_, clk);
  dff _88439_ (\oc8051_golden_model_1.TH1 [0], _43670_, clk);
  dff _88440_ (\oc8051_golden_model_1.TH1 [1], _43671_, clk);
  dff _88441_ (\oc8051_golden_model_1.TH1 [2], _43672_, clk);
  dff _88442_ (\oc8051_golden_model_1.TH1 [3], _43673_, clk);
  dff _88443_ (\oc8051_golden_model_1.TH1 [4], _43674_, clk);
  dff _88444_ (\oc8051_golden_model_1.TH1 [5], _43675_, clk);
  dff _88445_ (\oc8051_golden_model_1.TH1 [6], _43676_, clk);
  dff _88446_ (\oc8051_golden_model_1.TH1 [7], _40991_, clk);
  dff _88447_ (\oc8051_golden_model_1.TH0 [0], _43678_, clk);
  dff _88448_ (\oc8051_golden_model_1.TH0 [1], _43679_, clk);
  dff _88449_ (\oc8051_golden_model_1.TH0 [2], _43680_, clk);
  dff _88450_ (\oc8051_golden_model_1.TH0 [3], _43682_, clk);
  dff _88451_ (\oc8051_golden_model_1.TH0 [4], _43683_, clk);
  dff _88452_ (\oc8051_golden_model_1.TH0 [5], _43684_, clk);
  dff _88453_ (\oc8051_golden_model_1.TH0 [6], _43685_, clk);
  dff _88454_ (\oc8051_golden_model_1.TH0 [7], _40992_, clk);
  dff _88455_ (\oc8051_golden_model_1.PC [0], _43687_, clk);
  dff _88456_ (\oc8051_golden_model_1.PC [1], _43689_, clk);
  dff _88457_ (\oc8051_golden_model_1.PC [2], _43690_, clk);
  dff _88458_ (\oc8051_golden_model_1.PC [3], _43691_, clk);
  dff _88459_ (\oc8051_golden_model_1.PC [4], _43692_, clk);
  dff _88460_ (\oc8051_golden_model_1.PC [5], _43693_, clk);
  dff _88461_ (\oc8051_golden_model_1.PC [6], _43694_, clk);
  dff _88462_ (\oc8051_golden_model_1.PC [7], _43695_, clk);
  dff _88463_ (\oc8051_golden_model_1.PC [8], _43696_, clk);
  dff _88464_ (\oc8051_golden_model_1.PC [9], _43697_, clk);
  dff _88465_ (\oc8051_golden_model_1.PC [10], _43698_, clk);
  dff _88466_ (\oc8051_golden_model_1.PC [11], _43700_, clk);
  dff _88467_ (\oc8051_golden_model_1.PC [12], _43701_, clk);
  dff _88468_ (\oc8051_golden_model_1.PC [13], _43702_, clk);
  dff _88469_ (\oc8051_golden_model_1.PC [14], _43703_, clk);
  dff _88470_ (\oc8051_golden_model_1.PC [15], _40993_, clk);
  dff _88471_ (\oc8051_golden_model_1.P2 [0], _43705_, clk);
  dff _88472_ (\oc8051_golden_model_1.P2 [1], _43706_, clk);
  dff _88473_ (\oc8051_golden_model_1.P2 [2], _43707_, clk);
  dff _88474_ (\oc8051_golden_model_1.P2 [3], _43708_, clk);
  dff _88475_ (\oc8051_golden_model_1.P2 [4], _43709_, clk);
  dff _88476_ (\oc8051_golden_model_1.P2 [5], _43710_, clk);
  dff _88477_ (\oc8051_golden_model_1.P2 [6], _43711_, clk);
  dff _88478_ (\oc8051_golden_model_1.P2 [7], _40994_, clk);
  dff _88479_ (\oc8051_golden_model_1.P3 [0], _43713_, clk);
  dff _88480_ (\oc8051_golden_model_1.P3 [1], _43714_, clk);
  dff _88481_ (\oc8051_golden_model_1.P3 [2], _43715_, clk);
  dff _88482_ (\oc8051_golden_model_1.P3 [3], _43716_, clk);
  dff _88483_ (\oc8051_golden_model_1.P3 [4], _43717_, clk);
  dff _88484_ (\oc8051_golden_model_1.P3 [5], _43719_, clk);
  dff _88485_ (\oc8051_golden_model_1.P3 [6], _43720_, clk);
  dff _88486_ (\oc8051_golden_model_1.P3 [7], _40995_, clk);
  dff _88487_ (\oc8051_golden_model_1.P0 [0], _43721_, clk);
  dff _88488_ (\oc8051_golden_model_1.P0 [1], _43723_, clk);
  dff _88489_ (\oc8051_golden_model_1.P0 [2], _43724_, clk);
  dff _88490_ (\oc8051_golden_model_1.P0 [3], _43725_, clk);
  dff _88491_ (\oc8051_golden_model_1.P0 [4], _43726_, clk);
  dff _88492_ (\oc8051_golden_model_1.P0 [5], _43727_, clk);
  dff _88493_ (\oc8051_golden_model_1.P0 [6], _43728_, clk);
  dff _88494_ (\oc8051_golden_model_1.P0 [7], _40997_, clk);
  dff _88495_ (\oc8051_golden_model_1.P1 [0], _43730_, clk);
  dff _88496_ (\oc8051_golden_model_1.P1 [1], _43731_, clk);
  dff _88497_ (\oc8051_golden_model_1.P1 [2], _43732_, clk);
  dff _88498_ (\oc8051_golden_model_1.P1 [3], _43733_, clk);
  dff _88499_ (\oc8051_golden_model_1.P1 [4], _43734_, clk);
  dff _88500_ (\oc8051_golden_model_1.P1 [5], _43735_, clk);
  dff _88501_ (\oc8051_golden_model_1.P1 [6], _43736_, clk);
  dff _88502_ (\oc8051_golden_model_1.P1 [7], _40998_, clk);
  dff _88503_ (\oc8051_golden_model_1.IP [0], _43738_, clk);
  dff _88504_ (\oc8051_golden_model_1.IP [1], _43739_, clk);
  dff _88505_ (\oc8051_golden_model_1.IP [2], _43740_, clk);
  dff _88506_ (\oc8051_golden_model_1.IP [3], _43742_, clk);
  dff _88507_ (\oc8051_golden_model_1.IP [4], _43743_, clk);
  dff _88508_ (\oc8051_golden_model_1.IP [5], _43744_, clk);
  dff _88509_ (\oc8051_golden_model_1.IP [6], _43745_, clk);
  dff _88510_ (\oc8051_golden_model_1.IP [7], _40999_, clk);
  dff _88511_ (\oc8051_golden_model_1.IE [0], _43747_, clk);
  dff _88512_ (\oc8051_golden_model_1.IE [1], _43748_, clk);
  dff _88513_ (\oc8051_golden_model_1.IE [2], _43749_, clk);
  dff _88514_ (\oc8051_golden_model_1.IE [3], _43750_, clk);
  dff _88515_ (\oc8051_golden_model_1.IE [4], _43751_, clk);
  dff _88516_ (\oc8051_golden_model_1.IE [5], _43752_, clk);
  dff _88517_ (\oc8051_golden_model_1.IE [6], _43753_, clk);
  dff _88518_ (\oc8051_golden_model_1.IE [7], _41000_, clk);
  dff _88519_ (\oc8051_golden_model_1.SCON [0], _43755_, clk);
  dff _88520_ (\oc8051_golden_model_1.SCON [1], _43756_, clk);
  dff _88521_ (\oc8051_golden_model_1.SCON [2], _43757_, clk);
  dff _88522_ (\oc8051_golden_model_1.SCON [3], _43758_, clk);
  dff _88523_ (\oc8051_golden_model_1.SCON [4], _43759_, clk);
  dff _88524_ (\oc8051_golden_model_1.SCON [5], _43761_, clk);
  dff _88525_ (\oc8051_golden_model_1.SCON [6], _43762_, clk);
  dff _88526_ (\oc8051_golden_model_1.SCON [7], _41001_, clk);
  dff _88527_ (\oc8051_golden_model_1.SP [0], _43763_, clk);
  dff _88528_ (\oc8051_golden_model_1.SP [1], _43765_, clk);
  dff _88529_ (\oc8051_golden_model_1.SP [2], _43766_, clk);
  dff _88530_ (\oc8051_golden_model_1.SP [3], _43767_, clk);
  dff _88531_ (\oc8051_golden_model_1.SP [4], _43768_, clk);
  dff _88532_ (\oc8051_golden_model_1.SP [5], _43769_, clk);
  dff _88533_ (\oc8051_golden_model_1.SP [6], _43770_, clk);
  dff _88534_ (\oc8051_golden_model_1.SP [7], _41003_, clk);
  dff _88535_ (\oc8051_golden_model_1.SBUF [0], _43772_, clk);
  dff _88536_ (\oc8051_golden_model_1.SBUF [1], _43773_, clk);
  dff _88537_ (\oc8051_golden_model_1.SBUF [2], _43774_, clk);
  dff _88538_ (\oc8051_golden_model_1.SBUF [3], _43775_, clk);
  dff _88539_ (\oc8051_golden_model_1.SBUF [4], _43776_, clk);
  dff _88540_ (\oc8051_golden_model_1.SBUF [5], _43777_, clk);
  dff _88541_ (\oc8051_golden_model_1.SBUF [6], _43778_, clk);
  dff _88542_ (\oc8051_golden_model_1.SBUF [7], _41004_, clk);
  dff _88543_ (\oc8051_golden_model_1.PSW [0], _43779_, clk);
  dff _88544_ (\oc8051_golden_model_1.PSW [1], _43780_, clk);
  dff _88545_ (\oc8051_golden_model_1.PSW [2], _43781_, clk);
  dff _88546_ (\oc8051_golden_model_1.PSW [3], _43783_, clk);
  dff _88547_ (\oc8051_golden_model_1.PSW [4], _43784_, clk);
  dff _88548_ (\oc8051_golden_model_1.PSW [5], _43785_, clk);
  dff _88549_ (\oc8051_golden_model_1.PSW [6], _43786_, clk);
  dff _88550_ (\oc8051_golden_model_1.PSW [7], _41005_, clk);
  dff _88551_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02839_, clk);
  dff _88552_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02851_, clk);
  dff _88553_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02873_, clk);
  dff _88554_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02897_, clk);
  dff _88555_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02919_, clk);
  dff _88556_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00957_, clk);
  dff _88557_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02931_, clk);
  dff _88558_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00927_, clk);
  dff _88559_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02944_, clk);
  dff _88560_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02957_, clk);
  dff _88561_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02969_, clk);
  dff _88562_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02980_, clk);
  dff _88563_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _02994_, clk);
  dff _88564_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03006_, clk);
  dff _88565_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03020_, clk);
  dff _88566_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00976_, clk);
  dff _88567_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02359_, clk);
  dff _88568_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22218_, clk);
  dff _88569_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02546_, clk);
  dff _88570_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02703_, clk);
  dff _88571_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02884_, clk);
  dff _88572_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03126_, clk);
  dff _88573_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03363_, clk);
  dff _88574_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03564_, clk);
  dff _88575_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03763_, clk);
  dff _88576_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03958_, clk);
  dff _88577_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04057_, clk);
  dff _88578_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04156_, clk);
  dff _88579_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04250_, clk);
  dff _88580_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04349_, clk);
  dff _88581_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04447_, clk);
  dff _88582_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04546_, clk);
  dff _88583_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04645_, clk);
  dff _88584_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24376_, clk);
  dff _88585_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _39186_, clk);
  dff _88586_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _39188_, clk);
  dff _88587_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _39189_, clk);
  dff _88588_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _39190_, clk);
  dff _88589_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _39191_, clk);
  dff _88590_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _39192_, clk);
  dff _88591_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _39193_, clk);
  dff _88592_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _39173_, clk);
  dff _88593_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _39194_, clk);
  dff _88594_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _39195_, clk);
  dff _88595_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _39197_, clk);
  dff _88596_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _39198_, clk);
  dff _88597_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _39199_, clk);
  dff _88598_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _39200_, clk);
  dff _88599_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _39201_, clk);
  dff _88600_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _39174_, clk);
  dff _88601_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _39203_, clk);
  dff _88602_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _39204_, clk);
  dff _88603_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _39205_, clk);
  dff _88604_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _39206_, clk);
  dff _88605_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _39207_, clk);
  dff _88606_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _39209_, clk);
  dff _88607_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _39210_, clk);
  dff _88608_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _39176_, clk);
  dff _88609_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34279_, clk);
  dff _88610_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34282_, clk);
  dff _88611_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09718_, clk);
  dff _88612_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34284_, clk);
  dff _88613_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34286_, clk);
  dff _88614_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09721_, clk);
  dff _88615_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34288_, clk);
  dff _88616_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09724_, clk);
  dff _88617_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34290_, clk);
  dff _88618_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34292_, clk);
  dff _88619_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34294_, clk);
  dff _88620_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09727_, clk);
  dff _88621_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34296_, clk);
  dff _88622_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09730_, clk);
  dff _88623_ (\oc8051_top_1.oc8051_decoder1.wr , _09733_, clk);
  dff _88624_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09792_, clk);
  dff _88625_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09794_, clk);
  dff _88626_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09697_, clk);
  dff _88627_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09797_, clk);
  dff _88628_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09800_, clk);
  dff _88629_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09700_, clk);
  dff _88630_ (\oc8051_top_1.oc8051_decoder1.state [0], _09803_, clk);
  dff _88631_ (\oc8051_top_1.oc8051_decoder1.state [1], _09703_, clk);
  dff _88632_ (\oc8051_top_1.oc8051_decoder1.op [0], _09806_, clk);
  dff _88633_ (\oc8051_top_1.oc8051_decoder1.op [1], _09809_, clk);
  dff _88634_ (\oc8051_top_1.oc8051_decoder1.op [2], _09812_, clk);
  dff _88635_ (\oc8051_top_1.oc8051_decoder1.op [3], _09815_, clk);
  dff _88636_ (\oc8051_top_1.oc8051_decoder1.op [4], _09818_, clk);
  dff _88637_ (\oc8051_top_1.oc8051_decoder1.op [5], _09821_, clk);
  dff _88638_ (\oc8051_top_1.oc8051_decoder1.op [6], _09824_, clk);
  dff _88639_ (\oc8051_top_1.oc8051_decoder1.op [7], _09706_, clk);
  dff _88640_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09709_, clk);
  dff _88641_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34277_, clk);
  dff _88642_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09715_, clk);
  dff _88643_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09827_, clk);
  dff _88644_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09712_, clk);
  dff _88645_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39980_, clk);
  dff _88646_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _40013_, clk);
  dff _88647_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _40014_, clk);
  dff _88648_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _40015_, clk);
  dff _88649_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _40016_, clk);
  dff _88650_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _40017_, clk);
  dff _88651_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _40018_, clk);
  dff _88652_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _40019_, clk);
  dff _88653_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39981_, clk);
  dff _88654_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _40021_, clk);
  dff _88655_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _40022_, clk);
  dff _88656_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _40023_, clk);
  dff _88657_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _40024_, clk);
  dff _88658_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _40025_, clk);
  dff _88659_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _40026_, clk);
  dff _88660_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _40027_, clk);
  dff _88661_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39982_, clk);
  dff _88662_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _40028_, clk);
  dff _88663_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _40029_, clk);
  dff _88664_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _40030_, clk);
  dff _88665_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _40032_, clk);
  dff _88666_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _40033_, clk);
  dff _88667_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _40034_, clk);
  dff _88668_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _40035_, clk);
  dff _88669_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39983_, clk);
  dff _88670_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _40036_, clk);
  dff _88671_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _40037_, clk);
  dff _88672_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _40038_, clk);
  dff _88673_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _40039_, clk);
  dff _88674_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _40040_, clk);
  dff _88675_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _40041_, clk);
  dff _88676_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _40043_, clk);
  dff _88677_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39985_, clk);
  dff _88678_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39558_, clk);
  dff _88679_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39559_, clk);
  dff _88680_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39560_, clk);
  dff _88681_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39561_, clk);
  dff _88682_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _39275_, clk);
  dff _88683_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39347_, clk);
  dff _88684_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39348_, clk);
  dff _88685_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39349_, clk);
  dff _88686_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39350_, clk);
  dff _88687_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39351_, clk);
  dff _88688_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39353_, clk);
  dff _88689_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39354_, clk);
  dff _88690_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39355_, clk);
  dff _88691_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39356_, clk);
  dff _88692_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39357_, clk);
  dff _88693_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39358_, clk);
  dff _88694_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39359_, clk);
  dff _88695_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39360_, clk);
  dff _88696_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39361_, clk);
  dff _88697_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39362_, clk);
  dff _88698_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _39234_, clk);
  dff _88699_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39367_, clk);
  dff _88700_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39368_, clk);
  dff _88701_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39369_, clk);
  dff _88702_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39370_, clk);
  dff _88703_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39371_, clk);
  dff _88704_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39372_, clk);
  dff _88705_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39373_, clk);
  dff _88706_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39374_, clk);
  dff _88707_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39375_, clk);
  dff _88708_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39376_, clk);
  dff _88709_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39378_, clk);
  dff _88710_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39379_, clk);
  dff _88711_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39380_, clk);
  dff _88712_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39381_, clk);
  dff _88713_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39382_, clk);
  dff _88714_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _39235_, clk);
  dff _88715_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39562_, clk);
  dff _88716_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39563_, clk);
  dff _88717_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39564_, clk);
  dff _88718_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39565_, clk);
  dff _88719_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39567_, clk);
  dff _88720_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39568_, clk);
  dff _88721_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39569_, clk);
  dff _88722_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39570_, clk);
  dff _88723_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39571_, clk);
  dff _88724_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39572_, clk);
  dff _88725_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39573_, clk);
  dff _88726_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39574_, clk);
  dff _88727_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39575_, clk);
  dff _88728_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39576_, clk);
  dff _88729_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39578_, clk);
  dff _88730_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39579_, clk);
  dff _88731_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39580_, clk);
  dff _88732_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39581_, clk);
  dff _88733_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39582_, clk);
  dff _88734_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39583_, clk);
  dff _88735_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39584_, clk);
  dff _88736_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39585_, clk);
  dff _88737_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39586_, clk);
  dff _88738_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39587_, clk);
  dff _88739_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39589_, clk);
  dff _88740_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39590_, clk);
  dff _88741_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39591_, clk);
  dff _88742_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39592_, clk);
  dff _88743_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39593_, clk);
  dff _88744_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39594_, clk);
  dff _88745_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39595_, clk);
  dff _88746_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _39300_, clk);
  dff _88747_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _39273_, clk);
  dff _88748_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _88749_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39596_, clk);
  dff _88750_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39598_, clk);
  dff _88751_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39599_, clk);
  dff _88752_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39600_, clk);
  dff _88753_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39601_, clk);
  dff _88754_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39602_, clk);
  dff _88755_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39604_, clk);
  dff _88756_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _39276_, clk);
  dff _88757_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39605_, clk);
  dff _88758_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39606_, clk);
  dff _88759_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39607_, clk);
  dff _88760_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39608_, clk);
  dff _88761_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39609_, clk);
  dff _88762_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39610_, clk);
  dff _88763_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39611_, clk);
  dff _88764_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _39277_, clk);
  dff _88765_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39612_, clk);
  dff _88766_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39613_, clk);
  dff _88767_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39615_, clk);
  dff _88768_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39616_, clk);
  dff _88769_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39617_, clk);
  dff _88770_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39618_, clk);
  dff _88771_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39619_, clk);
  dff _88772_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _39279_, clk);
  dff _88773_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39280_, clk);
  dff _88774_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39281_, clk);
  dff _88775_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39620_, clk);
  dff _88776_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39621_, clk);
  dff _88777_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39622_, clk);
  dff _88778_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39623_, clk);
  dff _88779_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39624_, clk);
  dff _88780_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39626_, clk);
  dff _88781_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39627_, clk);
  dff _88782_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39282_, clk);
  dff _88783_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39628_, clk);
  dff _88784_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39629_, clk);
  dff _88785_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39630_, clk);
  dff _88786_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39631_, clk);
  dff _88787_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39632_, clk);
  dff _88788_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39633_, clk);
  dff _88789_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39634_, clk);
  dff _88790_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39635_, clk);
  dff _88791_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39636_, clk);
  dff _88792_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39637_, clk);
  dff _88793_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39638_, clk);
  dff _88794_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39639_, clk);
  dff _88795_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39640_, clk);
  dff _88796_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39641_, clk);
  dff _88797_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39642_, clk);
  dff _88798_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _39283_, clk);
  dff _88799_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39643_, clk);
  dff _88800_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39644_, clk);
  dff _88801_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39645_, clk);
  dff _88802_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39647_, clk);
  dff _88803_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39648_, clk);
  dff _88804_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39649_, clk);
  dff _88805_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39650_, clk);
  dff _88806_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39651_, clk);
  dff _88807_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39652_, clk);
  dff _88808_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39653_, clk);
  dff _88809_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39654_, clk);
  dff _88810_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39655_, clk);
  dff _88811_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39656_, clk);
  dff _88812_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39658_, clk);
  dff _88813_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39659_, clk);
  dff _88814_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _39285_, clk);
  dff _88815_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _39286_, clk);
  dff _88816_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39288_, clk);
  dff _88817_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _39287_, clk);
  dff _88818_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39660_, clk);
  dff _88819_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39661_, clk);
  dff _88820_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39662_, clk);
  dff _88821_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39663_, clk);
  dff _88822_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39664_, clk);
  dff _88823_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39665_, clk);
  dff _88824_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39666_, clk);
  dff _88825_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _39290_, clk);
  dff _88826_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39667_, clk);
  dff _88827_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39669_, clk);
  dff _88828_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _39291_, clk);
  dff _88829_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39670_, clk);
  dff _88830_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39671_, clk);
  dff _88831_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39672_, clk);
  dff _88832_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39673_, clk);
  dff _88833_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39674_, clk);
  dff _88834_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39675_, clk);
  dff _88835_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39676_, clk);
  dff _88836_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _39292_, clk);
  dff _88837_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39677_, clk);
  dff _88838_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39678_, clk);
  dff _88839_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39680_, clk);
  dff _88840_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39681_, clk);
  dff _88841_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39682_, clk);
  dff _88842_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39683_, clk);
  dff _88843_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39684_, clk);
  dff _88844_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _39293_, clk);
  dff _88845_ (\oc8051_top_1.oc8051_memory_interface1.reti , _39294_, clk);
  dff _88846_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39685_, clk);
  dff _88847_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39686_, clk);
  dff _88848_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39687_, clk);
  dff _88849_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39688_, clk);
  dff _88850_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39689_, clk);
  dff _88851_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39691_, clk);
  dff _88852_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39692_, clk);
  dff _88853_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _39295_, clk);
  dff _88854_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _39297_, clk);
  dff _88855_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _39298_, clk);
  dff _88856_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39693_, clk);
  dff _88857_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39694_, clk);
  dff _88858_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39695_, clk);
  dff _88859_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _39299_, clk);
  dff _88860_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39696_, clk);
  dff _88861_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39697_, clk);
  dff _88862_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39698_, clk);
  dff _88863_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39699_, clk);
  dff _88864_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39700_, clk);
  dff _88865_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39702_, clk);
  dff _88866_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39703_, clk);
  dff _88867_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39704_, clk);
  dff _88868_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39705_, clk);
  dff _88869_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39706_, clk);
  dff _88870_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39707_, clk);
  dff _88871_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39708_, clk);
  dff _88872_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39709_, clk);
  dff _88873_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39710_, clk);
  dff _88874_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39711_, clk);
  dff _88875_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39713_, clk);
  dff _88876_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39714_, clk);
  dff _88877_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39715_, clk);
  dff _88878_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39716_, clk);
  dff _88879_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39717_, clk);
  dff _88880_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39718_, clk);
  dff _88881_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39719_, clk);
  dff _88882_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39720_, clk);
  dff _88883_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39721_, clk);
  dff _88884_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39722_, clk);
  dff _88885_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39724_, clk);
  dff _88886_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39725_, clk);
  dff _88887_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39726_, clk);
  dff _88888_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39727_, clk);
  dff _88889_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39728_, clk);
  dff _88890_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39729_, clk);
  dff _88891_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _39301_, clk);
  dff _88892_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39730_, clk);
  dff _88893_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39731_, clk);
  dff _88894_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39732_, clk);
  dff _88895_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39733_, clk);
  dff _88896_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39735_, clk);
  dff _88897_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39736_, clk);
  dff _88898_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39737_, clk);
  dff _88899_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _39302_, clk);
  dff _88900_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _39303_, clk);
  dff _88901_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _39305_, clk);
  dff _88902_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39738_, clk);
  dff _88903_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39739_, clk);
  dff _88904_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39740_, clk);
  dff _88905_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39741_, clk);
  dff _88906_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39742_, clk);
  dff _88907_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39743_, clk);
  dff _88908_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39744_, clk);
  dff _88909_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39746_, clk);
  dff _88910_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39747_, clk);
  dff _88911_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39748_, clk);
  dff _88912_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39749_, clk);
  dff _88913_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39750_, clk);
  dff _88914_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39751_, clk);
  dff _88915_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39752_, clk);
  dff _88916_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39753_, clk);
  dff _88917_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _39306_, clk);
  dff _88918_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _39307_, clk);
  dff _88919_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _39308_, clk);
  dff _88920_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _39309_, clk);
  dff _88921_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39754_, clk);
  dff _88922_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39755_, clk);
  dff _88923_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39757_, clk);
  dff _88924_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39758_, clk);
  dff _88925_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39759_, clk);
  dff _88926_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39760_, clk);
  dff _88927_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39761_, clk);
  dff _88928_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39762_, clk);
  dff _88929_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39763_, clk);
  dff _88930_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39764_, clk);
  dff _88931_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39765_, clk);
  dff _88932_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39766_, clk);
  dff _88933_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39768_, clk);
  dff _88934_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39769_, clk);
  dff _88935_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39770_, clk);
  dff _88936_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _39310_, clk);
  dff _88937_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _39311_, clk);
  dff _88938_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _40237_, clk);
  dff _88939_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _40258_, clk);
  dff _88940_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _40259_, clk);
  dff _88941_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _40260_, clk);
  dff _88942_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _40261_, clk);
  dff _88943_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _40262_, clk);
  dff _88944_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _40263_, clk);
  dff _88945_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _40264_, clk);
  dff _88946_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _40239_, clk);
  dff _88947_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _40240_, clk);
  dff _88948_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _40265_, clk);
  dff _88949_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _40266_, clk);
  dff _88950_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _40241_, clk);
  dff _88951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03170_, clk);
  dff _88952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03173_, clk);
  dff _88953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03177_, clk);
  dff _88954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03181_, clk);
  dff _88955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03185_, clk);
  dff _88956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03189_, clk);
  dff _88957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03193_, clk);
  dff _88958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03196_, clk);
  dff _88959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03141_, clk);
  dff _88960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03145_, clk);
  dff _88961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03148_, clk);
  dff _88962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03152_, clk);
  dff _88963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03155_, clk);
  dff _88964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03159_, clk);
  dff _88965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03162_, clk);
  dff _88966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03165_, clk);
  dff _88967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02802_, clk);
  dff _88968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02807_, clk);
  dff _88969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02812_, clk);
  dff _88970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02817_, clk);
  dff _88971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02822_, clk);
  dff _88972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02827_, clk);
  dff _88973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02832_, clk);
  dff _88974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02834_, clk);
  dff _88975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02842_, clk);
  dff _88976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02845_, clk);
  dff _88977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02848_, clk);
  dff _88978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02853_, clk);
  dff _88979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02856_, clk);
  dff _88980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02859_, clk);
  dff _88981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02862_, clk);
  dff _88982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02865_, clk);
  dff _88983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02871_, clk);
  dff _88984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02875_, clk);
  dff _88985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02879_, clk);
  dff _88986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02882_, clk);
  dff _88987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02886_, clk);
  dff _88988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02889_, clk);
  dff _88989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02893_, clk);
  dff _88990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02895_, clk);
  dff _88991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02933_, clk);
  dff _88992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02937_, clk);
  dff _88993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02940_, clk);
  dff _88994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02945_, clk);
  dff _88995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02949_, clk);
  dff _88996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02952_, clk);
  dff _88997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02956_, clk);
  dff _88998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02959_, clk);
  dff _88999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02901_, clk);
  dff _89000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02904_, clk);
  dff _89001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02907_, clk);
  dff _89002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02910_, clk);
  dff _89003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02914_, clk);
  dff _89004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02917_, clk);
  dff _89005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02922_, clk);
  dff _89006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02925_, clk);
  dff _89007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03083_, clk);
  dff _89008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03086_, clk);
  dff _89009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03090_, clk);
  dff _89010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03094_, clk);
  dff _89011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03097_, clk);
  dff _89012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03101_, clk);
  dff _89013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03104_, clk);
  dff _89014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03107_, clk);
  dff _89015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03054_, clk);
  dff _89016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03058_, clk);
  dff _89017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03062_, clk);
  dff _89018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03065_, clk);
  dff _89019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03069_, clk);
  dff _89020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03072_, clk);
  dff _89021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03076_, clk);
  dff _89022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03078_, clk);
  dff _89023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03023_, clk);
  dff _89024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03027_, clk);
  dff _89025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03030_, clk);
  dff _89026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03034_, clk);
  dff _89027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03038_, clk);
  dff _89028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03041_, clk);
  dff _89029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03045_, clk);
  dff _89030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03047_, clk);
  dff _89031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02992_, clk);
  dff _89032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _02996_, clk);
  dff _89033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03000_, clk);
  dff _89034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03003_, clk);
  dff _89035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03008_, clk);
  dff _89036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03012_, clk);
  dff _89037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03015_, clk);
  dff _89038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03018_, clk);
  dff _89039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02963_, clk);
  dff _89040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02966_, clk);
  dff _89041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02971_, clk);
  dff _89042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02974_, clk);
  dff _89043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02977_, clk);
  dff _89044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02981_, clk);
  dff _89045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02985_, clk);
  dff _89046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02987_, clk);
  dff _89047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03111_, clk);
  dff _89048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03115_, clk);
  dff _89049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03119_, clk);
  dff _89050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03122_, clk);
  dff _89051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03127_, clk);
  dff _89052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03130_, clk);
  dff _89053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03134_, clk);
  dff _89054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03137_, clk);
  dff _89055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03265_, clk);
  dff _89056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03269_, clk);
  dff _89057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03273_, clk);
  dff _89058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03277_, clk);
  dff _89059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03281_, clk);
  dff _89060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03285_, clk);
  dff _89061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03289_, clk);
  dff _89062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02578_, clk);
  dff _89063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03233_, clk);
  dff _89064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03237_, clk);
  dff _89065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03241_, clk);
  dff _89066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03245_, clk);
  dff _89067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03249_, clk);
  dff _89068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03253_, clk);
  dff _89069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03257_, clk);
  dff _89070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03260_, clk);
  dff _89071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03201_, clk);
  dff _89072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03205_, clk);
  dff _89073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03209_, clk);
  dff _89074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03213_, clk);
  dff _89075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03217_, clk);
  dff _89076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03221_, clk);
  dff _89077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03225_, clk);
  dff _89078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03228_, clk);
  dff _89079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05085_, clk);
  dff _89080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05087_, clk);
  dff _89081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05089_, clk);
  dff _89082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05091_, clk);
  dff _89083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05093_, clk);
  dff _89084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05095_, clk);
  dff _89085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05097_, clk);
  dff _89086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02567_, clk);
  dff _89087_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0], clk);
  dff _89088_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1], clk);
  dff _89089_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2], clk);
  dff _89090_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3], clk);
  dff _89091_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4], clk);
  dff _89092_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5], clk);
  dff _89093_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6], clk);
  dff _89094_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7], clk);
  dff _89095_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8], clk);
  dff _89096_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9], clk);
  dff _89097_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10], clk);
  dff _89098_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11], clk);
  dff _89099_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12], clk);
  dff _89100_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13], clk);
  dff _89101_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14], clk);
  dff _89102_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15], clk);
  dff _89103_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16], clk);
  dff _89104_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17], clk);
  dff _89105_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18], clk);
  dff _89106_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19], clk);
  dff _89107_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20], clk);
  dff _89108_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21], clk);
  dff _89109_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22], clk);
  dff _89110_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23], clk);
  dff _89111_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24], clk);
  dff _89112_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25], clk);
  dff _89113_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26], clk);
  dff _89114_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27], clk);
  dff _89115_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28], clk);
  dff _89116_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29], clk);
  dff _89117_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30], clk);
  dff _89118_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31], clk);
  dff _89119_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _89120_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _40070_, clk);
  dff _89121_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _40156_, clk);
  dff _89122_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _40157_, clk);
  dff _89123_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _40158_, clk);
  dff _89124_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _40072_, clk);
  dff _89125_ (\oc8051_top_1.oc8051_sfr1.bit_out , _40073_, clk);
  dff _89126_ (\oc8051_top_1.oc8051_sfr1.wait_data , _40074_, clk);
  dff _89127_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _40159_, clk);
  dff _89128_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _40161_, clk);
  dff _89129_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _40162_, clk);
  dff _89130_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _40163_, clk);
  dff _89131_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _40164_, clk);
  dff _89132_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _40165_, clk);
  dff _89133_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _40166_, clk);
  dff _89134_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _40075_, clk);
  dff _89135_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _40076_, clk);
  dff _89136_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19851_, clk);
  dff _89137_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19863_, clk);
  dff _89138_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19875_, clk);
  dff _89139_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19886_, clk);
  dff _89140_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19898_, clk);
  dff _89141_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19910_, clk);
  dff _89142_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19922_, clk);
  dff _89143_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _18000_, clk);
  dff _89144_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08905_, clk);
  dff _89145_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08916_, clk);
  dff _89146_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08927_, clk);
  dff _89147_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08938_, clk);
  dff _89148_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08949_, clk);
  dff _89149_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08960_, clk);
  dff _89150_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08971_, clk);
  dff _89151_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06664_, clk);
  dff _89152_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13649_, clk);
  dff _89153_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13660_, clk);
  dff _89154_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13671_, clk);
  dff _89155_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13682_, clk);
  dff _89156_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13693_, clk);
  dff _89157_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13704_, clk);
  dff _89158_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13715_, clk);
  dff _89159_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12715_, clk);
  dff _89160_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13726_, clk);
  dff _89161_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13737_, clk);
  dff _89162_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13748_, clk);
  dff _89163_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13758_, clk);
  dff _89164_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13769_, clk);
  dff _89165_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13780_, clk);
  dff _89166_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13791_, clk);
  dff _89167_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12736_, clk);
  dff _89168_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _43104_, clk);
  dff _89169_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _43102_, clk);
  dff _89170_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _89171_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _43100_, clk);
  dff _89172_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00131_, clk);
  dff _89173_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00133_, clk);
  dff _89174_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00135_, clk);
  dff _89175_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00137_, clk);
  dff _89176_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00139_, clk);
  dff _89177_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00140_, clk);
  dff _89178_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00142_, clk);
  dff _89179_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _43098_, clk);
  dff _89180_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00144_, clk);
  dff _89181_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _43096_, clk);
  dff _89182_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _43094_, clk);
  dff _89183_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00146_, clk);
  dff _89184_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00148_, clk);
  dff _89185_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _43093_, clk);
  dff _89186_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00150_, clk);
  dff _89187_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00151_, clk);
  dff _89188_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _43091_, clk);
  dff _89189_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00153_, clk);
  dff _89190_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _43089_, clk);
  dff _89191_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00155_, clk);
  dff _89192_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _43087_, clk);
  dff _89193_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _43058_, clk);
  dff _89194_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _43056_, clk);
  dff _89195_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _43054_, clk);
  dff _89196_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _43052_, clk);
  dff _89197_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00157_, clk);
  dff _89198_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00159_, clk);
  dff _89199_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00161_, clk);
  dff _89200_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _43050_, clk);
  dff _89201_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00162_, clk);
  dff _89202_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00164_, clk);
  dff _89203_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00166_, clk);
  dff _89204_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00168_, clk);
  dff _89205_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00170_, clk);
  dff _89206_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00172_, clk);
  dff _89207_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00173_, clk);
  dff _89208_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _43048_, clk);
  dff _89209_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00175_, clk);
  dff _89210_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00177_, clk);
  dff _89211_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00179_, clk);
  dff _89212_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00181_, clk);
  dff _89213_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00183_, clk);
  dff _89214_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00184_, clk);
  dff _89215_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00186_, clk);
  dff _89216_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _43045_, clk);
  dff _89217_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40808_, clk);
  dff _89218_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40810_, clk);
  dff _89219_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40812_, clk);
  dff _89220_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40814_, clk);
  dff _89221_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40816_, clk);
  dff _89222_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40818_, clk);
  dff _89223_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40820_, clk);
  dff _89224_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31130_, clk);
  dff _89225_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40821_, clk);
  dff _89226_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40823_, clk);
  dff _89227_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40825_, clk);
  dff _89228_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40827_, clk);
  dff _89229_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40829_, clk);
  dff _89230_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40831_, clk);
  dff _89231_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40833_, clk);
  dff _89232_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31153_, clk);
  dff _89233_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40835_, clk);
  dff _89234_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40837_, clk);
  dff _89235_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40839_, clk);
  dff _89236_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40841_, clk);
  dff _89237_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40843_, clk);
  dff _89238_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40845_, clk);
  dff _89239_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40847_, clk);
  dff _89240_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31176_, clk);
  dff _89241_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40849_, clk);
  dff _89242_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40851_, clk);
  dff _89243_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40852_, clk);
  dff _89244_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40854_, clk);
  dff _89245_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40856_, clk);
  dff _89246_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40858_, clk);
  dff _89247_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40860_, clk);
  dff _89248_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31199_, clk);
  dff _89249_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17376_, clk);
  dff _89250_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17387_, clk);
  dff _89251_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17398_, clk);
  dff _89252_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17409_, clk);
  dff _89253_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17420_, clk);
  dff _89254_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17431_, clk);
  dff _89255_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15195_, clk);
  dff _89256_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09521_, clk);
  dff _89257_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10698_, clk);
  dff _89258_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10709_, clk);
  dff _89259_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10720_, clk);
  dff _89260_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10731_, clk);
  dff _89261_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10742_, clk);
  dff _89262_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10753_, clk);
  dff _89263_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10764_, clk);
  dff _89264_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09542_, clk);
  dff _89265_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _41311_, clk);
  dff _89266_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _41314_, clk);
  dff _89267_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41820_, clk);
  dff _89268_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41822_, clk);
  dff _89269_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41823_, clk);
  dff _89270_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41825_, clk);
  dff _89271_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41827_, clk);
  dff _89272_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41829_, clk);
  dff _89273_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41831_, clk);
  dff _89274_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _41317_, clk);
  dff _89275_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41833_, clk);
  dff _89276_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41835_, clk);
  dff _89277_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41837_, clk);
  dff _89278_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41839_, clk);
  dff _89279_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41840_, clk);
  dff _89280_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41842_, clk);
  dff _89281_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41844_, clk);
  dff _89282_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _41320_, clk);
  dff _89283_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _41323_, clk);
  dff _89284_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _41326_, clk);
  dff _89285_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41846_, clk);
  dff _89286_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41848_, clk);
  dff _89287_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41850_, clk);
  dff _89288_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41852_, clk);
  dff _89289_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41854_, clk);
  dff _89290_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41855_, clk);
  dff _89291_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41857_, clk);
  dff _89292_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _41329_, clk);
  dff _89293_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41859_, clk);
  dff _89294_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41861_, clk);
  dff _89295_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41863_, clk);
  dff _89296_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41865_, clk);
  dff _89297_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41867_, clk);
  dff _89298_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41869_, clk);
  dff _89299_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41870_, clk);
  dff _89300_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _41332_, clk);
  dff _89301_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _41335_, clk);
  dff _89302_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41872_, clk);
  dff _89303_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41874_, clk);
  dff _89304_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41876_, clk);
  dff _89305_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41877_, clk);
  dff _89306_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41879_, clk);
  dff _89307_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41881_, clk);
  dff _89308_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41883_, clk);
  dff _89309_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _41338_, clk);
  dff _89310_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01630_, clk);
  dff _89311_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01633_, clk);
  dff _89312_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01636_, clk);
  dff _89313_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01639_, clk);
  dff _89314_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02112_, clk);
  dff _89315_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02114_, clk);
  dff _89316_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02116_, clk);
  dff _89317_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02117_, clk);
  dff _89318_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02119_, clk);
  dff _89319_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02121_, clk);
  dff _89320_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02123_, clk);
  dff _89321_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01642_, clk);
  dff _89322_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02124_, clk);
  dff _89323_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02126_, clk);
  dff _89324_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02128_, clk);
  dff _89325_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02130_, clk);
  dff _89326_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02131_, clk);
  dff _89327_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02133_, clk);
  dff _89328_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02135_, clk);
  dff _89329_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01645_, clk);
  dff _89330_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01648_, clk);
  dff _89331_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02137_, clk);
  dff _89332_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02138_, clk);
  dff _89333_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02140_, clk);
  dff _89334_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02142_, clk);
  dff _89335_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02144_, clk);
  dff _89336_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02145_, clk);
  dff _89337_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02147_, clk);
  dff _89338_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01651_, clk);
  dff _89339_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02149_, clk);
  dff _89340_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02151_, clk);
  dff _89341_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02152_, clk);
  dff _89342_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02154_, clk);
  dff _89343_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02156_, clk);
  dff _89344_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02158_, clk);
  dff _89345_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02159_, clk);
  dff _89346_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01654_, clk);
  dff _89347_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01657_, clk);
  dff _89348_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02161_, clk);
  dff _89349_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02163_, clk);
  dff _89350_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02165_, clk);
  dff _89351_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02166_, clk);
  dff _89352_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02167_, clk);
  dff _89353_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02168_, clk);
  dff _89354_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02169_, clk);
  dff _89355_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01660_, clk);
  dff _89356_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01211_, clk);
  dff _89357_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01213_, clk);
  dff _89358_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01215_, clk);
  dff _89359_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01217_, clk);
  dff _89360_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01219_, clk);
  dff _89361_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01221_, clk);
  dff _89362_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01223_, clk);
  dff _89363_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01224_, clk);
  dff _89364_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01226_, clk);
  dff _89365_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01228_, clk);
  dff _89366_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01230_, clk);
  dff _89367_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00568_, clk);
  dff _89368_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00544_, clk);
  dff _89369_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00546_, clk);
  dff _89370_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00549_, clk);
  dff _89371_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00552_, clk);
  dff _89372_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00554_, clk);
  dff _89373_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00557_, clk);
  dff _89374_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01232_, clk);
  dff _89375_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00560_, clk);
  dff _89376_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01234_, clk);
  dff _89377_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01236_, clk);
  dff _89378_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01238_, clk);
  dff _89379_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00562_, clk);
  dff _89380_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01240_, clk);
  dff _89381_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01242_, clk);
  dff _89382_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01244_, clk);
  dff _89383_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01246_, clk);
  dff _89384_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01248_, clk);
  dff _89385_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01250_, clk);
  dff _89386_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01252_, clk);
  dff _89387_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00565_, clk);
  dff _89388_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00571_, clk);
  dff _89389_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00573_, clk);
  dff _89390_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00576_, clk);
  dff _89391_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00579_, clk);
  dff _89392_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00581_, clk);
  dff _89393_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01254_, clk);
  dff _89394_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01256_, clk);
  dff _89395_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01258_, clk);
  dff _89396_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00584_, clk);
  dff _89397_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01259_, clk);
  dff _89398_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01261_, clk);
  dff _89399_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01263_, clk);
  dff _89400_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01265_, clk);
  dff _89401_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01267_, clk);
  dff _89402_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01269_, clk);
  dff _89403_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01271_, clk);
  dff _89404_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01273_, clk);
  dff _89405_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01275_, clk);
  dff _89406_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01277_, clk);
  dff _89407_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00587_, clk);
  dff _89408_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01279_, clk);
  dff _89409_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01281_, clk);
  dff _89410_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01283_, clk);
  dff _89411_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01285_, clk);
  dff _89412_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01287_, clk);
  dff _89413_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01289_, clk);
  dff _89414_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01291_, clk);
  dff _89415_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00589_, clk);
  dff _89416_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01293_, clk);
  dff _89417_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01294_, clk);
  dff _89418_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01296_, clk);
  dff _89419_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01298_, clk);
  dff _89420_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01300_, clk);
  dff _89421_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01302_, clk);
  dff _89422_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01304_, clk);
  dff _89423_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00592_, clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [0], \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [1], \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [2], \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [3], \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [4], \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [5], \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [6], \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [7], \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [0], \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [1], \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [2], \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [3], \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [4], \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [5], \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [6], \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [7], \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [0], \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [1], \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [2], \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [3], \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [4], \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [5], \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [6], \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [7], \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [0], \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [1], \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [2], \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [3], \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [4], \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [5], \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [6], \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [7], \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1237 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1257 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1276 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1288 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1348 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1364 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1558 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1582 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1591 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1747 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1747 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1747 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1760 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1760 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1760 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1789 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1801 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1805 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1826 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1832 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1838 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1909 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1090 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1090 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1090 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1090 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1092 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1094 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1094 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1094 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1094 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1095 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1095 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1095 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1095 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1096 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1096 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1096 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1096 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1097 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1097 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1097 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1097 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1098 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1098 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1098 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1098 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1099 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1099 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1099 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1099 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1100 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1175 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1176 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1176 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1176 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1176 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1176 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1176 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1176 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1176 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1176 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1177 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1177 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1177 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1177 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1177 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1177 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1177 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1177 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1177 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1178 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1178 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1178 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1178 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1178 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1178 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1178 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1178 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1179 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1180 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1182 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1184 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1184 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1184 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1184 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1184 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1184 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1184 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1184 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1211 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1211 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1211 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1211 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1211 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1211 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1211 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1211 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1211 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1211 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1211 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1211 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n1211 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n1211 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n1211 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1213 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1213 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1213 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1213 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1213 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1213 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1213 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1213 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1215 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1215 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1215 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1215 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1215 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1215 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1215 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1215 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1215 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1219 [8], \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.n1220 , \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.n1221 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1221 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1221 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1221 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1222 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1222 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1222 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1222 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1222 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1226 [4], \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.n1227 , \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.n1228 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1228 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1228 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1228 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1228 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1228 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1228 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1228 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1228 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1236 , \oc8051_golden_model_1.n1237 [2]);
  buf(\oc8051_golden_model_1.n1237 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1237 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1237 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1237 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1237 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1241 [8], \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.n1242 , \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.n1247 [4], \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.n1248 , \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.n1256 , \oc8051_golden_model_1.n1257 [2]);
  buf(\oc8051_golden_model_1.n1257 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1257 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1257 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1257 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1257 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1259 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1259 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1259 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1259 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1259 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1259 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1259 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1259 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1259 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.n1262 , \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.n1263 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1263 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1263 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1263 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1268 [8], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1276 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1279 [8], \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.n1280 , \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.n1287 , \oc8051_golden_model_1.n1288 [2]);
  buf(\oc8051_golden_model_1.n1288 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1288 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1288 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1288 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1288 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1290 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1290 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1290 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1290 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1290 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n1290 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n1290 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n1290 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1290 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1292 [8], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1293 , \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1294 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1294 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1294 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1294 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1294 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1297 , \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1298 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1305 , \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.n1306 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1306 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1306 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.n1306 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1306 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1306 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1306 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1306 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1308 [4], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1309 , \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1310 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1310 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1310 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1310 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1310 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1310 [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1312 [8], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1313 , \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1320 , \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.n1321 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1321 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1321 [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.n1321 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1321 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1321 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1321 [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1322 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1322 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1322 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1322 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1322 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1325 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1325 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1325 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1325 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1325 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1325 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1325 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1325 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1326 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1326 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1326 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1326 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1326 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1326 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1326 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1326 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1326 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1327 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1327 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1327 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1327 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1327 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1327 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1327 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1327 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1328 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1329 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1329 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1329 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1329 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1329 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1329 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1329 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1329 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1330 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1330 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1333 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1335 [8], \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.n1336 , \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.n1337 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1337 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1339 [4], \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.n1340 , \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.n1348 [2]);
  buf(\oc8051_golden_model_1.n1348 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1348 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1348 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1348 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1348 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1352 [8], \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.n1355 [4], \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.n1356 , \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.n1363 , \oc8051_golden_model_1.n1364 [2]);
  buf(\oc8051_golden_model_1.n1364 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1364 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1364 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1364 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1364 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1368 [8], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.n1369 , \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.n1371 [4], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.n1372 , \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.n1379 , \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.n1380 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1380 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1380 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1380 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1380 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1384 [8], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.n1385 , \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.n1387 [4], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.n1388 , \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.n1395 , \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.n1396 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1396 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1396 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1396 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1396 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.n1558 [7]);
  buf(\oc8051_golden_model_1.n1557 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1557 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1557 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1557 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1557 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1557 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1557 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1558 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1558 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1558 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1558 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1558 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1558 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1558 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1581 , \oc8051_golden_model_1.n1582 [7]);
  buf(\oc8051_golden_model_1.n1582 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1582 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1582 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1582 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1582 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1582 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1582 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1589 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1589 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1589 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1589 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1590 , \oc8051_golden_model_1.n1591 [2]);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1591 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1591 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1591 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1591 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1591 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1738 , \oc8051_golden_model_1.n1747 [7]);
  buf(\oc8051_golden_model_1.n1740 , \oc8051_golden_model_1.n1747 [6]);
  buf(\oc8051_golden_model_1.n1746 , \oc8051_golden_model_1.n1747 [2]);
  buf(\oc8051_golden_model_1.n1747 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1751 , \oc8051_golden_model_1.n1760 [7]);
  buf(\oc8051_golden_model_1.n1753 , \oc8051_golden_model_1.n1760 [6]);
  buf(\oc8051_golden_model_1.n1759 , \oc8051_golden_model_1.n1760 [2]);
  buf(\oc8051_golden_model_1.n1760 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1760 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1760 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1760 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1760 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1764 , \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.n1766 , \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.n1772 , \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.n1773 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1773 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1773 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1773 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1773 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.n1779 , \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.n1785 , \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.n1786 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1786 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1786 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1786 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1786 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1788 , \oc8051_golden_model_1.n1789 [7]);
  buf(\oc8051_golden_model_1.n1789 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1789 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1789 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1789 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1789 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1789 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1789 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1794 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1794 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1794 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1794 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1794 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1794 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1794 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1794 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1794 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1800 , \oc8051_golden_model_1.n1801 [2]);
  buf(\oc8051_golden_model_1.n1801 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1801 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1801 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1801 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1801 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1801 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1801 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1804 , \oc8051_golden_model_1.n1805 [7]);
  buf(\oc8051_golden_model_1.n1805 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1825 , \oc8051_golden_model_1.n1826 [7]);
  buf(\oc8051_golden_model_1.n1826 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1826 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1826 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1826 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1826 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1826 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1826 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1831 , \oc8051_golden_model_1.n1832 [7]);
  buf(\oc8051_golden_model_1.n1832 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1832 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1832 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1832 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1832 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1832 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1832 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1837 , \oc8051_golden_model_1.n1838 [7]);
  buf(\oc8051_golden_model_1.n1838 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1838 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1838 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1838 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1838 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1838 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1838 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1843 , \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.n1844 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1844 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1844 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1844 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1844 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1844 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1844 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1849 , \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.n1850 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1850 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1850 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1850 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1850 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1850 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1850 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1851 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1851 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1851 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1851 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1851 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1851 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1851 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1851 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1852 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1853 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1853 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1853 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1889 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1889 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1889 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1889 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1889 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1889 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1889 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1889 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1908 , \oc8051_golden_model_1.n1909 [7]);
  buf(\oc8051_golden_model_1.n1909 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1909 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1909 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1909 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1909 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1909 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1909 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1913 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1913 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1913 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1913 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1914 [0], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1914 [1], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1914 [2], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1914 [3], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1915 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1915 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1915 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1915 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
