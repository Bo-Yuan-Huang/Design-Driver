
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [7:0] \uc8051golden_1.ACC ;
  wire [7:0] \uc8051golden_1.ACC_03 ;
  wire [7:0] \uc8051golden_1.ACC_13 ;
  wire [7:0] \uc8051golden_1.ACC_23 ;
  wire [7:0] \uc8051golden_1.ACC_33 ;
  wire [7:0] \uc8051golden_1.ACC_c4 ;
  wire [7:0] \uc8051golden_1.ACC_d6 ;
  wire [7:0] \uc8051golden_1.ACC_d7 ;
  wire [7:0] \uc8051golden_1.ACC_e4 ;
  wire [7:0] \uc8051golden_1.B ;
  wire [7:0] \uc8051golden_1.DPH ;
  wire [7:0] \uc8051golden_1.DPL ;
  wire [7:0] \uc8051golden_1.IE ;
  wire [7:0] \uc8051golden_1.IP ;
  wire [7:0] \uc8051golden_1.IRAM[0] ;
  wire [7:0] \uc8051golden_1.IRAM[10] ;
  wire [7:0] \uc8051golden_1.IRAM[11] ;
  wire [7:0] \uc8051golden_1.IRAM[12] ;
  wire [7:0] \uc8051golden_1.IRAM[13] ;
  wire [7:0] \uc8051golden_1.IRAM[14] ;
  wire [7:0] \uc8051golden_1.IRAM[15] ;
  wire [7:0] \uc8051golden_1.IRAM[1] ;
  wire [7:0] \uc8051golden_1.IRAM[2] ;
  wire [7:0] \uc8051golden_1.IRAM[3] ;
  wire [7:0] \uc8051golden_1.IRAM[4] ;
  wire [7:0] \uc8051golden_1.IRAM[5] ;
  wire [7:0] \uc8051golden_1.IRAM[6] ;
  wire [7:0] \uc8051golden_1.IRAM[7] ;
  wire [7:0] \uc8051golden_1.IRAM[8] ;
  wire [7:0] \uc8051golden_1.IRAM[9] ;
  wire [7:0] \uc8051golden_1.P0 ;
  wire [7:0] \uc8051golden_1.P1 ;
  wire [7:0] \uc8051golden_1.P2 ;
  wire [7:0] \uc8051golden_1.P3 ;
  wire [15:0] \uc8051golden_1.PC ;
  wire [7:0] \uc8051golden_1.PCON ;
  wire [15:0] \uc8051golden_1.PC_22 ;
  wire [15:0] \uc8051golden_1.PC_32 ;
  wire [7:0] \uc8051golden_1.PSW ;
  wire [7:0] \uc8051golden_1.PSW_13 ;
  wire [7:0] \uc8051golden_1.PSW_24 ;
  wire [7:0] \uc8051golden_1.PSW_25 ;
  wire [7:0] \uc8051golden_1.PSW_26 ;
  wire [7:0] \uc8051golden_1.PSW_27 ;
  wire [7:0] \uc8051golden_1.PSW_28 ;
  wire [7:0] \uc8051golden_1.PSW_29 ;
  wire [7:0] \uc8051golden_1.PSW_2a ;
  wire [7:0] \uc8051golden_1.PSW_2b ;
  wire [7:0] \uc8051golden_1.PSW_2c ;
  wire [7:0] \uc8051golden_1.PSW_2d ;
  wire [7:0] \uc8051golden_1.PSW_2e ;
  wire [7:0] \uc8051golden_1.PSW_2f ;
  wire [7:0] \uc8051golden_1.PSW_33 ;
  wire [7:0] \uc8051golden_1.PSW_34 ;
  wire [7:0] \uc8051golden_1.PSW_35 ;
  wire [7:0] \uc8051golden_1.PSW_36 ;
  wire [7:0] \uc8051golden_1.PSW_37 ;
  wire [7:0] \uc8051golden_1.PSW_38 ;
  wire [7:0] \uc8051golden_1.PSW_39 ;
  wire [7:0] \uc8051golden_1.PSW_3a ;
  wire [7:0] \uc8051golden_1.PSW_3b ;
  wire [7:0] \uc8051golden_1.PSW_3c ;
  wire [7:0] \uc8051golden_1.PSW_3d ;
  wire [7:0] \uc8051golden_1.PSW_3e ;
  wire [7:0] \uc8051golden_1.PSW_3f ;
  wire [7:0] \uc8051golden_1.PSW_72 ;
  wire [7:0] \uc8051golden_1.PSW_82 ;
  wire [7:0] \uc8051golden_1.PSW_84 ;
  wire [7:0] \uc8051golden_1.PSW_94 ;
  wire [7:0] \uc8051golden_1.PSW_95 ;
  wire [7:0] \uc8051golden_1.PSW_96 ;
  wire [7:0] \uc8051golden_1.PSW_97 ;
  wire [7:0] \uc8051golden_1.PSW_98 ;
  wire [7:0] \uc8051golden_1.PSW_99 ;
  wire [7:0] \uc8051golden_1.PSW_9a ;
  wire [7:0] \uc8051golden_1.PSW_9b ;
  wire [7:0] \uc8051golden_1.PSW_9c ;
  wire [7:0] \uc8051golden_1.PSW_9d ;
  wire [7:0] \uc8051golden_1.PSW_9e ;
  wire [7:0] \uc8051golden_1.PSW_9f ;
  wire [7:0] \uc8051golden_1.PSW_a0 ;
  wire [7:0] \uc8051golden_1.PSW_a2 ;
  wire [7:0] \uc8051golden_1.PSW_a4 ;
  wire [7:0] \uc8051golden_1.PSW_b0 ;
  wire [7:0] \uc8051golden_1.PSW_b3 ;
  wire [7:0] \uc8051golden_1.PSW_b4 ;
  wire [7:0] \uc8051golden_1.PSW_b5 ;
  wire [7:0] \uc8051golden_1.PSW_b6 ;
  wire [7:0] \uc8051golden_1.PSW_b7 ;
  wire [7:0] \uc8051golden_1.PSW_b8 ;
  wire [7:0] \uc8051golden_1.PSW_b9 ;
  wire [7:0] \uc8051golden_1.PSW_ba ;
  wire [7:0] \uc8051golden_1.PSW_bb ;
  wire [7:0] \uc8051golden_1.PSW_bc ;
  wire [7:0] \uc8051golden_1.PSW_bd ;
  wire [7:0] \uc8051golden_1.PSW_be ;
  wire [7:0] \uc8051golden_1.PSW_bf ;
  wire [7:0] \uc8051golden_1.PSW_c3 ;
  wire [7:0] \uc8051golden_1.PSW_d3 ;
  wire [7:0] \uc8051golden_1.PSW_d4 ;
  wire [7:0] \uc8051golden_1.RD_IRAM_0 ;
  wire [7:0] \uc8051golden_1.RD_IRAM_1 ;
  wire [15:0] \uc8051golden_1.RD_ROM_0_ADDR ;
  wire [7:0] \uc8051golden_1.SBUF ;
  wire [7:0] \uc8051golden_1.SCON ;
  wire [7:0] \uc8051golden_1.SP ;
  wire [7:0] \uc8051golden_1.TCON ;
  wire [7:0] \uc8051golden_1.TH0 ;
  wire [7:0] \uc8051golden_1.TH1 ;
  wire [7:0] \uc8051golden_1.TL0 ;
  wire [7:0] \uc8051golden_1.TL1 ;
  wire [7:0] \uc8051golden_1.TMOD ;
  wire \uc8051golden_1.clk ;
  wire [1:0] \uc8051golden_1.n0006 ;
  wire [7:0] \uc8051golden_1.n0007 ;
  wire [7:0] \uc8051golden_1.n0011 ;
  wire [7:0] \uc8051golden_1.n0019 ;
  wire [7:0] \uc8051golden_1.n0023 ;
  wire [7:0] \uc8051golden_1.n0027 ;
  wire [7:0] \uc8051golden_1.n0031 ;
  wire [7:0] \uc8051golden_1.n0035 ;
  wire [7:0] \uc8051golden_1.n0039 ;
  wire [7:0] \uc8051golden_1.n0561 ;
  wire [7:0] \uc8051golden_1.n0594 ;
  wire [15:0] \uc8051golden_1.n0701 ;
  wire [15:0] \uc8051golden_1.n0733 ;
  wire [7:0] \uc8051golden_1.n0994 ;
  wire [3:0] \uc8051golden_1.n1071 ;
  wire [3:0] \uc8051golden_1.n1073 ;
  wire [3:0] \uc8051golden_1.n1075 ;
  wire [3:0] \uc8051golden_1.n1076 ;
  wire [3:0] \uc8051golden_1.n1077 ;
  wire [3:0] \uc8051golden_1.n1078 ;
  wire [3:0] \uc8051golden_1.n1079 ;
  wire [3:0] \uc8051golden_1.n1080 ;
  wire [3:0] \uc8051golden_1.n1081 ;
  wire \uc8051golden_1.n1118 ;
  wire \uc8051golden_1.n1146 ;
  wire [8:0] \uc8051golden_1.n1147 ;
  wire [8:0] \uc8051golden_1.n1148 ;
  wire [7:0] \uc8051golden_1.n1149 ;
  wire \uc8051golden_1.n1150 ;
  wire \uc8051golden_1.n1151 ;
  wire [2:0] \uc8051golden_1.n1152 ;
  wire \uc8051golden_1.n1153 ;
  wire [1:0] \uc8051golden_1.n1154 ;
  wire [7:0] \uc8051golden_1.n1155 ;
  wire [15:0] \uc8051golden_1.n1181 ;
  wire [7:0] \uc8051golden_1.n1183 ;
  wire [8:0] \uc8051golden_1.n1185 ;
  wire [8:0] \uc8051golden_1.n1189 ;
  wire \uc8051golden_1.n1190 ;
  wire [3:0] \uc8051golden_1.n1191 ;
  wire [4:0] \uc8051golden_1.n1192 ;
  wire [4:0] \uc8051golden_1.n1196 ;
  wire \uc8051golden_1.n1197 ;
  wire [8:0] \uc8051golden_1.n1198 ;
  wire \uc8051golden_1.n1206 ;
  wire [7:0] \uc8051golden_1.n1207 ;
  wire [8:0] \uc8051golden_1.n1211 ;
  wire \uc8051golden_1.n1212 ;
  wire [4:0] \uc8051golden_1.n1217 ;
  wire \uc8051golden_1.n1218 ;
  wire \uc8051golden_1.n1226 ;
  wire [7:0] \uc8051golden_1.n1227 ;
  wire [8:0] \uc8051golden_1.n1229 ;
  wire [8:0] \uc8051golden_1.n1231 ;
  wire \uc8051golden_1.n1232 ;
  wire [3:0] \uc8051golden_1.n1233 ;
  wire [4:0] \uc8051golden_1.n1234 ;
  wire [4:0] \uc8051golden_1.n1236 ;
  wire \uc8051golden_1.n1237 ;
  wire [8:0] \uc8051golden_1.n1238 ;
  wire \uc8051golden_1.n1245 ;
  wire [7:0] \uc8051golden_1.n1246 ;
  wire [8:0] \uc8051golden_1.n1249 ;
  wire \uc8051golden_1.n1250 ;
  wire \uc8051golden_1.n1257 ;
  wire [7:0] \uc8051golden_1.n1258 ;
  wire [8:0] \uc8051golden_1.n1260 ;
  wire [8:0] \uc8051golden_1.n1262 ;
  wire \uc8051golden_1.n1263 ;
  wire [4:0] \uc8051golden_1.n1264 ;
  wire [4:0] \uc8051golden_1.n1266 ;
  wire \uc8051golden_1.n1267 ;
  wire [8:0] \uc8051golden_1.n1268 ;
  wire \uc8051golden_1.n1275 ;
  wire [7:0] \uc8051golden_1.n1276 ;
  wire [4:0] \uc8051golden_1.n1278 ;
  wire \uc8051golden_1.n1279 ;
  wire [7:0] \uc8051golden_1.n1280 ;
  wire [8:0] \uc8051golden_1.n1282 ;
  wire \uc8051golden_1.n1283 ;
  wire \uc8051golden_1.n1290 ;
  wire [7:0] \uc8051golden_1.n1291 ;
  wire [7:0] \uc8051golden_1.n1292 ;
  wire [8:0] \uc8051golden_1.n1295 ;
  wire [8:0] \uc8051golden_1.n1296 ;
  wire [7:0] \uc8051golden_1.n1297 ;
  wire \uc8051golden_1.n1298 ;
  wire [7:0] \uc8051golden_1.n1299 ;
  wire [7:0] \uc8051golden_1.n1300 ;
  wire [8:0] \uc8051golden_1.n1303 ;
  wire [8:0] \uc8051golden_1.n1305 ;
  wire \uc8051golden_1.n1306 ;
  wire [4:0] \uc8051golden_1.n1307 ;
  wire [4:0] \uc8051golden_1.n1309 ;
  wire \uc8051golden_1.n1310 ;
  wire \uc8051golden_1.n1317 ;
  wire [7:0] \uc8051golden_1.n1318 ;
  wire [8:0] \uc8051golden_1.n1322 ;
  wire \uc8051golden_1.n1323 ;
  wire [4:0] \uc8051golden_1.n1325 ;
  wire \uc8051golden_1.n1326 ;
  wire \uc8051golden_1.n1333 ;
  wire [7:0] \uc8051golden_1.n1334 ;
  wire [8:0] \uc8051golden_1.n1338 ;
  wire \uc8051golden_1.n1339 ;
  wire [4:0] \uc8051golden_1.n1341 ;
  wire \uc8051golden_1.n1342 ;
  wire \uc8051golden_1.n1349 ;
  wire [7:0] \uc8051golden_1.n1350 ;
  wire [8:0] \uc8051golden_1.n1354 ;
  wire \uc8051golden_1.n1355 ;
  wire [4:0] \uc8051golden_1.n1357 ;
  wire \uc8051golden_1.n1358 ;
  wire \uc8051golden_1.n1365 ;
  wire [7:0] \uc8051golden_1.n1366 ;
  wire \uc8051golden_1.n1520 ;
  wire [6:0] \uc8051golden_1.n1521 ;
  wire [7:0] \uc8051golden_1.n1522 ;
  wire \uc8051golden_1.n1545 ;
  wire [7:0] \uc8051golden_1.n1546 ;
  wire [3:0] \uc8051golden_1.n1553 ;
  wire \uc8051golden_1.n1554 ;
  wire [7:0] \uc8051golden_1.n1555 ;
  wire [7:0] \uc8051golden_1.n1680 ;
  wire \uc8051golden_1.n1683 ;
  wire \uc8051golden_1.n1685 ;
  wire \uc8051golden_1.n1691 ;
  wire [7:0] \uc8051golden_1.n1692 ;
  wire \uc8051golden_1.n1696 ;
  wire \uc8051golden_1.n1698 ;
  wire \uc8051golden_1.n1704 ;
  wire [7:0] \uc8051golden_1.n1705 ;
  wire \uc8051golden_1.n1709 ;
  wire \uc8051golden_1.n1711 ;
  wire \uc8051golden_1.n1717 ;
  wire [7:0] \uc8051golden_1.n1718 ;
  wire \uc8051golden_1.n1722 ;
  wire \uc8051golden_1.n1724 ;
  wire \uc8051golden_1.n1730 ;
  wire [7:0] \uc8051golden_1.n1731 ;
  wire \uc8051golden_1.n1733 ;
  wire [7:0] \uc8051golden_1.n1734 ;
  wire [7:0] \uc8051golden_1.n1735 ;
  wire [15:0] \uc8051golden_1.n1739 ;
  wire \uc8051golden_1.n1745 ;
  wire [7:0] \uc8051golden_1.n1746 ;
  wire \uc8051golden_1.n1749 ;
  wire [7:0] \uc8051golden_1.n1750 ;
  wire \uc8051golden_1.n1765 ;
  wire [7:0] \uc8051golden_1.n1766 ;
  wire \uc8051golden_1.n1771 ;
  wire [7:0] \uc8051golden_1.n1772 ;
  wire \uc8051golden_1.n1777 ;
  wire [7:0] \uc8051golden_1.n1778 ;
  wire \uc8051golden_1.n1783 ;
  wire [7:0] \uc8051golden_1.n1784 ;
  wire \uc8051golden_1.n1789 ;
  wire [7:0] \uc8051golden_1.n1790 ;
  wire [7:0] \uc8051golden_1.n1791 ;
  wire [3:0] \uc8051golden_1.n1792 ;
  wire [7:0] \uc8051golden_1.n1793 ;
  wire [7:0] \uc8051golden_1.n1828 ;
  wire \uc8051golden_1.n1847 ;
  wire [7:0] \uc8051golden_1.n1848 ;
  wire [7:0] \uc8051golden_1.n1852 ;
  wire [3:0] \uc8051golden_1.n1853 ;
  wire [7:0] \uc8051golden_1.n1854 ;
  wire \uc8051golden_1.rst ;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_42545_, rst);
  not (_18749_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_18770_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18771_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18770_);
  and (_18782_, _18771_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_18793_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18770_);
  and (_18804_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18770_);
  nor (_18815_, _18804_, _18793_);
  and (_18826_, _18815_, _18782_);
  nor (_18837_, _18826_, _18749_);
  and (_18848_, _18749_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18859_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_18870_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18859_);
  nor (_18881_, _18870_, _18848_);
  not (_18892_, _18881_);
  and (_18903_, _18892_, _18826_);
  or (_18914_, _18903_, _18837_);
  and (_22121_, _18914_, _42545_);
  nor (_18935_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18946_, _18935_);
  and (_18957_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_18968_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_18979_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_18990_, _18979_);
  not (_19001_, _18870_);
  nor (_19012_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_19023_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_19033_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _19023_);
  nor (_19044_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_19055_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_19066_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _19055_);
  nor (_19077_, _19066_, _19044_);
  nor (_19088_, _19077_, _19033_);
  not (_19099_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_19110_, _19033_, _19099_);
  nor (_19121_, _19110_, _19088_);
  and (_19132_, _19121_, _19012_);
  not (_19143_, _19132_);
  and (_19154_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_19165_, _19154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_19176_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_19187_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _19176_);
  and (_19198_, _19187_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_19209_, _19198_, _19165_);
  and (_19220_, _19209_, _19143_);
  nor (_19231_, _19220_, _19001_);
  not (_19242_, _18848_);
  nor (_19253_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_19264_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _19055_);
  nor (_19275_, _19264_, _19253_);
  nor (_19286_, _19275_, _19033_);
  not (_19297_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_19308_, _19033_, _19297_);
  nor (_19319_, _19308_, _19286_);
  and (_19330_, _19319_, _19012_);
  not (_19341_, _19330_);
  and (_19352_, _19154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_19362_, _19187_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_19373_, _19362_, _19352_);
  and (_19384_, _19373_, _19341_);
  nor (_19395_, _19384_, _19242_);
  nor (_19406_, _19395_, _19231_);
  nor (_19417_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_19428_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _19055_);
  nor (_19439_, _19428_, _19417_);
  nor (_19449_, _19439_, _19033_);
  not (_19460_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_19471_, _19033_, _19460_);
  nor (_19482_, _19471_, _19449_);
  and (_19493_, _19482_, _19012_);
  not (_19504_, _19493_);
  and (_19515_, _19154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_19526_, _19187_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_19536_, _19526_, _19515_);
  and (_19547_, _19536_, _19504_);
  nor (_19558_, _19547_, _18892_);
  nor (_19569_, _19558_, _18935_);
  and (_19580_, _19569_, _19406_);
  nor (_19591_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_19602_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _19055_);
  nor (_19613_, _19602_, _19591_);
  nor (_19623_, _19613_, _19033_);
  not (_19634_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_19645_, _19033_, _19634_);
  nor (_19656_, _19645_, _19623_);
  and (_19667_, _19656_, _19012_);
  not (_19678_, _19667_);
  and (_19689_, _19154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_19700_, _19187_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_19710_, _19700_, _19689_);
  and (_19721_, _19710_, _19678_);
  and (_19732_, _19721_, _18935_);
  nor (_19743_, _19732_, _19580_);
  not (_19765_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19777_, _19765_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19788_, _19777_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19800_, _19788_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_19812_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19824_, _19812_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19836_, _19824_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_19837_, _19836_, _19800_);
  not (_19848_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19859_, _19777_, _19848_);
  and (_19870_, _19859_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_19880_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19891_, _19880_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19902_, _19891_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_19913_, _19902_, _19870_);
  and (_19924_, _19913_, _19837_);
  and (_19935_, _19880_, _19765_);
  and (_19946_, _19935_, _19656_);
  and (_19957_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19967_, _19957_, _19848_);
  and (_19978_, _19967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_19989_, _19957_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_20000_, _19989_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_20011_, _20000_, _19978_);
  not (_20022_, _20011_);
  nor (_20033_, _20022_, _19946_);
  and (_20043_, _20033_, _19924_);
  not (_20054_, _20043_);
  and (_20065_, _20054_, _19743_);
  not (_20076_, _20065_);
  nor (_20087_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_20098_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _19055_);
  nor (_20109_, _20098_, _20087_);
  nor (_20120_, _20109_, _19033_);
  not (_20130_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_20141_, _19033_, _20130_);
  nor (_20152_, _20141_, _20120_);
  and (_20163_, _20152_, _19012_);
  not (_20174_, _20163_);
  and (_20185_, _19154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_20196_, _19187_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_20207_, _20196_, _20185_);
  and (_20217_, _20207_, _20174_);
  nor (_20228_, _20217_, _19001_);
  nor (_20239_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_20250_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _19055_);
  nor (_20261_, _20250_, _20239_);
  nor (_20272_, _20261_, _19033_);
  not (_20283_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_20294_, _19033_, _20283_);
  nor (_20304_, _20294_, _20272_);
  and (_20315_, _20304_, _19012_);
  not (_20326_, _20315_);
  and (_20337_, _19154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_20348_, _19187_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_20359_, _20348_, _20337_);
  and (_20370_, _20359_, _20326_);
  nor (_20381_, _20370_, _19242_);
  nor (_20391_, _20381_, _20228_);
  nor (_20402_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_20413_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _19055_);
  nor (_20424_, _20413_, _20402_);
  nor (_20435_, _20424_, _19033_);
  not (_20446_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_20457_, _19033_, _20446_);
  nor (_20467_, _20457_, _20435_);
  and (_20478_, _20467_, _19012_);
  not (_20489_, _20478_);
  and (_20500_, _19154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_20511_, _19187_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_20522_, _20511_, _20500_);
  and (_20533_, _20522_, _20489_);
  nor (_20544_, _20533_, _18892_);
  nor (_20554_, _20544_, _18935_);
  and (_20565_, _20554_, _20391_);
  nor (_20576_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_20587_, _19055_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_20598_, _20587_, _20576_);
  nor (_20609_, _20598_, _19033_);
  not (_20620_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_20631_, _19033_, _20620_);
  nor (_20641_, _20631_, _20609_);
  and (_20652_, _20641_, _19012_);
  not (_20673_, _20652_);
  and (_20684_, _19154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20685_, _19187_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_20696_, _20685_, _20684_);
  and (_20717_, _20696_, _20673_);
  and (_20728_, _20717_, _18935_);
  nor (_20729_, _20728_, _20565_);
  and (_20749_, _19788_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_20760_, _19824_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_20761_, _20760_, _20749_);
  and (_20772_, _19891_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_20783_, _19859_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_20794_, _20783_, _20772_);
  and (_20815_, _20794_, _20761_);
  and (_20816_, _20641_, _19935_);
  and (_20827_, _19967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_20837_, _19989_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_20848_, _20837_, _20827_);
  not (_20859_, _20848_);
  nor (_20870_, _20859_, _20816_);
  and (_20881_, _20870_, _20815_);
  not (_20892_, _20881_);
  and (_20903_, _20892_, _20729_);
  and (_20914_, _20903_, _20076_);
  not (_20924_, _20914_);
  and (_20945_, _19788_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_20946_, _19824_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_20957_, _20946_, _20945_);
  and (_20968_, _19891_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_20979_, _19859_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_20990_, _20979_, _20968_);
  and (_21001_, _20990_, _20957_);
  and (_21012_, _20304_, _19935_);
  and (_21022_, _19989_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_21033_, _19967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_21044_, _21033_, _21022_);
  not (_21055_, _21044_);
  nor (_21066_, _21055_, _21012_);
  and (_21077_, _21066_, _21001_);
  not (_21088_, _21077_);
  and (_21099_, _21088_, _20729_);
  and (_21119_, _19788_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_21120_, _19824_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_21131_, _21120_, _21119_);
  and (_21142_, _19891_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_21153_, _19859_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_21164_, _21153_, _21142_);
  and (_21175_, _21164_, _21131_);
  and (_21186_, _19935_, _19319_);
  and (_21197_, _19967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_21207_, _19989_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_21218_, _21207_, _21197_);
  not (_21229_, _21218_);
  nor (_21240_, _21229_, _21186_);
  and (_21251_, _21240_, _21175_);
  not (_21262_, _21251_);
  and (_21273_, _21262_, _19743_);
  and (_21284_, _21099_, _21273_);
  nor (_21294_, _21284_, _20065_);
  and (_21315_, _21284_, _20054_);
  nor (_21316_, _21315_, _21294_);
  and (_21327_, _21316_, _21099_);
  and (_21338_, _20903_, _20065_);
  and (_21349_, _20729_, _20054_);
  and (_21360_, _20892_, _19743_);
  nor (_21371_, _21360_, _21349_);
  nor (_21382_, _21371_, _21338_);
  and (_21392_, _21382_, _21327_);
  and (_21403_, _21382_, _21315_);
  nor (_21414_, _21403_, _21392_);
  nor (_21425_, _21414_, _20924_);
  and (_21436_, _21414_, _20924_);
  nor (_21447_, _21436_, _21425_);
  not (_21458_, _21447_);
  and (_21469_, _21262_, _20729_);
  and (_21480_, _19788_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_21490_, _19824_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_21501_, _21490_, _21480_);
  and (_21512_, _19891_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_21523_, _19859_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_21534_, _21523_, _21512_);
  and (_21545_, _21534_, _21501_);
  and (_21556_, _20152_, _19935_);
  and (_21567_, _19967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_21577_, _19989_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_21588_, _21577_, _21567_);
  not (_21599_, _21588_);
  nor (_21610_, _21599_, _21556_);
  and (_21621_, _21610_, _21545_);
  not (_21632_, _21621_);
  and (_21643_, _21632_, _19743_);
  and (_21664_, _21643_, _21469_);
  and (_21665_, _21088_, _19743_);
  nor (_21675_, _21665_, _21469_);
  nor (_21686_, _21675_, _21284_);
  and (_21697_, _21686_, _21664_);
  nor (_21708_, _21099_, _20065_);
  nor (_21719_, _21708_, _21327_);
  and (_21730_, _21719_, _21697_);
  nor (_21741_, _21382_, _21327_);
  nor (_21752_, _21741_, _21392_);
  nor (_21772_, _21752_, _21315_);
  nor (_21773_, _21772_, _21403_);
  and (_21784_, _21773_, _21730_);
  nor (_21795_, _21773_, _21730_);
  nor (_21806_, _21795_, _21784_);
  not (_21817_, _21806_);
  and (_21828_, _19788_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_21839_, _19824_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_21850_, _21839_, _21828_);
  and (_21860_, _19891_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_21871_, _19859_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_21882_, _21871_, _21860_);
  and (_21893_, _21882_, _21850_);
  and (_21904_, _20467_, _19935_);
  and (_21915_, _19989_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_21926_, _19967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_21936_, _21926_, _21915_);
  not (_21947_, _21936_);
  nor (_21958_, _21947_, _21904_);
  and (_21969_, _21958_, _21893_);
  not (_21980_, _21969_);
  and (_21991_, _21980_, _20729_);
  and (_22002_, _19788_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_22013_, _19824_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_22023_, _22013_, _22002_);
  and (_22034_, _19891_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_22045_, _19859_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_22056_, _22045_, _22034_);
  and (_22067_, _22056_, _22023_);
  and (_22078_, _19935_, _19121_);
  and (_22089_, _19967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_22100_, _19989_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_22110_, _22100_, _22089_);
  not (_22122_, _22110_);
  nor (_22133_, _22122_, _22078_);
  and (_22144_, _22133_, _22067_);
  not (_22155_, _22144_);
  and (_22166_, _22155_, _19743_);
  and (_22177_, _22166_, _21991_);
  and (_22188_, _21980_, _19743_);
  not (_22198_, _22188_);
  and (_22219_, _22155_, _20729_);
  and (_22220_, _22219_, _22198_);
  and (_22231_, _22220_, _21643_);
  nor (_22242_, _22231_, _22177_);
  and (_22253_, _21632_, _20729_);
  nor (_22264_, _22253_, _21273_);
  nor (_22275_, _22264_, _21664_);
  not (_22285_, _22275_);
  nor (_22296_, _22285_, _22242_);
  nor (_22307_, _21686_, _21664_);
  nor (_22318_, _22307_, _21697_);
  and (_22329_, _22318_, _22296_);
  nor (_22340_, _21719_, _21697_);
  nor (_22351_, _22340_, _21730_);
  and (_22362_, _22351_, _22329_);
  and (_22372_, _19788_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_22383_, _19824_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_22394_, _22383_, _22372_);
  and (_22405_, _19891_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_22416_, _19859_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_22427_, _22416_, _22405_);
  and (_22438_, _22427_, _22394_);
  and (_22448_, _19935_, _19482_);
  and (_22459_, _19989_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_22470_, _19967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_22481_, _22470_, _22459_);
  not (_22492_, _22481_);
  nor (_22513_, _22492_, _22448_);
  and (_22514_, _22513_, _22438_);
  not (_22525_, _22514_);
  and (_22535_, _22525_, _20729_);
  and (_22546_, _22535_, _22188_);
  nor (_22557_, _22166_, _21991_);
  nor (_22568_, _22557_, _22177_);
  and (_22579_, _22568_, _22546_);
  nor (_22590_, _22220_, _21643_);
  nor (_22601_, _22590_, _22231_);
  and (_22621_, _22601_, _22579_);
  and (_22622_, _22285_, _22242_);
  nor (_22633_, _22622_, _22296_);
  and (_22644_, _22633_, _22621_);
  nor (_22655_, _22318_, _22296_);
  nor (_22666_, _22655_, _22329_);
  and (_22677_, _22666_, _22644_);
  nor (_22688_, _22351_, _22329_);
  nor (_22698_, _22688_, _22362_);
  and (_22709_, _22698_, _22677_);
  nor (_22720_, _22709_, _22362_);
  nor (_22731_, _22720_, _21817_);
  nor (_22742_, _22731_, _21784_);
  nor (_22753_, _22742_, _21458_);
  or (_22764_, _22753_, _21338_);
  nor (_22775_, _22764_, _21425_);
  nor (_22785_, _22775_, _18990_);
  and (_22796_, _22775_, _18990_);
  nor (_22807_, _22796_, _22785_);
  not (_22818_, _22807_);
  and (_22839_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_22840_, _22742_, _21458_);
  nor (_22851_, _22840_, _22753_);
  and (_22862_, _22851_, _22839_);
  and (_22872_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_22883_, _22720_, _21817_);
  nor (_22894_, _22883_, _22731_);
  and (_22905_, _22894_, _22872_);
  nor (_22916_, _22894_, _22872_);
  nor (_22927_, _22916_, _22905_);
  and (_22938_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_22949_, _22698_, _22677_);
  nor (_22959_, _22949_, _22709_);
  and (_22970_, _22959_, _22938_);
  nor (_22981_, _22959_, _22938_);
  nor (_22992_, _22981_, _22970_);
  and (_23003_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_23014_, _22666_, _22644_);
  nor (_23025_, _23014_, _22677_);
  and (_23036_, _23025_, _23003_);
  nor (_23046_, _23025_, _23003_);
  nor (_23057_, _23046_, _23036_);
  not (_23068_, _23057_);
  and (_23079_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_23100_, _22633_, _22621_);
  nor (_23101_, _23100_, _22644_);
  and (_23112_, _23101_, _23079_);
  and (_23123_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_23134_, _22601_, _22579_);
  nor (_23144_, _23134_, _22621_);
  and (_23155_, _23144_, _23123_);
  and (_23166_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_23177_, _22568_, _22546_);
  nor (_23188_, _23177_, _22579_);
  and (_23199_, _23188_, _23166_);
  nor (_23210_, _23144_, _23123_);
  nor (_23221_, _23210_, _23155_);
  and (_23232_, _23221_, _23199_);
  nor (_23243_, _23232_, _23155_);
  not (_23254_, _23243_);
  nor (_23264_, _23101_, _23079_);
  nor (_23275_, _23264_, _23112_);
  and (_23286_, _23275_, _23254_);
  nor (_23297_, _23286_, _23112_);
  nor (_23308_, _23297_, _23068_);
  nor (_23319_, _23308_, _23036_);
  not (_23330_, _23319_);
  and (_23341_, _23330_, _22992_);
  nor (_23352_, _23341_, _22970_);
  not (_23363_, _23352_);
  and (_23383_, _23363_, _22927_);
  nor (_23384_, _23383_, _22905_);
  nor (_23395_, _22851_, _22839_);
  nor (_23406_, _23395_, _22862_);
  not (_23417_, _23406_);
  nor (_23428_, _23417_, _23384_);
  nor (_23439_, _23428_, _22862_);
  nor (_23450_, _23439_, _22818_);
  nor (_23461_, _23450_, _22785_);
  not (_23472_, _23461_);
  and (_23482_, _23472_, _18968_);
  and (_23493_, _23482_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_23504_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_23515_, _23504_, _23493_);
  and (_23526_, _23515_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_23537_, _23526_, _18957_);
  not (_23548_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or (_23559_, _18935_, _23548_);
  nor (_23570_, _23559_, _23537_);
  and (_23581_, _23537_, _23548_);
  or (_23591_, _23581_, _23570_);
  and (_24280_, _23591_, _42545_);
  nor (_23612_, _18826_, _18859_);
  and (_23623_, _18826_, _18859_);
  or (_23634_, _23623_, _23612_);
  and (_02351_, _23634_, _42545_);
  and (_23655_, _22525_, _19743_);
  and (_02542_, _23655_, _42545_);
  nor (_23676_, _22535_, _22188_);
  nor (_23687_, _23676_, _22546_);
  and (_02736_, _23687_, _42545_);
  nor (_23707_, _23188_, _23166_);
  nor (_23718_, _23707_, _23199_);
  and (_02964_, _23718_, _42545_);
  nor (_23739_, _23221_, _23199_);
  nor (_23750_, _23739_, _23232_);
  and (_03166_, _23750_, _42545_);
  nor (_23771_, _23275_, _23254_);
  nor (_23782_, _23771_, _23286_);
  and (_03371_, _23782_, _42545_);
  and (_23812_, _23297_, _23068_);
  nor (_23813_, _23812_, _23308_);
  and (_03603_, _23813_, _42545_);
  nor (_23834_, _23330_, _22992_);
  nor (_23845_, _23834_, _23341_);
  and (_03848_, _23845_, _42545_);
  nor (_23866_, _23363_, _22927_);
  nor (_23877_, _23866_, _23383_);
  and (_04074_, _23877_, _42545_);
  and (_23897_, _23417_, _23384_);
  nor (_23908_, _23897_, _23428_);
  and (_04170_, _23908_, _42545_);
  and (_23929_, _23439_, _22818_);
  nor (_23940_, _23929_, _23450_);
  and (_04270_, _23940_, _42545_);
  nor (_23961_, _23472_, _18968_);
  nor (_23971_, _23961_, _23482_);
  and (_04369_, _23971_, _42545_);
  and (_23992_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_24003_, _23992_, _23482_);
  nor (_24014_, _24003_, _23493_);
  and (_04468_, _24014_, _42545_);
  nor (_24035_, _23504_, _23493_);
  nor (_24046_, _24035_, _23515_);
  and (_04563_, _24046_, _42545_);
  and (_24066_, _18946_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_24077_, _24066_, _23515_);
  nor (_24088_, _24077_, _23526_);
  and (_04662_, _24088_, _42545_);
  nor (_24109_, _23526_, _18957_);
  nor (_24120_, _24109_, _23537_);
  and (_04760_, _24120_, _42545_);
  and (_24140_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18770_);
  nor (_24151_, _24140_, _18771_);
  not (_24162_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_24173_, _18793_, _24162_);
  and (_24184_, _24173_, _24151_);
  and (_24195_, _24184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24206_, _24195_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24216_, _24195_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24227_, _24216_, _24206_);
  and (_00925_, _24227_, _42545_);
  and (_00950_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _42545_);
  not (_24258_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_24269_, _20533_, _24258_);
  and (_24281_, _20217_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24292_, _24281_, _24269_);
  nor (_24302_, _24292_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24313_, _20370_, _24258_);
  and (_24324_, _20717_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24335_, _24324_, _24313_);
  and (_24346_, _24335_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24357_, _24346_, _24302_);
  nor (_24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24379_, _24368_, _20881_);
  nor (_24389_, _24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor (_24400_, _24389_, _24379_);
  not (_24411_, _24400_);
  and (_24422_, _19547_, _24258_);
  and (_24433_, _19220_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24444_, _24433_, _24422_);
  nor (_24455_, _24444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24465_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24476_, _19384_, _24258_);
  and (_24487_, _19721_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24498_, _24487_, _24476_);
  nor (_24519_, _24498_, _24465_);
  nor (_24520_, _24519_, _24455_);
  nor (_24531_, _24520_, _24411_);
  and (_24542_, _24520_, _24411_);
  nor (_24552_, _24542_, _24531_);
  nor (_24563_, _24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and (_24574_, _24368_, _20043_);
  nor (_24585_, _24574_, _24563_);
  not (_24596_, _24585_);
  nor (_24607_, _20533_, _24258_);
  nor (_24618_, _24607_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24629_, _20217_, _24258_);
  and (_24639_, _20370_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24650_, _24639_, _24629_);
  nor (_24661_, _24650_, _24465_);
  nor (_24672_, _24661_, _24618_);
  nor (_24683_, _24672_, _24596_);
  and (_24694_, _24672_, _24596_);
  nor (_24705_, _24694_, _24683_);
  not (_24715_, _24705_);
  nor (_24726_, _24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_24737_, _24368_, _21077_);
  nor (_24748_, _24737_, _24726_);
  not (_24759_, _24748_);
  nor (_24770_, _19547_, _24258_);
  nor (_24781_, _24770_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24792_, _19220_, _24258_);
  and (_24802_, _19384_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24813_, _24802_, _24792_);
  nor (_24824_, _24813_, _24465_);
  nor (_24835_, _24824_, _24781_);
  nor (_24846_, _24835_, _24759_);
  and (_24857_, _24835_, _24759_);
  and (_24868_, _24292_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24879_, _24868_);
  nor (_24889_, _24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_24900_, _24368_, _21251_);
  nor (_24911_, _24900_, _24889_);
  and (_24922_, _24911_, _24879_);
  and (_24933_, _24444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24944_, _24933_);
  and (_24955_, _24368_, _21621_);
  nor (_24966_, _24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_24976_, _24966_, _24955_);
  and (_24987_, _24976_, _24944_);
  nor (_24998_, _24976_, _24944_);
  nor (_25009_, _24998_, _24987_);
  not (_25020_, _25009_);
  and (_25031_, _24607_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_25042_, _25031_);
  and (_25063_, _24368_, _22144_);
  nor (_25064_, _24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_25075_, _25064_, _25063_);
  and (_25086_, _25075_, _25042_);
  and (_25097_, _24770_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_25108_, _25097_);
  nor (_25119_, _24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_25130_, _24368_, _21969_);
  nor (_25141_, _25130_, _25119_);
  nor (_25152_, _25141_, _25108_);
  not (_25163_, _25152_);
  nor (_25174_, _25075_, _25042_);
  nor (_25185_, _25174_, _25086_);
  and (_25196_, _25185_, _25163_);
  nor (_25207_, _25196_, _25086_);
  nor (_25218_, _25207_, _25020_);
  nor (_25229_, _25218_, _24987_);
  nor (_25239_, _24911_, _24879_);
  nor (_25250_, _25239_, _24922_);
  not (_25261_, _25250_);
  nor (_25272_, _25261_, _25229_);
  nor (_25283_, _25272_, _24922_);
  nor (_25294_, _25283_, _24857_);
  nor (_25305_, _25294_, _24846_);
  nor (_25326_, _25305_, _24715_);
  nor (_25327_, _25326_, _24683_);
  not (_25338_, _25327_);
  and (_25349_, _25338_, _24552_);
  or (_25360_, _25349_, _24531_);
  and (_25371_, _20717_, _19721_);
  or (_25382_, _25371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_25393_, _24498_);
  and (_25404_, _24335_, _25393_);
  nor (_25415_, _24813_, _24650_);
  and (_25426_, _25415_, _25404_);
  or (_25437_, _25426_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_25448_, _25437_, _25382_);
  and (_25459_, _25448_, _25360_);
  and (_25470_, _25459_, _24357_);
  nor (_25481_, _25338_, _24552_);
  or (_25492_, _25481_, _25349_);
  and (_25503_, _25492_, _25470_);
  nor (_25514_, _25470_, _24400_);
  nor (_25525_, _25514_, _25503_);
  not (_25536_, _25525_);
  and (_25547_, _25525_, _24357_);
  not (_25558_, _24520_);
  nor (_25569_, _25470_, _24596_);
  and (_25580_, _25305_, _24715_);
  nor (_25591_, _25580_, _25326_);
  and (_25602_, _25591_, _25470_);
  or (_25612_, _25602_, _25569_);
  and (_25633_, _25612_, _25558_);
  nor (_25634_, _25612_, _25558_);
  nor (_25645_, _25634_, _25633_);
  not (_25656_, _25645_);
  not (_25667_, _24672_);
  nor (_25678_, _25470_, _24759_);
  nor (_25689_, _24857_, _24846_);
  nor (_25700_, _25689_, _25283_);
  and (_25711_, _25689_, _25283_);
  or (_25722_, _25711_, _25700_);
  and (_25733_, _25722_, _25470_);
  or (_25744_, _25733_, _25678_);
  and (_25755_, _25744_, _25667_);
  nor (_25766_, _25744_, _25667_);
  not (_25777_, _24835_);
  and (_25788_, _25261_, _25229_);
  or (_25799_, _25788_, _25272_);
  and (_25810_, _25799_, _25470_);
  nor (_25821_, _25470_, _24911_);
  nor (_25832_, _25821_, _25810_);
  and (_25843_, _25832_, _25777_);
  and (_25854_, _25207_, _25020_);
  nor (_25865_, _25854_, _25218_);
  not (_25876_, _25865_);
  and (_25887_, _25876_, _25470_);
  nor (_25898_, _25470_, _24976_);
  nor (_25909_, _25898_, _25887_);
  and (_25920_, _25909_, _24879_);
  nor (_25931_, _25909_, _24879_);
  nor (_25942_, _25931_, _25920_);
  not (_25963_, _25942_);
  nor (_25964_, _25185_, _25163_);
  nor (_25974_, _25964_, _25196_);
  not (_25985_, _25974_);
  and (_25996_, _25985_, _25470_);
  nor (_26007_, _25470_, _25075_);
  nor (_26018_, _26007_, _25996_);
  and (_26029_, _26018_, _24944_);
  not (_26040_, _25141_);
  and (_26051_, _25470_, _25097_);
  or (_26062_, _26051_, _26040_);
  nand (_26073_, _25470_, _25097_);
  or (_26084_, _26073_, _25141_);
  and (_26095_, _26084_, _26062_);
  nor (_26106_, _26095_, _25031_);
  and (_26117_, _26095_, _25031_);
  nor (_26128_, _26117_, _26106_);
  and (_26139_, _24368_, _22514_);
  nor (_26150_, _24368_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_26161_, _26150_, _26139_);
  nor (_26172_, _26161_, _25108_);
  not (_26183_, _26172_);
  and (_26194_, _26183_, _26128_);
  nor (_26205_, _26194_, _26106_);
  nor (_26216_, _26018_, _24944_);
  nor (_26227_, _26216_, _26029_);
  not (_26238_, _26227_);
  nor (_26249_, _26238_, _26205_);
  nor (_26260_, _26249_, _26029_);
  nor (_26271_, _26260_, _25963_);
  nor (_26282_, _26271_, _25920_);
  nor (_26293_, _25832_, _25777_);
  nor (_26304_, _26293_, _25843_);
  not (_26314_, _26304_);
  nor (_26325_, _26314_, _26282_);
  nor (_26336_, _26325_, _25843_);
  nor (_26347_, _26336_, _25766_);
  nor (_26358_, _26347_, _25755_);
  nor (_26369_, _26358_, _25656_);
  or (_26380_, _26369_, _25633_);
  or (_26391_, _26380_, _25547_);
  and (_26402_, _26391_, _25448_);
  nor (_26413_, _26402_, _25536_);
  and (_26424_, _25547_, _25448_);
  and (_26445_, _26424_, _26380_);
  or (_26446_, _26445_, _26413_);
  and (_00968_, _26446_, _42545_);
  or (_26467_, _25525_, _24357_);
  and (_26478_, _26467_, _26402_);
  and (_02915_, _26478_, _42545_);
  and (_02928_, _25470_, _42545_);
  and (_02952_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _42545_);
  and (_02975_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _42545_);
  and (_02998_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _42545_);
  or (_26539_, _24184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_26550_, _24195_, rst);
  and (_03010_, _26550_, _26539_);
  not (_26571_, _26161_);
  and (_26582_, _26478_, _25097_);
  nor (_26593_, _26582_, _26571_);
  and (_26604_, _26582_, _26571_);
  or (_26615_, _26604_, _26593_);
  and (_03021_, _26615_, _42545_);
  nor (_26636_, _26478_, _26095_);
  nor (_26647_, _26183_, _26128_);
  nor (_26667_, _26647_, _26194_);
  and (_26668_, _26667_, _26478_);
  or (_26679_, _26668_, _26636_);
  and (_03034_, _26679_, _42545_);
  and (_26700_, _26238_, _26205_);
  or (_26711_, _26700_, _26249_);
  nand (_26722_, _26711_, _26478_);
  or (_26733_, _26478_, _26018_);
  and (_26744_, _26733_, _26722_);
  and (_03045_, _26744_, _42545_);
  and (_26765_, _26260_, _25963_);
  or (_26776_, _26765_, _26271_);
  nand (_26787_, _26776_, _26478_);
  or (_26798_, _26478_, _25909_);
  and (_26809_, _26798_, _26787_);
  and (_03058_, _26809_, _42545_);
  and (_26830_, _26314_, _26282_);
  or (_26841_, _26830_, _26325_);
  nand (_26852_, _26841_, _26478_);
  or (_26863_, _26478_, _25832_);
  and (_26874_, _26863_, _26852_);
  and (_03070_, _26874_, _42545_);
  or (_26895_, _25766_, _25755_);
  and (_26906_, _26895_, _26336_);
  nor (_26917_, _26895_, _26336_);
  or (_26928_, _26917_, _26906_);
  nand (_26939_, _26928_, _26478_);
  or (_26950_, _26478_, _25744_);
  and (_26961_, _26950_, _26939_);
  and (_03081_, _26961_, _42545_);
  and (_26982_, _26358_, _25656_);
  or (_26993_, _26982_, _26369_);
  nand (_27004_, _26993_, _26478_);
  or (_27014_, _26478_, _25612_);
  and (_27025_, _27014_, _27004_);
  and (_03091_, _27025_, _42545_);
  not (_27046_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27057_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18770_);
  and (_27068_, _27057_, _27046_);
  and (_27079_, _27068_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_27090_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_27101_, _27090_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_27112_, _27090_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_27123_, _27112_, _27101_);
  and (_27134_, _27123_, _27079_);
  not (_27145_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_27156_, _27068_, _27145_);
  and (_27167_, _27156_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_27178_, _27167_, _27134_);
  not (_27189_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_27200_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18770_);
  and (_27211_, _27200_, _27189_);
  and (_27222_, _27211_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27243_, _27222_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_27244_, _27211_, _27046_);
  and (_27255_, _27244_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_27266_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27277_, _27266_, _18770_);
  nor (_27288_, _27277_, _27200_);
  and (_27299_, _27288_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_27310_, _27299_, _27255_);
  nor (_27321_, _27310_, _27243_);
  and (_27332_, _27321_, _27178_);
  nor (_27343_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_27353_, _27343_, _27090_);
  and (_27364_, _27353_, _27079_);
  and (_27375_, _27156_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_27386_, _27375_, _27364_);
  and (_27397_, _27222_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_27408_, _27244_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_27419_, _27288_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_27430_, _27419_, _27408_);
  nor (_27441_, _27430_, _27397_);
  and (_27452_, _27441_, _27386_);
  and (_27463_, _27222_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_27474_, _27244_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_27485_, _27474_, _27463_);
  and (_27496_, _27156_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_27507_, _27496_);
  not (_27518_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_27529_, _27079_, _27518_);
  and (_27540_, _27288_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_27551_, _27540_, _27529_);
  and (_27562_, _27551_, _27507_);
  and (_27573_, _27562_, _27485_);
  and (_27584_, _27573_, _27452_);
  and (_27595_, _27584_, _27332_);
  and (_27606_, _27101_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_27617_, _27606_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_27628_, _27617_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_27639_, _27628_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_27650_, _27639_);
  not (_27661_, _27079_);
  nor (_27672_, _27628_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_27683_, _27672_, _27661_);
  and (_27694_, _27683_, _27650_);
  not (_27704_, _27694_);
  and (_27715_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27726_, _27715_, _27057_);
  and (_27737_, _27244_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_27748_, _27737_, _27726_);
  and (_27759_, _27156_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_27770_, _27222_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_27781_, _27770_, _27759_);
  and (_27792_, _27781_, _27748_);
  and (_27803_, _27792_, _27704_);
  nor (_27814_, _27617_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_27825_, _27814_);
  nor (_27836_, _27628_, _27661_);
  and (_27847_, _27836_, _27825_);
  not (_27858_, _27847_);
  and (_27879_, _27244_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_27880_, _27879_, _27726_);
  and (_27891_, _27156_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_27902_, _27222_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_27913_, _27902_, _27891_);
  and (_27924_, _27913_, _27880_);
  and (_27935_, _27924_, _27858_);
  nor (_27946_, _27935_, _27803_);
  not (_27957_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_27968_, _27639_, _27957_);
  and (_27979_, _27639_, _27957_);
  nor (_27990_, _27979_, _27968_);
  nor (_28001_, _27990_, _27661_);
  not (_28012_, _28001_);
  and (_28023_, _27156_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nor (_28033_, _27726_, _28023_);
  and (_28044_, _27222_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and (_28055_, _27244_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_28066_, _28055_, _28044_);
  and (_28077_, _28066_, _28033_);
  and (_28088_, _28077_, _28012_);
  not (_28099_, _28088_);
  not (_28110_, _27606_);
  nor (_28121_, _27101_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_28132_, _28121_, _27661_);
  and (_28143_, _28132_, _28110_);
  not (_28154_, _28143_);
  and (_28165_, _27288_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_28186_, _27156_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_28187_, _28186_, _28165_);
  and (_28198_, _27222_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_28209_, _27244_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_28220_, _28209_, _28198_);
  and (_28231_, _28220_, _28187_);
  and (_28242_, _28231_, _28154_);
  not (_28253_, _28242_);
  and (_28264_, _27222_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_28275_, _28264_);
  and (_28286_, _27156_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_28297_, _28286_, _27726_);
  and (_28308_, _28297_, _28275_);
  nor (_28319_, _27606_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_28330_, _28319_);
  nor (_28341_, _27617_, _27661_);
  and (_28351_, _28341_, _28330_);
  and (_28362_, _27288_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_28373_, _27244_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_28384_, _28373_, _28362_);
  not (_28395_, _28384_);
  nor (_28406_, _28395_, _28351_);
  and (_28417_, _28406_, _28308_);
  nor (_28428_, _28417_, _28253_);
  and (_28439_, _28428_, _28099_);
  and (_28450_, _28439_, _27946_);
  nand (_28461_, _28450_, _27595_);
  and (_28472_, _26446_, _24184_);
  and (_28483_, _23591_, _18826_);
  nor (_28494_, _20043_, _19721_);
  and (_28505_, _20043_, _19721_);
  nor (_28516_, _28505_, _28494_);
  not (_28537_, _28516_);
  nor (_28538_, _21077_, _20370_);
  nor (_28549_, _21251_, _19384_);
  and (_28560_, _21077_, _20370_);
  nor (_28571_, _28560_, _28538_);
  and (_28582_, _28571_, _28549_);
  nor (_28593_, _28582_, _28538_);
  nor (_28604_, _28593_, _28537_);
  and (_28615_, _21251_, _19384_);
  nor (_28626_, _28615_, _28549_);
  nor (_28637_, _21621_, _20217_);
  and (_28648_, _21621_, _20217_);
  nor (_28658_, _28648_, _28637_);
  nor (_28669_, _22144_, _19220_);
  and (_28680_, _22144_, _19220_);
  nor (_28691_, _28680_, _28669_);
  not (_28702_, _28691_);
  nor (_28713_, _21969_, _20533_);
  nor (_28724_, _22514_, _19547_);
  and (_28735_, _21969_, _20533_);
  nor (_28746_, _28735_, _28713_);
  and (_28757_, _28746_, _28724_);
  nor (_28768_, _28757_, _28713_);
  nor (_28779_, _28768_, _28702_);
  nor (_28790_, _28779_, _28669_);
  nor (_28801_, _28790_, _28658_);
  and (_28812_, _28790_, _28658_);
  nor (_28823_, _28812_, _28801_);
  not (_28834_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_28845_, _19033_, _28834_);
  not (_28856_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_28867_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28878_, _28867_, _20598_);
  nor (_28889_, _28878_, _28856_);
  nor (_28910_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28911_, _28910_, _19275_);
  not (_28922_, _28911_);
  not (_28933_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_28944_, _28933_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28955_, _28944_, _19613_);
  not (_28965_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28976_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _28965_);
  and (_28987_, _28976_, _20261_);
  nor (_28998_, _28987_, _28955_);
  and (_29009_, _28998_, _28922_);
  and (_29020_, _29009_, _28889_);
  and (_29031_, _28867_, _20109_);
  nor (_29042_, _29031_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_29053_, _28976_, _20424_);
  not (_29064_, _29053_);
  and (_29075_, _28944_, _19077_);
  and (_29086_, _28910_, _19439_);
  nor (_29097_, _29086_, _29075_);
  and (_29108_, _29097_, _29064_);
  and (_29119_, _29108_, _29042_);
  nor (_29130_, _29119_, _29020_);
  nor (_29141_, _29130_, _19033_);
  nor (_29152_, _29141_, _28845_);
  and (_29163_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_29174_, _29163_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_29185_, _29174_);
  and (_29196_, _29185_, _29152_);
  and (_29207_, _29185_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_29218_, _29207_, _29196_);
  and (_29229_, _22514_, _19547_);
  nor (_29240_, _29229_, _28724_);
  not (_29251_, _29240_);
  nor (_29262_, _29251_, _29218_);
  and (_29272_, _29262_, _28746_);
  and (_29283_, _28768_, _28702_);
  nor (_29294_, _29283_, _28779_);
  and (_29305_, _29294_, _29272_);
  not (_29316_, _29305_);
  nor (_29327_, _29316_, _28823_);
  nor (_29338_, _28790_, _28648_);
  or (_29349_, _29338_, _28637_);
  or (_29360_, _29349_, _29327_);
  and (_29371_, _29360_, _28626_);
  nor (_29382_, _28571_, _28549_);
  nor (_29393_, _29382_, _28582_);
  and (_29404_, _29393_, _29371_);
  and (_29415_, _28593_, _28537_);
  nor (_29436_, _29415_, _28604_);
  and (_29437_, _29436_, _29404_);
  or (_29448_, _29437_, _28604_);
  nor (_29459_, _29448_, _28494_);
  nor (_29470_, _20881_, _20717_);
  and (_29481_, _20881_, _20717_);
  nor (_29492_, _29481_, _29470_);
  not (_29503_, _29492_);
  nor (_29514_, _29503_, _29459_);
  not (_29525_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_29536_, _24140_, _29525_);
  and (_29547_, _29536_, _18815_);
  nand (_29558_, _29503_, _29459_);
  nand (_29569_, _29558_, _29547_);
  nor (_29579_, _29569_, _29514_);
  not (_29590_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_29601_, _18771_, _29590_);
  and (_29612_, _29601_, _18815_);
  not (_29623_, _29612_);
  not (_29634_, _19721_);
  nor (_29645_, _20043_, _29634_);
  and (_29656_, _21088_, _20370_);
  not (_29667_, _19384_);
  and (_29678_, _21251_, _29667_);
  nor (_29689_, _29678_, _28571_);
  nor (_29710_, _29689_, _29656_);
  nor (_29711_, _29710_, _28516_);
  nor (_29722_, _29711_, _29645_);
  and (_29733_, _29710_, _28516_);
  nor (_29744_, _29733_, _29711_);
  not (_29755_, _29744_);
  and (_29766_, _29678_, _28571_);
  nor (_29777_, _29766_, _29689_);
  not (_29788_, _29777_);
  not (_29799_, _28626_);
  not (_29810_, _19547_);
  and (_29821_, _22514_, _29810_);
  nor (_29832_, _29821_, _28746_);
  not (_29843_, _20533_);
  nor (_29854_, _21969_, _29843_);
  nor (_29865_, _29854_, _29832_);
  nor (_29876_, _29865_, _28691_);
  not (_29886_, _19220_);
  nor (_29897_, _22144_, _29886_);
  nor (_29908_, _29897_, _29876_);
  nor (_29919_, _29908_, _28658_);
  and (_29930_, _29908_, _28658_);
  nor (_29941_, _29930_, _29919_);
  not (_29952_, _29941_);
  and (_29963_, _29865_, _28691_);
  nor (_29974_, _29963_, _29876_);
  not (_29984_, _29974_);
  and (_29995_, _29821_, _28746_);
  nor (_30006_, _29995_, _29832_);
  not (_30017_, _30006_);
  nor (_30028_, _29240_, _29218_);
  and (_30039_, _30028_, _30017_);
  and (_30050_, _30039_, _29984_);
  and (_30061_, _30050_, _29952_);
  not (_30072_, _20217_);
  or (_30083_, _21621_, _30072_);
  and (_30094_, _21621_, _30072_);
  or (_30104_, _29908_, _30094_);
  and (_30115_, _30104_, _30083_);
  or (_30126_, _30115_, _30061_);
  and (_30137_, _30126_, _29799_);
  and (_30148_, _30137_, _29788_);
  and (_30159_, _30148_, _29755_);
  nor (_30170_, _30159_, _29722_);
  nor (_30181_, _30170_, _29492_);
  and (_30192_, _30170_, _29492_);
  nor (_30203_, _30192_, _30181_);
  nor (_30213_, _30203_, _29623_);
  and (_30224_, _18804_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30235_, _30224_, _29601_);
  nor (_30246_, _22514_, _21969_);
  and (_30257_, _30246_, _22155_);
  and (_30268_, _30257_, _21632_);
  and (_30279_, _30268_, _21262_);
  and (_30290_, _30279_, _21088_);
  and (_30301_, _30290_, _20054_);
  and (_30312_, _30301_, _29218_);
  not (_30332_, _29218_);
  and (_30333_, _21077_, _20043_);
  and (_30344_, _22514_, _21969_);
  and (_30355_, _30344_, _22144_);
  and (_30366_, _30355_, _21621_);
  and (_30377_, _30366_, _21251_);
  and (_30388_, _30377_, _30333_);
  and (_30399_, _30388_, _30332_);
  nor (_30410_, _30399_, _30312_);
  and (_30421_, _30410_, _20881_);
  nor (_30431_, _30410_, _20881_);
  nor (_30442_, _30431_, _30421_);
  and (_30453_, _30442_, _30235_);
  not (_30464_, _20717_);
  nor (_30475_, _29218_, _30464_);
  not (_30486_, _30475_);
  and (_30497_, _29218_, _20881_);
  and (_30508_, _30224_, _18782_);
  not (_30519_, _30508_);
  nor (_30530_, _30519_, _30497_);
  and (_30540_, _30530_, _30486_);
  nor (_30551_, _30540_, _30453_);
  and (_30562_, _29536_, _24173_);
  and (_30573_, _22144_, _21969_);
  nor (_30584_, _30573_, _21621_);
  and (_30595_, _30584_, _30562_);
  and (_30606_, _30595_, _21262_);
  nor (_30617_, _30606_, _21088_);
  and (_30628_, _30617_, _20043_);
  nor (_30639_, _30333_, _20881_);
  nor (_30650_, _30639_, _30595_);
  and (_30660_, _30650_, _29218_);
  nor (_30671_, _30660_, _30628_);
  and (_30682_, _30671_, _20881_);
  nor (_30693_, _30671_, _20881_);
  or (_30704_, _30693_, _30682_);
  and (_30715_, _30704_, _30562_);
  and (_30726_, _30224_, _29536_);
  not (_30737_, _30726_);
  nor (_30748_, _30737_, _29218_);
  not (_30758_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30769_, _18804_, _30758_);
  and (_30780_, _30769_, _29536_);
  not (_30791_, _30780_);
  nor (_30802_, _30791_, _29481_);
  and (_30813_, _30769_, _24151_);
  and (_30824_, _30813_, _29492_);
  nor (_30835_, _30824_, _30802_);
  and (_30846_, _24173_, _18782_);
  and (_30857_, _30846_, _29470_);
  and (_30868_, _29601_, _24173_);
  and (_30878_, _30868_, _20881_);
  nor (_30889_, _30878_, _30857_);
  and (_30900_, _30224_, _24151_);
  not (_30911_, _30900_);
  nor (_30922_, _30911_, _22514_);
  and (_30933_, _24151_, _18815_);
  not (_30944_, _30933_);
  nor (_30955_, _30944_, _20881_);
  and (_30966_, _30769_, _18771_);
  not (_30977_, _30966_);
  nor (_30987_, _30977_, _20043_);
  or (_30998_, _30987_, _30955_);
  nor (_31009_, _30998_, _30922_);
  and (_31020_, _31009_, _30889_);
  nand (_31042_, _31020_, _30835_);
  or (_31043_, _31042_, _30748_);
  nor (_31065_, _31043_, _30715_);
  nand (_31066_, _31065_, _30551_);
  or (_31088_, _31066_, _30213_);
  or (_31089_, _31088_, _29579_);
  or (_31110_, _31089_, _28483_);
  or (_31111_, _31110_, _28472_);
  or (_31122_, _31111_, _28461_);
  not (_31133_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31144_, \oc8051_top_1.oc8051_decoder1.wr , _18770_);
  not (_31165_, _31144_);
  nor (_31166_, _31165_, _27068_);
  and (_31187_, _31166_, _31133_);
  not (_31188_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_31208_, _28461_, _31188_);
  and (_31209_, _31208_, _31187_);
  and (_31230_, _31209_, _31122_);
  nor (_31231_, _31166_, _31188_);
  not (_31252_, _29547_);
  nor (_31253_, _29514_, _29470_);
  nor (_31274_, _31253_, _31252_);
  not (_31275_, _31274_);
  and (_31296_, _20881_, _30464_);
  nor (_31297_, _31296_, _30181_);
  nor (_31317_, _31297_, _29623_);
  and (_31318_, _29218_, _20043_);
  and (_31339_, _31318_, _30617_);
  nor (_31340_, _31339_, _30497_);
  not (_31361_, _30562_);
  nor (_31362_, _29218_, _20881_);
  not (_31383_, _31362_);
  nor (_31384_, _31383_, _30628_);
  nor (_31405_, _31384_, _31361_);
  and (_31406_, _31405_, _31340_);
  and (_31427_, _29174_, _29152_);
  and (_31428_, _30769_, _29601_);
  and (_31448_, _30846_, _29152_);
  nor (_31449_, _31448_, _31428_);
  nor (_31470_, _31449_, _31427_);
  nor (_31471_, _30944_, _29218_);
  and (_31492_, _30769_, _18782_);
  not (_31493_, _31492_);
  nor (_31514_, _31493_, _20881_);
  nor (_31515_, _30737_, _22514_);
  or (_31535_, _31515_, _30595_);
  or (_31536_, _31535_, _31514_);
  or (_31557_, _31536_, _31471_);
  nor (_31558_, _29207_, _29152_);
  not (_31579_, _30813_);
  nor (_31580_, _31579_, _29196_);
  nor (_31601_, _31580_, _30780_);
  nor (_31602_, _31601_, _31558_);
  nor (_31623_, _30911_, _29152_);
  or (_31624_, _31623_, _29218_);
  or (_31645_, _30868_, _30332_);
  and (_31646_, _31645_, _31624_);
  or (_31666_, _31646_, _31602_);
  or (_31667_, _31666_, _31557_);
  or (_31688_, _31667_, _31470_);
  nor (_31689_, _31688_, _31406_);
  not (_31710_, _31689_);
  nor (_31711_, _31710_, _31317_);
  and (_31732_, _31711_, _31275_);
  not (_31733_, _27332_);
  nor (_31754_, _27573_, _27452_);
  and (_31755_, _31754_, _31733_);
  and (_31765_, _31755_, _28450_);
  nand (_31776_, _31765_, _31732_);
  or (_31787_, _31765_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_31798_, _31166_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31809_, _31798_, _31787_);
  and (_31820_, _31809_, _31776_);
  or (_31831_, _31820_, _31231_);
  or (_31842_, _31831_, _31230_);
  and (_06624_, _31842_, _42545_);
  and (_31863_, _26615_, _24184_);
  not (_31873_, _31863_);
  and (_31884_, _23908_, _18826_);
  and (_31895_, _29251_, _29218_);
  nor (_31906_, _31895_, _29262_);
  nor (_31917_, _29612_, _29547_);
  not (_31928_, _31917_);
  and (_31939_, _31928_, _31906_);
  not (_31950_, _31939_);
  nor (_31961_, _31493_, _29218_);
  not (_31972_, _31961_);
  nor (_31982_, _31579_, _28724_);
  nor (_31993_, _31982_, _30780_);
  or (_32004_, _31993_, _29229_);
  and (_32015_, _30846_, _28724_);
  and (_32026_, _30868_, _22514_);
  nor (_32037_, _32026_, _32015_);
  nor (_32048_, _30519_, _19547_);
  and (_32059_, _30235_, _22514_);
  nor (_32070_, _32059_, _32048_);
  and (_32081_, _30224_, _29525_);
  not (_32093_, _32081_);
  nor (_32112_, _32093_, _21969_);
  not (_32123_, _32112_);
  and (_32134_, _31428_, _20892_);
  nor (_32145_, _30933_, _30562_);
  nor (_32156_, _32145_, _22514_);
  nor (_32167_, _32156_, _32134_);
  and (_32178_, _32167_, _32123_);
  and (_32189_, _32178_, _32070_);
  and (_32200_, _32189_, _32037_);
  and (_32211_, _32200_, _32004_);
  and (_32221_, _32211_, _31972_);
  and (_32232_, _32221_, _31950_);
  not (_32243_, _32232_);
  nor (_32254_, _32243_, _31884_);
  and (_32265_, _32254_, _31873_);
  not (_32276_, _32265_);
  or (_32287_, _32276_, _28461_);
  not (_32298_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_32309_, _28461_, _32298_);
  and (_32319_, _32309_, _31187_);
  and (_32330_, _32319_, _32287_);
  nor (_32341_, _31166_, _32298_);
  not (_32352_, _31732_);
  or (_32363_, _32352_, _28461_);
  and (_32374_, _32309_, _31798_);
  and (_32385_, _32374_, _32363_);
  or (_32396_, _32385_, _32341_);
  or (_32407_, _32396_, _32330_);
  and (_08891_, _32407_, _42545_);
  and (_32427_, _23940_, _18826_);
  not (_32438_, _32427_);
  and (_32449_, _26679_, _24184_);
  nor (_32460_, _30519_, _20533_);
  nor (_32471_, _30344_, _30246_);
  not (_32482_, _32471_);
  nor (_32493_, _32482_, _29218_);
  and (_32504_, _32482_, _29218_);
  nor (_32515_, _32504_, _32493_);
  and (_32526_, _32515_, _30235_);
  nor (_32537_, _32526_, _32460_);
  nor (_32547_, _30944_, _21969_);
  nor (_32558_, _32093_, _22144_);
  nor (_32569_, _30977_, _22514_);
  or (_32580_, _32569_, _32558_);
  nor (_32591_, _32580_, _32547_);
  and (_32602_, _30846_, _28713_);
  and (_32613_, _30868_, _21969_);
  nor (_32624_, _32613_, _32602_);
  and (_32635_, _32624_, _32591_);
  nor (_32646_, _30584_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_32656_, _32646_, _21980_);
  nor (_32667_, _32646_, _21980_);
  nor (_32678_, _32667_, _32656_);
  nor (_32689_, _32678_, _31361_);
  and (_32700_, _30813_, _28746_);
  nor (_32711_, _30791_, _28735_);
  or (_32722_, _32711_, _32700_);
  nor (_32733_, _32722_, _32689_);
  and (_32744_, _32733_, _32635_);
  and (_32755_, _32744_, _32537_);
  nor (_32765_, _28746_, _28724_);
  or (_32776_, _32765_, _28757_);
  and (_32787_, _32776_, _29262_);
  nor (_32798_, _32776_, _29262_);
  or (_32809_, _32798_, _32787_);
  and (_32820_, _32809_, _29547_);
  nor (_32831_, _30028_, _30017_);
  nor (_32842_, _32831_, _30039_);
  nor (_32853_, _32842_, _29623_);
  nor (_32864_, _32853_, _32820_);
  and (_32874_, _32864_, _32755_);
  not (_32885_, _32874_);
  nor (_32896_, _32885_, _32449_);
  and (_32907_, _32896_, _32438_);
  not (_32918_, _32907_);
  or (_32929_, _32918_, _28461_);
  not (_32940_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_32951_, _28461_, _32940_);
  and (_32962_, _32951_, _31187_);
  and (_32973_, _32962_, _32929_);
  nor (_32983_, _31166_, _32940_);
  not (_32994_, _27452_);
  nor (_33005_, _27573_, _32994_);
  and (_33016_, _33005_, _27332_);
  and (_33027_, _33016_, _28450_);
  nand (_33038_, _33027_, _31732_);
  or (_33049_, _33027_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_33060_, _33049_, _31798_);
  and (_33071_, _33060_, _33038_);
  or (_33082_, _33071_, _32983_);
  or (_33092_, _33082_, _32973_);
  and (_08902_, _33092_, _42545_);
  and (_33113_, _23971_, _18826_);
  not (_33124_, _33113_);
  and (_33135_, _26744_, _24184_);
  nor (_33146_, _30519_, _19220_);
  and (_33157_, _30344_, _30332_);
  and (_33168_, _30246_, _29218_);
  nor (_33179_, _33168_, _33157_);
  nor (_33190_, _33179_, _22144_);
  not (_33200_, _30235_);
  and (_33211_, _33179_, _22144_);
  or (_33222_, _33211_, _33200_);
  nor (_33233_, _33222_, _33190_);
  nor (_33244_, _33233_, _33146_);
  nor (_33255_, _30039_, _29984_);
  nor (_33266_, _33255_, _30050_);
  nor (_33277_, _33266_, _29623_);
  not (_33288_, _33277_);
  nor (_33299_, _32093_, _21621_);
  and (_33310_, _30846_, _28669_);
  and (_33320_, _30868_, _22144_);
  nor (_33331_, _33320_, _33310_);
  nor (_33342_, _30791_, _28680_);
  and (_33353_, _30813_, _28691_);
  nor (_33364_, _33353_, _33342_);
  nor (_33375_, _30977_, _21969_);
  nor (_33386_, _30944_, _22144_);
  nor (_33397_, _33386_, _33375_);
  and (_33408_, _33397_, _33364_);
  nand (_33419_, _33408_, _33331_);
  nor (_33429_, _33419_, _33299_);
  and (_33440_, _33429_, _33288_);
  nor (_33451_, _29294_, _29272_);
  nor (_33462_, _33451_, _31252_);
  and (_33473_, _33462_, _29316_);
  nor (_33484_, _32667_, _22144_);
  and (_33495_, _30573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_33506_, _33495_, _33484_);
  nor (_33517_, _33506_, _31361_);
  nor (_33528_, _33517_, _33473_);
  and (_33538_, _33528_, _33440_);
  and (_33549_, _33538_, _33244_);
  not (_33560_, _33549_);
  nor (_33571_, _33560_, _33135_);
  and (_33582_, _33571_, _33124_);
  not (_33593_, _33582_);
  or (_33604_, _33593_, _28461_);
  not (_33615_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_33626_, _28461_, _33615_);
  and (_33637_, _33626_, _31187_);
  and (_33647_, _33637_, _33604_);
  nor (_33658_, _31166_, _33615_);
  nand (_33669_, _28450_, _27332_);
  or (_33680_, _31754_, _33669_);
  and (_33691_, _33680_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_33702_, _27332_, _27573_);
  and (_33713_, _33702_, _32994_);
  not (_33724_, _33713_);
  nor (_33735_, _33724_, _31732_);
  and (_33746_, _27332_, _27452_);
  and (_33756_, _33746_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_33767_, _33756_, _33735_);
  and (_33778_, _33767_, _28450_);
  or (_33789_, _33778_, _33691_);
  and (_33800_, _33789_, _31798_);
  or (_33811_, _33800_, _33658_);
  or (_33822_, _33811_, _33647_);
  and (_08913_, _33822_, _42545_);
  and (_33843_, _24014_, _18826_);
  not (_33854_, _33843_);
  and (_33864_, _26809_, _24184_);
  nor (_33875_, _30050_, _29952_);
  nor (_33886_, _33875_, _30061_);
  nor (_33897_, _33886_, _29623_);
  not (_33908_, _33897_);
  nor (_33919_, _30791_, _28648_);
  and (_33930_, _30813_, _28658_);
  nor (_33941_, _33930_, _33919_);
  and (_33952_, _29316_, _28823_);
  or (_33963_, _33952_, _31252_);
  nor (_33973_, _33963_, _29327_);
  nor (_33984_, _30519_, _20217_);
  nor (_33995_, _30355_, _29218_);
  nor (_34006_, _30257_, _30332_);
  nor (_34017_, _34006_, _33995_);
  and (_34028_, _34017_, _21632_);
  not (_34039_, _34028_);
  nor (_34050_, _34017_, _21632_);
  nor (_34061_, _34050_, _33200_);
  and (_34072_, _34061_, _34039_);
  nor (_34083_, _34072_, _33984_);
  nor (_34093_, _30977_, _22144_);
  nor (_34104_, _30944_, _21621_);
  nor (_34115_, _34104_, _34093_);
  not (_34126_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_34137_, _30573_, _34126_);
  nor (_34148_, _34137_, _21632_);
  or (_34159_, _34148_, _31361_);
  nor (_34170_, _34159_, _30584_);
  and (_34181_, _30846_, _28637_);
  and (_34192_, _30868_, _21621_);
  nor (_34202_, _34192_, _34181_);
  nor (_34213_, _32093_, _21251_);
  not (_34224_, _34213_);
  nand (_34235_, _34224_, _34202_);
  nor (_34246_, _34235_, _34170_);
  and (_34257_, _34246_, _34115_);
  nand (_34268_, _34257_, _34083_);
  nor (_34279_, _34268_, _33973_);
  and (_34290_, _34279_, _33941_);
  and (_34301_, _34290_, _33908_);
  not (_34311_, _34301_);
  nor (_34322_, _34311_, _33864_);
  and (_34333_, _34322_, _33854_);
  not (_34344_, _34333_);
  or (_34355_, _34344_, _28461_);
  not (_34366_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_34377_, _28461_, _34366_);
  and (_34388_, _34377_, _31187_);
  and (_34399_, _34388_, _34355_);
  nor (_34410_, _31166_, _34366_);
  and (_34420_, _33669_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_34431_, _31754_, _27332_);
  not (_34442_, _34431_);
  nor (_34453_, _34442_, _31732_);
  nor (_34464_, _33746_, _33702_);
  nor (_34475_, _34464_, _34366_);
  or (_34486_, _34475_, _34453_);
  and (_34497_, _34486_, _28450_);
  or (_34508_, _34497_, _34420_);
  and (_34519_, _34508_, _31798_);
  or (_34529_, _34519_, _34410_);
  or (_34540_, _34529_, _34399_);
  and (_08924_, _34540_, _42545_);
  and (_34561_, _26874_, _24184_);
  not (_34572_, _34561_);
  and (_34583_, _24046_, _18826_);
  nor (_34594_, _30126_, _28626_);
  and (_34605_, _30126_, _28626_);
  nor (_34616_, _34605_, _34594_);
  and (_34627_, _34616_, _29612_);
  not (_34637_, _34627_);
  nor (_34648_, _29360_, _28626_);
  not (_34659_, _34648_);
  nor (_34670_, _31252_, _29371_);
  and (_34681_, _34670_, _34659_);
  and (_34692_, _29218_, _21262_);
  nor (_34703_, _29218_, _19384_);
  or (_34714_, _34703_, _34692_);
  and (_34725_, _34714_, _30508_);
  and (_34736_, _30268_, _29218_);
  and (_34746_, _30366_, _30332_);
  nor (_34757_, _34746_, _34736_);
  nor (_34768_, _34757_, _21251_);
  not (_34779_, _34768_);
  and (_34790_, _34757_, _21251_);
  nor (_34801_, _34790_, _33200_);
  and (_34812_, _34801_, _34779_);
  nor (_34823_, _34812_, _34725_);
  nor (_34834_, _30595_, _21262_);
  not (_34845_, _34834_);
  nor (_34856_, _30606_, _31361_);
  and (_34866_, _34856_, _34845_);
  not (_34877_, _34866_);
  and (_34888_, _30813_, _28626_);
  nor (_34899_, _30791_, _28615_);
  not (_34910_, _34899_);
  and (_34921_, _30846_, _28549_);
  and (_34932_, _30868_, _21251_);
  nor (_34943_, _34932_, _34921_);
  nand (_34954_, _34943_, _34910_);
  nor (_34965_, _34954_, _34888_);
  nor (_34975_, _32093_, _21077_);
  not (_34986_, _34975_);
  nor (_34997_, _30944_, _21251_);
  nor (_35008_, _30977_, _21621_);
  nor (_35019_, _35008_, _34997_);
  and (_35030_, _35019_, _34986_);
  and (_35041_, _35030_, _34965_);
  and (_35052_, _35041_, _34877_);
  and (_35063_, _35052_, _34823_);
  not (_35074_, _35063_);
  nor (_35084_, _35074_, _34681_);
  and (_35095_, _35084_, _34637_);
  not (_35106_, _35095_);
  nor (_35117_, _35106_, _34583_);
  and (_35128_, _35117_, _34572_);
  not (_35139_, _35128_);
  or (_35150_, _35139_, _28461_);
  not (_35161_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_35172_, _28461_, _35161_);
  and (_35183_, _35172_, _31187_);
  and (_35193_, _35183_, _35150_);
  nor (_35204_, _31166_, _35161_);
  not (_35215_, _28450_);
  and (_35226_, _27584_, _31733_);
  nor (_35237_, _27584_, _31733_);
  nor (_35248_, _35237_, _35226_);
  or (_35259_, _35248_, _35215_);
  and (_35270_, _35259_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_35281_, _35226_, _32352_);
  and (_35292_, _35237_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_35302_, _35292_, _35281_);
  and (_35313_, _35302_, _28450_);
  or (_35324_, _35313_, _35270_);
  and (_35335_, _35324_, _31798_);
  or (_35346_, _35335_, _35204_);
  or (_35357_, _35346_, _35193_);
  and (_08935_, _35357_, _42545_);
  and (_35378_, _26961_, _24184_);
  not (_35388_, _35378_);
  and (_35399_, _24088_, _18826_);
  nor (_35410_, _29393_, _29371_);
  nor (_35421_, _35410_, _29404_);
  and (_35432_, _35421_, _29547_);
  not (_35443_, _35432_);
  nor (_35454_, _30137_, _29788_);
  nor (_35465_, _35454_, _30148_);
  nor (_35476_, _35465_, _29623_);
  nor (_35487_, _29218_, _20370_);
  and (_35497_, _29218_, _21088_);
  nor (_35508_, _35497_, _35487_);
  nor (_35519_, _35508_, _30519_);
  nor (_35530_, _30279_, _30332_);
  nor (_35541_, _30377_, _29218_);
  nor (_35552_, _35541_, _35530_);
  nor (_35563_, _35552_, _21088_);
  not (_35574_, _35563_);
  and (_35585_, _35552_, _21088_);
  nor (_35596_, _35585_, _33200_);
  and (_35607_, _35596_, _35574_);
  nor (_35617_, _35607_, _35519_);
  not (_35628_, _30660_);
  and (_35639_, _35628_, _30617_);
  nor (_35650_, _30660_, _30606_);
  nor (_35661_, _35650_, _21077_);
  nor (_35672_, _35661_, _35639_);
  nor (_35683_, _35672_, _31361_);
  and (_35694_, _30813_, _28571_);
  not (_35705_, _35694_);
  nor (_35716_, _30791_, _28560_);
  not (_35727_, _35716_);
  and (_35737_, _30846_, _28538_);
  and (_35748_, _30868_, _21077_);
  nor (_35759_, _35748_, _35737_);
  and (_35770_, _35759_, _35727_);
  and (_35781_, _35770_, _35705_);
  nor (_35792_, _32093_, _20043_);
  not (_35803_, _35792_);
  nor (_35814_, _30944_, _21077_);
  nor (_35825_, _30977_, _21251_);
  nor (_35836_, _35825_, _35814_);
  and (_35847_, _35836_, _35803_);
  and (_35858_, _35847_, _35781_);
  not (_35868_, _35858_);
  nor (_35879_, _35868_, _35683_);
  and (_35890_, _35879_, _35617_);
  not (_35901_, _35890_);
  nor (_35912_, _35901_, _35476_);
  and (_35923_, _35912_, _35443_);
  not (_35934_, _35923_);
  nor (_35945_, _35934_, _35399_);
  and (_35956_, _35945_, _35388_);
  not (_35967_, _35956_);
  or (_35978_, _35967_, _28461_);
  not (_35988_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_35999_, _28461_, _35988_);
  and (_36010_, _35999_, _31187_);
  and (_36021_, _36010_, _35978_);
  nor (_36032_, _31166_, _35988_);
  and (_36043_, _33005_, _31733_);
  and (_36054_, _36043_, _28450_);
  nand (_36065_, _36054_, _31732_);
  or (_36076_, _36054_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_36087_, _36076_, _31798_);
  and (_36098_, _36087_, _36065_);
  or (_36109_, _36098_, _36032_);
  or (_36119_, _36109_, _36021_);
  and (_08946_, _36119_, _42545_);
  and (_36140_, _27025_, _24184_);
  not (_36151_, _36140_);
  and (_36162_, _24120_, _18826_);
  nor (_36173_, _29436_, _29404_);
  not (_36184_, _36173_);
  nor (_36194_, _31252_, _29437_);
  and (_36205_, _36194_, _36184_);
  not (_36216_, _36205_);
  nor (_36227_, _30148_, _29755_);
  nor (_36238_, _36227_, _30159_);
  nor (_36249_, _36238_, _29623_);
  nor (_36260_, _29218_, _29634_);
  or (_36271_, _36260_, _30519_);
  nor (_36281_, _36271_, _31318_);
  nor (_36292_, _29218_, _21088_);
  nand (_36303_, _36292_, _30377_);
  nand (_36314_, _30290_, _29218_);
  and (_36325_, _36314_, _36303_);
  and (_36336_, _36325_, _20043_);
  nor (_36347_, _36325_, _20043_);
  or (_36358_, _36347_, _33200_);
  nor (_36368_, _36358_, _36336_);
  nor (_36379_, _36368_, _36281_);
  nor (_36390_, _35639_, _20043_);
  and (_36401_, _35639_, _20043_);
  nor (_36412_, _36401_, _36390_);
  nor (_36423_, _36412_, _31361_);
  and (_36434_, _30813_, _28516_);
  nor (_36445_, _30791_, _28505_);
  not (_36455_, _36445_);
  and (_36466_, _30846_, _28494_);
  and (_36477_, _30868_, _20043_);
  nor (_36488_, _36477_, _36466_);
  nand (_36499_, _36488_, _36455_);
  nor (_36510_, _36499_, _36434_);
  nor (_36521_, _32093_, _20881_);
  not (_36531_, _36521_);
  nor (_36542_, _30944_, _20043_);
  nor (_36553_, _30977_, _21077_);
  nor (_36564_, _36553_, _36542_);
  and (_36575_, _36564_, _36531_);
  and (_36586_, _36575_, _36510_);
  not (_36597_, _36586_);
  nor (_36608_, _36597_, _36423_);
  and (_36618_, _36608_, _36379_);
  not (_36629_, _36618_);
  nor (_36640_, _36629_, _36249_);
  and (_36651_, _36640_, _36216_);
  not (_36662_, _36651_);
  nor (_36673_, _36662_, _36162_);
  and (_36684_, _36673_, _36151_);
  not (_36695_, _36684_);
  or (_36705_, _36695_, _28461_);
  not (_36716_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_36727_, _28461_, _36716_);
  and (_36738_, _36727_, _31187_);
  and (_36749_, _36738_, _36705_);
  nor (_36760_, _31166_, _36716_);
  nor (_36771_, _27332_, _27452_);
  and (_36782_, _36771_, _27573_);
  and (_36793_, _36782_, _28450_);
  nand (_36804_, _36793_, _31732_);
  or (_36814_, _36793_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_36825_, _36814_, _31798_);
  and (_36836_, _36825_, _36804_);
  or (_36847_, _36836_, _36760_);
  or (_36858_, _36847_, _36749_);
  and (_08957_, _36858_, _42545_);
  and (_36879_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36890_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_36901_, _36890_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_36912_, _36901_);
  not (_36922_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_36933_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_36944_, _36933_, _36922_);
  and (_36955_, _36890_, _18770_);
  and (_36966_, _36955_, _36944_);
  not (_36977_, _36966_);
  not (_36988_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_36999_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37010_, _36999_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_37021_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  not (_37032_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_37043_, _36999_, _37032_);
  and (_37054_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_37065_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37076_, _37065_, _37032_);
  and (_37087_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_37098_, _37087_, _37054_);
  or (_37109_, _37098_, _37021_);
  and (_37120_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_37131_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_37142_, _37131_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37153_, _37142_, _37032_);
  and (_37163_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_37174_, _37163_, _37120_);
  nor (_37185_, _36999_, _37032_);
  and (_37196_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_37207_, _37131_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37218_, _37207_, _37032_);
  and (_37229_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_37240_, _37229_, _37196_);
  nand (_37251_, _37240_, _37174_);
  nor (_37262_, _37251_, _37109_);
  and (_37272_, _37262_, _36988_);
  nor (_37283_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _36988_);
  or (_37294_, _37283_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37305_, _37294_, _37272_);
  and (_37316_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_37327_, _37316_, _37305_);
  nor (_37338_, _37327_, _36977_);
  not (_37349_, _37338_);
  not (_37360_, _36944_);
  nor (_37371_, _36955_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_37382_, _37371_, _37360_);
  and (_37392_, _37382_, _37349_);
  not (_37403_, _37392_);
  and (_37414_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_37425_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_37436_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_37447_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_37458_, _37447_, _37436_);
  and (_37469_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_37480_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_37491_, _37480_, _37469_);
  and (_37501_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_37512_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_37523_, _37512_, _37501_);
  and (_37534_, _37523_, _37491_);
  and (_37545_, _37534_, _37458_);
  nor (_37556_, _37545_, _37120_);
  and (_37567_, _37556_, _36988_);
  nor (_37578_, _37567_, _37425_);
  nor (_37589_, _37578_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37600_, _37589_, _37414_);
  and (_37611_, _37600_, _36966_);
  not (_37622_, _37611_);
  nor (_37633_, _36955_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_37644_, _37633_, _37360_);
  and (_37655_, _37644_, _37622_);
  and (_37666_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37675_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37686_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_37697_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_37708_, _37697_, _37686_);
  and (_37719_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_37730_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_37741_, _37730_, _37719_);
  and (_37746_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_37747_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_37748_, _37747_, _37746_);
  and (_37749_, _37748_, _37741_);
  and (_37750_, _37749_, _37708_);
  nor (_37751_, _37750_, _37120_);
  and (_37752_, _37751_, _36988_);
  nor (_37753_, _37752_, _37675_);
  nor (_37754_, _37753_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37755_, _37754_, _37666_);
  and (_37756_, _37755_, _36966_);
  not (_37757_, _37756_);
  nor (_37758_, _36955_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_37759_, _37758_, _37360_);
  and (_37760_, _37759_, _37757_);
  not (_37761_, _37760_);
  and (_37762_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37763_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_37764_, _37120_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37765_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_37766_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_37767_, _37766_, _37765_);
  and (_37768_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_37769_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_37770_, _37769_, _37768_);
  and (_37771_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_37772_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_37773_, _37772_, _37771_);
  and (_37774_, _37773_, _37770_);
  and (_37775_, _37774_, _37767_);
  nor (_37776_, _37775_, _37764_);
  nor (_37777_, _37776_, _37763_);
  nor (_37778_, _37777_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37779_, _37778_, _37762_);
  nor (_37780_, _37779_, _36977_);
  and (_37781_, _36977_, \oc8051_top_1.oc8051_decoder1.op [6]);
  or (_37782_, _37781_, _37780_);
  and (_37783_, _37782_, _36944_);
  nor (_37784_, _37783_, _37761_);
  and (_37785_, _37784_, _37655_);
  and (_37786_, _37785_, _37403_);
  and (_37787_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37788_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37789_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_37790_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_37791_, _37790_, _37789_);
  and (_37792_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_37793_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_37794_, _37793_, _37792_);
  and (_37795_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_37796_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_37797_, _37796_, _37795_);
  and (_37798_, _37797_, _37794_);
  and (_37799_, _37798_, _37791_);
  nor (_37800_, _37799_, _37120_);
  and (_37801_, _37800_, _36988_);
  nor (_37802_, _37801_, _37788_);
  nor (_37803_, _37802_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37804_, _37803_, _37787_);
  and (_37805_, _37804_, _36966_);
  not (_37806_, _37805_);
  nor (_37807_, _36955_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_37808_, _37807_, _37360_);
  and (_37809_, _37808_, _37806_);
  and (_37810_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_37811_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_37812_, _37811_, _37810_);
  and (_37813_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_37814_, _37813_, _37120_);
  and (_37815_, _37814_, _37812_);
  and (_37816_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not (_37817_, _37816_);
  and (_37818_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_37819_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_37820_, _37819_, _37818_);
  and (_37821_, _37820_, _37817_);
  and (_37822_, _37821_, _37815_);
  and (_37823_, _37822_, _36988_);
  nor (_37824_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _36988_);
  or (_37825_, _37824_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37826_, _37825_, _37823_);
  and (_37827_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_37828_, _37827_, _37826_);
  nor (_37829_, _37828_, _36977_);
  not (_37830_, _37829_);
  nor (_37831_, _36955_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_37832_, _37831_, _37360_);
  and (_37833_, _37832_, _37830_);
  and (_37834_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_37835_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37836_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37837_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_37838_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_37839_, _37838_, _37837_);
  and (_37840_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_37841_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_37842_, _37841_, _37840_);
  and (_37843_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_37844_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_37845_, _37844_, _37843_);
  and (_37846_, _37845_, _37842_);
  and (_37847_, _37846_, _37839_);
  nor (_37848_, _37847_, _37120_);
  and (_37849_, _37848_, _36988_);
  or (_37850_, _37849_, _37836_);
  and (_37851_, _37850_, _37835_);
  nor (_37852_, _37851_, _37834_);
  and (_37853_, _37852_, _36966_);
  not (_37854_, _37853_);
  nor (_37855_, _36955_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_37856_, _37855_, _37360_);
  and (_37857_, _37856_, _37854_);
  and (_37858_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37859_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37860_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_37861_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_37862_, _37861_, _37860_);
  and (_37863_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_37864_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_37865_, _37864_, _37863_);
  and (_37866_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_37867_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_37868_, _37867_, _37866_);
  and (_37869_, _37868_, _37865_);
  and (_37870_, _37869_, _37862_);
  nor (_37871_, _37870_, _37120_);
  and (_37872_, _37871_, _36988_);
  or (_37873_, _37872_, _37859_);
  and (_37874_, _37873_, _37835_);
  nor (_37875_, _37874_, _37858_);
  and (_37876_, _37875_, _36966_);
  not (_37877_, _37876_);
  nor (_37878_, _36955_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_37879_, _37878_, _37360_);
  and (_37880_, _37879_, _37877_);
  nor (_37881_, _37880_, _37857_);
  and (_37882_, _37881_, _37833_);
  and (_37883_, _37882_, _37809_);
  and (_37884_, _37883_, _37786_);
  not (_37885_, _37883_);
  nor (_37886_, _37783_, _37760_);
  and (_37887_, _37886_, _37655_);
  and (_37888_, _37887_, _37392_);
  not (_37889_, _37655_);
  and (_37890_, _37783_, _37760_);
  and (_37891_, _37890_, _37889_);
  and (_37892_, _37891_, _37392_);
  nor (_37893_, _37892_, _37888_);
  nor (_37894_, _37893_, _37885_);
  nor (_37895_, _37894_, _37884_);
  and (_37896_, _37887_, _37403_);
  not (_37897_, _37857_);
  and (_37898_, _37880_, _37897_);
  nor (_37899_, _37833_, _37809_);
  and (_37900_, _37899_, _37898_);
  and (_37901_, _37900_, _37896_);
  and (_37902_, _37900_, _37786_);
  nor (_37903_, _37902_, _37901_);
  and (_37904_, _37903_, _37895_);
  nor (_37905_, _37904_, _36912_);
  not (_37906_, _37905_);
  and (_37907_, _37783_, _37889_);
  and (_37908_, _37899_, _37881_);
  not (_37909_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_37910_, _18770_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_37911_, _37910_, _37909_);
  and (_37912_, _37911_, _37908_);
  and (_37913_, _37912_, _37907_);
  and (_37914_, _37902_, _18770_);
  and (_37915_, _37901_, _18770_);
  nor (_37916_, _37915_, _37914_);
  nor (_37917_, _37916_, _36890_);
  nor (_37918_, _37917_, _37913_);
  and (_37919_, _37918_, _37906_);
  nor (_37920_, _37919_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37921_, _37920_, _36879_);
  and (_37922_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_37923_, _37809_);
  and (_37924_, _37882_, _37923_);
  and (_37925_, _37888_, _37924_);
  not (_37926_, _37833_);
  and (_37927_, _37926_, _37809_);
  and (_37928_, _37927_, _37898_);
  and (_37929_, _37896_, _37928_);
  nor (_37930_, _37929_, _37925_);
  nor (_37931_, _37783_, _37655_);
  and (_37932_, _37931_, _37760_);
  and (_37933_, _37932_, _37924_);
  and (_37934_, _37880_, _37833_);
  and (_37935_, _37934_, _37897_);
  and (_37936_, _37935_, _37786_);
  nor (_37937_, _37936_, _37933_);
  and (_37938_, _37937_, _37930_);
  and (_37939_, _37891_, _37403_);
  and (_37940_, _37939_, _37928_);
  and (_37941_, _37783_, _37761_);
  and (_37942_, _37941_, _37655_);
  and (_37943_, _37942_, _37403_);
  and (_37944_, _37943_, _37928_);
  nor (_37945_, _37944_, _37940_);
  and (_37946_, _37896_, _37924_);
  and (_37947_, _37941_, _37889_);
  and (_37948_, _37947_, _37392_);
  and (_37949_, _37948_, _37882_);
  nor (_37950_, _37949_, _37946_);
  and (_37951_, _37950_, _37945_);
  and (_37952_, _37951_, _37938_);
  and (_37953_, _37932_, _37403_);
  and (_37954_, _37908_, _37953_);
  not (_37955_, _37954_);
  and (_37956_, _37932_, _37392_);
  and (_37957_, _37956_, _37908_);
  and (_37958_, _37931_, _37761_);
  and (_37959_, _37958_, _37392_);
  and (_37960_, _37959_, _37908_);
  nor (_37961_, _37960_, _37957_);
  and (_37962_, _37961_, _37955_);
  and (_37963_, _37786_, _37857_);
  not (_37964_, _37963_);
  and (_37965_, _37890_, _37655_);
  and (_37966_, _37965_, _37403_);
  and (_37967_, _37966_, _37928_);
  and (_37968_, _37958_, _37403_);
  and (_37969_, _37968_, _37928_);
  nor (_37970_, _37969_, _37967_);
  and (_37971_, _37970_, _37964_);
  and (_37972_, _37971_, _37962_);
  and (_37973_, _37972_, _37952_);
  and (_37974_, _37942_, _37392_);
  and (_37975_, _37974_, _37928_);
  and (_37976_, _37959_, _37928_);
  nor (_37977_, _37976_, _37975_);
  and (_37978_, _37908_, _37785_);
  and (_37979_, _37947_, _37403_);
  and (_37980_, _37979_, _37928_);
  nor (_37981_, _37980_, _37978_);
  and (_37982_, _37981_, _37977_);
  and (_37983_, _37785_, _37392_);
  and (_37984_, _37983_, _37924_);
  and (_37985_, _37943_, _37924_);
  nor (_37986_, _37985_, _37984_);
  and (_37987_, _37892_, _37924_);
  and (_37988_, _37979_, _37882_);
  nor (_37989_, _37988_, _37987_);
  and (_37990_, _37989_, _37986_);
  and (_37991_, _37990_, _37982_);
  and (_37992_, _37939_, _37882_);
  and (_37993_, _37908_, _37942_);
  nor (_37994_, _37993_, _37992_);
  not (_37995_, _37994_);
  not (_37996_, _37928_);
  nor (_37997_, _37983_, _37888_);
  nor (_37998_, _37997_, _37996_);
  nor (_37999_, _37998_, _37995_);
  nor (_38000_, _37948_, _37932_);
  nor (_38001_, _38000_, _37996_);
  and (_38002_, _37974_, _37924_);
  and (_38003_, _37786_, _37924_);
  nor (_38004_, _38003_, _38002_);
  not (_38005_, _38004_);
  nor (_38006_, _38005_, _38001_);
  and (_38007_, _38006_, _37999_);
  and (_38008_, _38007_, _37991_);
  and (_38009_, _38008_, _37973_);
  nor (_38010_, _38009_, _36912_);
  and (_38011_, \oc8051_top_1.oc8051_decoder1.state [0], _18770_);
  and (_38012_, _38011_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_38013_, _38012_, _37933_);
  nor (_38014_, _37913_, _38013_);
  not (_38015_, _38014_);
  nor (_38016_, _38015_, _38010_);
  nor (_38017_, _38016_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38018_, _38017_, _37922_);
  and (_38019_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38020_, _37403_, _37857_);
  and (_38021_, _38020_, _37934_);
  and (_38022_, _38021_, _37947_);
  and (_38023_, _37935_, _37932_);
  or (_38024_, _38023_, _38022_);
  and (_38025_, _38021_, _37785_);
  and (_38026_, _37958_, _37935_);
  nor (_38027_, _38026_, _38025_);
  not (_38028_, _38027_);
  nor (_38029_, _38028_, _38024_);
  and (_38030_, _37935_, _37403_);
  and (_38031_, _38030_, _37965_);
  and (_38032_, _38030_, _37941_);
  and (_38033_, _38032_, _37889_);
  nor (_38034_, _38033_, _38031_);
  and (_38035_, _37935_, _37896_);
  and (_38036_, _37939_, _37935_);
  nor (_38037_, _38036_, _38035_);
  and (_38038_, _38037_, _38034_);
  and (_38039_, _38038_, _38029_);
  and (_38040_, _37942_, _37935_);
  and (_38041_, _38021_, _37887_);
  nor (_38042_, _38041_, _38040_);
  and (_38043_, _37974_, _37908_);
  nor (_38044_, _38043_, _37933_);
  and (_38045_, _38044_, _38042_);
  and (_38046_, _38045_, _37895_);
  and (_38047_, _38046_, _38039_);
  nor (_38048_, _38047_, _36912_);
  and (_38049_, _37913_, _37760_);
  or (_38050_, _38049_, _38013_);
  nor (_38051_, _38050_, _38048_);
  nor (_38052_, _38051_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38053_, _38052_, _38019_);
  nor (_38054_, _38053_, _38018_);
  and (_38055_, _38054_, _37921_);
  and (_09507_, _38055_, _42545_);
  and (_38056_, _28417_, _27935_);
  not (_38057_, _27803_);
  nor (_38058_, _38057_, _28088_);
  and (_38059_, _38058_, _38056_);
  and (_38060_, _38059_, _33005_);
  and (_38061_, _31187_, _28242_);
  and (_38062_, _38061_, _27332_);
  and (_38063_, _38062_, _38060_);
  not (_38064_, _38063_);
  and (_38065_, _38064_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_38066_, _38060_, _27332_);
  and (_38067_, _38066_, _38061_);
  not (_38068_, _38067_);
  or (_38069_, _24184_, _18826_);
  and (_38070_, _29536_, _24162_);
  or (_38071_, _30966_, _30933_);
  or (_38072_, _38071_, _38070_);
  or (_38073_, _38072_, _38069_);
  nor (_38074_, _38073_, _32081_);
  nor (_38075_, _38074_, _20043_);
  not (_38076_, _38075_);
  and (_38077_, _38076_, _36510_);
  and (_38078_, _38077_, _36379_);
  nor (_38079_, _38078_, _38068_);
  nor (_38080_, _38079_, _38065_);
  and (_38081_, _38064_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38082_, _38074_, _21077_);
  not (_38083_, _38082_);
  and (_38084_, _38083_, _35781_);
  and (_38085_, _38084_, _35617_);
  nor (_38086_, _38085_, _38068_);
  nor (_38087_, _38086_, _38081_);
  and (_38088_, _38064_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38089_, _38074_, _21251_);
  not (_38090_, _38089_);
  and (_38091_, _38090_, _34965_);
  and (_38092_, _38091_, _34823_);
  nor (_38093_, _38092_, _38068_);
  nor (_38094_, _38093_, _38088_);
  and (_38095_, _38064_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38096_, _38074_, _21621_);
  not (_38097_, _38096_);
  and (_38098_, _38097_, _34202_);
  and (_38099_, _38098_, _33941_);
  and (_38100_, _38099_, _34083_);
  nor (_38101_, _38100_, _38068_);
  nor (_38102_, _38101_, _38095_);
  and (_38103_, _38064_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38104_, _38074_, _22144_);
  not (_38105_, _38104_);
  and (_38106_, _38105_, _33331_);
  and (_38107_, _38106_, _33364_);
  and (_38108_, _38107_, _33244_);
  nor (_38109_, _38108_, _38068_);
  nor (_38110_, _38109_, _38103_);
  and (_38111_, _38064_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38112_, _38074_, _21969_);
  nor (_38113_, _38112_, _32722_);
  and (_38114_, _38113_, _32624_);
  and (_38115_, _38114_, _32537_);
  nor (_38116_, _38115_, _38068_);
  nor (_38117_, _38116_, _38111_);
  nor (_38118_, _38063_, _27518_);
  nor (_38119_, _38074_, _22514_);
  not (_38120_, _38119_);
  and (_38121_, _38120_, _32070_);
  and (_38122_, _38121_, _32037_);
  and (_38123_, _38122_, _32004_);
  not (_38124_, _38123_);
  and (_38125_, _38124_, _38067_);
  nor (_38126_, _38125_, _38118_);
  and (_38127_, _38126_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38128_, _38127_, _38117_);
  and (_38129_, _38128_, _38110_);
  and (_38130_, _38129_, _38102_);
  and (_38131_, _38130_, _38094_);
  and (_38132_, _38131_, _38087_);
  and (_38133_, _38132_, _38080_);
  nor (_38134_, _38063_, _27957_);
  and (_38135_, _38134_, _38133_);
  nor (_38136_, _38134_, _38133_);
  nor (_38137_, _38136_, _38135_);
  and (_38138_, _38137_, _27661_);
  nor (_38139_, _38063_, _28001_);
  not (_38140_, _38139_);
  nor (_38141_, _38140_, _38138_);
  nor (_38142_, _38074_, _20881_);
  not (_38143_, _38142_);
  and (_38144_, _38143_, _30889_);
  and (_38145_, _38144_, _30835_);
  and (_38146_, _38145_, _30551_);
  and (_38147_, _38146_, _38067_);
  nor (_38148_, _38147_, _38141_);
  and (_09528_, _38148_, _42545_);
  not (_38149_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38150_, _38126_, _38149_);
  nor (_38151_, _38126_, _38149_);
  nor (_38152_, _38151_, _38150_);
  and (_38153_, _38152_, _27661_);
  nor (_38154_, _38153_, _27529_);
  nor (_38155_, _38154_, _38067_);
  nor (_38156_, _38155_, _38125_);
  nand (_10658_, _38156_, _42545_);
  nor (_38157_, _38127_, _38117_);
  nor (_38158_, _38157_, _38128_);
  nor (_38159_, _38158_, _27079_);
  nor (_38160_, _38159_, _27364_);
  nor (_38161_, _38160_, _38067_);
  nor (_38162_, _38161_, _38116_);
  nand (_10669_, _38162_, _42545_);
  nor (_38163_, _38128_, _38110_);
  nor (_38164_, _38163_, _38129_);
  nor (_38165_, _38164_, _27079_);
  nor (_38166_, _38165_, _27134_);
  nor (_38167_, _38166_, _38067_);
  nor (_38168_, _38167_, _38109_);
  nand (_10680_, _38168_, _42545_);
  nor (_38169_, _38129_, _38102_);
  nor (_38170_, _38169_, _38130_);
  nor (_38171_, _38170_, _27079_);
  nor (_38172_, _38171_, _28143_);
  nor (_38173_, _38172_, _38067_);
  nor (_38174_, _38173_, _38101_);
  nor (_10691_, _38174_, rst);
  nor (_38175_, _38130_, _38094_);
  nor (_38176_, _38175_, _38131_);
  nor (_38177_, _38176_, _27079_);
  nor (_38178_, _38177_, _28351_);
  nor (_38179_, _38178_, _38067_);
  nor (_38180_, _38179_, _38093_);
  nor (_10702_, _38180_, rst);
  nor (_38181_, _38131_, _38087_);
  nor (_38182_, _38181_, _38132_);
  nor (_38183_, _38182_, _27079_);
  nor (_38184_, _38183_, _27847_);
  nor (_38185_, _38184_, _38067_);
  nor (_38186_, _38185_, _38086_);
  nor (_10713_, _38186_, rst);
  nor (_38187_, _38132_, _38080_);
  nor (_38188_, _38187_, _38133_);
  nor (_38189_, _38188_, _27079_);
  nor (_38190_, _38189_, _27694_);
  nor (_38191_, _38190_, _38067_);
  nor (_38192_, _38191_, _38079_);
  nor (_10724_, _38192_, rst);
  and (_38193_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18770_);
  and (_38194_, _38193_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38195_, _38059_, _34431_);
  nand (_38196_, _38195_, _38061_);
  or (_38197_, _38196_, _31111_);
  not (_38198_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand (_38199_, _38196_, _38198_);
  and (_38200_, _38199_, _38197_);
  or (_38201_, _38200_, _38194_);
  not (_38202_, _38194_);
  nor (_38203_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38204_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38205_, _38204_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38206_, _38205_, _38203_);
  nor (_38207_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38208_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38209_, _38208_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38210_, _38209_, _38207_);
  not (_38211_, _38210_);
  nor (_38212_, _38211_, _31253_);
  nor (_38213_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38214_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38215_, _38214_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38216_, _38215_, _38213_);
  and (_38217_, _38216_, _38212_);
  nor (_38218_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38219_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38220_, _38219_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38221_, _38220_, _38218_);
  and (_38222_, _38221_, _38217_);
  and (_38223_, _38222_, _38206_);
  nor (_38224_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38225_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38226_, _38225_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38227_, _38226_, _38224_);
  and (_38228_, _38227_, _38223_);
  nor (_38229_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38230_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38231_, _38230_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38232_, _38231_, _38229_);
  and (_38233_, _38232_, _38228_);
  nor (_38234_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38235_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38236_, _38235_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38237_, _38236_, _38234_);
  and (_38238_, _38237_, _38233_);
  nor (_38239_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38240_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38241_, _38240_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38242_, _38241_, _38239_);
  or (_38243_, _38242_, _38238_);
  nand (_38244_, _38242_, _38238_);
  and (_38245_, _38244_, _29547_);
  and (_38246_, _38245_, _38243_);
  and (_38247_, _23877_, _18826_);
  and (_38248_, _29218_, _20370_);
  not (_38249_, _38248_);
  and (_38250_, _30301_, _20892_);
  and (_38251_, _38250_, _29810_);
  and (_38252_, _38251_, _29843_);
  and (_38253_, _38252_, _29886_);
  and (_38254_, _38253_, _30072_);
  nor (_38255_, _38254_, _30332_);
  and (_38256_, _29218_, _19384_);
  nor (_38257_, _38256_, _38255_);
  and (_38258_, _38257_, _38249_);
  and (_38259_, _30388_, _20881_);
  and (_38260_, _20217_, _19220_);
  and (_38261_, _20533_, _19547_);
  and (_38262_, _38261_, _38260_);
  and (_38263_, _38262_, _38259_);
  and (_38264_, _20370_, _19384_);
  and (_38265_, _38264_, _38263_);
  nor (_38266_, _38265_, _29218_);
  not (_38267_, _38266_);
  and (_38268_, _38267_, _38258_);
  nor (_38269_, _29218_, _19721_);
  and (_38270_, _29218_, _19721_);
  nor (_38271_, _38270_, _38269_);
  and (_38272_, _38271_, _38268_);
  nand (_38273_, _38272_, _30464_);
  or (_38274_, _38272_, _30464_);
  and (_38275_, _38274_, _38273_);
  and (_38276_, _38275_, _30235_);
  and (_38277_, _29218_, _30464_);
  or (_38278_, _38277_, _31362_);
  and (_38279_, _38278_, _30508_);
  nor (_38280_, _31493_, _21621_);
  nor (_38281_, _30944_, _20717_);
  and (_38282_, _24184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  or (_38283_, _38282_, _38281_);
  or (_38284_, _38283_, _38280_);
  or (_38285_, _38284_, _38279_);
  or (_38286_, _38285_, _38276_);
  or (_38287_, _38286_, _38247_);
  or (_38288_, _38287_, _38246_);
  or (_38289_, _38288_, _38202_);
  and (_38290_, _38289_, _42545_);
  and (_12675_, _38290_, _38201_);
  and (_38291_, _38059_, _33713_);
  and (_38292_, _38291_, _38061_);
  nor (_38293_, _38292_, _38194_);
  or (_38294_, _38293_, _31111_);
  not (_38295_, _38293_);
  or (_38296_, _38295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38297_, _38296_, _42545_);
  and (_12696_, _38297_, _38294_);
  nor (_38298_, _38196_, _32265_);
  and (_38299_, _38196_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38300_, _38299_, _38194_);
  or (_38301_, _38300_, _38298_);
  and (_38302_, _26478_, _24184_);
  not (_38303_, _38302_);
  and (_38304_, _38211_, _31253_);
  nor (_38305_, _38304_, _38212_);
  and (_38306_, _38305_, _29547_);
  nor (_38307_, _31362_, _30497_);
  not (_38308_, _38307_);
  nor (_38309_, _38308_, _30410_);
  nor (_38310_, _38309_, _29810_);
  and (_38311_, _38309_, _29810_);
  nor (_38312_, _38311_, _38310_);
  and (_38313_, _38312_, _30235_);
  nor (_38314_, _30944_, _19547_);
  and (_38315_, _23655_, _18826_);
  nor (_38316_, _31493_, _21251_);
  nor (_38317_, _30519_, _22514_);
  or (_38318_, _38317_, _38316_);
  or (_38319_, _38318_, _38315_);
  nor (_38320_, _38319_, _38314_);
  not (_38321_, _38320_);
  nor (_38322_, _38321_, _38313_);
  not (_38323_, _38322_);
  nor (_38324_, _38323_, _38306_);
  and (_38325_, _38324_, _38303_);
  nand (_38326_, _38325_, _38194_);
  and (_38327_, _38326_, _42545_);
  and (_13611_, _38327_, _38301_);
  nor (_38328_, _38196_, _32907_);
  and (_38329_, _38196_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38330_, _38329_, _38194_);
  or (_38331_, _38330_, _38328_);
  nor (_38332_, _38216_, _38212_);
  nor (_38333_, _38332_, _38217_);
  and (_38334_, _38333_, _29547_);
  not (_38335_, _38334_);
  and (_38336_, _25470_, _24184_);
  nor (_38337_, _38251_, _30332_);
  and (_38338_, _38259_, _19547_);
  nor (_38339_, _38338_, _29218_);
  or (_38340_, _38339_, _38337_);
  nor (_38341_, _38340_, _29843_);
  and (_38342_, _38340_, _29843_);
  or (_38343_, _38342_, _38341_);
  and (_38344_, _38343_, _30235_);
  nor (_38345_, _30944_, _20533_);
  and (_38346_, _23687_, _18826_);
  nor (_38347_, _31493_, _21077_);
  nor (_38348_, _30519_, _21969_);
  or (_38349_, _38348_, _38347_);
  or (_38350_, _38349_, _38346_);
  nor (_38351_, _38350_, _38345_);
  not (_38352_, _38351_);
  nor (_38353_, _38352_, _38344_);
  not (_38354_, _38353_);
  nor (_38355_, _38354_, _38336_);
  and (_38356_, _38355_, _38335_);
  nand (_38357_, _38356_, _38194_);
  and (_38358_, _38357_, _42545_);
  and (_13622_, _38358_, _38331_);
  nor (_38359_, _38196_, _33582_);
  and (_38360_, _38196_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38361_, _38360_, _38194_);
  or (_38362_, _38361_, _38359_);
  nor (_38363_, _38221_, _38217_);
  nor (_38364_, _38363_, _38222_);
  and (_38365_, _38364_, _29547_);
  not (_38366_, _38365_);
  and (_38367_, _38338_, _20533_);
  and (_38368_, _38367_, _30332_);
  and (_38369_, _38252_, _29218_);
  nor (_38370_, _38369_, _38368_);
  and (_38371_, _38370_, _19220_);
  nor (_38372_, _38370_, _19220_);
  nor (_38373_, _38372_, _38371_);
  and (_38374_, _38373_, _30235_);
  not (_38375_, _38374_);
  nor (_38376_, _30519_, _22144_);
  and (_38377_, _24184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38378_, _38377_, _38376_);
  and (_38379_, _23718_, _18826_);
  nor (_38380_, _31493_, _20043_);
  nor (_38381_, _30944_, _19220_);
  or (_38382_, _38381_, _38380_);
  nor (_38383_, _38382_, _38379_);
  and (_38384_, _38383_, _38378_);
  and (_38385_, _38384_, _38375_);
  and (_38386_, _38385_, _38366_);
  nand (_38387_, _38386_, _38194_);
  and (_38390_, _38387_, _42545_);
  and (_13633_, _38390_, _38362_);
  nor (_38392_, _38196_, _34333_);
  and (_38393_, _38196_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38394_, _38393_, _38194_);
  or (_38395_, _38394_, _38392_);
  nor (_38396_, _38222_, _38206_);
  nor (_38397_, _38396_, _38223_);
  and (_38398_, _38397_, _29547_);
  not (_38399_, _38398_);
  nor (_38400_, _38253_, _30072_);
  not (_38402_, _38400_);
  and (_38411_, _38402_, _38255_);
  and (_38417_, _38367_, _19220_);
  nor (_38423_, _38417_, _20217_);
  nor (_38426_, _38423_, _38263_);
  nor (_38427_, _38426_, _29218_);
  nor (_38428_, _38427_, _38411_);
  nor (_38429_, _38428_, _33200_);
  nor (_38430_, _30944_, _20217_);
  or (_38431_, _38430_, _31514_);
  nor (_38432_, _38431_, _38429_);
  and (_38433_, _23750_, _18826_);
  nor (_38434_, _30519_, _21621_);
  and (_38435_, _24184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_38436_, _38435_, _38434_);
  nor (_38437_, _38436_, _38433_);
  and (_38438_, _38437_, _38432_);
  and (_38439_, _38438_, _38399_);
  nand (_38440_, _38439_, _38194_);
  and (_38441_, _38440_, _42545_);
  and (_13644_, _38441_, _38395_);
  nor (_38442_, _38196_, _35128_);
  and (_38443_, _38196_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38444_, _38443_, _38194_);
  or (_38445_, _38444_, _38442_);
  nor (_38446_, _38227_, _38223_);
  nor (_38447_, _38446_, _38228_);
  and (_38448_, _38447_, _29547_);
  not (_38449_, _38448_);
  and (_38452_, _23782_, _18826_);
  nor (_38453_, _38263_, _29218_);
  nor (_38454_, _38453_, _38255_);
  nor (_38455_, _38454_, _29667_);
  and (_38456_, _38454_, _29667_);
  nor (_38457_, _38456_, _38455_);
  and (_38458_, _38457_, _30235_);
  and (_38459_, _24184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38460_, _29218_, _21262_);
  or (_38461_, _38460_, _30519_);
  nor (_38462_, _38461_, _38256_);
  nor (_38463_, _31493_, _22514_);
  nor (_38464_, _30944_, _19384_);
  or (_38465_, _38464_, _38463_);
  or (_38466_, _38465_, _38462_);
  nor (_38467_, _38466_, _38459_);
  not (_38468_, _38467_);
  nor (_38469_, _38468_, _38458_);
  not (_38470_, _38469_);
  nor (_38471_, _38470_, _38452_);
  and (_38472_, _38471_, _38449_);
  nand (_38473_, _38472_, _38194_);
  and (_38474_, _38473_, _42545_);
  and (_13655_, _38474_, _38445_);
  nor (_38475_, _38196_, _35956_);
  and (_38476_, _38196_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38477_, _38476_, _38194_);
  or (_38478_, _38477_, _38475_);
  nor (_38479_, _38232_, _38228_);
  nor (_38480_, _38479_, _38233_);
  and (_38481_, _38480_, _29547_);
  not (_38482_, _38481_);
  and (_38483_, _23813_, _18826_);
  and (_38484_, _38263_, _19384_);
  nor (_38485_, _38484_, _29218_);
  not (_38486_, _38485_);
  and (_38487_, _38486_, _38257_);
  and (_38488_, _38487_, _20370_);
  nor (_38490_, _38487_, _20370_);
  nor (_38494_, _38490_, _38488_);
  nor (_38500_, _38494_, _33200_);
  and (_38505_, _24184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_38512_, _36292_, _30519_);
  and (_38520_, _38512_, _38249_);
  nor (_38528_, _31493_, _21969_);
  nor (_38529_, _30944_, _20370_);
  or (_38530_, _38529_, _38528_);
  or (_38531_, _38530_, _38520_);
  nor (_38532_, _38531_, _38505_);
  not (_38533_, _38532_);
  nor (_38534_, _38533_, _38500_);
  not (_38535_, _38534_);
  nor (_38536_, _38535_, _38483_);
  and (_38537_, _38536_, _38482_);
  nand (_38538_, _38537_, _38194_);
  and (_38539_, _38538_, _42545_);
  and (_13665_, _38539_, _38478_);
  nor (_38540_, _38196_, _36684_);
  and (_38541_, _38196_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38542_, _38541_, _38194_);
  or (_38543_, _38542_, _38540_);
  nor (_38544_, _38237_, _38233_);
  nor (_38545_, _38544_, _38238_);
  and (_38546_, _38545_, _29547_);
  and (_38547_, _23845_, _18826_);
  and (_38548_, _38268_, _19721_);
  nor (_38549_, _38268_, _19721_);
  or (_38550_, _38549_, _38548_);
  and (_38551_, _38550_, _30235_);
  or (_38552_, _29218_, _20054_);
  nor (_38553_, _38270_, _30519_);
  and (_38554_, _38553_, _38552_);
  nor (_38555_, _31493_, _22144_);
  nor (_38556_, _30944_, _19721_);
  and (_38557_, _24184_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or (_38558_, _38557_, _38556_);
  or (_38559_, _38558_, _38555_);
  or (_38560_, _38559_, _38554_);
  or (_38561_, _38560_, _38551_);
  or (_38562_, _38561_, _38547_);
  or (_38563_, _38562_, _38546_);
  or (_38564_, _38563_, _38202_);
  and (_38570_, _38564_, _42545_);
  and (_13676_, _38570_, _38543_);
  nand (_38581_, _38295_, _32265_);
  or (_38582_, _38295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_38583_, _38582_, _42545_);
  and (_13687_, _38583_, _38581_);
  nand (_38599_, _38295_, _32907_);
  or (_38600_, _38295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38601_, _38600_, _42545_);
  and (_13698_, _38601_, _38599_);
  nand (_38602_, _38295_, _33582_);
  or (_38603_, _38295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38604_, _38603_, _42545_);
  and (_13709_, _38604_, _38602_);
  nand (_38605_, _38295_, _34333_);
  or (_38606_, _38295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38607_, _38606_, _42545_);
  and (_13720_, _38607_, _38605_);
  nand (_38608_, _38295_, _35128_);
  or (_38609_, _38295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38610_, _38609_, _42545_);
  and (_13731_, _38610_, _38608_);
  nand (_38611_, _38295_, _35956_);
  or (_38612_, _38295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38613_, _38612_, _42545_);
  and (_13742_, _38613_, _38611_);
  nand (_38614_, _38295_, _36684_);
  or (_38615_, _38295_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38616_, _38615_, _42545_);
  and (_13753_, _38616_, _38614_);
  not (_38617_, _27935_);
  nor (_38618_, _38617_, _27803_);
  and (_38619_, _38618_, _31798_);
  and (_38620_, _38619_, _28439_);
  and (_38621_, _31755_, _32352_);
  not (_38622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38623_, _31755_, _38622_);
  or (_38624_, _38623_, _38621_);
  and (_38625_, _38624_, _38620_);
  nor (_38626_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_38627_, _38626_);
  nand (_38628_, _38627_, _31732_);
  and (_38629_, _38626_, _38622_);
  nor (_38630_, _38629_, _38620_);
  and (_38631_, _38630_, _38628_);
  nor (_38632_, _28417_, _38617_);
  nor (_38633_, _27803_, _28088_);
  and (_38634_, _38061_, _27595_);
  and (_38635_, _38634_, _38633_);
  and (_38636_, _38635_, _38632_);
  or (_38637_, _38636_, _38631_);
  or (_38638_, _38637_, _38625_);
  nand (_38639_, _38636_, _38146_);
  and (_38640_, _38639_, _42545_);
  and (_15156_, _38640_, _38638_);
  and (_38641_, _38632_, _38633_);
  and (_38642_, _38641_, _38634_);
  and (_38643_, _38620_, _33016_);
  nand (_38644_, _38643_, _31732_);
  or (_38645_, _38643_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_38646_, _38645_, _38644_);
  or (_38647_, _38646_, _38642_);
  nand (_38648_, _38636_, _38115_);
  and (_38649_, _38648_, _42545_);
  and (_17337_, _38649_, _38647_);
  or (_38650_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_38651_, _23940_, _23908_);
  or (_38652_, _38651_, _23971_);
  or (_38653_, _38652_, _24014_);
  or (_38654_, _38653_, _24046_);
  or (_38655_, _38654_, _24088_);
  or (_38656_, _38655_, _24120_);
  or (_38657_, _38656_, _23591_);
  and (_38658_, _38657_, _18826_);
  or (_38659_, _31297_, _30170_);
  not (_38660_, _31296_);
  nand (_38661_, _38660_, _30170_);
  and (_38662_, _38661_, _29612_);
  and (_38663_, _38662_, _38659_);
  not (_38664_, _29470_);
  nand (_38665_, _29459_, _38664_);
  or (_38666_, _29481_, _29459_);
  and (_38667_, _29547_, _38666_);
  and (_38668_, _38667_, _38665_);
  and (_38669_, _38264_, _25371_);
  and (_38670_, _38262_, _24184_);
  nand (_38671_, _38670_, _38669_);
  nand (_38672_, _38671_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_38673_, _38672_, _38668_);
  or (_38674_, _38673_, _38663_);
  or (_38675_, _38674_, _38658_);
  and (_38676_, _38675_, _38650_);
  or (_38677_, _38676_, _38620_);
  not (_38678_, _38620_);
  and (_38679_, _33724_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_38680_, _38679_, _33735_);
  or (_38681_, _38680_, _38678_);
  and (_38682_, _38681_, _38677_);
  or (_38683_, _38682_, _38636_);
  nand (_38684_, _38636_, _38108_);
  and (_38685_, _38684_, _42545_);
  and (_17348_, _38685_, _38683_);
  and (_38686_, _38620_, _34431_);
  nand (_38687_, _38686_, _31732_);
  not (_38688_, _38636_);
  or (_38689_, _38686_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_38690_, _38689_, _38688_);
  and (_38691_, _38690_, _38687_);
  nor (_38692_, _38688_, _38100_);
  or (_38693_, _38692_, _38691_);
  and (_17359_, _38693_, _42545_);
  or (_38694_, _38678_, _35248_);
  not (_38695_, _38642_);
  and (_38696_, _38695_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_38697_, _38695_, _38092_);
  nor (_38698_, _38697_, _38696_);
  nor (_38491_, _38698_, rst);
  and (_38699_, _38491_, _38694_);
  and (_38700_, _35237_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_38701_, _38700_, _35281_);
  nor (_38702_, _38636_, rst);
  and (_38703_, _38702_, _38620_);
  and (_38704_, _38703_, _38701_);
  or (_17370_, _38704_, _38699_);
  and (_38705_, _38620_, _36043_);
  nand (_38706_, _38705_, _31732_);
  or (_38707_, _38705_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_38708_, _38707_, _38706_);
  or (_38709_, _38708_, _38642_);
  nand (_38710_, _38636_, _38085_);
  and (_38711_, _38710_, _42545_);
  and (_17381_, _38711_, _38709_);
  and (_38712_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_38713_, _29547_, _29360_);
  and (_38714_, _30126_, _29612_);
  or (_38715_, _38714_, _38713_);
  and (_38716_, _38715_, _38712_);
  nand (_38717_, _38712_, _30944_);
  and (_38718_, _38717_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_38719_, _38718_, _38620_);
  or (_38720_, _38719_, _38716_);
  not (_38721_, _36782_);
  nor (_38722_, _38721_, _31732_);
  or (_38723_, _36782_, _34126_);
  nand (_38724_, _38723_, _38620_);
  or (_38725_, _38724_, _38722_);
  and (_38726_, _38725_, _38720_);
  or (_38727_, _38726_, _38636_);
  nand (_38728_, _38636_, _38078_);
  and (_38729_, _38728_, _42545_);
  and (_17392_, _38729_, _38727_);
  not (_38730_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38731_, _38193_, _38730_);
  not (_38732_, _38731_);
  or (_38733_, _38732_, _38288_);
  nor (_38734_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38735_, _38734_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38736_, _27332_, _28242_);
  and (_38737_, _38736_, _27584_);
  and (_38738_, _28417_, _38617_);
  and (_38739_, _38738_, _38633_);
  and (_38740_, _38739_, _38737_);
  and (_38741_, _38740_, _31187_);
  nor (_38742_, _38741_, _38735_);
  not (_38743_, _38742_);
  and (_38744_, _38743_, _31111_);
  and (_38745_, _28417_, _28242_);
  and (_38746_, _38745_, _27946_);
  not (_38747_, _31798_);
  nor (_38748_, _38747_, _28088_);
  and (_38749_, _38748_, _38746_);
  and (_38750_, _38749_, _31755_);
  or (_38751_, _38750_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_38752_, _38742_, _38732_);
  nand (_38753_, _38750_, _31732_);
  and (_38754_, _38753_, _38752_);
  and (_38755_, _38754_, _38751_);
  or (_38756_, _38755_, _38731_);
  or (_38757_, _38756_, _38744_);
  and (_38758_, _38757_, _38733_);
  and (_17961_, _38758_, _42545_);
  nor (_38759_, _38732_, _38325_);
  and (_38760_, _38743_, _32265_);
  not (_38761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38762_, _38749_, _38761_);
  nor (_38763_, _38762_, _38743_);
  and (_38764_, _38745_, _28099_);
  and (_38765_, _31798_, _27946_);
  and (_38766_, _38765_, _38764_);
  and (_38767_, _32352_, _27595_);
  nor (_38768_, _27595_, _38761_);
  nor (_38769_, _38768_, _38767_);
  not (_38770_, _38769_);
  nand (_38771_, _38770_, _38766_);
  and (_38780_, _38771_, _38763_);
  nor (_38791_, _38780_, _38731_);
  not (_38802_, _38791_);
  nor (_38811_, _38802_, _38760_);
  nor (_38817_, _38811_, _38759_);
  nor (_19754_, _38817_, rst);
  nor (_38838_, _38732_, _38356_);
  and (_38849_, _38743_, _32907_);
  not (_38860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_38871_, _38749_, _38860_);
  nor (_38882_, _38871_, _38743_);
  not (_38893_, _33016_);
  nor (_38904_, _38893_, _31732_);
  nor (_38915_, _33016_, _38860_);
  nor (_38926_, _38915_, _38904_);
  not (_38937_, _38926_);
  and (_38948_, _38752_, _38766_);
  nand (_38959_, _38948_, _38937_);
  and (_38970_, _38959_, _38882_);
  nor (_38981_, _38970_, _38731_);
  not (_38985_, _38981_);
  nor (_38986_, _38985_, _38849_);
  nor (_38987_, _38986_, _38838_);
  nor (_19766_, _38987_, rst);
  nor (_38988_, _38732_, _38386_);
  and (_38989_, _38743_, _33582_);
  not (_38990_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_38991_, _38749_, _38990_);
  nor (_38992_, _38991_, _38743_);
  not (_38993_, _38766_);
  nor (_38994_, _33713_, _38990_);
  nor (_38995_, _38994_, _33735_);
  or (_38996_, _38995_, _38993_);
  and (_38997_, _38996_, _38992_);
  nor (_38998_, _38997_, _38731_);
  not (_38999_, _38998_);
  nor (_39000_, _38999_, _38989_);
  nor (_39001_, _39000_, _38988_);
  nor (_19778_, _39001_, rst);
  nor (_39002_, _38742_, _34333_);
  not (_39003_, _38749_);
  and (_39004_, _38752_, _39003_);
  and (_39005_, _39004_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  not (_39006_, _38948_);
  and (_39007_, _34442_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39008_, _39007_, _34453_);
  nor (_39009_, _39008_, _39006_);
  nor (_39010_, _39009_, _39005_);
  and (_39011_, _39010_, _38732_);
  not (_39012_, _39011_);
  nor (_39013_, _39012_, _39002_);
  and (_39014_, _38731_, _38439_);
  or (_39015_, _39014_, _39013_);
  nor (_19789_, _39015_, rst);
  nor (_39016_, _38742_, _35128_);
  and (_39017_, _38749_, _35226_);
  and (_39018_, _39017_, _31732_);
  nor (_39019_, _39017_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_39020_, _39019_);
  and (_39021_, _39020_, _38752_);
  not (_39022_, _39021_);
  nor (_39023_, _39022_, _39018_);
  or (_39024_, _39023_, _39016_);
  and (_39025_, _39024_, _38732_);
  nor (_39026_, _38732_, _38472_);
  or (_39027_, _39026_, _39025_);
  and (_19801_, _39027_, _42545_);
  nor (_39028_, _38742_, _35956_);
  and (_39029_, _38749_, _36043_);
  and (_39030_, _39029_, _31732_);
  nor (_39031_, _39029_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_39032_, _39031_);
  and (_39033_, _39032_, _38752_);
  not (_39034_, _39033_);
  nor (_39035_, _39034_, _39030_);
  or (_39036_, _39035_, _39028_);
  and (_39037_, _39036_, _38732_);
  nor (_39038_, _38732_, _38537_);
  or (_39039_, _39038_, _39037_);
  and (_19813_, _39039_, _42545_);
  nor (_39040_, _38732_, _38563_);
  nor (_39041_, _38742_, _36684_);
  and (_39042_, _38749_, _36782_);
  nor (_39043_, _39042_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not (_39044_, _39043_);
  not (_39045_, _38752_);
  and (_39046_, _39042_, _31732_);
  nor (_39047_, _39046_, _39045_);
  and (_39048_, _39047_, _39044_);
  nor (_39049_, _39048_, _38731_);
  not (_39050_, _39049_);
  nor (_39051_, _39050_, _39041_);
  nor (_39052_, _39051_, _39040_);
  and (_19825_, _39052_, _42545_);
  and (_39053_, _27935_, _27803_);
  and (_39054_, _38764_, _39053_);
  and (_39055_, _39054_, _31755_);
  nand (_39056_, _39055_, _31732_);
  or (_39057_, _39055_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39058_, _39057_, _31798_);
  and (_39059_, _39058_, _39056_);
  and (_39060_, _38059_, _38737_);
  nand (_39061_, _39060_, _38146_);
  or (_39062_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39063_, _39062_, _31187_);
  and (_39064_, _39063_, _39061_);
  not (_39065_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_39066_, _31166_, _39065_);
  or (_39067_, _39066_, rst);
  or (_39068_, _39067_, _39064_);
  or (_31031_, _39068_, _39059_);
  and (_39069_, _39053_, _28439_);
  and (_39070_, _39069_, _31755_);
  nand (_39071_, _39070_, _31732_);
  or (_39072_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39073_, _39072_, _31798_);
  and (_39074_, _39073_, _39071_);
  and (_39075_, _38632_, _38058_);
  and (_39076_, _39075_, _38737_);
  nand (_39077_, _39076_, _38146_);
  or (_39078_, _39076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39079_, _39078_, _31187_);
  and (_39080_, _39079_, _39077_);
  not (_39081_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_39082_, _31166_, _39081_);
  or (_39083_, _39082_, rst);
  or (_39084_, _39083_, _39080_);
  or (_31054_, _39084_, _39074_);
  and (_39085_, _38617_, _27803_);
  and (_39086_, _39085_, _38764_);
  and (_39087_, _39086_, _31755_);
  nand (_39088_, _39087_, _31732_);
  or (_39089_, _39087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39090_, _39089_, _31798_);
  and (_39091_, _39090_, _39088_);
  and (_39092_, _38738_, _38058_);
  and (_39093_, _39092_, _38737_);
  not (_39094_, _39093_);
  nor (_39095_, _39094_, _38146_);
  not (_39096_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_39097_, _39093_, _39096_);
  or (_39098_, _39097_, _39095_);
  and (_39099_, _39098_, _31187_);
  nor (_39100_, _31166_, _39096_);
  or (_39101_, _39100_, rst);
  or (_39102_, _39101_, _39099_);
  or (_31077_, _39102_, _39091_);
  and (_39103_, _39085_, _28439_);
  nand (_39104_, _39103_, _31755_);
  or (_39105_, _39104_, _32352_);
  not (_39106_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nand (_39107_, _39104_, _39106_);
  and (_39108_, _39107_, _31798_);
  and (_39109_, _39108_, _39105_);
  nor (_39110_, _28417_, _27935_);
  and (_39111_, _38058_, _39110_);
  and (_39112_, _39111_, _38737_);
  not (_39113_, _39112_);
  nor (_39114_, _39113_, _38146_);
  nor (_39115_, _39112_, _39106_);
  or (_39116_, _39115_, _39114_);
  and (_39117_, _39116_, _31187_);
  nor (_39118_, _31166_, _39106_);
  or (_39119_, _39118_, rst);
  or (_39120_, _39119_, _39117_);
  or (_31099_, _39120_, _39109_);
  or (_39121_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_39122_, _39121_, _31798_);
  and (_39123_, _39054_, _27595_);
  nand (_39124_, _39123_, _31732_);
  and (_39125_, _39124_, _39122_);
  nand (_39126_, _39060_, _38123_);
  and (_39127_, _39126_, _31187_);
  and (_39128_, _39127_, _39121_);
  not (_39129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39130_, _31166_, _39129_);
  or (_39131_, _39130_, rst);
  or (_39132_, _39131_, _39128_);
  or (_40232_, _39132_, _39125_);
  and (_39133_, _33005_, _38736_);
  and (_39134_, _39133_, _38059_);
  nand (_39135_, _39134_, _31732_);
  or (_39136_, _39134_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39137_, _39136_, _31798_);
  and (_39138_, _39137_, _39135_);
  nand (_39139_, _39060_, _38115_);
  or (_39140_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39141_, _39140_, _31187_);
  and (_39142_, _39141_, _39139_);
  not (_39143_, _31166_);
  and (_39144_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_39145_, _39144_, rst);
  or (_39146_, _39145_, _39142_);
  or (_40234_, _39146_, _39138_);
  not (_39147_, _34464_);
  nand (_39148_, _39054_, _39147_);
  and (_39149_, _39148_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39150_, _33746_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39151_, _39150_, _33735_);
  and (_39152_, _39151_, _39054_);
  or (_39153_, _39152_, _39149_);
  and (_39154_, _39153_, _31798_);
  nand (_39155_, _39060_, _38108_);
  or (_39156_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39157_, _39156_, _31187_);
  and (_39158_, _39157_, _39155_);
  and (_39159_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39160_, _39159_, rst);
  or (_39161_, _39160_, _39158_);
  or (_40236_, _39161_, _39154_);
  nand (_39162_, _39054_, _27332_);
  and (_39163_, _39162_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39164_, _39147_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39165_, _39164_, _34453_);
  and (_39166_, _39165_, _39054_);
  or (_39167_, _39166_, _39163_);
  and (_39168_, _39167_, _31798_);
  nand (_39169_, _39060_, _38100_);
  or (_39170_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39171_, _39170_, _31187_);
  and (_39172_, _39171_, _39169_);
  and (_39173_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39174_, _39173_, rst);
  or (_39175_, _39174_, _39172_);
  or (_40238_, _39175_, _39168_);
  not (_39176_, _39054_);
  or (_39177_, _39176_, _35248_);
  and (_39178_, _39177_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39179_, _35237_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39180_, _39179_, _35281_);
  and (_39181_, _39180_, _39054_);
  or (_39182_, _39181_, _39178_);
  and (_39183_, _39182_, _31798_);
  nand (_39184_, _39060_, _38092_);
  or (_39185_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39186_, _39185_, _31187_);
  and (_39187_, _39186_, _39184_);
  and (_39188_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39189_, _39188_, rst);
  or (_39190_, _39189_, _39187_);
  or (_40240_, _39190_, _39183_);
  and (_39191_, _39054_, _36043_);
  nand (_39192_, _39191_, _31732_);
  or (_39193_, _39191_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39194_, _39193_, _31798_);
  and (_39195_, _39194_, _39192_);
  nand (_39196_, _39060_, _38085_);
  or (_39197_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39198_, _39197_, _31187_);
  and (_39199_, _39198_, _39196_);
  and (_39200_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39201_, _39200_, rst);
  or (_39202_, _39201_, _39199_);
  or (_40242_, _39202_, _39195_);
  and (_39203_, _39054_, _36782_);
  nand (_39208_, _39203_, _31732_);
  or (_39214_, _39203_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39215_, _39214_, _31798_);
  and (_39216_, _39215_, _39208_);
  nand (_39217_, _39060_, _38078_);
  or (_39218_, _39060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39219_, _39218_, _31187_);
  and (_39220_, _39219_, _39217_);
  and (_39221_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39222_, _39221_, rst);
  or (_39223_, _39222_, _39220_);
  or (_40243_, _39223_, _39216_);
  and (_39224_, _39069_, _27595_);
  nand (_39225_, _39224_, _31732_);
  or (_39226_, _39076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39227_, _39226_, _31798_);
  and (_39228_, _39227_, _39225_);
  nand (_39229_, _39076_, _38123_);
  and (_39230_, _39229_, _31187_);
  and (_39231_, _39230_, _39226_);
  not (_39232_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_39233_, _31166_, _39232_);
  or (_39234_, _39233_, rst);
  or (_39235_, _39234_, _39231_);
  or (_40245_, _39235_, _39228_);
  and (_39236_, _39069_, _33016_);
  nand (_39237_, _39236_, _31732_);
  or (_39238_, _39236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39239_, _39238_, _31798_);
  and (_39240_, _39239_, _39237_);
  nand (_39241_, _39076_, _38115_);
  or (_39242_, _39076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39243_, _39242_, _31187_);
  and (_39244_, _39243_, _39241_);
  and (_39245_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39246_, _39245_, rst);
  or (_39247_, _39246_, _39244_);
  or (_40247_, _39247_, _39240_);
  and (_39248_, _39069_, _33713_);
  nand (_39249_, _39248_, _31732_);
  or (_39250_, _39248_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39251_, _39250_, _31798_);
  and (_39252_, _39251_, _39249_);
  nand (_39253_, _39076_, _38108_);
  or (_39254_, _39076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39255_, _39254_, _31187_);
  and (_39256_, _39255_, _39253_);
  and (_39257_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39258_, _39257_, rst);
  or (_39259_, _39258_, _39256_);
  or (_40249_, _39259_, _39252_);
  and (_39260_, _39069_, _34431_);
  nand (_39261_, _39260_, _31732_);
  or (_39262_, _39260_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39263_, _39262_, _31798_);
  and (_39264_, _39263_, _39261_);
  nand (_39265_, _39076_, _38100_);
  or (_39266_, _39076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39267_, _39266_, _31187_);
  and (_39268_, _39267_, _39265_);
  and (_39269_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39270_, _39269_, rst);
  or (_39271_, _39270_, _39268_);
  or (_40251_, _39271_, _39264_);
  and (_39272_, _39069_, _35226_);
  nand (_39273_, _39272_, _31732_);
  or (_39274_, _39272_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39275_, _39274_, _31798_);
  and (_39276_, _39275_, _39273_);
  nand (_39277_, _39076_, _38092_);
  or (_39278_, _39076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39279_, _39278_, _31187_);
  and (_39280_, _39279_, _39277_);
  and (_39281_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39282_, _39281_, rst);
  or (_39283_, _39282_, _39280_);
  or (_40253_, _39283_, _39276_);
  and (_39284_, _39069_, _36043_);
  nand (_39285_, _39284_, _31732_);
  or (_39286_, _39284_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39287_, _39286_, _31798_);
  and (_39288_, _39287_, _39285_);
  nand (_39289_, _39076_, _38085_);
  or (_39290_, _39076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39291_, _39290_, _31187_);
  and (_39292_, _39291_, _39289_);
  and (_39293_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39294_, _39293_, rst);
  or (_39295_, _39294_, _39292_);
  or (_40255_, _39295_, _39288_);
  and (_39296_, _39069_, _36782_);
  nand (_39297_, _39296_, _31732_);
  or (_39298_, _39296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39299_, _39298_, _31798_);
  and (_39300_, _39299_, _39297_);
  nand (_39301_, _39076_, _38078_);
  or (_39302_, _39076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39303_, _39302_, _31187_);
  and (_39314_, _39303_, _39301_);
  and (_39325_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39336_, _39325_, rst);
  or (_39347_, _39336_, _39314_);
  or (_40257_, _39347_, _39300_);
  nand (_39364_, _39093_, _31732_);
  or (_39365_, _39093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39366_, _39365_, _31798_);
  and (_39367_, _39366_, _39364_);
  nand (_39368_, _39093_, _38123_);
  and (_39369_, _39365_, _31187_);
  and (_39370_, _39369_, _39368_);
  not (_39371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_39372_, _31166_, _39371_);
  or (_39373_, _39372_, rst);
  or (_39374_, _39373_, _39370_);
  or (_40259_, _39374_, _39367_);
  and (_39375_, _39086_, _33016_);
  nand (_39376_, _39375_, _31732_);
  or (_39377_, _39375_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39378_, _39377_, _31798_);
  and (_39379_, _39378_, _39376_);
  nor (_39380_, _39094_, _38115_);
  and (_39381_, _39094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39382_, _39381_, _39380_);
  and (_39383_, _39382_, _31187_);
  and (_39384_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39385_, _39384_, rst);
  or (_39386_, _39385_, _39383_);
  or (_40261_, _39386_, _39379_);
  and (_39387_, _39086_, _33713_);
  nand (_39388_, _39387_, _31732_);
  or (_39389_, _39387_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39390_, _39389_, _31798_);
  and (_39391_, _39390_, _39388_);
  nor (_39392_, _39094_, _38108_);
  and (_39393_, _39094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39394_, _39393_, _39392_);
  and (_39395_, _39394_, _31187_);
  and (_39396_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39397_, _39396_, rst);
  or (_39398_, _39397_, _39395_);
  or (_40263_, _39398_, _39391_);
  and (_39399_, _39086_, _34431_);
  nand (_39400_, _39399_, _31732_);
  or (_39401_, _39399_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39402_, _39401_, _31798_);
  and (_39403_, _39402_, _39400_);
  nor (_39404_, _39094_, _38100_);
  and (_39405_, _39094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39406_, _39405_, _39404_);
  and (_39407_, _39406_, _31187_);
  and (_39408_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39409_, _39408_, rst);
  or (_39410_, _39409_, _39407_);
  or (_40265_, _39410_, _39403_);
  and (_39411_, _39086_, _35226_);
  nand (_39412_, _39411_, _31732_);
  or (_39413_, _39411_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39414_, _39413_, _31798_);
  and (_39415_, _39414_, _39412_);
  nor (_39416_, _39094_, _38092_);
  and (_39417_, _39094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39418_, _39417_, _39416_);
  and (_39419_, _39418_, _31187_);
  and (_39420_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39421_, _39420_, rst);
  or (_39422_, _39421_, _39419_);
  or (_40267_, _39422_, _39415_);
  and (_39424_, _39086_, _36043_);
  nand (_39430_, _39424_, _31732_);
  or (_39431_, _39424_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39432_, _39431_, _31798_);
  and (_39433_, _39432_, _39430_);
  nor (_39434_, _39094_, _38085_);
  and (_39435_, _39094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39436_, _39435_, _39434_);
  and (_39437_, _39436_, _31187_);
  and (_39438_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39439_, _39438_, rst);
  or (_39440_, _39439_, _39437_);
  or (_40269_, _39440_, _39433_);
  and (_39441_, _39086_, _36782_);
  nand (_39442_, _39441_, _31732_);
  or (_39443_, _39441_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39444_, _39443_, _31798_);
  and (_39445_, _39444_, _39442_);
  nor (_39446_, _39094_, _38078_);
  and (_39447_, _39094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39448_, _39447_, _39446_);
  and (_39449_, _39448_, _31187_);
  and (_39450_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39451_, _39450_, rst);
  or (_39452_, _39451_, _39449_);
  or (_40271_, _39452_, _39445_);
  and (_39453_, _39103_, _27595_);
  nand (_39454_, _39453_, _31732_);
  or (_39455_, _39112_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39456_, _39455_, _31798_);
  and (_39457_, _39456_, _39454_);
  nand (_39458_, _39112_, _38123_);
  and (_39459_, _39455_, _31187_);
  and (_39460_, _39459_, _39458_);
  not (_39461_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_39462_, _31166_, _39461_);
  or (_39463_, _39462_, rst);
  or (_39464_, _39463_, _39460_);
  or (_40272_, _39464_, _39457_);
  and (_39465_, _39103_, _33016_);
  nand (_39466_, _39465_, _31732_);
  or (_39467_, _39465_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39468_, _39467_, _31798_);
  and (_39469_, _39468_, _39466_);
  nor (_39470_, _39113_, _38115_);
  and (_39471_, _39113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39472_, _39471_, _39470_);
  and (_39473_, _39472_, _31187_);
  and (_39474_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39475_, _39474_, rst);
  or (_39476_, _39475_, _39473_);
  or (_40274_, _39476_, _39469_);
  and (_39477_, _39103_, _33713_);
  nand (_39478_, _39477_, _31732_);
  or (_39479_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39480_, _39479_, _31798_);
  and (_39481_, _39480_, _39478_);
  nor (_39482_, _39113_, _38108_);
  and (_39483_, _39113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39484_, _39483_, _39482_);
  and (_39485_, _39484_, _31187_);
  and (_39486_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39487_, _39486_, rst);
  or (_39488_, _39487_, _39485_);
  or (_40276_, _39488_, _39481_);
  and (_39489_, _39103_, _34431_);
  nand (_39490_, _39489_, _31732_);
  or (_39491_, _39489_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39492_, _39491_, _31798_);
  and (_39493_, _39492_, _39490_);
  nor (_39494_, _39113_, _38100_);
  and (_39495_, _39113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39496_, _39495_, _39494_);
  and (_39497_, _39496_, _31187_);
  and (_39498_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39499_, _39498_, rst);
  or (_39500_, _39499_, _39497_);
  or (_40278_, _39500_, _39493_);
  and (_39501_, _39103_, _35226_);
  nand (_39502_, _39501_, _31732_);
  or (_39503_, _39501_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39504_, _39503_, _31798_);
  and (_39508_, _39504_, _39502_);
  nor (_39516_, _39113_, _38092_);
  and (_39517_, _39113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39518_, _39517_, _39516_);
  and (_39519_, _39518_, _31187_);
  and (_39520_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39521_, _39520_, rst);
  or (_39522_, _39521_, _39519_);
  or (_40280_, _39522_, _39508_);
  and (_39523_, _39103_, _36043_);
  nand (_39524_, _39523_, _31732_);
  or (_39525_, _39523_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39526_, _39525_, _31798_);
  and (_39527_, _39526_, _39524_);
  nor (_39528_, _39113_, _38085_);
  and (_39529_, _39113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39530_, _39529_, _39528_);
  and (_39531_, _39530_, _31187_);
  and (_39532_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39533_, _39532_, rst);
  or (_39534_, _39533_, _39531_);
  or (_40282_, _39534_, _39527_);
  and (_39535_, _39103_, _36782_);
  nand (_39536_, _39535_, _31732_);
  or (_39537_, _39535_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39538_, _39537_, _31798_);
  and (_39539_, _39538_, _39536_);
  nor (_39540_, _39113_, _38078_);
  and (_39541_, _39113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39542_, _39541_, _39540_);
  and (_39543_, _39542_, _31187_);
  and (_39544_, _39143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39545_, _39544_, rst);
  or (_39546_, _39545_, _39543_);
  or (_40284_, _39546_, _39539_);
  and (_40734_, t0_i, _42545_);
  and (_40737_, t1_i, _42545_);
  not (_39547_, _31187_);
  nor (_39548_, _39547_, _28242_);
  and (_39549_, _39548_, _34431_);
  and (_39550_, _39549_, _38059_);
  nand (_39551_, _39550_, _38146_);
  nor (_39552_, _27332_, _28242_);
  and (_39553_, _39552_, _38060_);
  and (_39554_, _39553_, _31187_);
  not (_39555_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_39556_, _39555_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_39558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _39557_);
  nor (_39559_, _39558_, _39556_);
  or (_39560_, _39559_, _39554_);
  and (_39561_, _39560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_39562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_39563_, t1_i);
  and (_39564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _39563_);
  nor (_39565_, _39564_, _39562_);
  not (_39566_, _39565_);
  not (_39567_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_39568_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39567_);
  nor (_39569_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_39570_, _39569_);
  and (_39571_, _39570_, _39568_);
  and (_39572_, _39571_, _39566_);
  not (_39573_, _39572_);
  nand (_39574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_39575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_39576_, _39575_, _39574_);
  nor (_39577_, _39576_, _39573_);
  and (_39578_, _39577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_39579_, _39578_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_39580_, _39579_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_39581_, _39580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_39582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_39583_, _39576_, _39582_);
  and (_39588_, _39583_, _39572_);
  and (_39589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_39590_, _39589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_39591_, _39590_, _39588_);
  nor (_39592_, _39591_, _39559_);
  and (_39593_, _39592_, _39581_);
  and (_39594_, _39591_, _39556_);
  and (_39595_, _39594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39596_, _39595_, _39593_);
  nor (_39597_, _39596_, _39554_);
  or (_39598_, _39597_, _39561_);
  or (_39599_, _39550_, _39598_);
  and (_39600_, _39599_, _42545_);
  and (_40740_, _39600_, _39551_);
  not (_39601_, _39554_);
  nor (_39602_, _39601_, _38146_);
  and (_39603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39612_, _39603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39614_, _39612_, _39588_);
  and (_39615_, _39614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_39616_, _39615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39617_, _39616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_39618_, _39617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_39619_, _39618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39621_, _39620_);
  and (_39622_, _39618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39623_, _39622_, _39621_);
  and (_39624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not (_39625_, _39558_);
  and (_39626_, _39622_, _39590_);
  nor (_39627_, _39626_, _39625_);
  or (_39628_, _39627_, _39624_);
  or (_39629_, _39590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_39630_, _39629_, _39628_);
  or (_39631_, _39630_, _39623_);
  and (_39632_, _39631_, _39619_);
  and (_39633_, _39548_, _38195_);
  nor (_39634_, _39633_, _39554_);
  and (_39635_, _39634_, _39632_);
  and (_39636_, _39633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_39637_, _39636_, _39635_);
  or (_39638_, _39637_, _39602_);
  and (_40743_, _39638_, _42545_);
  and (_39639_, _39573_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_39640_, _39639_, _39626_);
  and (_39641_, _39640_, _39558_);
  or (_39642_, _39639_, _39622_);
  and (_39643_, _39642_, _39620_);
  nand (_39644_, _39572_, _39555_);
  and (_39645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_39646_, _39645_, _39644_);
  or (_39647_, _39646_, _39594_);
  or (_39648_, _39647_, _39643_);
  or (_39649_, _39648_, _39641_);
  and (_39650_, _39649_, _42545_);
  and (_40746_, _39650_, _39634_);
  and (_39651_, _39548_, _35226_);
  and (_39652_, _39651_, _38059_);
  nor (_39653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_39654_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_39655_, t0_i);
  and (_39656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _39655_);
  nor (_39657_, _39656_, _39654_);
  not (_39658_, _39657_);
  not (_39659_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_39660_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_39661_, _39660_, _39659_);
  and (_39662_, _39661_, _39658_);
  not (_39663_, _39662_);
  and (_39664_, _39663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_39665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_39666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_39667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_39668_, _39667_, _39666_);
  and (_39669_, _39668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_39670_, _39669_, _39662_);
  and (_39671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_39672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_39673_, _39672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_39674_, _39673_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_39675_, _39674_, _39671_);
  and (_39676_, _39675_, _39670_);
  and (_39677_, _39676_, _39665_);
  or (_39678_, _39677_, _39664_);
  and (_39679_, _39678_, _39653_);
  and (_39680_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_39681_, _39680_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_39682_, _39681_, _39670_);
  not (_39683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _39683_);
  and (_39685_, _39675_, _39665_);
  and (_39686_, _39685_, _39684_);
  or (_39687_, _39686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39688_, _39687_, _39682_);
  not (_39689_, _39653_);
  and (_39690_, _39664_, _39689_);
  or (_39691_, _39690_, _39688_);
  or (_39692_, _39691_, _39679_);
  nand (_39693_, _39692_, _42545_);
  nor (_39694_, _39693_, _39652_);
  and (_39695_, _39548_, _33713_);
  and (_39696_, _39695_, _38059_);
  not (_39697_, _39696_);
  and (_40749_, _39697_, _39694_);
  nand (_39698_, _39696_, _38146_);
  not (_39699_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand (_39700_, _39652_, _39699_);
  and (_39701_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_39702_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_39703_, _39702_, _39670_);
  or (_39704_, _39703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_39705_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_39706_, _39705_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand (_39707_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_39708_, _39707_, _39682_);
  and (_39709_, _39708_, _39689_);
  or (_39710_, _39709_, _39652_);
  and (_39711_, _39710_, _39704_);
  or (_39712_, _39711_, _39701_);
  and (_39713_, _39712_, _39700_);
  or (_39714_, _39713_, _39696_);
  and (_39715_, _39714_, _42545_);
  and (_40752_, _39715_, _39698_);
  or (_39716_, _39706_, _39684_);
  not (_39717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_39718_, _39681_, _39669_);
  and (_39719_, _39662_, _39683_);
  and (_39720_, _39719_, _39718_);
  and (_39721_, _39720_, _39675_);
  and (_39722_, _39721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_39723_, _39722_, _39717_);
  and (_39724_, _39722_, _39717_);
  or (_39725_, _39724_, _39723_);
  and (_39726_, _39725_, _39716_);
  and (_39727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39728_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_39729_, _39728_, _39674_);
  and (_39730_, _39729_, _39671_);
  and (_39731_, _39730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_39732_, _39731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_39733_, _39728_, _39685_);
  and (_39734_, _39733_, _39732_);
  and (_39735_, _39734_, _39727_);
  and (_39736_, _39676_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_39737_, _39736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_39738_, _39677_, _39689_);
  and (_39739_, _39738_, _39737_);
  or (_39740_, _39739_, _39735_);
  or (_39741_, _39740_, _39726_);
  or (_39742_, _39741_, _39652_);
  nand (_39743_, _39652_, _38146_);
  and (_39744_, _39743_, _39742_);
  or (_39745_, _39744_, _39696_);
  nand (_39746_, _39696_, _39717_);
  and (_39747_, _39746_, _42545_);
  and (_40755_, _39747_, _39745_);
  not (_39748_, _39728_);
  or (_39749_, _39748_, _39685_);
  or (_39750_, _39728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_39751_, _39727_, _42545_);
  and (_39752_, _39751_, _39750_);
  nand (_39753_, _39752_, _39749_);
  nor (_39754_, _39753_, _39652_);
  and (_40758_, _39754_, _39697_);
  and (_39755_, _39548_, _38066_);
  or (_39756_, _39755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_39757_, _39756_, _42545_);
  nand (_39758_, _39755_, _38146_);
  and (_40761_, _39758_, _39757_);
  not (_39759_, _39550_);
  not (_39760_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_39761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_39762_, _39761_, _39554_);
  and (_39763_, _39762_, _39572_);
  and (_39764_, _39763_, _39760_);
  nor (_39765_, _39763_, _39760_);
  or (_39766_, _39765_, _39764_);
  and (_39767_, _39766_, _39759_);
  and (_39768_, _39550_, _38124_);
  nor (_39769_, _39550_, _39554_);
  and (_39770_, _39590_, _39583_);
  and (_39771_, _39770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39772_, _39771_, _39556_);
  and (_39773_, _39772_, _39769_);
  or (_39774_, _39773_, _39768_);
  or (_39775_, _39774_, _39767_);
  and (_41247_, _39775_, _42545_);
  not (_39776_, _39633_);
  nand (_39777_, _39776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_39778_, _39777_, _39762_);
  not (_39779_, _39761_);
  and (_39780_, _39572_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_39781_, _39780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_39782_, _39780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_39783_, _39782_, _39781_);
  and (_39784_, _39783_, _39779_);
  and (_39785_, _39594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_39786_, _39785_, _39784_);
  and (_39787_, _39786_, _39634_);
  nor (_39788_, _39759_, _38115_);
  or (_39789_, _39788_, _39787_);
  or (_39790_, _39789_, _39778_);
  and (_41249_, _39790_, _42545_);
  nor (_39791_, _39782_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_39792_, _39782_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_39793_, _39792_, _39791_);
  and (_39794_, _39793_, _39779_);
  and (_39795_, _39594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_39796_, _39795_, _39794_);
  and (_39797_, _39796_, _39634_);
  nand (_39798_, _39776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_39799_, _39798_, _39762_);
  or (_39800_, _39799_, _39797_);
  nor (_39801_, _39776_, _38108_);
  or (_39802_, _39801_, _39800_);
  and (_41251_, _39802_, _42545_);
  or (_39803_, _39792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_39804_, _39761_, _39577_);
  and (_39805_, _39804_, _39803_);
  and (_39806_, _39594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_39807_, _39806_, _39805_);
  and (_39808_, _39807_, _39634_);
  nand (_39809_, _39776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_39810_, _39809_, _39762_);
  or (_39811_, _39810_, _39808_);
  nor (_39812_, _39776_, _38100_);
  or (_39813_, _39812_, _39811_);
  and (_41253_, _39813_, _42545_);
  or (_39814_, _39577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_39815_, _39761_, _39588_);
  and (_39816_, _39815_, _39814_);
  and (_39817_, _39594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_39818_, _39817_, _39816_);
  and (_39819_, _39818_, _39634_);
  or (_39820_, _39633_, _39582_);
  nor (_39821_, _39820_, _39762_);
  or (_39822_, _39821_, _39819_);
  nor (_39823_, _39776_, _38092_);
  or (_39824_, _39823_, _39822_);
  and (_41254_, _39824_, _42545_);
  or (_39825_, _39588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_39826_, _39588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_39827_, _39826_, _39559_);
  and (_39828_, _39827_, _39825_);
  and (_39829_, _39594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_39830_, _39829_, _39828_);
  and (_39831_, _39830_, _39634_);
  and (_39832_, _39776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_39833_, _39832_, _39560_);
  or (_39834_, _39833_, _39831_);
  nor (_39835_, _39776_, _38085_);
  or (_39836_, _39835_, _39834_);
  and (_41256_, _39836_, _42545_);
  and (_39837_, _39556_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_39838_, _39837_, _39572_);
  and (_39839_, _39838_, _39770_);
  nor (_39840_, _39826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_39841_, _39840_, _39559_);
  nor (_39842_, _39841_, _39580_);
  or (_39843_, _39842_, _39839_);
  and (_39844_, _39843_, _39634_);
  and (_39845_, _39776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_39846_, _39845_, _39560_);
  or (_39847_, _39846_, _39844_);
  nor (_39848_, _39776_, _38078_);
  or (_39849_, _39848_, _39847_);
  and (_41258_, _39849_, _42545_);
  and (_39850_, _39554_, _38124_);
  and (_39851_, _39633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39852_, _39588_, _39557_);
  nor (_39853_, _39590_, _39555_);
  not (_39854_, _39853_);
  and (_39855_, _39854_, _39852_);
  nand (_39856_, _39855_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_39857_, _39855_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39858_, _39857_, _39856_);
  and (_39859_, _39858_, _39634_);
  or (_39860_, _39859_, _39851_);
  or (_39861_, _39860_, _39850_);
  and (_41260_, _39861_, _42545_);
  nor (_39862_, _39601_, _38115_);
  and (_39863_, _39633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not (_39864_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_39865_, _39591_, _39625_);
  not (_39866_, _39865_);
  not (_39867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_39868_, _39852_, _39558_);
  nor (_39869_, _39868_, _39867_);
  and (_39870_, _39869_, _39866_);
  nor (_39871_, _39870_, _39864_);
  and (_39872_, _39870_, _39864_);
  or (_39873_, _39872_, _39871_);
  and (_39874_, _39873_, _39634_);
  or (_39875_, _39874_, _39863_);
  or (_39876_, _39875_, _39862_);
  and (_41262_, _39876_, _42545_);
  nor (_39877_, _39601_, _38108_);
  nand (_39878_, _39614_, _39557_);
  nand (_39879_, _39854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_39880_, _39879_, _39878_);
  and (_39881_, _39620_, _39583_);
  and (_39882_, _39770_, _39558_);
  or (_39883_, _39882_, _39881_);
  and (_39884_, _39603_, _39572_);
  and (_39885_, _39884_, _39883_);
  or (_39886_, _39885_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39887_, _39886_, _39880_);
  and (_39888_, _39887_, _39634_);
  and (_39889_, _39633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_39890_, _39889_, _39888_);
  or (_39891_, _39890_, _39877_);
  and (_41264_, _39891_, _42545_);
  nand (_39892_, _39554_, _38100_);
  and (_39893_, _39615_, _39590_);
  and (_39894_, _39614_, _39590_);
  or (_39895_, _39894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_39896_, _39895_, _39558_);
  nor (_39897_, _39896_, _39893_);
  and (_39898_, _39878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_39899_, _39878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_39900_, _39899_, _39898_);
  and (_39901_, _39900_, _39625_);
  or (_39902_, _39901_, _39897_);
  or (_39903_, _39902_, _39554_);
  and (_39904_, _39903_, _39759_);
  and (_39905_, _39904_, _39892_);
  and (_39906_, _39550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_39907_, _39906_, _39905_);
  and (_41266_, _39907_, _42545_);
  nor (_39908_, _39601_, _38092_);
  and (_39909_, _39633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_39910_, _39893_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_39911_, _39910_, _39558_);
  and (_39912_, _39893_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_39913_, _39912_, _39911_);
  and (_39914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39915_, _39603_, _39583_);
  and (_39916_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39917_, _39916_, _39572_);
  and (_39918_, _39917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_39919_, _39918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_39920_, _39918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39921_, _39920_, _39919_);
  and (_39922_, _39921_, _39620_);
  or (_39923_, _39922_, _39914_);
  or (_39924_, _39923_, _39913_);
  and (_39925_, _39924_, _39634_);
  or (_39926_, _39925_, _39909_);
  or (_39927_, _39926_, _39908_);
  and (_41268_, _39927_, _42545_);
  nand (_39928_, _39554_, _38085_);
  and (_39929_, _39616_, _39620_);
  and (_39930_, _39912_, _39558_);
  nor (_39931_, _39930_, _39929_);
  and (_39932_, _39931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_39933_, _39931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_39934_, _39933_, _39932_);
  or (_39935_, _39934_, _39554_);
  and (_39936_, _39935_, _39759_);
  and (_39937_, _39936_, _39928_);
  and (_39938_, _39550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_39939_, _39938_, _39937_);
  and (_41270_, _39939_, _42545_);
  nand (_39940_, _39554_, _38078_);
  nor (_39941_, _39853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_39942_, _39941_, _39617_);
  or (_39943_, _39942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_39944_, _39942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_39945_, _39944_, _39943_);
  or (_39946_, _39945_, _39554_);
  and (_39947_, _39946_, _39759_);
  and (_39948_, _39947_, _39940_);
  and (_39949_, _39550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_39950_, _39949_, _39948_);
  and (_41271_, _39950_, _42545_);
  and (_39951_, _39548_, _38291_);
  nor (_39952_, _39663_, _39652_);
  or (_39953_, _39952_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_39954_, _39662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_39955_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_39956_, _39955_, _39718_);
  nand (_39957_, _39956_, _39954_);
  or (_39958_, _39957_, _39652_);
  and (_39959_, _39958_, _39953_);
  or (_39960_, _39959_, _39951_);
  nand (_39961_, _39696_, _38123_);
  and (_39962_, _39961_, _42545_);
  and (_41273_, _39962_, _39960_);
  nor (_39963_, _39954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_39964_, _39954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_39965_, _39964_, _39963_);
  and (_39966_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_39967_, _39966_, _39682_);
  nor (_39968_, _39967_, _39965_);
  nor (_39969_, _39968_, _39652_);
  and (_39970_, _39652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_39971_, _39970_, _39969_);
  and (_39972_, _39971_, _39697_);
  nor (_39973_, _39697_, _38115_);
  or (_39974_, _39973_, _39972_);
  and (_41275_, _39974_, _42545_);
  nand (_39975_, _39951_, _38108_);
  and (_39976_, _39652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_39977_, _39964_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_39978_, _39954_, _39666_);
  nor (_39979_, _39978_, _39977_);
  and (_39980_, _39706_, _39682_);
  and (_39981_, _39980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_39982_, _39981_, _39979_);
  nor (_39983_, _39982_, _39652_);
  or (_39984_, _39983_, _39976_);
  or (_39985_, _39984_, _39951_);
  and (_39986_, _39985_, _42545_);
  and (_41277_, _39986_, _39975_);
  nand (_39987_, _39951_, _38100_);
  and (_39988_, _39652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_39989_, _39668_, _39662_);
  nor (_39990_, _39978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_39991_, _39990_, _39989_);
  and (_39992_, _39980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_39993_, _39992_, _39991_);
  nor (_39994_, _39993_, _39652_);
  or (_39995_, _39994_, _39988_);
  or (_39996_, _39995_, _39951_);
  and (_39997_, _39996_, _42545_);
  and (_41279_, _39997_, _39987_);
  nand (_39998_, _39951_, _38092_);
  and (_39999_, _39652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40000_, _39989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40001_, _40000_, _39670_);
  and (_40002_, _39980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_40003_, _40002_, _40001_);
  nor (_40004_, _40003_, _39652_);
  or (_40005_, _40004_, _39999_);
  or (_40006_, _40005_, _39951_);
  and (_40007_, _40006_, _42545_);
  and (_41281_, _40007_, _39998_);
  nand (_40008_, _39951_, _38085_);
  and (_40009_, _39652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_40010_, _39670_, _39689_);
  and (_40011_, _40010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_40012_, _40010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_40013_, _40012_, _40011_);
  and (_40014_, _39980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_40015_, _40014_, _40013_);
  nor (_40016_, _40015_, _39652_);
  or (_40017_, _40016_, _40009_);
  or (_40018_, _40017_, _39951_);
  and (_40019_, _40018_, _42545_);
  and (_41283_, _40019_, _40008_);
  and (_40020_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_40021_, _40020_, _39662_);
  and (_40022_, _40021_, _39718_);
  not (_40023_, _40011_);
  nor (_40024_, _40023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_40025_, _40024_, _40022_);
  nor (_40026_, _40025_, _39652_);
  or (_40027_, _40023_, _39652_);
  and (_40028_, _40027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_40029_, _40028_, _40026_);
  and (_40030_, _40029_, _39697_);
  nor (_40031_, _39697_, _38078_);
  or (_40032_, _40031_, _40030_);
  and (_41285_, _40032_, _42545_);
  or (_40033_, _39720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40034_, _40033_, _39716_);
  and (_40035_, _39720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_40036_, _40035_, _40034_);
  and (_40037_, _39728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40038_, _39728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40039_, _40038_, _39727_);
  nor (_40040_, _40039_, _40037_);
  and (_40041_, _39670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40042_, _39670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40043_, _40042_, _39653_);
  nor (_40044_, _40043_, _40041_);
  or (_40045_, _40044_, _40040_);
  or (_40046_, _40045_, _40036_);
  or (_40047_, _40046_, _39652_);
  nand (_40048_, _39652_, _38123_);
  and (_40049_, _40048_, _40047_);
  or (_40050_, _40049_, _39696_);
  or (_40051_, _39697_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_40052_, _40051_, _42545_);
  and (_41287_, _40052_, _40050_);
  nand (_40053_, _39652_, _38115_);
  or (_40054_, _40035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40055_, _39718_, _39662_);
  and (_40056_, _40055_, _39672_);
  not (_40057_, _40056_);
  or (_40058_, _40057_, _39706_);
  and (_40059_, _40058_, _39716_);
  and (_40060_, _40059_, _40054_);
  and (_40061_, _39728_, _39672_);
  or (_40062_, _40037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_40063_, _40062_, _39727_);
  nor (_40064_, _40063_, _40061_);
  or (_40065_, _40041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40066_, _40041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_40067_, _40066_, _39689_);
  and (_40068_, _40067_, _40065_);
  or (_40069_, _40068_, _40064_);
  or (_40070_, _40069_, _40060_);
  or (_40071_, _40070_, _39652_);
  and (_40072_, _40071_, _40053_);
  or (_40073_, _40072_, _39696_);
  or (_40074_, _39697_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40075_, _40074_, _42545_);
  and (_41288_, _40075_, _40073_);
  nand (_40076_, _39652_, _38108_);
  and (_40077_, _39672_, _39662_);
  and (_40078_, _40077_, _39669_);
  or (_40079_, _40078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40080_, _39673_, _39670_);
  nor (_40081_, _40080_, _39689_);
  and (_40082_, _40081_, _40079_);
  or (_40083_, _40056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40084_, _40055_, _39673_);
  not (_40085_, _40084_);
  and (_40086_, _40085_, _39684_);
  and (_40087_, _40086_, _40083_);
  and (_40088_, _40061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_40089_, _40088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40090_, _39728_, _39673_);
  nand (_40091_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40092_, _40091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40093_, _40092_, _40089_);
  or (_40094_, _40093_, _40087_);
  or (_40095_, _40094_, _40082_);
  or (_40096_, _40095_, _39652_);
  and (_40097_, _40096_, _40076_);
  or (_40098_, _40097_, _39696_);
  or (_40099_, _39697_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40100_, _40099_, _42545_);
  and (_41290_, _40100_, _40098_);
  nand (_40101_, _39652_, _38100_);
  not (_40102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40103_, _40084_, _39683_);
  nor (_40104_, _40103_, _40102_);
  and (_40105_, _40103_, _40102_);
  or (_40106_, _40105_, _40104_);
  and (_40107_, _40106_, _39716_);
  or (_40108_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_40109_, _39729_);
  and (_40110_, _40109_, _39727_);
  and (_40111_, _40110_, _40108_);
  or (_40112_, _40080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40113_, _39674_, _39670_);
  nor (_40114_, _40113_, _39689_);
  and (_40115_, _40114_, _40112_);
  or (_40116_, _40115_, _40111_);
  or (_40117_, _40116_, _40107_);
  or (_40118_, _40117_, _39652_);
  and (_40119_, _40118_, _40101_);
  or (_40120_, _40119_, _39696_);
  nand (_40121_, _39696_, _40102_);
  and (_40122_, _40121_, _42545_);
  and (_41292_, _40122_, _40120_);
  nand (_40123_, _39652_, _38092_);
  or (_40124_, _40113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40125_, _40078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40126_, _40125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40127_, _40126_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_40128_, _40127_, _39689_);
  and (_40129_, _40128_, _40124_);
  and (_40130_, _40055_, _39674_);
  or (_40131_, _40130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_40132_, _40130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40133_, _40132_, _39684_);
  and (_40134_, _40133_, _40131_);
  and (_40135_, _39729_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_40136_, _40135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40137_, _40136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40138_, _39729_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_40139_, _40138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40140_, _40139_, _40137_);
  or (_40141_, _40140_, _40134_);
  or (_40142_, _40141_, _40129_);
  or (_40143_, _40142_, _39652_);
  and (_40144_, _40143_, _40123_);
  or (_40145_, _40144_, _39696_);
  or (_40146_, _39697_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40147_, _40146_, _42545_);
  and (_41294_, _40147_, _40145_);
  nand (_40148_, _39652_, _38085_);
  not (_40149_, _40127_);
  nor (_40150_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40151_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_40152_, _40151_, _40150_);
  and (_40153_, _40152_, _39653_);
  nor (_40154_, _40132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_40155_, _40154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_40156_, _40154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40157_, _40156_, _39716_);
  and (_40158_, _40157_, _40155_);
  not (_40159_, _39730_);
  and (_40160_, _40159_, _39727_);
  or (_40161_, _40138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40162_, _40161_, _40160_);
  or (_40163_, _40162_, _40158_);
  or (_40164_, _40163_, _40153_);
  nor (_40165_, _40164_, _39652_);
  nor (_40166_, _40165_, _39951_);
  and (_40167_, _40166_, _40148_);
  and (_40168_, _39696_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_40169_, _40168_, _40167_);
  and (_41296_, _40169_, _42545_);
  or (_40170_, _39721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_40171_, _40170_, _39716_);
  nor (_40172_, _40171_, _39722_);
  or (_40173_, _39730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_40174_, _39731_);
  and (_40175_, _40174_, _39727_);
  and (_40176_, _40175_, _40173_);
  or (_40177_, _39676_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_40178_, _39736_, _39689_);
  and (_40179_, _40178_, _40177_);
  or (_40180_, _40179_, _40176_);
  nor (_40181_, _40180_, _40172_);
  nor (_40182_, _40181_, _39652_);
  not (_40183_, _38078_);
  and (_40184_, _39652_, _40183_);
  or (_40185_, _40184_, _40182_);
  and (_40186_, _40185_, _39697_);
  and (_40187_, _39696_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40188_, _40187_, _40186_);
  and (_41298_, _40188_, _42545_);
  nor (_40189_, _39755_, _39705_);
  and (_40190_, _39755_, _38124_);
  or (_40191_, _40190_, _40189_);
  and (_41300_, _40191_, _42545_);
  or (_40192_, _39755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40193_, _40192_, _42545_);
  nand (_40194_, _39755_, _38115_);
  and (_41302_, _40194_, _40193_);
  or (_40195_, _39755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_40196_, _40195_, _42545_);
  nand (_40197_, _39755_, _38108_);
  and (_41304_, _40197_, _40196_);
  or (_40198_, _39755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_40199_, _40198_, _42545_);
  nand (_40200_, _39755_, _38100_);
  and (_41305_, _40200_, _40199_);
  or (_40201_, _39755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_40202_, _40201_, _42545_);
  nand (_40203_, _39755_, _38092_);
  and (_41307_, _40203_, _40202_);
  or (_40204_, _39755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_40205_, _40204_, _42545_);
  nand (_40206_, _39755_, _38085_);
  and (_41309_, _40206_, _40205_);
  or (_40207_, _39755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_40208_, _40207_, _42545_);
  nand (_40209_, _39755_, _38078_);
  and (_41311_, _40209_, _40208_);
  and (_40210_, _38061_, _31755_);
  and (_40211_, _40210_, _39111_);
  not (_40212_, _28417_);
  nor (_40213_, _38747_, _28242_);
  nand (_40214_, _40213_, _40212_);
  nor (_40215_, _40214_, _28088_);
  and (_40216_, _40215_, _39085_);
  and (_40217_, _40216_, _31755_);
  nand (_40218_, _40217_, _31732_);
  or (_40219_, _40217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_40220_, _40219_, _40218_);
  or (_40221_, _40220_, _40211_);
  nand (_40222_, _40211_, _38146_);
  and (_40223_, _40222_, _42545_);
  and (_42479_, _40223_, _40221_);
  and (_40224_, _39548_, _27595_);
  and (_40225_, _40224_, _39092_);
  not (_40226_, _40225_);
  and (_40227_, _28417_, _28253_);
  and (_40228_, _40227_, _38748_);
  and (_40229_, _40228_, _39085_);
  and (_40230_, _40229_, _31755_);
  or (_40231_, _40230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40233_, _40231_, _40226_);
  nand (_40235_, _40230_, _31732_);
  and (_40237_, _40235_, _40233_);
  nor (_40239_, _40226_, _38146_);
  or (_40241_, _40239_, _40237_);
  and (_42482_, _40241_, _42545_);
  and (_40244_, _40224_, _38059_);
  and (_40246_, _40213_, _28417_);
  and (_40248_, _40246_, _28099_);
  and (_40250_, _40248_, _39053_);
  nand (_40252_, _40250_, _27573_);
  and (_40254_, _40252_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40256_, _40254_, _40244_);
  or (_40258_, _27584_, _33702_);
  and (_40260_, _40258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40262_, _40260_, _38722_);
  and (_40264_, _40262_, _40250_);
  or (_40266_, _40264_, _40256_);
  nand (_40268_, _40244_, _38078_);
  and (_40270_, _40268_, _42545_);
  and (_42484_, _40270_, _40266_);
  not (_40273_, _40244_);
  nor (_40275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_40277_, _40275_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_40279_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_40281_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_40283_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40285_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40283_);
  and (_40286_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40287_, _40286_, _40285_);
  nor (_40288_, _40287_, _40281_);
  or (_40289_, _40288_, _40279_);
  and (_40290_, _40283_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40291_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_40292_, _40291_, _40290_);
  nor (_40293_, _40292_, _40281_);
  and (_40294_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40283_);
  and (_40295_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40296_, _40295_, _40294_);
  nand (_40297_, _40296_, _40293_);
  or (_40298_, _40297_, _40289_);
  and (_40299_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_40300_, _40299_, _40277_);
  and (_40301_, _38059_, _31755_);
  and (_40302_, _40301_, _40213_);
  or (_40303_, _40302_, _40300_);
  and (_40304_, _40303_, _40273_);
  nand (_40305_, _40302_, _31732_);
  and (_40306_, _40305_, _40304_);
  nor (_40307_, _40273_, _38146_);
  or (_40308_, _40307_, _40306_);
  and (_42487_, _40308_, _42545_);
  and (_40309_, _39553_, _31798_);
  nand (_40310_, _40309_, _31732_);
  not (_40311_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_40312_, _40311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_40313_, _40296_, _40281_);
  not (_40314_, _40313_);
  or (_40315_, _40314_, _40293_);
  or (_40316_, _40315_, _40289_);
  and (_40317_, _40316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_40318_, _40317_, _40312_);
  or (_40319_, _40318_, _40309_);
  and (_40320_, _40319_, _40273_);
  and (_40321_, _40320_, _40310_);
  nor (_40327_, _40273_, _38085_);
  or (_40333_, _40327_, _40321_);
  and (_42489_, _40333_, _42545_);
  not (_40344_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_40348_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40344_);
  nand (_40349_, _40288_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_40350_, _40313_, _40293_);
  or (_40351_, _40350_, _40349_);
  and (_40352_, _40351_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_40353_, _40352_, _40348_);
  and (_40354_, _40213_, _38066_);
  or (_40355_, _40354_, _40353_);
  and (_40356_, _40355_, _40273_);
  nand (_40357_, _40354_, _31732_);
  and (_40358_, _40357_, _40356_);
  nor (_40359_, _40273_, _38115_);
  or (_40360_, _40359_, _40358_);
  and (_42491_, _40360_, _42545_);
  and (_40365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_40369_, _40349_, _40315_);
  and (_40371_, _40369_, _40365_);
  and (_40372_, _40213_, _38195_);
  or (_40373_, _40372_, _40371_);
  and (_40377_, _40373_, _40273_);
  nand (_40383_, _40372_, _31732_);
  and (_40384_, _40383_, _40377_);
  nor (_40385_, _40273_, _38100_);
  or (_40386_, _40385_, _40384_);
  and (_42493_, _40386_, _42545_);
  nand (_40395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_40396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40283_);
  and (_40397_, _40396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40402_, _40397_, _40395_);
  or (_40407_, _40402_, _40281_);
  and (_40408_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40409_, _40408_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_40411_, _40409_);
  and (_40417_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40420_, _40417_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_40421_, _40420_);
  and (_40422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40428_, _40422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_40433_, _40432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_40434_, _40433_, _40428_);
  and (_40440_, _40434_, _40421_);
  and (_40444_, _40440_, _40411_);
  not (_40445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_40450_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_40451_, _40450_, _40445_);
  nand (_40456_, _40451_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_40457_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_40459_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_40460_, _40459_, _40457_);
  and (_40466_, _40460_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_40469_, _40466_);
  and (_40470_, _40469_, _40456_);
  nand (_40471_, _40470_, _40444_);
  and (_40477_, _40471_, _40407_);
  and (_40481_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_40482_, _40481_, _40283_);
  and (_40483_, _40482_, _40477_);
  not (_40489_, _40483_);
  not (_40493_, _40482_);
  and (_40494_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40281_);
  not (_40499_, _40494_);
  not (_40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40505_, _40417_, _40500_);
  not (_40506_, _40505_);
  not (_40507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40511_, _40422_, _40507_);
  not (_40517_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40518_, _40432_, _40517_);
  nor (_40519_, _40518_, _40511_);
  and (_40522_, _40519_, _40506_);
  nor (_40529_, _40522_, _40499_);
  not (_40530_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40531_, _40451_, _40530_);
  not (_40534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40540_, _40460_, _40534_);
  nor (_40542_, _40540_, _40531_);
  not (_40543_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40546_, _40408_, _40543_);
  not (_40552_, _40546_);
  and (_40553_, _40552_, _40542_);
  nor (_40554_, _40553_, _40499_);
  nor (_40555_, _40554_, _40529_);
  or (_40556_, _40555_, _40493_);
  and (_40557_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42545_);
  and (_40558_, _40557_, _40556_);
  and (_42531_, _40558_, _40489_);
  nor (_40559_, _40481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40560_, _40559_);
  not (_40561_, _40477_);
  and (_40562_, _40555_, _40561_);
  nor (_40563_, _40562_, _40560_);
  nand (_40564_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42545_);
  nor (_42533_, _40564_, _40563_);
  and (_40565_, _40470_, _40411_);
  nand (_40566_, _40565_, _40477_);
  or (_40567_, _40554_, _40477_);
  and (_40568_, _40567_, _40482_);
  and (_40569_, _40568_, _40566_);
  or (_40570_, _40569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_40571_, _40489_, _40440_);
  nor (_40572_, _40493_, _40477_);
  nand (_40573_, _40572_, _40529_);
  and (_40574_, _40573_, _42545_);
  and (_40575_, _40574_, _40571_);
  and (_42535_, _40575_, _40570_);
  and (_40576_, _40566_, _40559_);
  or (_40577_, _40576_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40578_, _40559_, _40477_);
  not (_40579_, _40578_);
  or (_40580_, _40579_, _40440_);
  or (_40581_, _40554_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_40582_, _40559_, _40529_);
  and (_40583_, _40582_, _40581_);
  or (_40584_, _40583_, _40477_);
  and (_40585_, _40584_, _42545_);
  and (_40586_, _40585_, _40580_);
  and (_42537_, _40586_, _40577_);
  nand (_40587_, _40562_, _40281_);
  nor (_40588_, _40283_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_40589_, _40588_, _40481_);
  and (_40590_, _40589_, _42545_);
  and (_42539_, _40590_, _40587_);
  and (_40591_, _40562_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_40592_, _40283_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_40593_, _40592_, _40588_);
  nor (_40594_, _40593_, _40561_);
  or (_40595_, _40594_, _40481_);
  or (_40596_, _40595_, _40591_);
  not (_40597_, _40481_);
  or (_40598_, _40593_, _40597_);
  and (_40599_, _40598_, _42545_);
  and (_42541_, _40599_, _40596_);
  and (_40600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42545_);
  and (_42543_, _40600_, _40481_);
  nor (_42548_, _40275_, rst);
  and (_42549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _42545_);
  nor (_40601_, _40562_, _40481_);
  and (_40602_, _40481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_40603_, _40602_, _40601_);
  and (_00130_, _40603_, _42545_);
  and (_40604_, _40481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_40605_, _40604_, _40601_);
  and (_00132_, _40605_, _42545_);
  and (_40606_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42545_);
  and (_00134_, _40606_, _40481_);
  nor (_40607_, _40555_, _40477_);
  not (_40608_, _40518_);
  nor (_40609_, _40540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_40610_, _40609_, _40531_);
  or (_40611_, _40610_, _40546_);
  and (_40612_, _40611_, _40608_);
  or (_40613_, _40612_, _40511_);
  and (_40614_, _40613_, _40506_);
  and (_40615_, _40614_, _40607_);
  not (_40616_, _40433_);
  or (_40617_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40618_, _40617_, _40456_);
  or (_40619_, _40618_, _40409_);
  and (_40620_, _40619_, _40616_);
  or (_40621_, _40620_, _40428_);
  and (_40622_, _40477_, _40421_);
  and (_40623_, _40622_, _40621_);
  or (_40624_, _40623_, _40481_);
  or (_40625_, _40624_, _40615_);
  or (_40626_, _40597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40627_, _40626_, _42545_);
  and (_00136_, _40627_, _40625_);
  not (_40628_, _40428_);
  or (_40629_, _40433_, _40409_);
  and (_40630_, _40470_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_40631_, _40630_, _40629_);
  and (_40632_, _40631_, _40628_);
  and (_40633_, _40632_, _40622_);
  nor (_40634_, _40511_, _40505_);
  or (_40635_, _40546_, _40518_);
  and (_40636_, _40542_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_40637_, _40636_, _40635_);
  and (_40638_, _40637_, _40634_);
  and (_40639_, _40638_, _40607_);
  or (_40640_, _40639_, _40481_);
  or (_40641_, _40640_, _40633_);
  or (_40642_, _40597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_40643_, _40642_, _42545_);
  and (_00138_, _40643_, _40641_);
  and (_40644_, _40552_, _40494_);
  nand (_40645_, _40644_, _40522_);
  or (_40646_, _40645_, _40542_);
  nor (_40647_, _40646_, _40477_);
  nand (_40648_, _40444_, _40407_);
  nor (_40649_, _40648_, _40470_);
  or (_40650_, _40649_, _40481_);
  or (_40651_, _40650_, _40647_);
  or (_40652_, _40597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_40653_, _40652_, _42545_);
  and (_00140_, _40653_, _40651_);
  and (_40654_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42545_);
  and (_00141_, _40654_, _40481_);
  and (_40655_, _40481_, _40283_);
  or (_40656_, _40655_, _40563_);
  or (_40657_, _40656_, _40572_);
  and (_00143_, _40657_, _42545_);
  not (_40658_, _40601_);
  and (_40659_, _40658_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_40660_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40283_);
  or (_40661_, _40660_, _40421_);
  and (_40662_, _40661_, _40477_);
  not (_40663_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_40664_, _40466_, _40283_);
  or (_40665_, _40664_, _40663_);
  nor (_40666_, _40456_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40667_, _40666_, _40409_);
  nand (_40668_, _40667_, _40665_);
  or (_40669_, _40411_, _40286_);
  and (_40670_, _40669_, _40668_);
  or (_40671_, _40670_, _40433_);
  or (_40672_, _40660_, _40616_);
  and (_40673_, _40672_, _40628_);
  and (_40674_, _40673_, _40671_);
  and (_40675_, _40428_, _40286_);
  or (_40676_, _40675_, _40420_);
  or (_40677_, _40676_, _40674_);
  and (_40678_, _40677_, _40662_);
  or (_40679_, _40660_, _40506_);
  and (_40680_, _40540_, _40283_);
  or (_40681_, _40680_, _40663_);
  and (_40682_, _40531_, _40283_);
  nor (_40683_, _40682_, _40546_);
  nand (_40684_, _40683_, _40681_);
  or (_40685_, _40552_, _40286_);
  and (_40686_, _40685_, _40684_);
  or (_40687_, _40686_, _40518_);
  not (_40688_, _40511_);
  or (_40689_, _40660_, _40608_);
  and (_40690_, _40689_, _40688_);
  and (_40691_, _40690_, _40687_);
  and (_40692_, _40511_, _40286_);
  or (_40693_, _40692_, _40505_);
  or (_40694_, _40693_, _40691_);
  and (_40695_, _40694_, _40607_);
  and (_40696_, _40695_, _40679_);
  or (_40697_, _40696_, _40678_);
  and (_40698_, _40697_, _40597_);
  or (_40699_, _40698_, _40659_);
  and (_00145_, _40699_, _42545_);
  and (_40700_, _40658_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40701_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40283_);
  and (_40702_, _40701_, _40421_);
  or (_40703_, _40702_, _40440_);
  or (_40704_, _40664_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40705_, _40704_, _40667_);
  nand (_40706_, _40409_, _40295_);
  nand (_40707_, _40706_, _40434_);
  or (_40708_, _40707_, _40705_);
  and (_40709_, _40708_, _40703_);
  and (_40710_, _40420_, _40295_);
  or (_40711_, _40710_, _40709_);
  and (_40712_, _40711_, _40477_);
  and (_40713_, _40505_, _40295_);
  and (_40714_, _40701_, _40506_);
  or (_40715_, _40714_, _40522_);
  and (_40716_, _40546_, _40295_);
  not (_40717_, _40519_);
  or (_40718_, _40680_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40719_, _40718_, _40683_);
  or (_40720_, _40719_, _40717_);
  or (_40721_, _40720_, _40716_);
  and (_40722_, _40721_, _40715_);
  or (_40723_, _40722_, _40713_);
  and (_40724_, _40723_, _40607_);
  or (_40725_, _40724_, _40712_);
  and (_40726_, _40725_, _40597_);
  or (_40727_, _40726_, _40700_);
  and (_00147_, _40727_, _42545_);
  and (_40728_, _40658_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_40729_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40730_, _40729_, _40421_);
  and (_40731_, _40730_, _40477_);
  not (_40732_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_40733_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40735_, _40733_, _40732_);
  nor (_40736_, _40456_, _40283_);
  nor (_40738_, _40736_, _40409_);
  nand (_40739_, _40738_, _40735_);
  or (_40741_, _40411_, _40285_);
  and (_40742_, _40741_, _40739_);
  or (_40744_, _40742_, _40433_);
  or (_40745_, _40729_, _40616_);
  and (_40747_, _40745_, _40628_);
  and (_40748_, _40747_, _40744_);
  and (_40750_, _40428_, _40285_);
  or (_40751_, _40750_, _40420_);
  or (_40753_, _40751_, _40748_);
  and (_40754_, _40753_, _40731_);
  or (_40756_, _40729_, _40506_);
  and (_40757_, _40540_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40759_, _40757_, _40732_);
  and (_40760_, _40531_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40762_, _40760_, _40546_);
  nand (_40763_, _40762_, _40759_);
  or (_40764_, _40552_, _40285_);
  and (_40765_, _40764_, _40763_);
  or (_40766_, _40765_, _40518_);
  or (_40767_, _40729_, _40608_);
  and (_40768_, _40767_, _40688_);
  and (_40769_, _40768_, _40766_);
  and (_40770_, _40511_, _40285_);
  or (_40771_, _40770_, _40505_);
  or (_40772_, _40771_, _40769_);
  and (_40773_, _40772_, _40607_);
  and (_40774_, _40773_, _40756_);
  or (_40775_, _40774_, _40754_);
  and (_40776_, _40775_, _40597_);
  or (_40777_, _40776_, _40728_);
  and (_00149_, _40777_, _42545_);
  and (_40778_, _40505_, _40294_);
  or (_40779_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40780_, _40779_, _40506_);
  or (_40781_, _40780_, _40522_);
  and (_40782_, _40546_, _40294_);
  or (_40783_, _40757_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40784_, _40783_, _40762_);
  or (_40785_, _40784_, _40717_);
  or (_40786_, _40785_, _40782_);
  and (_40787_, _40786_, _40781_);
  or (_40788_, _40787_, _40778_);
  and (_40789_, _40788_, _40607_);
  or (_40790_, _40733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40791_, _40790_, _40738_);
  and (_40792_, _40409_, _40294_);
  or (_40793_, _40792_, _40791_);
  and (_40794_, _40793_, _40434_);
  not (_40795_, _40434_);
  and (_40796_, _40779_, _40795_);
  or (_40797_, _40796_, _40420_);
  or (_40798_, _40797_, _40794_);
  or (_40799_, _40421_, _40294_);
  and (_40800_, _40799_, _40477_);
  and (_40801_, _40800_, _40798_);
  and (_40802_, _40562_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40803_, _40802_, _40481_);
  or (_40804_, _40803_, _40801_);
  or (_40805_, _40804_, _40789_);
  or (_40806_, _40597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40807_, _40806_, _42545_);
  and (_00151_, _40807_, _40805_);
  or (_40808_, _40560_, _40555_);
  and (_40809_, _40808_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_40810_, _40809_, _40578_);
  and (_00152_, _40810_, _42545_);
  and (_40811_, _40556_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_40812_, _40811_, _40483_);
  and (_00154_, _40812_, _42545_);
  and (_40813_, _40250_, _27595_);
  or (_40814_, _40813_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_40815_, _40814_, _40273_);
  nand (_40816_, _40813_, _31732_);
  and (_40817_, _40816_, _40815_);
  and (_40818_, _40244_, _38124_);
  or (_40819_, _40818_, _40817_);
  and (_00156_, _40819_, _42545_);
  not (_40820_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand (_40821_, _40250_, _33713_);
  nand (_40822_, _40821_, _40820_);
  and (_40823_, _40822_, _40273_);
  or (_40824_, _40821_, _32352_);
  and (_40825_, _40824_, _40823_);
  nor (_40826_, _40273_, _38108_);
  or (_40827_, _40826_, _40825_);
  and (_00158_, _40827_, _42545_);
  nand (_40828_, _40250_, _35226_);
  nand (_40829_, _40828_, _39659_);
  and (_40830_, _40829_, _40273_);
  or (_40831_, _40828_, _32352_);
  and (_40832_, _40831_, _40830_);
  nor (_40833_, _40273_, _38092_);
  or (_40834_, _40833_, _40832_);
  and (_00160_, _40834_, _42545_);
  and (_40835_, _40229_, _27595_);
  or (_40836_, _40835_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40837_, _40836_, _40226_);
  nand (_40838_, _40835_, _31732_);
  and (_40839_, _40838_, _40837_);
  and (_40840_, _40225_, _38124_);
  or (_40841_, _40840_, _40839_);
  and (_00162_, _40841_, _42545_);
  and (_40842_, _40229_, _33016_);
  or (_40843_, _40842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40844_, _40843_, _40226_);
  nand (_40845_, _40842_, _31732_);
  and (_40846_, _40845_, _40844_);
  nor (_40847_, _40226_, _38115_);
  or (_40848_, _40847_, _40846_);
  and (_00163_, _40848_, _42545_);
  nand (_40849_, _40229_, _39147_);
  and (_40850_, _40849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40851_, _40850_, _40225_);
  and (_40852_, _33746_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40853_, _40852_, _33735_);
  and (_40854_, _40853_, _40229_);
  or (_40855_, _40854_, _40851_);
  nand (_40856_, _40225_, _38108_);
  and (_40857_, _40856_, _42545_);
  and (_00165_, _40857_, _40855_);
  and (_40858_, _40229_, _34431_);
  or (_40859_, _40858_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40860_, _40859_, _40226_);
  nand (_40861_, _40858_, _31732_);
  and (_40862_, _40861_, _40860_);
  nor (_40863_, _40226_, _38100_);
  or (_40864_, _40863_, _40862_);
  and (_00167_, _40864_, _42545_);
  and (_40865_, _40229_, _35226_);
  or (_40866_, _40865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_40867_, _40866_, _40226_);
  nand (_40868_, _40865_, _31732_);
  and (_40869_, _40868_, _40867_);
  nor (_40870_, _40226_, _38092_);
  or (_40871_, _40870_, _40869_);
  and (_00169_, _40871_, _42545_);
  and (_40872_, _40229_, _36043_);
  or (_40873_, _40872_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_40874_, _40873_, _40226_);
  nand (_40875_, _40872_, _31732_);
  and (_40876_, _40875_, _40874_);
  nor (_40877_, _40226_, _38085_);
  or (_40878_, _40877_, _40876_);
  and (_00171_, _40878_, _42545_);
  and (_40879_, _40229_, _36782_);
  or (_40880_, _40879_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_40881_, _40880_, _40226_);
  nand (_40882_, _40879_, _31732_);
  and (_40883_, _40882_, _40881_);
  nor (_40884_, _40226_, _38078_);
  or (_40885_, _40884_, _40883_);
  and (_00173_, _40885_, _42545_);
  and (_40886_, _40216_, _27595_);
  nand (_40887_, _40886_, _31732_);
  or (_40888_, _40886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40889_, _40888_, _40887_);
  or (_40890_, _40889_, _40211_);
  nand (_40891_, _40211_, _38123_);
  and (_40892_, _40891_, _42545_);
  and (_00174_, _40892_, _40890_);
  and (_40893_, _40216_, _33016_);
  nand (_40894_, _40893_, _31732_);
  not (_40895_, _40211_);
  or (_40896_, _40893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40897_, _40896_, _40895_);
  and (_40898_, _40897_, _40894_);
  nor (_40899_, _40895_, _38115_);
  or (_40900_, _40899_, _40898_);
  and (_00176_, _40900_, _42545_);
  and (_40901_, _33746_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40902_, _40901_, _33735_);
  and (_40903_, _40902_, _40216_);
  nand (_40904_, _40216_, _39147_);
  and (_40905_, _40904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40906_, _40905_, _40211_);
  or (_40907_, _40906_, _40903_);
  nand (_40908_, _40211_, _38108_);
  and (_40909_, _40908_, _42545_);
  and (_00178_, _40909_, _40907_);
  and (_40910_, _40216_, _34431_);
  nand (_40911_, _40910_, _31732_);
  or (_40912_, _40910_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40913_, _40912_, _40895_);
  and (_40914_, _40913_, _40911_);
  nor (_40915_, _40895_, _38100_);
  or (_40916_, _40915_, _40914_);
  and (_00180_, _40916_, _42545_);
  and (_40917_, _40216_, _35226_);
  nand (_40918_, _40917_, _31732_);
  or (_40919_, _40917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40920_, _40919_, _40895_);
  and (_40921_, _40920_, _40918_);
  nor (_40922_, _40895_, _38092_);
  or (_40923_, _40922_, _40921_);
  and (_00182_, _40923_, _42545_);
  and (_40924_, _40216_, _36043_);
  nand (_40925_, _40924_, _31732_);
  or (_40926_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40927_, _40926_, _40925_);
  or (_40928_, _40927_, _40211_);
  nand (_40929_, _40211_, _38085_);
  and (_40930_, _40929_, _42545_);
  and (_00184_, _40930_, _40928_);
  and (_40931_, _40216_, _36782_);
  nand (_40932_, _40931_, _31732_);
  or (_40933_, _40931_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_40934_, _40933_, _40895_);
  and (_40935_, _40934_, _40932_);
  nor (_40936_, _40895_, _38078_);
  or (_40937_, _40936_, _40935_);
  and (_00185_, _40937_, _42545_);
  and (_40938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_40939_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_40940_, _40275_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_40941_, _40940_, _40939_);
  not (_40942_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_40943_, _40942_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_40944_, _40943_, _40941_);
  nor (_40945_, _40944_, _40938_);
  or (_40946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_40947_, _40946_, _42545_);
  nor (_00546_, _40947_, _40945_);
  nor (_40948_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_40949_, _40948_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_40950_, _40948_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_40951_, _40950_, _42545_);
  and (_00548_, _40951_, _40949_);
  not (_40952_, rxd_i);
  and (_40953_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _40952_);
  nor (_40954_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_40955_, _40954_);
  and (_40956_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_40957_, _40956_, _40955_);
  and (_40958_, _40957_, _40953_);
  not (_40959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_40960_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _40959_);
  and (_40961_, _40960_, _40954_);
  or (_40962_, _40961_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or (_40963_, _40962_, _40958_);
  and (_40964_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _42545_);
  and (_00551_, _40964_, _40963_);
  and (_40965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_40966_, _40965_, _40955_);
  not (_40967_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_40968_, _40954_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_40969_, _40968_, _40967_);
  nor (_40970_, _40969_, _40966_);
  not (_40971_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_40972_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _40971_);
  not (_40973_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_40974_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _40973_);
  and (_40975_, _40974_, _40972_);
  not (_40976_, _40975_);
  or (_40977_, _40976_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and (_40978_, _40975_, _40966_);
  and (_40979_, _40966_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_40980_, _40979_, _40978_);
  and (_40981_, _40980_, _40977_);
  or (_40982_, _40981_, _40970_);
  not (_40983_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand (_40984_, _40954_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_40985_, _40984_, _40983_);
  not (_40986_, _40985_);
  or (_40987_, _40986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_40988_, _40987_, _40982_);
  nand (_00554_, _40988_, _40964_);
  not (_40989_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_40990_, _40966_);
  nor (_40991_, _40967_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_40992_, _40991_);
  not (_40993_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_40994_, _40954_, _40993_);
  and (_40995_, _40994_, _40992_);
  and (_40996_, _40995_, _40990_);
  nor (_40997_, _40996_, _40989_);
  and (_40998_, _40996_, rxd_i);
  or (_40999_, _40998_, rst);
  or (_00556_, _40999_, _40997_);
  nor (_41000_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41001_, _41000_, _40972_);
  and (_41002_, _41001_, _40979_);
  nand (_41003_, _41002_, _40952_);
  or (_41004_, _41002_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_41005_, _41004_, _42545_);
  and (_00559_, _41005_, _41003_);
  and (_41006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41007_, _41006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41008_, _41007_, _40971_);
  and (_41009_, _41008_, _40979_);
  and (_41010_, _40957_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41011_, _41010_, _40979_);
  nor (_41012_, _41007_, _40990_);
  or (_41013_, _41012_, _41011_);
  and (_41014_, _41013_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_41015_, _41014_, _41009_);
  and (_00562_, _41015_, _42545_);
  and (_41016_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _42545_);
  nand (_41017_, _41016_, _40993_);
  nand (_41018_, _40964_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_00564_, _41018_, _41017_);
  and (_41019_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _40993_);
  not (_41020_, _40957_);
  nand (_41021_, _40961_, _40983_);
  and (_41022_, _41021_, _41020_);
  and (_41023_, _41022_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_41024_, _41023_, _40966_);
  or (_41025_, _40975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_41026_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41027_, _41026_, _40978_);
  and (_41028_, _41027_, _41025_);
  and (_41029_, _41028_, _41024_);
  or (_41030_, _41029_, _40985_);
  nand (_41031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41032_, _41031_, _40966_);
  or (_41033_, _41032_, _40976_);
  and (_41034_, _41033_, _40986_);
  or (_41035_, _41034_, rxd_i);
  and (_41036_, _41035_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41037_, _41036_, _41030_);
  or (_41038_, _41037_, _41019_);
  and (_00567_, _41038_, _42545_);
  and (_41039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_41041_, _40940_, _41040_);
  or (_41042_, _41041_, _40943_);
  nor (_41043_, _41042_, _41039_);
  or (_41044_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41045_, _41044_, _42545_);
  nor (_00570_, _41045_, _41043_);
  nor (_41046_, _41043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41047_, _41046_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41048_, _41046_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_41049_, _41048_, _42545_);
  and (_00572_, _41049_, _41047_);
  not (_41050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  nor (_41051_, _31733_, _28242_);
  and (_41052_, _41051_, _33005_);
  and (_41053_, _41052_, _31187_);
  and (_41054_, _41053_, _39075_);
  and (_41055_, _41054_, _42545_);
  nand (_41056_, _41055_, _41050_);
  nor (_41057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_41058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_41059_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41060_, _41059_, _41058_);
  and (_41061_, _41060_, _41057_);
  not (_41062_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_41063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_41064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41065_, _41064_, _41063_);
  and (_41066_, _41065_, _41062_);
  and (_41067_, _41066_, _41061_);
  not (_41068_, _41067_);
  or (_41069_, _41068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  or (_41070_, _41067_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not (_41071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_41072_, _40984_, _41071_);
  and (_41073_, _41072_, _41070_);
  and (_41074_, _41073_, _41069_);
  nor (_41075_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41076_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41077_, _41076_, _41075_);
  and (_41078_, _40955_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_41079_, _41078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41080_, _41079_, _41077_);
  not (_41081_, _41080_);
  or (_41082_, _41081_, _41070_);
  and (_41083_, _41077_, _41078_);
  or (_41084_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _41071_);
  nor (_41085_, _41084_, _41083_);
  nor (_41086_, _41085_, _41072_);
  and (_41087_, _41086_, _41082_);
  nor (_41088_, _41087_, _41074_);
  nor (_41089_, _41054_, rst);
  nand (_41090_, _41089_, _41088_);
  and (_00575_, _41090_, _41056_);
  nor (_41091_, _41068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_41092_, _41083_, _41091_);
  and (_41093_, _41072_, _41067_);
  or (_41094_, _41071_, rst);
  nor (_41095_, _41094_, _41093_);
  and (_41096_, _41095_, _41092_);
  or (_00578_, _41096_, _41055_);
  or (_41097_, _41081_, _41091_);
  or (_41098_, _41083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41099_, _40984_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41100_, _41099_, _41098_);
  and (_41101_, _41100_, _41097_);
  or (_41102_, _41101_, _41093_);
  and (_00580_, _41102_, _41089_);
  and (_41103_, _41079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_41104_, _41103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_41105_, _41104_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nand (_41106_, _41105_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or (_41107_, _41105_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41108_, _41107_, _41106_);
  and (_00583_, _41108_, _41089_);
  nor (_41109_, _41080_, _41072_);
  and (_41110_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41111_, _41110_, _41089_);
  and (_41112_, _41055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_00586_, _41112_, _41111_);
  and (_41113_, _40210_, _38059_);
  or (_41114_, _41113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_41115_, _41114_, _42545_);
  nand (_41116_, _41113_, _38146_);
  and (_00588_, _41116_, _41115_);
  and (_41117_, _40215_, _39053_);
  and (_41118_, _41117_, _31755_);
  nand (_41119_, _41118_, _31732_);
  and (_41120_, _40224_, _39075_);
  not (_41121_, _41120_);
  or (_41122_, _41118_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_41123_, _41122_, _41121_);
  and (_41124_, _41123_, _41119_);
  nor (_41125_, _41121_, _38146_);
  or (_41126_, _41125_, _41124_);
  and (_00591_, _41126_, _42545_);
  nor (_41127_, _40985_, _40978_);
  not (_41128_, _41127_);
  nor (_41129_, _41022_, _40966_);
  nor (_41130_, _41129_, _41128_);
  nor (_41131_, _41130_, _40993_);
  or (_41132_, _41131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_41133_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _40993_);
  or (_41134_, _41133_, _41127_);
  and (_41135_, _41134_, _42545_);
  and (_01207_, _41135_, _41132_);
  or (_41136_, _41131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_41137_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _40993_);
  or (_41138_, _41137_, _41127_);
  and (_41139_, _41138_, _42545_);
  and (_01208_, _41139_, _41136_);
  or (_41140_, _41131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_41141_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _40993_);
  or (_41142_, _41141_, _41127_);
  and (_41143_, _41142_, _42545_);
  and (_01209_, _41143_, _41140_);
  or (_41144_, _41131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_41145_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _40993_);
  or (_41146_, _41145_, _41127_);
  and (_41147_, _41146_, _42545_);
  and (_01210_, _41147_, _41144_);
  or (_41148_, _41131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_41149_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _40993_);
  or (_41150_, _41149_, _41127_);
  and (_41151_, _41150_, _42545_);
  and (_01211_, _41151_, _41148_);
  or (_41152_, _41131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_41153_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _40993_);
  or (_41154_, _41153_, _41127_);
  and (_41155_, _41154_, _42545_);
  and (_01213_, _41155_, _41152_);
  or (_41156_, _41131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_41157_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _40993_);
  or (_41158_, _41157_, _41127_);
  and (_41159_, _41158_, _42545_);
  and (_01215_, _41159_, _41156_);
  or (_41160_, _41131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_41161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _40993_);
  or (_41162_, _41161_, _41127_);
  and (_41163_, _41162_, _42545_);
  and (_01217_, _41163_, _41160_);
  nor (_41164_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_41165_, _41164_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_41166_, _40976_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_41167_, _40975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41168_, _41167_, _40966_);
  and (_41169_, _41168_, _41166_);
  or (_41170_, _40957_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41171_, _41170_, _41021_);
  and (_41172_, _41171_, _40990_);
  or (_41173_, _41172_, _41169_);
  or (_41174_, _41173_, _40985_);
  or (_41175_, _40986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41176_, _41175_, _40964_);
  and (_41177_, _41176_, _41174_);
  or (_01219_, _41177_, _41165_);
  and (_41178_, _40975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_41179_, _41178_, _41022_);
  or (_41180_, _41179_, _41130_);
  and (_41181_, _41180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41182_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _40993_);
  nand (_41183_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41184_, _41183_, _41127_);
  or (_41185_, _41184_, _41182_);
  or (_41186_, _41185_, _41181_);
  and (_01221_, _41186_, _42545_);
  not (_41187_, _41131_);
  and (_41188_, _41187_, _41016_);
  or (_41189_, _41179_, _41128_);
  and (_41190_, _40964_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_41191_, _41190_, _41189_);
  or (_01223_, _41191_, _41188_);
  or (_41192_, _41009_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_41193_, _41009_, _40952_);
  and (_41194_, _41193_, _42545_);
  and (_01225_, _41194_, _41192_);
  or (_41195_, _41011_, _40973_);
  or (_41196_, _40979_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41197_, _41196_, _42545_);
  and (_01227_, _41197_, _41195_);
  and (_41198_, _41011_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_41199_, _41000_, _41006_);
  and (_41200_, _41199_, _40979_);
  or (_41201_, _41200_, _41198_);
  and (_01229_, _41201_, _42545_);
  and (_41202_, _41013_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41203_, _41006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41204_, _41203_, _41012_);
  or (_41205_, _41204_, _41202_);
  and (_01231_, _41205_, _42545_);
  and (_41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _40993_);
  and (_41207_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41208_, _41207_, _41206_);
  and (_01233_, _41208_, _42545_);
  and (_41209_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _40993_);
  and (_41210_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41211_, _41210_, _41209_);
  and (_01235_, _41211_, _42545_);
  and (_41212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _40993_);
  and (_41213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41214_, _41213_, _41212_);
  and (_01237_, _41214_, _42545_);
  and (_41215_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _40993_);
  and (_41216_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41217_, _41216_, _41215_);
  and (_01239_, _41217_, _42545_);
  and (_41218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _40993_);
  and (_41219_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41220_, _41219_, _41218_);
  and (_01241_, _41220_, _42545_);
  and (_41221_, _40964_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01243_, _41221_, _41165_);
  and (_41222_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41223_, _41222_, _41182_);
  and (_01245_, _41223_, _42545_);
  nor (_41224_, _41079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41225_, _41224_, _41103_);
  and (_01246_, _41225_, _41089_);
  nor (_41226_, _41103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_41227_, _41226_, _41104_);
  and (_01248_, _41227_, _41089_);
  nor (_41228_, _41104_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_41229_, _41228_, _41105_);
  and (_01250_, _41229_, _41089_);
  and (_41230_, _41067_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41231_, _41230_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41232_, _41231_, _41072_);
  or (_41233_, _41080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41234_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41235_, _41234_, _41233_);
  nor (_41236_, _41235_, _41232_);
  nor (_41237_, _41236_, _41054_);
  nor (_41238_, _40955_, _38123_);
  and (_41239_, _41238_, _41054_);
  or (_41240_, _41239_, _41237_);
  and (_01252_, _41240_, _42545_);
  not (_41241_, _41109_);
  and (_41242_, _41241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_41243_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_41244_, _41243_, _41242_);
  and (_41245_, _41244_, _41089_);
  nand (_41246_, _40954_, _38115_);
  nand (_41248_, _40955_, _38123_);
  and (_41250_, _41248_, _41055_);
  and (_41252_, _41250_, _41246_);
  or (_01254_, _41252_, _41245_);
  nor (_41255_, _41109_, _41062_);
  and (_41257_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_41259_, _41257_, _41255_);
  and (_41261_, _41259_, _41089_);
  nand (_41263_, _40954_, _38108_);
  nand (_41265_, _40955_, _38115_);
  and (_41267_, _41265_, _41055_);
  and (_41269_, _41267_, _41263_);
  or (_01256_, _41269_, _41261_);
  nand (_41272_, _41109_, _41062_);
  or (_41274_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_41276_, _41274_, _41272_);
  and (_41278_, _41276_, _41089_);
  nand (_41280_, _40955_, _38108_);
  nand (_41282_, _40954_, _38100_);
  and (_41284_, _41282_, _41055_);
  and (_41286_, _41284_, _41280_);
  or (_01258_, _41286_, _41278_);
  nand (_41289_, _41109_, _41058_);
  or (_41291_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41293_, _41291_, _41289_);
  and (_41295_, _41293_, _41089_);
  nand (_41297_, _40955_, _38100_);
  nand (_41299_, _40954_, _38092_);
  and (_41301_, _41299_, _41055_);
  and (_41303_, _41301_, _41297_);
  or (_01260_, _41303_, _41295_);
  or (_41306_, _41241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_41308_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_41310_, _41308_, _41306_);
  and (_41312_, _41310_, _41089_);
  nand (_41313_, _40954_, _38085_);
  nand (_41314_, _40955_, _38092_);
  and (_41315_, _41314_, _41055_);
  and (_41316_, _41315_, _41313_);
  or (_01262_, _41316_, _41312_);
  or (_41317_, _41241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or (_41318_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41319_, _41318_, _41317_);
  and (_41320_, _41319_, _41089_);
  nand (_41321_, _40954_, _38078_);
  nand (_41322_, _40955_, _38085_);
  and (_41323_, _41322_, _41055_);
  and (_41324_, _41323_, _41321_);
  or (_01264_, _41324_, _41320_);
  or (_41325_, _41241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_41326_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41327_, _41326_, _41325_);
  and (_41328_, _41327_, _41089_);
  nand (_41329_, _40954_, _38146_);
  nand (_41330_, _40955_, _38078_);
  and (_41331_, _41330_, _41055_);
  and (_41332_, _41331_, _41329_);
  or (_01266_, _41332_, _41328_);
  and (_41333_, _41054_, _40955_);
  nand (_41334_, _41333_, _38146_);
  and (_41335_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41336_, _41241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41337_, _41336_, _41335_);
  or (_41338_, _41337_, _41054_);
  and (_41339_, _41338_, _42545_);
  and (_01268_, _41339_, _41334_);
  or (_41340_, _41241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41341_, _41109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41342_, _41341_, _41340_);
  and (_41343_, _41342_, _41089_);
  or (_41344_, _40942_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41345_, _41344_, _40955_);
  and (_41346_, _41345_, _41055_);
  or (_01270_, _41346_, _41343_);
  nand (_41347_, _41113_, _38123_);
  or (_41348_, _41113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_41349_, _41348_, _42545_);
  and (_01272_, _41349_, _41347_);
  or (_41350_, _41113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_41351_, _41350_, _42545_);
  nand (_41352_, _41113_, _38115_);
  and (_01274_, _41352_, _41351_);
  or (_41353_, _41113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_41354_, _41353_, _42545_);
  nand (_41355_, _41113_, _38108_);
  and (_01276_, _41355_, _41354_);
  or (_41356_, _41113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_41357_, _41356_, _42545_);
  nand (_41358_, _41113_, _38100_);
  and (_01278_, _41358_, _41357_);
  or (_41359_, _41113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_41360_, _41359_, _42545_);
  nand (_41361_, _41113_, _38092_);
  and (_01280_, _41361_, _41360_);
  or (_41362_, _41113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_41363_, _41362_, _42545_);
  nand (_41364_, _41113_, _38085_);
  and (_01281_, _41364_, _41363_);
  or (_41365_, _41113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_41366_, _41365_, _42545_);
  nand (_41367_, _41113_, _38078_);
  and (_01283_, _41367_, _41366_);
  not (_41368_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_41369_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41368_);
  or (_41370_, _41369_, _40954_);
  nor (_41371_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41372_, _41371_, _41370_);
  or (_41373_, _41372_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_41374_, _41373_, _41117_);
  or (_41375_, _27595_, _40959_);
  nand (_41376_, _41375_, _41117_);
  or (_41377_, _41376_, _38767_);
  and (_41378_, _41377_, _41374_);
  or (_41379_, _41378_, _41120_);
  nand (_41380_, _41120_, _38123_);
  and (_41381_, _41380_, _42545_);
  and (_01285_, _41381_, _41379_);
  or (_41382_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_41383_, _41382_, _41117_);
  nand (_41384_, _38893_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_41385_, _41384_, _41117_);
  or (_41386_, _41385_, _38904_);
  and (_41387_, _41386_, _41383_);
  or (_41388_, _41387_, _41120_);
  nand (_41389_, _41120_, _38115_);
  and (_41390_, _41389_, _42545_);
  and (_01287_, _41390_, _41388_);
  not (_41391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41392_, _40968_, _41391_);
  and (_41393_, _41392_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_41394_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_41395_, _41392_, _41394_);
  or (_41396_, _41395_, _41393_);
  or (_41397_, _41396_, _41117_);
  or (_41398_, _33713_, _41394_);
  nand (_41399_, _41398_, _41117_);
  or (_41400_, _41399_, _33735_);
  and (_41401_, _41400_, _41397_);
  or (_41402_, _41401_, _41120_);
  nand (_41403_, _41120_, _38108_);
  and (_41404_, _41403_, _42545_);
  and (_01289_, _41404_, _41402_);
  and (_41405_, _41117_, _34431_);
  nand (_41406_, _41405_, _31732_);
  or (_41407_, _41405_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41408_, _41407_, _41121_);
  and (_41409_, _41408_, _41406_);
  nor (_41410_, _41121_, _38100_);
  or (_41411_, _41410_, _41409_);
  and (_01291_, _41411_, _42545_);
  and (_41412_, _41117_, _35226_);
  nand (_41413_, _41412_, _31732_);
  or (_41414_, _41412_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_41415_, _41414_, _41121_);
  and (_41416_, _41415_, _41413_);
  nor (_41417_, _41121_, _38092_);
  or (_41418_, _41417_, _41416_);
  and (_01293_, _41418_, _42545_);
  and (_41419_, _41117_, _36043_);
  nand (_41420_, _41419_, _31732_);
  or (_41421_, _41419_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_41422_, _41421_, _41121_);
  and (_41423_, _41422_, _41420_);
  nor (_41424_, _41121_, _38085_);
  or (_41425_, _41424_, _41423_);
  and (_01295_, _41425_, _42545_);
  and (_41426_, _41117_, _36782_);
  nand (_41427_, _41426_, _31732_);
  or (_41428_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_41429_, _41428_, _41427_);
  or (_41430_, _41429_, _41120_);
  nand (_41431_, _41120_, _38078_);
  and (_41432_, _41431_, _42545_);
  and (_01297_, _41432_, _41430_);
  and (_01622_, t2_i, _42545_);
  nor (_41433_, t2_i, rst);
  and (_01625_, _41433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand (_41434_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _42545_);
  nor (_01628_, _41434_, t2ex_i);
  and (_01631_, t2ex_i, _42545_);
  not (_41435_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_41436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_41437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_41438_, _41437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41439_, _41438_, _41436_);
  nor (_41440_, _41439_, _41435_);
  and (_41441_, _41439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_41442_, _41441_, _41440_);
  and (_41443_, _38056_, _38633_);
  and (_41444_, _41443_, _39695_);
  nor (_41445_, _41444_, _41442_);
  and (_41446_, _27573_, _32994_);
  and (_41447_, _41051_, _41446_);
  and (_41448_, _41443_, _41447_);
  and (_41449_, _41448_, _31187_);
  not (_41450_, _41449_);
  nor (_41451_, _41450_, _38146_);
  or (_41452_, _41451_, _41445_);
  and (_41453_, _41443_, _39549_);
  not (_41454_, _41453_);
  and (_41455_, _41454_, _41452_);
  and (_41456_, _41453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_41457_, _41456_, _41455_);
  and (_01634_, _41457_, _42545_);
  nand (_41458_, _41453_, _38146_);
  not (_41459_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_41460_, _41439_);
  nor (_41461_, _41444_, _41460_);
  nor (_41462_, _41461_, _41459_);
  and (_41463_, _41461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_41464_, _41463_, _41462_);
  or (_41465_, _41464_, _41453_);
  and (_41466_, _41465_, _42545_);
  and (_01637_, _41466_, _41458_);
  and (_41467_, _41443_, _39651_);
  and (_41468_, _39548_, _36043_);
  and (_41469_, _41468_, _41443_);
  nor (_41470_, _41469_, _41467_);
  not (_41471_, _41437_);
  or (_41472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_41473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_41474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _41473_);
  and (_41475_, _41474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_41476_, _41475_, _41472_);
  and (_41477_, _41476_, _41471_);
  and (_41478_, _41477_, _41470_);
  or (_41479_, _41478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_41480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41481_, _41480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_41482_, _41481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_41483_, _41482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_41484_, _41483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_41485_, _41484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_41486_, _41485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_41487_, _41486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_41488_, _41487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_41489_, _41488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_41490_, _41489_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_41491_, _41490_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_41492_, _41491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_41493_, _41492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_41494_, _41493_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_41495_, _41494_);
  nand (_41496_, _41495_, _41478_);
  and (_41497_, _41496_, _42545_);
  and (_01640_, _41497_, _41479_);
  nand (_41498_, _41467_, _38146_);
  and (_41499_, _41443_, _36043_);
  and (_41500_, _41499_, _39548_);
  not (_41501_, _41500_);
  not (_41502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41503_, _41436_, _41502_);
  and (_41504_, _41503_, _41437_);
  and (_41505_, _41504_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not (_41506_, _41504_);
  nor (_41507_, _41438_, _41435_);
  and (_41508_, _41494_, _41476_);
  and (_41509_, _41508_, _41507_);
  and (_41510_, _41485_, _41476_);
  or (_41511_, _41510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_41512_, _41510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_41513_, _41512_, _41511_);
  or (_41514_, _41513_, _41509_);
  and (_41515_, _41514_, _41506_);
  or (_41516_, _41515_, _41505_);
  or (_41517_, _41516_, _41467_);
  and (_41518_, _41517_, _41501_);
  and (_41519_, _41518_, _41498_);
  and (_41520_, _41500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_41521_, _41520_, _41519_);
  and (_01643_, _41521_, _42545_);
  and (_41522_, _41493_, _41476_);
  or (_41523_, _41522_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_41524_, _41438_, _41459_);
  nand (_41525_, _41524_, _41508_);
  and (_41526_, _41525_, _41523_);
  or (_41527_, _41526_, _41504_);
  nand (_41528_, _41504_, _41459_);
  and (_41529_, _41528_, _41470_);
  and (_41530_, _41529_, _41527_);
  and (_41531_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_41532_, _41531_, _41530_);
  not (_41533_, _38146_);
  and (_41534_, _41469_, _41533_);
  or (_41535_, _41534_, _41532_);
  and (_01646_, _41535_, _42545_);
  and (_41536_, _41506_, _41476_);
  and (_41537_, _41536_, _41437_);
  nand (_41538_, _41537_, _41494_);
  nand (_41539_, _41538_, _41470_);
  or (_41540_, _41470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41541_, _41540_, _42545_);
  and (_01649_, _41541_, _41539_);
  or (_41542_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41543_, _40228_, _38618_);
  or (_41544_, _41543_, _41542_);
  not (_41545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_41546_, _31755_, _41545_);
  nand (_41547_, _41546_, _41543_);
  or (_41548_, _41547_, _38621_);
  and (_41549_, _41548_, _41544_);
  and (_41550_, _41443_, _40224_);
  or (_41551_, _41550_, _41549_);
  nand (_41552_, _41550_, _38146_);
  and (_41553_, _41552_, _42545_);
  and (_01652_, _41553_, _41551_);
  or (_41554_, _41439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not (_41555_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_41556_, _41439_, _41555_);
  and (_41557_, _41556_, _41554_);
  or (_41558_, _41557_, _41444_);
  nand (_41559_, _41444_, _38123_);
  and (_41560_, _41559_, _41558_);
  or (_41561_, _41560_, _41453_);
  not (_41562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_41563_, _41453_, _41562_);
  and (_41564_, _41563_, _42545_);
  and (_02115_, _41564_, _41561_);
  nand (_41565_, _41444_, _38115_);
  and (_41566_, _41460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41567_, _41439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_41568_, _41567_, _41566_);
  or (_41569_, _41568_, _41444_);
  and (_41570_, _41569_, _41565_);
  or (_41571_, _41570_, _41453_);
  or (_41572_, _41454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41573_, _41572_, _42545_);
  and (_02117_, _41573_, _41571_);
  nand (_41574_, _41444_, _38108_);
  and (_41575_, _41460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41576_, _41439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_41577_, _41576_, _41575_);
  or (_41578_, _41577_, _41444_);
  and (_41579_, _41578_, _41574_);
  or (_41580_, _41579_, _41453_);
  or (_41581_, _41454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41582_, _41581_, _42545_);
  and (_02118_, _41582_, _41580_);
  nand (_41583_, _41444_, _38100_);
  and (_41584_, _41460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41585_, _41439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_41586_, _41585_, _41584_);
  or (_41587_, _41586_, _41444_);
  and (_41588_, _41587_, _41583_);
  or (_41589_, _41588_, _41453_);
  or (_41590_, _41454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41591_, _41590_, _42545_);
  and (_02120_, _41591_, _41589_);
  nand (_41592_, _41444_, _38092_);
  and (_41593_, _41460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_41594_, _41439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_41595_, _41594_, _41593_);
  or (_41596_, _41595_, _41444_);
  and (_41597_, _41596_, _41592_);
  or (_41598_, _41597_, _41453_);
  or (_41599_, _41454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_41600_, _41599_, _42545_);
  and (_02122_, _41600_, _41598_);
  and (_41601_, _41460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41602_, _41439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_41603_, _41602_, _41601_);
  nor (_41604_, _41603_, _41444_);
  nor (_41605_, _41450_, _38085_);
  or (_41606_, _41605_, _41604_);
  and (_41607_, _41606_, _41454_);
  and (_41608_, _41453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_41609_, _41608_, _41607_);
  and (_02124_, _41609_, _42545_);
  and (_41610_, _41460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_41611_, _41439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_41612_, _41611_, _41610_);
  nor (_41613_, _41612_, _41444_);
  nor (_41614_, _41450_, _38078_);
  or (_41615_, _41614_, _41613_);
  and (_41616_, _41615_, _41454_);
  and (_41617_, _41453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_41618_, _41617_, _41616_);
  and (_02125_, _41618_, _42545_);
  or (_41619_, _41461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_41620_, _41461_);
  or (_41621_, _41620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_41622_, _41621_, _41619_);
  or (_41623_, _41622_, _41453_);
  nand (_41624_, _41453_, _38123_);
  and (_41625_, _41624_, _42545_);
  and (_02127_, _41625_, _41623_);
  or (_41626_, _41461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  not (_41627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_41628_, _41461_, _41627_);
  and (_41629_, _41628_, _41626_);
  or (_41630_, _41629_, _41453_);
  nand (_41631_, _41453_, _38115_);
  and (_41632_, _41631_, _42545_);
  and (_02129_, _41632_, _41630_);
  nand (_41633_, _41453_, _38108_);
  and (_41634_, _41620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_41635_, _41461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_41636_, _41635_, _41634_);
  or (_41637_, _41636_, _41453_);
  and (_41638_, _41637_, _42545_);
  and (_02131_, _41638_, _41633_);
  nand (_41639_, _41453_, _38100_);
  and (_41640_, _41620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_41641_, _41461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41642_, _41641_, _41640_);
  or (_41643_, _41642_, _41453_);
  and (_41644_, _41643_, _42545_);
  and (_02132_, _41644_, _41639_);
  nand (_41645_, _41453_, _38092_);
  and (_41646_, _41620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_41647_, _41461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41648_, _41647_, _41646_);
  or (_41649_, _41648_, _41453_);
  and (_41650_, _41649_, _42545_);
  and (_02134_, _41650_, _41645_);
  and (_41651_, _41620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_41652_, _41461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41653_, _41652_, _41651_);
  and (_41654_, _41653_, _41454_);
  nor (_41655_, _41454_, _38085_);
  or (_41656_, _41655_, _41654_);
  and (_02136_, _41656_, _42545_);
  nand (_41657_, _41453_, _38078_);
  and (_41658_, _41620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_41659_, _41461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_41660_, _41659_, _41658_);
  or (_41661_, _41660_, _41453_);
  and (_41662_, _41661_, _42545_);
  and (_02138_, _41662_, _41657_);
  or (_41663_, _41476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41664_, _41476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_41665_, _41438_, _41562_);
  nand (_41666_, _41665_, _41494_);
  nand (_41667_, _41666_, _41664_);
  and (_41668_, _41667_, _41663_);
  or (_41669_, _41668_, _41504_);
  and (_41670_, _41504_, _41562_);
  nor (_41671_, _41670_, _41467_);
  and (_41672_, _41671_, _41669_);
  and (_41673_, _41467_, _38124_);
  or (_41674_, _41673_, _41500_);
  or (_41675_, _41674_, _41672_);
  nand (_41676_, _41469_, _41555_);
  and (_41677_, _41676_, _42545_);
  and (_02139_, _41677_, _41675_);
  not (_41678_, _41438_);
  and (_41679_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41680_, _41679_, _41536_);
  and (_41681_, _41680_, _41494_);
  and (_41682_, _41504_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_41683_, _41664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_41684_, _41480_, _41476_);
  and (_41685_, _41684_, _41506_);
  and (_41686_, _41685_, _41683_);
  nor (_41687_, _41686_, _41682_);
  nand (_41688_, _41687_, _41470_);
  or (_41689_, _41688_, _41681_);
  nand (_41690_, _41467_, _38115_);
  or (_41691_, _41501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_41692_, _41691_, _42545_);
  and (_41693_, _41692_, _41690_);
  and (_02141_, _41693_, _41689_);
  and (_41694_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41695_, _41694_, _41508_);
  and (_41696_, _41684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_41697_, _41684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_41698_, _41697_, _41504_);
  or (_41699_, _41698_, _41696_);
  or (_41700_, _41699_, _41695_);
  nor (_41701_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor (_41702_, _41701_, _41467_);
  and (_41703_, _41702_, _41700_);
  not (_41704_, _41467_);
  nor (_41705_, _41704_, _38108_);
  or (_41706_, _41705_, _41703_);
  or (_41707_, _41706_, _41500_);
  or (_41708_, _41501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_41709_, _41708_, _42545_);
  and (_02143_, _41709_, _41707_);
  and (_41710_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41711_, _41710_, _41508_);
  nand (_41712_, _41481_, _41476_);
  and (_41713_, _41712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_41714_, _41712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_41715_, _41714_, _41504_);
  or (_41716_, _41715_, _41713_);
  or (_41717_, _41716_, _41711_);
  nor (_41718_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor (_41719_, _41718_, _41467_);
  and (_41720_, _41719_, _41717_);
  nor (_41721_, _41704_, _38100_);
  or (_41722_, _41721_, _41720_);
  or (_41723_, _41722_, _41500_);
  or (_41724_, _41501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_41725_, _41724_, _42545_);
  and (_02145_, _41725_, _41723_);
  and (_41726_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_41727_, _41726_, _41508_);
  nand (_41728_, _41482_, _41476_);
  and (_41729_, _41728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_41730_, _41728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_41731_, _41730_, _41504_);
  or (_41732_, _41731_, _41729_);
  or (_41733_, _41732_, _41727_);
  nor (_41734_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_41735_, _41734_, _41467_);
  and (_41736_, _41735_, _41733_);
  nor (_41737_, _41704_, _38092_);
  or (_41738_, _41737_, _41736_);
  or (_41739_, _41738_, _41500_);
  or (_41740_, _41501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_41741_, _41740_, _42545_);
  and (_02146_, _41741_, _41739_);
  or (_41742_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41743_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41744_, _41743_, _41508_);
  nand (_41745_, _41483_, _41476_);
  and (_41746_, _41745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_41747_, _41745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_41748_, _41747_, _41504_);
  or (_41749_, _41748_, _41746_);
  or (_41750_, _41749_, _41744_);
  nand (_41751_, _41750_, _41742_);
  nand (_41752_, _41751_, _41704_);
  nand (_41753_, _41467_, _38085_);
  and (_41754_, _41753_, _41752_);
  or (_41755_, _41754_, _41469_);
  or (_41756_, _41501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_41757_, _41756_, _42545_);
  and (_02148_, _41757_, _41755_);
  nor (_41758_, _41704_, _38078_);
  and (_41759_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_41760_, _41759_, _41508_);
  and (_41761_, _41484_, _41476_);
  nor (_41762_, _41761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_41763_, _41762_, _41510_);
  or (_41764_, _41763_, _41504_);
  or (_41765_, _41764_, _41760_);
  nor (_41766_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_41767_, _41766_, _41467_);
  and (_41768_, _41767_, _41765_);
  or (_41769_, _41768_, _41500_);
  or (_41770_, _41769_, _41758_);
  or (_41771_, _41501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_41772_, _41771_, _42545_);
  and (_02150_, _41772_, _41770_);
  not (_41773_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_41774_, _41438_, _41773_);
  and (_41775_, _41774_, _41508_);
  and (_41776_, _41486_, _41476_);
  or (_41777_, _41776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_41778_, _41487_, _41476_);
  and (_41779_, _41778_, _41777_);
  or (_41780_, _41779_, _41504_);
  or (_41781_, _41780_, _41775_);
  and (_41782_, _41504_, _41773_);
  nor (_41783_, _41782_, _41467_);
  and (_41784_, _41783_, _41781_);
  and (_41785_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_41786_, _41785_, _41500_);
  or (_41787_, _41786_, _41784_);
  nand (_41788_, _41469_, _38123_);
  and (_41789_, _41788_, _42545_);
  and (_02152_, _41789_, _41787_);
  and (_41790_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_41791_, _41790_, _41508_);
  nand (_41792_, _41778_, _41627_);
  or (_41793_, _41778_, _41627_);
  and (_41794_, _41793_, _41792_);
  or (_41795_, _41794_, _41504_);
  or (_41796_, _41795_, _41791_);
  nor (_41797_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_41798_, _41797_, _41467_);
  and (_41799_, _41798_, _41796_);
  and (_41800_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_41801_, _41800_, _41500_);
  or (_41802_, _41801_, _41799_);
  nand (_41803_, _41500_, _38115_);
  and (_41804_, _41803_, _42545_);
  and (_02153_, _41804_, _41802_);
  and (_41805_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_41806_, _41805_, _41508_);
  nand (_41807_, _41488_, _41476_);
  and (_41808_, _41807_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_41809_, _41807_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_41810_, _41809_, _41504_);
  or (_41811_, _41810_, _41808_);
  or (_41812_, _41811_, _41806_);
  nor (_41813_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_41814_, _41813_, _41467_);
  and (_41815_, _41814_, _41812_);
  and (_41816_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_41817_, _41816_, _41500_);
  or (_41818_, _41817_, _41815_);
  nand (_41819_, _41500_, _38108_);
  and (_41820_, _41819_, _42545_);
  and (_02155_, _41820_, _41818_);
  and (_41821_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_41822_, _41821_, _41508_);
  nand (_41823_, _41489_, _41476_);
  and (_41824_, _41823_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_41825_, _41823_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41826_, _41825_, _41504_);
  or (_41827_, _41826_, _41824_);
  or (_41828_, _41827_, _41822_);
  nor (_41829_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_41830_, _41829_, _41467_);
  and (_41831_, _41830_, _41828_);
  and (_41832_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41833_, _41832_, _41500_);
  or (_41834_, _41833_, _41831_);
  nand (_41835_, _41500_, _38100_);
  and (_41836_, _41835_, _42545_);
  and (_02157_, _41836_, _41834_);
  and (_41837_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_41838_, _41837_, _41508_);
  nand (_41839_, _41490_, _41476_);
  and (_41840_, _41839_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_41841_, _41839_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41842_, _41841_, _41504_);
  or (_41843_, _41842_, _41840_);
  or (_41844_, _41843_, _41838_);
  nor (_41845_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_41846_, _41845_, _41467_);
  and (_41847_, _41846_, _41844_);
  and (_41848_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41849_, _41848_, _41500_);
  or (_41850_, _41849_, _41847_);
  nand (_41851_, _41500_, _38092_);
  and (_41852_, _41851_, _42545_);
  and (_02159_, _41852_, _41850_);
  and (_41853_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_41854_, _41853_, _41508_);
  nand (_41855_, _41491_, _41476_);
  and (_41856_, _41855_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_41857_, _41855_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41858_, _41857_, _41504_);
  or (_41859_, _41858_, _41856_);
  or (_41860_, _41859_, _41854_);
  nor (_41861_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_41862_, _41861_, _41467_);
  and (_41863_, _41862_, _41860_);
  and (_41864_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41865_, _41864_, _41500_);
  or (_41866_, _41865_, _41863_);
  nand (_41867_, _41500_, _38085_);
  and (_41868_, _41867_, _42545_);
  and (_02160_, _41868_, _41866_);
  and (_41869_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_41870_, _41869_, _41508_);
  and (_41871_, _41492_, _41476_);
  nor (_41872_, _41871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_41873_, _41872_, _41522_);
  or (_41874_, _41873_, _41504_);
  or (_41875_, _41874_, _41870_);
  nor (_41876_, _41506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_41877_, _41876_, _41467_);
  and (_41878_, _41877_, _41875_);
  and (_41879_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_41880_, _41879_, _41500_);
  or (_41881_, _41880_, _41878_);
  nand (_41882_, _41500_, _38078_);
  and (_41883_, _41882_, _42545_);
  and (_02162_, _41883_, _41881_);
  not (_41884_, _41550_);
  and (_41885_, _41543_, _27595_);
  or (_41886_, _41885_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41887_, _41886_, _41884_);
  nand (_41888_, _41885_, _31732_);
  and (_41889_, _41888_, _41887_);
  and (_41890_, _41550_, _38124_);
  or (_41891_, _41890_, _41889_);
  and (_02164_, _41891_, _42545_);
  and (_41892_, _41543_, _33016_);
  or (_41893_, _41892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_41894_, _41893_, _41884_);
  nand (_41895_, _41892_, _31732_);
  and (_41896_, _41895_, _41894_);
  nor (_41897_, _41884_, _38115_);
  or (_41898_, _41897_, _41896_);
  and (_02166_, _41898_, _42545_);
  nand (_41899_, _41543_, _39147_);
  and (_41900_, _41899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_41901_, _41900_, _41550_);
  and (_41902_, _33746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_41903_, _41902_, _33735_);
  and (_41904_, _41903_, _41543_);
  or (_41905_, _41904_, _41901_);
  nand (_41906_, _41550_, _38108_);
  and (_41907_, _41906_, _42545_);
  and (_02167_, _41907_, _41905_);
  and (_41908_, _41543_, _34431_);
  or (_41909_, _41908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_41910_, _41909_, _41884_);
  nand (_41911_, _41908_, _31732_);
  and (_41912_, _41911_, _41910_);
  nor (_41913_, _41884_, _38100_);
  or (_41914_, _41913_, _41912_);
  and (_02169_, _41914_, _42545_);
  and (_41915_, _41543_, _35226_);
  or (_41916_, _41915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_41917_, _41916_, _41884_);
  nand (_41918_, _41915_, _31732_);
  and (_41919_, _41918_, _41917_);
  nor (_41920_, _41884_, _38092_);
  or (_41921_, _41920_, _41919_);
  and (_02171_, _41921_, _42545_);
  and (_41922_, _41543_, _36043_);
  or (_41923_, _41922_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_41924_, _41923_, _41884_);
  nand (_41925_, _41922_, _31732_);
  and (_41926_, _41925_, _41924_);
  nor (_41927_, _41884_, _38085_);
  or (_41928_, _41927_, _41926_);
  and (_02173_, _41928_, _42545_);
  not (_41929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41930_, _41436_, _41929_);
  or (_41931_, _41930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_41932_, _41931_, _41543_);
  nand (_41933_, _38721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_41934_, _41933_, _41543_);
  or (_41935_, _41934_, _38722_);
  and (_41936_, _41935_, _41932_);
  or (_41937_, _41936_, _41550_);
  nand (_41938_, _41550_, _38078_);
  and (_41939_, _41938_, _42545_);
  and (_02174_, _41939_, _41937_);
  and (_41940_, _28088_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41941_, _41940_, _28253_);
  nor (_41942_, _27573_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_41943_, _41942_, _41941_);
  nor (_41944_, _28088_, _27068_);
  nor (_41945_, _41944_, _31165_);
  not (_41946_, _41945_);
  nor (_41947_, _41946_, _41943_);
  and (_41948_, _41940_, _40212_);
  nor (_41949_, _27452_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_41950_, _41949_, _41948_);
  nor (_41951_, _41950_, _41946_);
  and (_41952_, _41951_, _41947_);
  and (_41953_, _41940_, _38057_);
  nor (_41954_, _41940_, _28242_);
  nor (_41955_, _41954_, _41953_);
  nor (_41956_, _41955_, _41946_);
  and (_41957_, _41940_, _38617_);
  nor (_41958_, _27332_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_41959_, _41958_, _41957_);
  nor (_41960_, _41959_, _41946_);
  and (_41961_, _41960_, _41956_);
  and (_41962_, _41961_, _41952_);
  and (_41963_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_41964_, _41963_, _28867_);
  nor (_41965_, _41964_, _31732_);
  nand (_41966_, _28867_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41967_, _20598_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41968_, _41967_, _41966_);
  nor (_41969_, _38146_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_41970_, _41969_, _41968_);
  or (_41971_, _41970_, _41965_);
  and (_41972_, _41971_, _41945_);
  and (_41973_, _41972_, _41962_);
  not (_41974_, _41962_);
  and (_41975_, _41974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_02565_, _41975_, _41973_);
  and (_41976_, _38148_, _38055_);
  not (_41977_, _41976_);
  not (_41978_, _38053_);
  and (_41979_, _41978_, _38018_);
  and (_41980_, _38695_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_41981_, _41980_, _38692_);
  nor (_41982_, _41981_, _28253_);
  and (_41983_, _41981_, _28253_);
  or (_41984_, _41983_, _41982_);
  not (_41985_, _41984_);
  and (_41986_, _37809_, _27573_);
  not (_41987_, _41986_);
  nor (_41988_, _37809_, _27573_);
  not (_41989_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_41990_, _31144_, _41989_);
  not (_41991_, _41990_);
  and (_41992_, _27803_, _28088_);
  and (_41993_, _41992_, _38056_);
  and (_41994_, _41993_, _41052_);
  not (_41995_, _41994_);
  and (_41996_, _41993_, _38737_);
  and (_41997_, _41993_, _39133_);
  nor (_41998_, _41997_, _41996_);
  and (_41999_, _27595_, _28253_);
  and (_42000_, _41993_, _41999_);
  not (_42001_, _42000_);
  and (_42002_, _42001_, _41998_);
  and (_42003_, _42002_, _41995_);
  not (_42004_, _42003_);
  and (_42005_, _41992_, _38632_);
  and (_42006_, _42005_, _41999_);
  and (_42007_, _42005_, _38737_);
  and (_42008_, _42005_, _39133_);
  nor (_42009_, _42008_, _42007_);
  not (_42010_, _42009_);
  or (_42011_, _42010_, _42006_);
  nor (_42012_, _42011_, _42004_);
  nor (_42013_, _42012_, _41991_);
  and (_42014_, _42005_, _41052_);
  and (_42015_, _42014_, _41990_);
  nor (_42016_, _42015_, _42013_);
  nor (_42017_, _42016_, _41988_);
  and (_42018_, _42017_, _41987_);
  and (_42019_, _38698_, _40212_);
  nor (_42020_, _38698_, _40212_);
  nor (_42021_, _42020_, _42019_);
  and (_42022_, _42021_, _42018_);
  and (_42023_, _42022_, _41985_);
  nor (_42024_, _41981_, _37923_);
  and (_42025_, _42024_, _38698_);
  and (_42026_, _42025_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_42027_, _41981_, _37809_);
  and (_42028_, _42027_, _38698_);
  and (_42029_, _42028_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_42030_, _42029_, _42026_);
  not (_42031_, _38698_);
  and (_42032_, _42024_, _42031_);
  and (_42033_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_42034_, _41981_, _37923_);
  and (_42035_, _42034_, _42031_);
  and (_42036_, _42035_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_42037_, _42036_, _42033_);
  and (_42038_, _42037_, _42030_);
  and (_42039_, _42034_, _38698_);
  and (_42040_, _42039_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_42041_, _41981_, _37809_);
  and (_42042_, _42041_, _42031_);
  and (_42043_, _42042_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_42044_, _42043_, _42040_);
  and (_42045_, _42041_, _38698_);
  and (_42046_, _42045_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_42047_, _42027_, _42031_);
  and (_42048_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_42049_, _42048_, _42046_);
  and (_42050_, _42049_, _42044_);
  and (_42051_, _42050_, _42038_);
  nor (_42052_, _42051_, _42023_);
  and (_42053_, _42023_, _41533_);
  nor (_42054_, _42053_, _42052_);
  not (_42055_, _42054_);
  and (_42056_, _42055_, _41979_);
  not (_42057_, _42056_);
  not (_42058_, _37921_);
  nor (_42059_, _41978_, _38018_);
  not (_42060_, _36955_);
  and (_42061_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_42062_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_42063_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_42064_, _42063_, _42062_);
  and (_42065_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_42066_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_42067_, _42066_, _42065_);
  and (_42068_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_42069_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_42070_, _42069_, _42068_);
  and (_42071_, _42070_, _42067_);
  and (_42072_, _42071_, _42064_);
  nor (_42073_, _37120_, _42060_);
  not (_42074_, _42073_);
  nor (_42075_, _42074_, _42072_);
  nor (_42076_, _42075_, _42061_);
  not (_42077_, _42076_);
  and (_42078_, _42077_, _42059_);
  nor (_42079_, _42078_, _42058_);
  and (_42080_, _42079_, _42057_);
  and (_42081_, _42080_, _41977_);
  and (_42082_, _37908_, _37786_);
  nor (_42083_, _42082_, _37987_);
  and (_42084_, _37983_, _37908_);
  nor (_42085_, _42084_, _37946_);
  and (_42086_, _42085_, _38004_);
  and (_42087_, _42086_, _42083_);
  not (_42088_, _37925_);
  and (_42089_, _37986_, _42088_);
  and (_42090_, _42089_, _37962_);
  and (_42091_, _42090_, _42087_);
  nor (_42092_, _42091_, _36912_);
  not (_42093_, _37911_);
  nor (_42094_, _42093_, _37961_);
  nor (_42095_, _42094_, _42092_);
  not (_42096_, _42095_);
  and (_42097_, _42096_, _42081_);
  and (_42098_, _41979_, _37921_);
  and (_42099_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_42100_, _42035_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_42101_, _42100_, _42099_);
  and (_42102_, _42045_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_42103_, _42039_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_42104_, _42103_, _42102_);
  and (_42105_, _42104_, _42101_);
  and (_42106_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_42107_, _42028_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_42108_, _42107_, _42106_);
  and (_42109_, _42042_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_42110_, _42025_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_42111_, _42110_, _42109_);
  and (_42112_, _42111_, _42108_);
  and (_42113_, _42112_, _42105_);
  nor (_42114_, _42113_, _42023_);
  not (_42115_, _38092_);
  and (_42116_, _42023_, _42115_);
  nor (_42117_, _42116_, _42114_);
  not (_42118_, _42117_);
  and (_42119_, _42118_, _42098_);
  not (_42120_, _42119_);
  and (_42121_, _42058_, _38053_);
  not (_42122_, _38180_);
  and (_42123_, _42122_, _38055_);
  nor (_42124_, _42123_, _42121_);
  and (_42125_, _37921_, _38053_);
  and (_42126_, _42125_, _38018_);
  and (_42127_, _42126_, _42031_);
  and (_42128_, _42059_, _37921_);
  and (_42129_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_42130_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42131_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_42132_, _42131_, _42130_);
  and (_42133_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_42134_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_42135_, _42134_, _42133_);
  and (_42136_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_42137_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_42138_, _42137_, _42136_);
  and (_42139_, _42138_, _42135_);
  and (_42140_, _42139_, _42132_);
  nor (_42141_, _42140_, _42074_);
  nor (_42142_, _42141_, _42129_);
  not (_42143_, _42142_);
  and (_42144_, _42143_, _42128_);
  nor (_42145_, _42144_, _42127_);
  and (_42146_, _42145_, _42124_);
  and (_42147_, _42146_, _42120_);
  not (_42148_, _42147_);
  and (_42149_, _42148_, _42097_);
  and (_42150_, _42045_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_42151_, _42039_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_42152_, _42151_, _42150_);
  and (_42153_, _42035_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_42154_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_42155_, _42154_, _42153_);
  and (_42156_, _42155_, _42152_);
  and (_42157_, _42025_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_42158_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_42159_, _42158_, _42157_);
  and (_42160_, _42042_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_42161_, _42028_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_42162_, _42161_, _42160_);
  and (_42163_, _42162_, _42159_);
  and (_42164_, _42163_, _42156_);
  nor (_42165_, _42164_, _42023_);
  not (_42166_, _38115_);
  and (_42167_, _42023_, _42166_);
  nor (_42168_, _42167_, _42165_);
  not (_42169_, _42168_);
  and (_42170_, _42169_, _42098_);
  not (_42171_, _42170_);
  and (_42172_, _41979_, _42058_);
  not (_42173_, _38162_);
  and (_42174_, _42173_, _38055_);
  nor (_42175_, _42174_, _42172_);
  and (_42176_, _42126_, _37833_);
  and (_42177_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_42178_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42179_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_42180_, _42179_, _42178_);
  and (_42181_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_42182_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_42183_, _42182_, _42181_);
  and (_42184_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_42185_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_42186_, _42185_, _42184_);
  and (_42187_, _42186_, _42183_);
  and (_42188_, _42187_, _42180_);
  nor (_42189_, _42188_, _42074_);
  nor (_42190_, _42189_, _42177_);
  not (_42191_, _42190_);
  and (_42192_, _42191_, _42128_);
  nor (_42193_, _42192_, _42176_);
  and (_42194_, _42193_, _42175_);
  and (_42195_, _42194_, _42171_);
  nor (_42196_, _42195_, _42096_);
  nor (_42197_, _42196_, _42149_);
  nand (_42198_, _42197_, _41950_);
  or (_42199_, _42197_, _41950_);
  and (_42200_, _42199_, _42198_);
  not (_42201_, _42200_);
  not (_42202_, _41943_);
  and (_42203_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_42204_, _42039_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_42205_, _42204_, _42203_);
  and (_42206_, _42045_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_42207_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_42208_, _42207_, _42206_);
  and (_42209_, _42208_, _42205_);
  and (_42210_, _42035_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_42211_, _42028_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_42212_, _42211_, _42210_);
  and (_42213_, _42042_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_42214_, _42025_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_42215_, _42214_, _42213_);
  and (_42216_, _42215_, _42212_);
  and (_42217_, _42216_, _42209_);
  nor (_42218_, _42217_, _42023_);
  not (_42219_, _38100_);
  and (_42220_, _42023_, _42219_);
  nor (_42221_, _42220_, _42218_);
  not (_42222_, _42221_);
  and (_42223_, _42222_, _42098_);
  not (_42224_, _42223_);
  and (_42225_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_42226_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_42227_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_42228_, _42227_, _42226_);
  and (_42229_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_42230_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_42231_, _42230_, _42229_);
  and (_42232_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_42233_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_42234_, _42233_, _42232_);
  and (_42235_, _42234_, _42231_);
  and (_42236_, _42235_, _42228_);
  nor (_42237_, _42236_, _42074_);
  nor (_42238_, _42237_, _42225_);
  not (_42239_, _42238_);
  and (_42240_, _42239_, _42128_);
  not (_42241_, _42240_);
  not (_42242_, _38174_);
  and (_42243_, _42242_, _38055_);
  not (_42244_, _41981_);
  and (_42245_, _42126_, _42244_);
  nor (_42246_, _42245_, _42243_);
  and (_42247_, _42246_, _42241_);
  and (_42248_, _42247_, _42224_);
  not (_42249_, _42248_);
  and (_42250_, _42249_, _42097_);
  and (_42251_, _42045_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_42252_, _42039_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_42253_, _42252_, _42251_);
  and (_42254_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_42255_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_42256_, _42255_, _42254_);
  and (_42257_, _42256_, _42253_);
  and (_42258_, _42025_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_42259_, _42035_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_42260_, _42259_, _42258_);
  and (_42261_, _42042_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_42262_, _42028_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_42263_, _42262_, _42261_);
  and (_42264_, _42263_, _42260_);
  and (_42265_, _42264_, _42257_);
  nor (_42266_, _42265_, _42023_);
  and (_42267_, _42023_, _38124_);
  nor (_42268_, _42267_, _42266_);
  not (_42269_, _42268_);
  and (_42270_, _42269_, _42098_);
  not (_42271_, _42270_);
  and (_42272_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_42273_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_42274_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42275_, _42274_, _42273_);
  and (_42276_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42277_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_42278_, _42277_, _42276_);
  and (_42279_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_42280_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_42281_, _42280_, _42279_);
  and (_42282_, _42281_, _42278_);
  and (_42283_, _42282_, _42275_);
  nor (_42284_, _42283_, _42074_);
  nor (_42285_, _42284_, _42272_);
  not (_42286_, _42285_);
  and (_42287_, _42286_, _42128_);
  not (_42288_, _42287_);
  not (_42289_, _38156_);
  and (_42290_, _42289_, _38055_);
  and (_42291_, _42126_, _37809_);
  nor (_42292_, _42291_, _42290_);
  and (_42293_, _42292_, _42288_);
  and (_42294_, _42293_, _42271_);
  nor (_42295_, _42294_, _42096_);
  nor (_42296_, _42295_, _42250_);
  and (_42297_, _42296_, _42202_);
  nor (_42298_, _42296_, _42202_);
  nor (_42299_, _42298_, _42297_);
  and (_42300_, _42299_, _42201_);
  not (_42301_, _38192_);
  and (_42302_, _42301_, _38055_);
  not (_42303_, _42302_);
  and (_42304_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_42305_, _42045_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_42306_, _42305_, _42304_);
  and (_42307_, _42042_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_42308_, _42028_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_42309_, _42308_, _42307_);
  and (_42310_, _42309_, _42306_);
  and (_42311_, _42025_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_42312_, _42039_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_42313_, _42312_, _42311_);
  and (_42314_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_42315_, _42035_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_42316_, _42315_, _42314_);
  and (_42317_, _42316_, _42313_);
  and (_42318_, _42317_, _42310_);
  nor (_42319_, _42318_, _42023_);
  and (_42320_, _42023_, _40183_);
  nor (_42321_, _42320_, _42319_);
  not (_42322_, _42321_);
  and (_42323_, _42322_, _42098_);
  not (_42324_, _42323_);
  nor (_42325_, _41979_, _37921_);
  and (_42326_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_42327_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42328_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_42329_, _42328_, _42327_);
  and (_42330_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_42331_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42332_, _42331_, _42330_);
  and (_42333_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_42334_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_42335_, _42334_, _42333_);
  and (_42336_, _42335_, _42332_);
  and (_42337_, _42336_, _42329_);
  nor (_42338_, _42337_, _42074_);
  nor (_42339_, _42338_, _42326_);
  not (_42340_, _42339_);
  and (_42341_, _42340_, _42059_);
  nor (_42342_, _42341_, _42325_);
  and (_42343_, _42342_, _42324_);
  and (_42344_, _42343_, _42303_);
  and (_42345_, _42344_, _42097_);
  nor (_42346_, _42249_, _42097_);
  nor (_42347_, _42346_, _42345_);
  nor (_42348_, _42347_, _41955_);
  and (_42349_, _42347_, _41955_);
  nor (_42350_, _42349_, _42348_);
  not (_42351_, _41959_);
  and (_42352_, _38054_, _42058_);
  not (_42353_, _42352_);
  and (_42354_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_42355_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42356_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_42357_, _42356_, _42355_);
  and (_42358_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_42359_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_42360_, _42359_, _42358_);
  and (_42361_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_42362_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_42363_, _42362_, _42361_);
  and (_42364_, _42363_, _42360_);
  and (_42365_, _42364_, _42357_);
  nor (_42366_, _42365_, _42074_);
  nor (_42367_, _42366_, _42354_);
  not (_42368_, _42367_);
  and (_42369_, _42368_, _42128_);
  and (_42370_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_42371_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_42372_, _42371_, _42370_);
  and (_42373_, _42028_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_42374_, _42025_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_42375_, _42374_, _42373_);
  and (_42376_, _42375_, _42372_);
  and (_42377_, _42035_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_42378_, _42039_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_42379_, _42378_, _42377_);
  and (_42380_, _42045_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_42381_, _42042_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_42382_, _42381_, _42380_);
  and (_42383_, _42382_, _42379_);
  and (_42384_, _42383_, _42376_);
  nor (_42385_, _42384_, _42023_);
  not (_42386_, _38085_);
  and (_42387_, _42023_, _42386_);
  nor (_42388_, _42387_, _42385_);
  not (_42389_, _42388_);
  and (_42390_, _42389_, _42098_);
  nor (_42391_, _42390_, _42369_);
  and (_42392_, _42121_, _38018_);
  not (_42393_, _38186_);
  and (_42394_, _42393_, _38055_);
  nor (_42395_, _42394_, _42392_);
  and (_42396_, _42395_, _42391_);
  and (_42397_, _42396_, _42353_);
  not (_42398_, _42397_);
  and (_42399_, _42398_, _42097_);
  and (_42400_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_42401_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_42402_, _42401_, _42400_);
  and (_42403_, _42028_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_42404_, _42025_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_42405_, _42404_, _42403_);
  and (_42406_, _42405_, _42402_);
  and (_42407_, _42045_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_42408_, _42039_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_42409_, _42408_, _42407_);
  and (_42410_, _42035_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_42411_, _42042_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_42412_, _42411_, _42410_);
  and (_42413_, _42412_, _42409_);
  and (_42414_, _42413_, _42406_);
  nor (_42415_, _42414_, _42023_);
  not (_42416_, _38108_);
  and (_42417_, _42023_, _42416_);
  nor (_42418_, _42417_, _42415_);
  not (_42419_, _42418_);
  and (_42420_, _42419_, _42098_);
  not (_42421_, _42420_);
  and (_42422_, _42126_, _37880_);
  and (_42423_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_42424_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_42425_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_42426_, _42425_, _42424_);
  and (_42427_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_42428_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_42429_, _42428_, _42427_);
  and (_42430_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_42431_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_42432_, _42431_, _42430_);
  and (_42433_, _42432_, _42429_);
  and (_42434_, _42433_, _42426_);
  nor (_42435_, _42434_, _42074_);
  nor (_42436_, _42435_, _42423_);
  not (_42437_, _42436_);
  and (_42438_, _42437_, _42128_);
  not (_42439_, _38168_);
  and (_42440_, _42439_, _38055_);
  or (_42441_, _42440_, _42438_);
  nor (_42442_, _42441_, _42422_);
  and (_42443_, _42442_, _42421_);
  nor (_42444_, _42443_, _42096_);
  nor (_42445_, _42444_, _42399_);
  and (_42446_, _42445_, _42351_);
  nor (_42447_, _42445_, _42351_);
  nor (_42448_, _42447_, _42446_);
  and (_42449_, _42448_, _42350_);
  and (_42450_, _42449_, _42300_);
  and (_42451_, _42450_, _41945_);
  nor (_42452_, _42147_, _42097_);
  nor (_42453_, _41940_, _28417_);
  not (_42454_, _42453_);
  and (_42455_, _42454_, _42452_);
  nor (_42456_, _42454_, _42452_);
  nor (_42457_, _42456_, _42455_);
  nor (_42458_, _42398_, _42097_);
  nor (_42459_, _41940_, _38617_);
  not (_42460_, _42459_);
  nor (_42461_, _42460_, _42458_);
  and (_42462_, _42460_, _42458_);
  nor (_42463_, _42462_, _42461_);
  and (_42464_, _42463_, _42457_);
  nor (_42465_, _42081_, _28099_);
  and (_42466_, _42081_, _28099_);
  nor (_42467_, _42466_, _42465_);
  nor (_42468_, _42344_, _42097_);
  nor (_42469_, _41940_, _27803_);
  not (_42470_, _42469_);
  and (_42471_, _42470_, _42468_);
  nor (_42472_, _42470_, _42468_);
  nor (_42473_, _42472_, _42471_);
  and (_42474_, _42473_, _42467_);
  and (_42475_, _42474_, _42464_);
  and (_42476_, _42475_, _42451_);
  not (_42477_, _42445_);
  not (_42478_, _42296_);
  and (_42480_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_42481_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_42483_, _42481_, _42197_);
  or (_42485_, _42483_, _42480_);
  and (_42486_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_42488_, _42197_);
  and (_42490_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_42492_, _42490_, _42488_);
  or (_42494_, _42492_, _42486_);
  and (_42495_, _42494_, _42485_);
  or (_42496_, _42495_, _42477_);
  not (_42497_, _42347_);
  and (_42498_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_42499_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_42500_, _42499_, _42197_);
  or (_42501_, _42500_, _42498_);
  and (_42502_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_42503_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_42504_, _42503_, _42488_);
  or (_42505_, _42504_, _42502_);
  and (_42506_, _42505_, _42501_);
  or (_42507_, _42506_, _42445_);
  and (_42508_, _42507_, _42497_);
  and (_42509_, _42508_, _42496_);
  or (_42510_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_42511_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_42512_, _42511_, _42510_);
  or (_42513_, _42512_, _42488_);
  or (_42514_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_42515_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_42516_, _42515_, _42514_);
  or (_42517_, _42516_, _42197_);
  and (_42518_, _42517_, _42513_);
  or (_42519_, _42518_, _42477_);
  or (_42520_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_42521_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_42522_, _42521_, _42520_);
  or (_42523_, _42522_, _42488_);
  or (_42524_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_42525_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_42526_, _42525_, _42524_);
  or (_42527_, _42526_, _42197_);
  and (_42528_, _42527_, _42523_);
  or (_42529_, _42528_, _42445_);
  and (_42530_, _42529_, _42347_);
  and (_42532_, _42530_, _42519_);
  or (_42534_, _42532_, _42509_);
  or (_42536_, _42534_, _42476_);
  not (_42538_, _42476_);
  or (_42540_, _42538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_42542_, _42538_, _42451_);
  nor (_42544_, _42542_, rst);
  and (_42546_, _42544_, _42540_);
  and (_42547_, _42546_, _42536_);
  and (_39585_, _41971_, _42545_);
  and (_42550_, _39585_, _42542_);
  or (_02573_, _42550_, _42547_);
  nor (_42551_, _41960_, _41956_);
  nor (_42552_, _41951_, _41947_);
  and (_42553_, _42552_, _41945_);
  and (_42554_, _42553_, _42551_);
  and (_42555_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _28856_);
  and (_42556_, _42555_, _28910_);
  nand (_42557_, _42556_, _31732_);
  not (_42558_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42559_, _38123_, _42558_);
  or (_42560_, _19439_, _42558_);
  and (_42561_, _42560_, _42559_);
  or (_42562_, _42561_, _42556_);
  and (_42563_, _42562_, _42557_);
  and (_42564_, _42563_, _42554_);
  not (_42565_, _42554_);
  and (_42566_, _42565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_02617_, _42566_, _42564_);
  nand (_42567_, _42555_, _28976_);
  nor (_42568_, _42567_, _31732_);
  nor (_42569_, _38115_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42570_, _42555_, _28933_);
  and (_42571_, _42555_, _28867_);
  or (_42572_, _42571_, _41963_);
  or (_42573_, _42572_, _42570_);
  and (_42574_, _42573_, _20424_);
  or (_42575_, _42574_, _42569_);
  or (_42576_, _42575_, _42568_);
  and (_42577_, _42576_, _42554_);
  and (_42578_, _42565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_02623_, _42578_, _42577_);
  and (_42579_, _42565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_42580_, _42555_, _28944_);
  nor (_42581_, _42580_, _31732_);
  nor (_42582_, _38108_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42583_, _42555_, _28965_);
  or (_42584_, _42583_, _42572_);
  and (_42585_, _42584_, _19077_);
  or (_42586_, _42585_, _42582_);
  or (_42587_, _42586_, _42581_);
  and (_42588_, _42587_, _42554_);
  or (_02628_, _42588_, _42579_);
  and (_42589_, _42571_, _32352_);
  nor (_42590_, _38100_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42591_, _42570_, _41963_);
  or (_42592_, _42591_, _42583_);
  and (_42593_, _42592_, _20109_);
  or (_42594_, _42593_, _42590_);
  or (_42595_, _42594_, _42589_);
  and (_42596_, _42595_, _42554_);
  and (_42597_, _42565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_02634_, _42597_, _42596_);
  nand (_42598_, _41963_, _28910_);
  nor (_42599_, _42598_, _31732_);
  nor (_42600_, _38092_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42601_, _28910_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42602_, _19275_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42603_, _42602_, _42601_);
  or (_42604_, _42603_, _42600_);
  or (_42605_, _42604_, _42599_);
  and (_42606_, _42605_, _42554_);
  and (_42607_, _42565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_02638_, _42607_, _42606_);
  nand (_42608_, _41963_, _28976_);
  nor (_42609_, _42608_, _31732_);
  nor (_42610_, _38085_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42611_, _28976_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42612_, _20261_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42613_, _42612_, _42611_);
  or (_42614_, _42613_, _42610_);
  or (_42615_, _42614_, _42609_);
  and (_42616_, _42615_, _42554_);
  and (_42617_, _42565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_02642_, _42617_, _42616_);
  nand (_42618_, _41963_, _28944_);
  nor (_42619_, _42618_, _31732_);
  nor (_42620_, _38078_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42621_, _28944_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42622_, _19613_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42623_, _42622_, _42621_);
  or (_42624_, _42623_, _42620_);
  or (_42625_, _42624_, _42619_);
  and (_42626_, _42625_, _42554_);
  and (_42627_, _42565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_02647_, _42627_, _42626_);
  and (_42628_, _42565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_42629_, _42554_, _41971_);
  or (_02649_, _42629_, _42628_);
  and (_42630_, _42563_, _41945_);
  and (_42631_, _41950_, _41947_);
  and (_42632_, _42631_, _42551_);
  and (_42633_, _42632_, _42630_);
  not (_42634_, _42632_);
  and (_42635_, _42634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_02655_, _42635_, _42633_);
  and (_42636_, _42576_, _41945_);
  and (_42637_, _42632_, _42636_);
  and (_42638_, _42634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_02658_, _42638_, _42637_);
  and (_42639_, _42587_, _41945_);
  and (_42640_, _42632_, _42639_);
  and (_42641_, _42634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_02662_, _42641_, _42640_);
  and (_42642_, _42595_, _41945_);
  and (_42643_, _42632_, _42642_);
  and (_42644_, _42634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_02665_, _42644_, _42643_);
  and (_42645_, _42605_, _41945_);
  and (_42646_, _42632_, _42645_);
  and (_42647_, _42634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_02669_, _42647_, _42646_);
  and (_42648_, _42615_, _41945_);
  and (_42649_, _42632_, _42648_);
  and (_42650_, _42634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_02672_, _42650_, _42649_);
  and (_42651_, _42625_, _41945_);
  and (_42652_, _42632_, _42651_);
  and (_42653_, _42634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_02675_, _42653_, _42652_);
  and (_42654_, _42632_, _41972_);
  and (_42655_, _42634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_02677_, _42655_, _42654_);
  and (_42656_, _41951_, _41943_);
  and (_42657_, _42656_, _42551_);
  and (_42658_, _42657_, _42630_);
  not (_42659_, _42657_);
  and (_42660_, _42659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_02684_, _42660_, _42658_);
  and (_42661_, _42657_, _42636_);
  and (_42662_, _42659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_02687_, _42662_, _42661_);
  and (_42663_, _42657_, _42639_);
  and (_42664_, _42659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_02690_, _42664_, _42663_);
  and (_42665_, _42657_, _42642_);
  and (_42666_, _42659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_02692_, _42666_, _42665_);
  and (_42667_, _42657_, _42645_);
  and (_42668_, _42659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_02694_, _42668_, _42667_);
  and (_42669_, _42657_, _42648_);
  and (_42670_, _42659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_02697_, _42670_, _42669_);
  and (_42671_, _42657_, _42651_);
  and (_42672_, _42659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_02701_, _42672_, _42671_);
  and (_42673_, _42657_, _41972_);
  and (_42674_, _42659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_02703_, _42674_, _42673_);
  and (_42675_, _42551_, _41952_);
  and (_42676_, _42675_, _42630_);
  not (_42677_, _42675_);
  and (_42678_, _42677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_02708_, _42678_, _42676_);
  and (_42679_, _42675_, _42636_);
  and (_42680_, _42677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_02711_, _42680_, _42679_);
  and (_42681_, _42675_, _42639_);
  and (_42682_, _42677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_02714_, _42682_, _42681_);
  and (_42683_, _42675_, _42642_);
  and (_42684_, _42677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_02718_, _42684_, _42683_);
  and (_42685_, _42675_, _42645_);
  and (_42686_, _42677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_02721_, _42686_, _42685_);
  and (_42687_, _42675_, _42648_);
  and (_42688_, _42677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_02724_, _42688_, _42687_);
  and (_42689_, _42675_, _42651_);
  and (_42690_, _42677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_02727_, _42690_, _42689_);
  and (_42691_, _42675_, _41972_);
  and (_42692_, _42677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_02730_, _42692_, _42691_);
  and (_42693_, _41960_, _41955_);
  and (_42694_, _42693_, _42552_);
  and (_42695_, _42694_, _42630_);
  not (_42696_, _42694_);
  and (_42697_, _42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_02737_, _42697_, _42695_);
  and (_42698_, _42694_, _42636_);
  and (_42699_, _42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_02740_, _42699_, _42698_);
  and (_42700_, _42694_, _42639_);
  and (_42701_, _42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_02744_, _42701_, _42700_);
  and (_42702_, _42694_, _42642_);
  and (_42703_, _42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_02747_, _42703_, _42702_);
  and (_42704_, _42694_, _42645_);
  and (_42705_, _42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_02750_, _42705_, _42704_);
  and (_42706_, _42694_, _42648_);
  and (_42707_, _42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_02753_, _42707_, _42706_);
  and (_42708_, _42694_, _42651_);
  and (_42709_, _42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_02757_, _42709_, _42708_);
  and (_42710_, _42694_, _41972_);
  and (_42711_, _42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_02759_, _42711_, _42710_);
  and (_42712_, _42693_, _42631_);
  and (_42713_, _42712_, _42630_);
  not (_42714_, _42712_);
  and (_42715_, _42714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_02763_, _42715_, _42713_);
  and (_42716_, _42712_, _42636_);
  and (_42717_, _42714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_02766_, _42717_, _42716_);
  and (_42718_, _42712_, _42639_);
  and (_42719_, _42714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_02770_, _42719_, _42718_);
  and (_42720_, _42712_, _42642_);
  and (_42721_, _42714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_02773_, _42721_, _42720_);
  and (_42722_, _42712_, _42645_);
  and (_42723_, _42714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_02776_, _42723_, _42722_);
  and (_42724_, _42712_, _42648_);
  and (_42725_, _42714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_02779_, _42725_, _42724_);
  and (_42726_, _42712_, _42651_);
  and (_42727_, _42714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_02783_, _42727_, _42726_);
  and (_42728_, _42712_, _41972_);
  and (_42729_, _42714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_02785_, _42729_, _42728_);
  and (_42730_, _42693_, _42656_);
  and (_42731_, _42730_, _42630_);
  not (_42732_, _42730_);
  and (_42733_, _42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_02789_, _42733_, _42731_);
  and (_42734_, _42730_, _42636_);
  and (_42735_, _42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_02792_, _42735_, _42734_);
  and (_42736_, _42730_, _42639_);
  and (_42737_, _42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_02796_, _42737_, _42736_);
  and (_42738_, _42730_, _42642_);
  and (_42739_, _42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_02799_, _42739_, _42738_);
  and (_42740_, _42730_, _42645_);
  and (_42741_, _42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_02802_, _42741_, _42740_);
  and (_42742_, _42730_, _42648_);
  and (_42743_, _42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_02805_, _42743_, _42742_);
  and (_42744_, _42730_, _42651_);
  and (_42745_, _42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_02809_, _42745_, _42744_);
  and (_42746_, _42730_, _41972_);
  and (_42747_, _42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_02811_, _42747_, _42746_);
  and (_42748_, _42693_, _41952_);
  and (_42749_, _42748_, _42630_);
  not (_42750_, _42748_);
  and (_42751_, _42750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_02815_, _42751_, _42749_);
  and (_42752_, _42748_, _42636_);
  and (_42753_, _42750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_02818_, _42753_, _42752_);
  and (_42754_, _42748_, _42639_);
  and (_42755_, _42750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_02822_, _42755_, _42754_);
  and (_42756_, _42748_, _42642_);
  and (_42757_, _42750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_02825_, _42757_, _42756_);
  and (_42758_, _42748_, _42645_);
  and (_42759_, _42750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_02828_, _42759_, _42758_);
  and (_42760_, _42748_, _42648_);
  and (_42761_, _42750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_02831_, _42761_, _42760_);
  and (_42762_, _42748_, _42651_);
  and (_42763_, _42750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_02835_, _42763_, _42762_);
  and (_42764_, _42748_, _41972_);
  and (_42765_, _42750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_02837_, _42765_, _42764_);
  and (_42766_, _41959_, _41956_);
  and (_42767_, _42766_, _42552_);
  and (_42768_, _42767_, _42630_);
  not (_42769_, _42767_);
  and (_42770_, _42769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_02843_, _42770_, _42768_);
  and (_42771_, _42767_, _42636_);
  and (_42772_, _42769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_02847_, _42772_, _42771_);
  and (_42773_, _42767_, _42639_);
  and (_42774_, _42769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_02850_, _42774_, _42773_);
  and (_42775_, _42767_, _42642_);
  and (_42776_, _42769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_02853_, _42776_, _42775_);
  and (_42777_, _42767_, _42645_);
  and (_42778_, _42769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_02856_, _42778_, _42777_);
  and (_42779_, _42767_, _42648_);
  and (_42780_, _42769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_02860_, _42780_, _42779_);
  and (_42781_, _42767_, _42651_);
  and (_42782_, _42769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_02864_, _42782_, _42781_);
  and (_42783_, _42767_, _41972_);
  and (_42784_, _42769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_02866_, _42784_, _42783_);
  and (_42785_, _42766_, _42631_);
  and (_42786_, _42785_, _42630_);
  not (_42787_, _42785_);
  and (_42788_, _42787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_02871_, _42788_, _42786_);
  and (_42789_, _42785_, _42636_);
  and (_42790_, _42787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_02874_, _42790_, _42789_);
  and (_42791_, _42785_, _42639_);
  and (_42792_, _42787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_02878_, _42792_, _42791_);
  and (_42793_, _42785_, _42642_);
  and (_42794_, _42787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_02881_, _42794_, _42793_);
  and (_42795_, _42785_, _42645_);
  and (_42796_, _42787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_02885_, _42796_, _42795_);
  and (_42797_, _42785_, _42648_);
  and (_42798_, _42787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_02889_, _42798_, _42797_);
  and (_42799_, _42785_, _42651_);
  and (_42800_, _42787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_02892_, _42800_, _42799_);
  and (_42801_, _42785_, _41972_);
  and (_42802_, _42787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_02895_, _42802_, _42801_);
  and (_42803_, _42766_, _42656_);
  and (_42804_, _42803_, _42630_);
  not (_42805_, _42803_);
  and (_42806_, _42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_02899_, _42806_, _42804_);
  and (_42807_, _42803_, _42636_);
  and (_42808_, _42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_02903_, _42808_, _42807_);
  and (_42809_, _42803_, _42639_);
  and (_42810_, _42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_02906_, _42810_, _42809_);
  and (_42811_, _42803_, _42642_);
  and (_42812_, _42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_02910_, _42812_, _42811_);
  and (_42813_, _42803_, _42645_);
  and (_42814_, _42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_02914_, _42814_, _42813_);
  and (_42815_, _42803_, _42648_);
  and (_42816_, _42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_02918_, _42816_, _42815_);
  and (_42817_, _42803_, _42651_);
  and (_42818_, _42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_02922_, _42818_, _42817_);
  and (_42819_, _42803_, _41972_);
  and (_42820_, _42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_02924_, _42820_, _42819_);
  and (_42821_, _42766_, _41952_);
  and (_42822_, _42821_, _42630_);
  not (_42823_, _42821_);
  and (_42824_, _42823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_02930_, _42824_, _42822_);
  and (_42825_, _42821_, _42636_);
  and (_42826_, _42823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_02933_, _42826_, _42825_);
  and (_42827_, _42821_, _42639_);
  and (_42828_, _42823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_02936_, _42828_, _42827_);
  and (_42829_, _42821_, _42642_);
  and (_42830_, _42823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_02940_, _42830_, _42829_);
  and (_42831_, _42821_, _42645_);
  and (_42832_, _42823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_02943_, _42832_, _42831_);
  and (_42833_, _42821_, _42648_);
  and (_42834_, _42823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_02947_, _42834_, _42833_);
  and (_42835_, _42821_, _42651_);
  and (_42836_, _42823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_02950_, _42836_, _42835_);
  and (_42837_, _42821_, _41972_);
  and (_42838_, _42823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_02954_, _42838_, _42837_);
  and (_42839_, _42552_, _41961_);
  and (_42840_, _42839_, _42630_);
  not (_42841_, _42839_);
  and (_42842_, _42841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_02959_, _42842_, _42840_);
  and (_42843_, _42839_, _42636_);
  and (_42844_, _42841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_02962_, _42844_, _42843_);
  and (_42845_, _42839_, _42639_);
  and (_42846_, _42841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_02966_, _42846_, _42845_);
  and (_42847_, _42839_, _42642_);
  and (_42848_, _42841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_02970_, _42848_, _42847_);
  and (_42849_, _42839_, _42645_);
  and (_42850_, _42841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_02973_, _42850_, _42849_);
  and (_42851_, _42839_, _42648_);
  and (_42852_, _42841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_02977_, _42852_, _42851_);
  and (_42853_, _42839_, _42651_);
  and (_42854_, _42841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_02980_, _42854_, _42853_);
  and (_42855_, _42839_, _41972_);
  and (_42856_, _42841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_02983_, _42856_, _42855_);
  and (_42857_, _42631_, _41961_);
  and (_42858_, _42857_, _42630_);
  not (_42859_, _42857_);
  and (_42860_, _42859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_02987_, _42860_, _42858_);
  and (_42861_, _42857_, _42636_);
  and (_42862_, _42859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_02990_, _42862_, _42861_);
  and (_42863_, _42857_, _42639_);
  and (_42864_, _42859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_02993_, _42864_, _42863_);
  and (_42865_, _42857_, _42642_);
  and (_42866_, _42859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_02997_, _42866_, _42865_);
  and (_42867_, _42857_, _42645_);
  and (_42868_, _42859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_03001_, _42868_, _42867_);
  and (_42869_, _42857_, _42648_);
  and (_42870_, _42859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_03004_, _42870_, _42869_);
  and (_42871_, _42857_, _42651_);
  and (_42872_, _42859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_03007_, _42872_, _42871_);
  and (_42873_, _42857_, _41972_);
  and (_42874_, _42859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_03011_, _42874_, _42873_);
  and (_42875_, _42656_, _41961_);
  and (_42876_, _42875_, _42630_);
  not (_42877_, _42875_);
  and (_42878_, _42877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_03015_, _42878_, _42876_);
  and (_42879_, _42875_, _42636_);
  and (_42880_, _42877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_03018_, _42880_, _42879_);
  and (_42881_, _42875_, _42639_);
  and (_42882_, _42877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_03022_, _42882_, _42881_);
  and (_42883_, _42875_, _42642_);
  and (_42884_, _42877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_03026_, _42884_, _42883_);
  and (_42885_, _42875_, _42645_);
  and (_42886_, _42877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_03029_, _42886_, _42885_);
  and (_42887_, _42875_, _42648_);
  and (_42888_, _42877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_03032_, _42888_, _42887_);
  and (_42897_, _42875_, _42651_);
  and (_42904_, _42877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_03036_, _42904_, _42897_);
  and (_42915_, _42875_, _41972_);
  and (_42920_, _42877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_03038_, _42920_, _42915_);
  and (_42933_, _42630_, _41962_);
  and (_42937_, _41974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_03042_, _42937_, _42933_);
  and (_42951_, _42636_, _41962_);
  and (_42955_, _41974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_03047_, _42955_, _42951_);
  and (_42967_, _42639_, _41962_);
  and (_42973_, _41974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_03051_, _42973_, _42967_);
  and (_42979_, _42642_, _41962_);
  and (_42990_, _41974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_03054_, _42990_, _42979_);
  and (_43000_, _42645_, _41962_);
  and (_43008_, _41974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_03059_, _43008_, _43000_);
  and (_43016_, _42648_, _41962_);
  and (_43024_, _41974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_03063_, _43024_, _43016_);
  and (_43033_, _42651_, _41962_);
  and (_43040_, _41974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_03066_, _43040_, _43033_);
  and (_43051_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_43056_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_43064_, _43056_, _42197_);
  or (_43070_, _43064_, _43051_);
  and (_43073_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_43074_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_43075_, _43074_, _42488_);
  or (_43076_, _43075_, _43073_);
  and (_43077_, _43076_, _43070_);
  or (_43078_, _43077_, _42477_);
  and (_43079_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_43080_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_43081_, _43080_, _42197_);
  or (_43082_, _43081_, _43079_);
  and (_43083_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_43084_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_43085_, _43084_, _42488_);
  or (_43086_, _43085_, _43083_);
  and (_43087_, _43086_, _43082_);
  or (_43088_, _43087_, _42445_);
  and (_43089_, _43088_, _42497_);
  and (_43090_, _43089_, _43078_);
  or (_43091_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_43092_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_43093_, _43092_, _43091_);
  or (_43094_, _43093_, _42488_);
  or (_43095_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_43096_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_43097_, _43096_, _43095_);
  or (_43098_, _43097_, _42197_);
  and (_43099_, _43098_, _43094_);
  or (_43100_, _43099_, _42477_);
  or (_43101_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_43102_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_43103_, _43102_, _43101_);
  or (_43104_, _43103_, _42488_);
  or (_43105_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_43106_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_43107_, _43106_, _43105_);
  or (_43108_, _43107_, _42197_);
  and (_43109_, _43108_, _43104_);
  or (_43110_, _43109_, _42445_);
  and (_43111_, _43110_, _42347_);
  and (_43112_, _43111_, _43100_);
  or (_43113_, _43112_, _43090_);
  or (_43114_, _43113_, _42476_);
  or (_43115_, _42538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_43116_, _43115_, _42544_);
  and (_43117_, _43116_, _43114_);
  and (_39604_, _42563_, _42545_);
  and (_43118_, _39604_, _42542_);
  or (_03193_, _43118_, _43117_);
  and (_43119_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_43120_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_43121_, _43120_, _42197_);
  or (_43122_, _43121_, _43119_);
  and (_43123_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_43124_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_43125_, _43124_, _42488_);
  or (_43126_, _43125_, _43123_);
  and (_43127_, _43126_, _43122_);
  or (_43128_, _43127_, _42477_);
  and (_43129_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_43130_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_43131_, _43130_, _42197_);
  or (_43132_, _43131_, _43129_);
  and (_43133_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_43134_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_43135_, _43134_, _42488_);
  or (_43136_, _43135_, _43133_);
  and (_43137_, _43136_, _43132_);
  or (_43138_, _43137_, _42445_);
  and (_43139_, _43138_, _42497_);
  and (_43140_, _43139_, _43128_);
  or (_43141_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_43142_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_43143_, _43142_, _43141_);
  or (_43144_, _43143_, _42488_);
  or (_43145_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_43146_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_43147_, _43146_, _43145_);
  or (_43148_, _43147_, _42197_);
  and (_43149_, _43148_, _43144_);
  or (_43150_, _43149_, _42477_);
  or (_43151_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_43152_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_43153_, _43152_, _43151_);
  or (_43154_, _43153_, _42488_);
  or (_43155_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_43156_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_43157_, _43156_, _43155_);
  or (_43158_, _43157_, _42197_);
  and (_43159_, _43158_, _43154_);
  or (_43160_, _43159_, _42445_);
  and (_43161_, _43160_, _42347_);
  and (_43162_, _43161_, _43150_);
  or (_43163_, _43162_, _43140_);
  or (_43164_, _43163_, _42476_);
  or (_43165_, _42538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_43166_, _43165_, _42544_);
  and (_43167_, _43166_, _43164_);
  and (_39605_, _42576_, _42545_);
  and (_43168_, _39605_, _42542_);
  or (_03194_, _43168_, _43167_);
  and (_43169_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and (_43170_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_43171_, _43170_, _42197_);
  or (_43172_, _43171_, _43169_);
  and (_43173_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_43174_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_43175_, _43174_, _42488_);
  or (_43176_, _43175_, _43173_);
  and (_43177_, _43176_, _43172_);
  or (_43178_, _43177_, _42477_);
  and (_43179_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_43180_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_43181_, _43180_, _42197_);
  or (_43182_, _43181_, _43179_);
  and (_43183_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_43184_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_43185_, _43184_, _42488_);
  or (_43186_, _43185_, _43183_);
  and (_43187_, _43186_, _43182_);
  or (_43188_, _43187_, _42445_);
  and (_43189_, _43188_, _42497_);
  and (_43190_, _43189_, _43178_);
  or (_43191_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_43192_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_43193_, _43192_, _43191_);
  or (_43194_, _43193_, _42488_);
  or (_43195_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_43196_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_43197_, _43196_, _43195_);
  or (_43198_, _43197_, _42197_);
  and (_43199_, _43198_, _43194_);
  or (_43200_, _43199_, _42477_);
  or (_43201_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_43202_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_43203_, _43202_, _43201_);
  or (_43204_, _43203_, _42488_);
  or (_43205_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_43206_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_43207_, _43206_, _43205_);
  or (_43208_, _43207_, _42197_);
  and (_43209_, _43208_, _43204_);
  or (_43210_, _43209_, _42445_);
  and (_43211_, _43210_, _42347_);
  and (_43212_, _43211_, _43200_);
  or (_43213_, _43212_, _43190_);
  or (_43214_, _43213_, _42476_);
  or (_43215_, _42538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_43216_, _43215_, _42544_);
  and (_43217_, _43216_, _43214_);
  and (_39606_, _42587_, _42545_);
  and (_43218_, _39606_, _42542_);
  or (_03196_, _43218_, _43217_);
  and (_43219_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_43220_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_43221_, _43220_, _42197_);
  or (_43222_, _43221_, _43219_);
  and (_43223_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_43224_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_43225_, _43224_, _42488_);
  or (_43226_, _43225_, _43223_);
  and (_43227_, _43226_, _43222_);
  or (_43228_, _43227_, _42477_);
  and (_43229_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_43230_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_43231_, _43230_, _42197_);
  or (_43232_, _43231_, _43229_);
  and (_43233_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_43234_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_43235_, _43234_, _42488_);
  or (_43236_, _43235_, _43233_);
  and (_43237_, _43236_, _43232_);
  or (_43238_, _43237_, _42445_);
  and (_43239_, _43238_, _42497_);
  and (_43240_, _43239_, _43228_);
  or (_43241_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_43242_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_43243_, _43242_, _43241_);
  or (_43244_, _43243_, _42488_);
  or (_43245_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_43246_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_43247_, _43246_, _43245_);
  or (_43248_, _43247_, _42197_);
  and (_43249_, _43248_, _43244_);
  or (_43250_, _43249_, _42477_);
  or (_43251_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_43252_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_43253_, _43252_, _43251_);
  or (_43254_, _43253_, _42488_);
  or (_43255_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_43256_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_43257_, _43256_, _43255_);
  or (_43258_, _43257_, _42197_);
  and (_43259_, _43258_, _43254_);
  or (_43260_, _43259_, _42445_);
  and (_43261_, _43260_, _42347_);
  and (_43262_, _43261_, _43250_);
  or (_43263_, _43262_, _43240_);
  and (_43264_, _43263_, _42538_);
  and (_43265_, _42476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_43266_, _43265_, _42542_);
  or (_43267_, _43266_, _43264_);
  and (_39607_, _42595_, _42545_);
  or (_43268_, _39607_, _42544_);
  and (_03198_, _43268_, _43267_);
  and (_43269_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_43270_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_43271_, _43270_, _42197_);
  or (_43272_, _43271_, _43269_);
  and (_43273_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_43274_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_43275_, _43274_, _42488_);
  or (_43276_, _43275_, _43273_);
  and (_43277_, _43276_, _43272_);
  or (_43278_, _43277_, _42477_);
  and (_43279_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_43280_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_43281_, _43280_, _42197_);
  or (_43282_, _43281_, _43279_);
  and (_43283_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_43284_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_43285_, _43284_, _42488_);
  or (_43286_, _43285_, _43283_);
  and (_43287_, _43286_, _43282_);
  or (_43288_, _43287_, _42445_);
  and (_43289_, _43288_, _42497_);
  and (_43290_, _43289_, _43278_);
  or (_43291_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_43292_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_43293_, _43292_, _43291_);
  or (_43294_, _43293_, _42488_);
  or (_43295_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_43296_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_43297_, _43296_, _43295_);
  or (_43298_, _43297_, _42197_);
  and (_43299_, _43298_, _43294_);
  or (_43300_, _43299_, _42477_);
  or (_43301_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_43302_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_43303_, _43302_, _43301_);
  or (_43304_, _43303_, _42488_);
  or (_43305_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_43306_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_43307_, _43306_, _43305_);
  or (_43308_, _43307_, _42197_);
  and (_43309_, _43308_, _43304_);
  or (_43310_, _43309_, _42445_);
  and (_43311_, _43310_, _42347_);
  and (_43312_, _43311_, _43300_);
  or (_43313_, _43312_, _43290_);
  or (_43314_, _43313_, _42476_);
  or (_43315_, _42538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_43316_, _43315_, _42544_);
  and (_43317_, _43316_, _43314_);
  and (_39608_, _42605_, _42545_);
  and (_43318_, _39608_, _42542_);
  or (_03200_, _43318_, _43317_);
  and (_43319_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_43320_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_43321_, _43320_, _42197_);
  or (_43322_, _43321_, _43319_);
  and (_43323_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_43324_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_43325_, _43324_, _42488_);
  or (_43326_, _43325_, _43323_);
  and (_43327_, _43326_, _43322_);
  or (_43328_, _43327_, _42477_);
  and (_43329_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_43330_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_43331_, _43330_, _42197_);
  or (_43332_, _43331_, _43329_);
  and (_43333_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_43334_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_43335_, _43334_, _42488_);
  or (_43336_, _43335_, _43333_);
  and (_43337_, _43336_, _43332_);
  or (_43338_, _43337_, _42445_);
  and (_43339_, _43338_, _42497_);
  and (_43340_, _43339_, _43328_);
  or (_43341_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_43342_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_43343_, _43342_, _43341_);
  or (_43344_, _43343_, _42488_);
  or (_43345_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_43346_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_43347_, _43346_, _43345_);
  or (_43348_, _43347_, _42197_);
  and (_43349_, _43348_, _43344_);
  or (_43350_, _43349_, _42477_);
  or (_43351_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_43352_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_43353_, _43352_, _43351_);
  or (_43354_, _43353_, _42488_);
  or (_43355_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_43356_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_43357_, _43356_, _43355_);
  or (_43358_, _43357_, _42197_);
  and (_43359_, _43358_, _43354_);
  or (_43360_, _43359_, _42445_);
  and (_43361_, _43360_, _42347_);
  and (_43362_, _43361_, _43350_);
  or (_43363_, _43362_, _43340_);
  or (_43364_, _43363_, _42476_);
  or (_43365_, _42538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_43366_, _43365_, _42544_);
  and (_43367_, _43366_, _43364_);
  and (_39609_, _42615_, _42545_);
  and (_43368_, _39609_, _42542_);
  or (_03201_, _43368_, _43367_);
  and (_43369_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_43370_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_43371_, _43370_, _42197_);
  or (_43372_, _43371_, _43369_);
  and (_43373_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_43374_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_43375_, _43374_, _42488_);
  or (_43376_, _43375_, _43373_);
  and (_43377_, _43376_, _43372_);
  or (_43378_, _43377_, _42477_);
  and (_43379_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_43380_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_43381_, _43380_, _42197_);
  or (_43382_, _43381_, _43379_);
  and (_43383_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_43384_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_43385_, _43384_, _42488_);
  or (_43386_, _43385_, _43383_);
  and (_43387_, _43386_, _43382_);
  or (_43388_, _43387_, _42445_);
  and (_43389_, _43388_, _42497_);
  and (_43390_, _43389_, _43378_);
  or (_43391_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_43392_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_43393_, _43392_, _43391_);
  or (_43394_, _43393_, _42488_);
  or (_43395_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_43396_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_43397_, _43396_, _43395_);
  or (_43398_, _43397_, _42197_);
  and (_43399_, _43398_, _43394_);
  or (_43400_, _43399_, _42477_);
  or (_43401_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_43402_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_43403_, _43402_, _43401_);
  or (_43404_, _43403_, _42488_);
  or (_43405_, _42296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_43406_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_43407_, _43406_, _43405_);
  or (_43408_, _43407_, _42197_);
  and (_43409_, _43408_, _43404_);
  or (_43410_, _43409_, _42445_);
  and (_43411_, _43410_, _42347_);
  and (_43412_, _43411_, _43400_);
  or (_43413_, _43412_, _43390_);
  and (_43414_, _43413_, _42538_);
  and (_43415_, _42476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or (_43416_, _43415_, _42542_);
  or (_43417_, _43416_, _43414_);
  and (_39610_, _42625_, _42545_);
  or (_43418_, _39610_, _42544_);
  and (_03203_, _43418_, _43417_);
  or (_43419_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_43420_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_43421_, _43420_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_43422_, _43421_, _43419_);
  nand (_43423_, _43422_, _42545_);
  or (_43424_, \oc8051_gm_cxrom_1.cell0.data [7], _42545_);
  and (_03209_, _43424_, _43423_);
  or (_43425_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43426_, \oc8051_gm_cxrom_1.cell0.data [0], _43420_);
  nand (_43427_, _43426_, _43425_);
  nand (_43428_, _43427_, _42545_);
  or (_43429_, \oc8051_gm_cxrom_1.cell0.data [0], _42545_);
  and (_03215_, _43429_, _43428_);
  or (_43430_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43431_, \oc8051_gm_cxrom_1.cell0.data [1], _43420_);
  nand (_43432_, _43431_, _43430_);
  nand (_43433_, _43432_, _42545_);
  or (_43434_, \oc8051_gm_cxrom_1.cell0.data [1], _42545_);
  and (_03218_, _43434_, _43433_);
  or (_43435_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43436_, \oc8051_gm_cxrom_1.cell0.data [2], _43420_);
  nand (_43437_, _43436_, _43435_);
  nand (_43438_, _43437_, _42545_);
  or (_43439_, \oc8051_gm_cxrom_1.cell0.data [2], _42545_);
  and (_03222_, _43439_, _43438_);
  or (_43440_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43441_, \oc8051_gm_cxrom_1.cell0.data [3], _43420_);
  nand (_43442_, _43441_, _43440_);
  nand (_43443_, _43442_, _42545_);
  or (_43444_, \oc8051_gm_cxrom_1.cell0.data [3], _42545_);
  and (_03225_, _43444_, _43443_);
  or (_43445_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43446_, \oc8051_gm_cxrom_1.cell0.data [4], _43420_);
  nand (_43447_, _43446_, _43445_);
  nand (_43448_, _43447_, _42545_);
  or (_43449_, \oc8051_gm_cxrom_1.cell0.data [4], _42545_);
  and (_03228_, _43449_, _43448_);
  or (_43450_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43451_, \oc8051_gm_cxrom_1.cell0.data [5], _43420_);
  nand (_43452_, _43451_, _43450_);
  nand (_43453_, _43452_, _42545_);
  or (_43454_, \oc8051_gm_cxrom_1.cell0.data [5], _42545_);
  and (_03232_, _43454_, _43453_);
  or (_43455_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43456_, \oc8051_gm_cxrom_1.cell0.data [6], _43420_);
  nand (_43457_, _43456_, _43455_);
  nand (_43458_, _43457_, _42545_);
  or (_43459_, \oc8051_gm_cxrom_1.cell0.data [6], _42545_);
  and (_03235_, _43459_, _43458_);
  or (_00001_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_00002_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_00003_, _00002_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_00004_, _00003_, _00001_);
  nand (_00005_, _00004_, _42545_);
  or (_00006_, \oc8051_gm_cxrom_1.cell1.data [7], _42545_);
  and (_03254_, _00006_, _00005_);
  or (_00007_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00008_, \oc8051_gm_cxrom_1.cell1.data [0], _00002_);
  nand (_00009_, _00008_, _00007_);
  nand (_00010_, _00009_, _42545_);
  or (_00011_, \oc8051_gm_cxrom_1.cell1.data [0], _42545_);
  and (_03260_, _00011_, _00010_);
  or (_00012_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00013_, \oc8051_gm_cxrom_1.cell1.data [1], _00002_);
  nand (_00014_, _00013_, _00012_);
  nand (_00015_, _00014_, _42545_);
  or (_00016_, \oc8051_gm_cxrom_1.cell1.data [1], _42545_);
  and (_03263_, _00016_, _00015_);
  or (_00017_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00018_, \oc8051_gm_cxrom_1.cell1.data [2], _00002_);
  nand (_00019_, _00018_, _00017_);
  nand (_00020_, _00019_, _42545_);
  or (_00021_, \oc8051_gm_cxrom_1.cell1.data [2], _42545_);
  and (_03267_, _00021_, _00020_);
  or (_00022_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00023_, \oc8051_gm_cxrom_1.cell1.data [3], _00002_);
  nand (_00024_, _00023_, _00022_);
  nand (_00025_, _00024_, _42545_);
  or (_00026_, \oc8051_gm_cxrom_1.cell1.data [3], _42545_);
  and (_03270_, _00026_, _00025_);
  or (_00027_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00028_, \oc8051_gm_cxrom_1.cell1.data [4], _00002_);
  nand (_00029_, _00028_, _00027_);
  nand (_00030_, _00029_, _42545_);
  or (_00031_, \oc8051_gm_cxrom_1.cell1.data [4], _42545_);
  and (_03274_, _00031_, _00030_);
  or (_00032_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00033_, \oc8051_gm_cxrom_1.cell1.data [5], _00002_);
  nand (_00034_, _00033_, _00032_);
  nand (_00035_, _00034_, _42545_);
  or (_00036_, \oc8051_gm_cxrom_1.cell1.data [5], _42545_);
  and (_03277_, _00036_, _00035_);
  or (_00037_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00038_, \oc8051_gm_cxrom_1.cell1.data [6], _00002_);
  nand (_00039_, _00038_, _00037_);
  nand (_00040_, _00039_, _42545_);
  or (_00041_, \oc8051_gm_cxrom_1.cell1.data [6], _42545_);
  and (_03280_, _00041_, _00040_);
  or (_00042_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_00043_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_00044_, _00043_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_00045_, _00044_, _00042_);
  nand (_00046_, _00045_, _42545_);
  or (_00047_, \oc8051_gm_cxrom_1.cell2.data [7], _42545_);
  and (_03297_, _00047_, _00046_);
  or (_00048_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00049_, \oc8051_gm_cxrom_1.cell2.data [0], _00043_);
  nand (_00050_, _00049_, _00048_);
  nand (_00051_, _00050_, _42545_);
  or (_00052_, \oc8051_gm_cxrom_1.cell2.data [0], _42545_);
  and (_03304_, _00052_, _00051_);
  or (_00053_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00054_, \oc8051_gm_cxrom_1.cell2.data [1], _00043_);
  nand (_00055_, _00054_, _00053_);
  nand (_00056_, _00055_, _42545_);
  or (_00057_, \oc8051_gm_cxrom_1.cell2.data [1], _42545_);
  and (_03307_, _00057_, _00056_);
  or (_00058_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00059_, \oc8051_gm_cxrom_1.cell2.data [2], _00043_);
  nand (_00060_, _00059_, _00058_);
  nand (_00061_, _00060_, _42545_);
  or (_00062_, \oc8051_gm_cxrom_1.cell2.data [2], _42545_);
  and (_03311_, _00062_, _00061_);
  or (_00063_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00064_, \oc8051_gm_cxrom_1.cell2.data [3], _00043_);
  nand (_00065_, _00064_, _00063_);
  nand (_00066_, _00065_, _42545_);
  or (_00067_, \oc8051_gm_cxrom_1.cell2.data [3], _42545_);
  and (_03314_, _00067_, _00066_);
  or (_00068_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00069_, \oc8051_gm_cxrom_1.cell2.data [4], _00043_);
  nand (_00070_, _00069_, _00068_);
  nand (_00071_, _00070_, _42545_);
  or (_00072_, \oc8051_gm_cxrom_1.cell2.data [4], _42545_);
  and (_03318_, _00072_, _00071_);
  or (_00073_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00074_, \oc8051_gm_cxrom_1.cell2.data [5], _00043_);
  nand (_00075_, _00074_, _00073_);
  nand (_00076_, _00075_, _42545_);
  or (_00077_, \oc8051_gm_cxrom_1.cell2.data [5], _42545_);
  and (_03321_, _00077_, _00076_);
  or (_00078_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00079_, \oc8051_gm_cxrom_1.cell2.data [6], _00043_);
  nand (_00080_, _00079_, _00078_);
  nand (_00081_, _00080_, _42545_);
  or (_00082_, \oc8051_gm_cxrom_1.cell2.data [6], _42545_);
  and (_03325_, _00082_, _00081_);
  or (_00083_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_00084_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_00085_, _00084_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_00086_, _00085_, _00083_);
  nand (_00087_, _00086_, _42545_);
  or (_00088_, \oc8051_gm_cxrom_1.cell3.data [7], _42545_);
  and (_03344_, _00088_, _00087_);
  or (_00089_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00090_, \oc8051_gm_cxrom_1.cell3.data [0], _00084_);
  nand (_00091_, _00090_, _00089_);
  nand (_00092_, _00091_, _42545_);
  or (_00093_, \oc8051_gm_cxrom_1.cell3.data [0], _42545_);
  and (_03350_, _00093_, _00092_);
  or (_00094_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00095_, \oc8051_gm_cxrom_1.cell3.data [1], _00084_);
  nand (_00096_, _00095_, _00094_);
  nand (_00097_, _00096_, _42545_);
  or (_00098_, \oc8051_gm_cxrom_1.cell3.data [1], _42545_);
  and (_03354_, _00098_, _00097_);
  or (_00099_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00100_, \oc8051_gm_cxrom_1.cell3.data [2], _00084_);
  nand (_00101_, _00100_, _00099_);
  nand (_00102_, _00101_, _42545_);
  or (_00103_, \oc8051_gm_cxrom_1.cell3.data [2], _42545_);
  and (_03357_, _00103_, _00102_);
  or (_00104_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00105_, \oc8051_gm_cxrom_1.cell3.data [3], _00084_);
  nand (_00106_, _00105_, _00104_);
  nand (_00107_, _00106_, _42545_);
  or (_00108_, \oc8051_gm_cxrom_1.cell3.data [3], _42545_);
  and (_03361_, _00108_, _00107_);
  or (_00109_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00110_, \oc8051_gm_cxrom_1.cell3.data [4], _00084_);
  nand (_00111_, _00110_, _00109_);
  nand (_00112_, _00111_, _42545_);
  or (_00113_, \oc8051_gm_cxrom_1.cell3.data [4], _42545_);
  and (_03364_, _00113_, _00112_);
  or (_00114_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00115_, \oc8051_gm_cxrom_1.cell3.data [5], _00084_);
  nand (_00116_, _00115_, _00114_);
  nand (_00117_, _00116_, _42545_);
  or (_00118_, \oc8051_gm_cxrom_1.cell3.data [5], _42545_);
  and (_03368_, _00118_, _00117_);
  or (_00119_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00120_, \oc8051_gm_cxrom_1.cell3.data [6], _00084_);
  nand (_00121_, _00120_, _00119_);
  nand (_00122_, _00121_, _42545_);
  or (_00123_, \oc8051_gm_cxrom_1.cell3.data [6], _42545_);
  and (_03373_, _00123_, _00122_);
  or (_00124_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_00125_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_00126_, _00125_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_00127_, _00126_, _00124_);
  nand (_00128_, _00127_, _42545_);
  or (_00129_, \oc8051_gm_cxrom_1.cell4.data [7], _42545_);
  and (_03391_, _00129_, _00128_);
  or (_00131_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00133_, \oc8051_gm_cxrom_1.cell4.data [0], _00125_);
  nand (_00135_, _00133_, _00131_);
  nand (_00137_, _00135_, _42545_);
  or (_00139_, \oc8051_gm_cxrom_1.cell4.data [0], _42545_);
  and (_03397_, _00139_, _00137_);
  or (_00142_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00144_, \oc8051_gm_cxrom_1.cell4.data [1], _00125_);
  nand (_00146_, _00144_, _00142_);
  nand (_00148_, _00146_, _42545_);
  or (_00150_, \oc8051_gm_cxrom_1.cell4.data [1], _42545_);
  and (_03400_, _00150_, _00148_);
  or (_00153_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00155_, \oc8051_gm_cxrom_1.cell4.data [2], _00125_);
  nand (_00157_, _00155_, _00153_);
  nand (_00159_, _00157_, _42545_);
  or (_00161_, \oc8051_gm_cxrom_1.cell4.data [2], _42545_);
  and (_03404_, _00161_, _00159_);
  or (_00164_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00166_, \oc8051_gm_cxrom_1.cell4.data [3], _00125_);
  nand (_00168_, _00166_, _00164_);
  nand (_00170_, _00168_, _42545_);
  or (_00172_, \oc8051_gm_cxrom_1.cell4.data [3], _42545_);
  and (_03407_, _00172_, _00170_);
  or (_00175_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00177_, \oc8051_gm_cxrom_1.cell4.data [4], _00125_);
  nand (_00179_, _00177_, _00175_);
  nand (_00181_, _00179_, _42545_);
  or (_00183_, \oc8051_gm_cxrom_1.cell4.data [4], _42545_);
  and (_03411_, _00183_, _00181_);
  or (_00186_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00187_, \oc8051_gm_cxrom_1.cell4.data [5], _00125_);
  nand (_00188_, _00187_, _00186_);
  nand (_00189_, _00188_, _42545_);
  or (_00190_, \oc8051_gm_cxrom_1.cell4.data [5], _42545_);
  and (_03415_, _00190_, _00189_);
  or (_00191_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00192_, \oc8051_gm_cxrom_1.cell4.data [6], _00125_);
  nand (_00193_, _00192_, _00191_);
  nand (_00194_, _00193_, _42545_);
  or (_00195_, \oc8051_gm_cxrom_1.cell4.data [6], _42545_);
  and (_03419_, _00195_, _00194_);
  or (_00196_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_00197_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_00198_, _00197_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_00199_, _00198_, _00196_);
  nand (_00200_, _00199_, _42545_);
  or (_00201_, \oc8051_gm_cxrom_1.cell5.data [7], _42545_);
  and (_03441_, _00201_, _00200_);
  or (_00202_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00203_, \oc8051_gm_cxrom_1.cell5.data [0], _00197_);
  nand (_00204_, _00203_, _00202_);
  nand (_00205_, _00204_, _42545_);
  or (_00206_, \oc8051_gm_cxrom_1.cell5.data [0], _42545_);
  and (_03448_, _00206_, _00205_);
  or (_00207_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00208_, \oc8051_gm_cxrom_1.cell5.data [1], _00197_);
  nand (_00209_, _00208_, _00207_);
  nand (_00210_, _00209_, _42545_);
  or (_00211_, \oc8051_gm_cxrom_1.cell5.data [1], _42545_);
  and (_03452_, _00211_, _00210_);
  or (_00212_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00213_, \oc8051_gm_cxrom_1.cell5.data [2], _00197_);
  nand (_00214_, _00213_, _00212_);
  nand (_00215_, _00214_, _42545_);
  or (_00216_, \oc8051_gm_cxrom_1.cell5.data [2], _42545_);
  and (_03456_, _00216_, _00215_);
  or (_00217_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00218_, \oc8051_gm_cxrom_1.cell5.data [3], _00197_);
  nand (_00219_, _00218_, _00217_);
  nand (_00220_, _00219_, _42545_);
  or (_00221_, \oc8051_gm_cxrom_1.cell5.data [3], _42545_);
  and (_03460_, _00221_, _00220_);
  or (_00222_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00223_, \oc8051_gm_cxrom_1.cell5.data [4], _00197_);
  nand (_00224_, _00223_, _00222_);
  nand (_00225_, _00224_, _42545_);
  or (_00226_, \oc8051_gm_cxrom_1.cell5.data [4], _42545_);
  and (_03464_, _00226_, _00225_);
  or (_00227_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00228_, \oc8051_gm_cxrom_1.cell5.data [5], _00197_);
  nand (_00229_, _00228_, _00227_);
  nand (_00230_, _00229_, _42545_);
  or (_00231_, \oc8051_gm_cxrom_1.cell5.data [5], _42545_);
  and (_03468_, _00231_, _00230_);
  or (_00232_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00233_, \oc8051_gm_cxrom_1.cell5.data [6], _00197_);
  nand (_00234_, _00233_, _00232_);
  nand (_00235_, _00234_, _42545_);
  or (_00236_, \oc8051_gm_cxrom_1.cell5.data [6], _42545_);
  and (_03472_, _00236_, _00235_);
  or (_00237_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_00238_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_00239_, _00238_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_00240_, _00239_, _00237_);
  nand (_00241_, _00240_, _42545_);
  or (_00242_, \oc8051_gm_cxrom_1.cell6.data [7], _42545_);
  and (_03494_, _00242_, _00241_);
  or (_00243_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00244_, \oc8051_gm_cxrom_1.cell6.data [0], _00238_);
  nand (_00245_, _00244_, _00243_);
  nand (_00246_, _00245_, _42545_);
  or (_00247_, \oc8051_gm_cxrom_1.cell6.data [0], _42545_);
  and (_03501_, _00247_, _00246_);
  or (_00248_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00249_, \oc8051_gm_cxrom_1.cell6.data [1], _00238_);
  nand (_00250_, _00249_, _00248_);
  nand (_00251_, _00250_, _42545_);
  or (_00252_, \oc8051_gm_cxrom_1.cell6.data [1], _42545_);
  and (_03505_, _00252_, _00251_);
  or (_00253_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00254_, \oc8051_gm_cxrom_1.cell6.data [2], _00238_);
  nand (_00255_, _00254_, _00253_);
  nand (_00256_, _00255_, _42545_);
  or (_00257_, \oc8051_gm_cxrom_1.cell6.data [2], _42545_);
  and (_03509_, _00257_, _00256_);
  or (_00258_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00259_, \oc8051_gm_cxrom_1.cell6.data [3], _00238_);
  nand (_00260_, _00259_, _00258_);
  nand (_00261_, _00260_, _42545_);
  or (_00262_, \oc8051_gm_cxrom_1.cell6.data [3], _42545_);
  and (_03513_, _00262_, _00261_);
  or (_00263_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00264_, \oc8051_gm_cxrom_1.cell6.data [4], _00238_);
  nand (_00265_, _00264_, _00263_);
  nand (_00266_, _00265_, _42545_);
  or (_00267_, \oc8051_gm_cxrom_1.cell6.data [4], _42545_);
  and (_03517_, _00267_, _00266_);
  or (_00268_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00269_, \oc8051_gm_cxrom_1.cell6.data [5], _00238_);
  nand (_00270_, _00269_, _00268_);
  nand (_00271_, _00270_, _42545_);
  or (_00272_, \oc8051_gm_cxrom_1.cell6.data [5], _42545_);
  and (_03521_, _00272_, _00271_);
  or (_00273_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00274_, \oc8051_gm_cxrom_1.cell6.data [6], _00238_);
  nand (_00275_, _00274_, _00273_);
  nand (_00276_, _00275_, _42545_);
  or (_00277_, \oc8051_gm_cxrom_1.cell6.data [6], _42545_);
  and (_03525_, _00277_, _00276_);
  or (_00278_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_00279_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_00280_, _00279_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_00281_, _00280_, _00278_);
  nand (_00282_, _00281_, _42545_);
  or (_00283_, \oc8051_gm_cxrom_1.cell7.data [7], _42545_);
  and (_03547_, _00283_, _00282_);
  or (_00284_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00285_, \oc8051_gm_cxrom_1.cell7.data [0], _00279_);
  nand (_00286_, _00285_, _00284_);
  nand (_00287_, _00286_, _42545_);
  or (_00288_, \oc8051_gm_cxrom_1.cell7.data [0], _42545_);
  and (_03554_, _00288_, _00287_);
  or (_00289_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00290_, \oc8051_gm_cxrom_1.cell7.data [1], _00279_);
  nand (_00291_, _00290_, _00289_);
  nand (_00292_, _00291_, _42545_);
  or (_00293_, \oc8051_gm_cxrom_1.cell7.data [1], _42545_);
  and (_03558_, _00293_, _00292_);
  or (_00294_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00295_, \oc8051_gm_cxrom_1.cell7.data [2], _00279_);
  nand (_00296_, _00295_, _00294_);
  nand (_00297_, _00296_, _42545_);
  or (_00298_, \oc8051_gm_cxrom_1.cell7.data [2], _42545_);
  and (_03562_, _00298_, _00297_);
  or (_00299_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00300_, \oc8051_gm_cxrom_1.cell7.data [3], _00279_);
  nand (_00301_, _00300_, _00299_);
  nand (_00302_, _00301_, _42545_);
  or (_00303_, \oc8051_gm_cxrom_1.cell7.data [3], _42545_);
  and (_03566_, _00303_, _00302_);
  or (_00304_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00305_, \oc8051_gm_cxrom_1.cell7.data [4], _00279_);
  nand (_00306_, _00305_, _00304_);
  nand (_00307_, _00306_, _42545_);
  or (_00308_, \oc8051_gm_cxrom_1.cell7.data [4], _42545_);
  and (_03570_, _00308_, _00307_);
  or (_00309_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00310_, \oc8051_gm_cxrom_1.cell7.data [5], _00279_);
  nand (_00311_, _00310_, _00309_);
  nand (_00312_, _00311_, _42545_);
  or (_00313_, \oc8051_gm_cxrom_1.cell7.data [5], _42545_);
  and (_03574_, _00313_, _00312_);
  or (_00314_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00315_, \oc8051_gm_cxrom_1.cell7.data [6], _00279_);
  nand (_00316_, _00315_, _00314_);
  nand (_00317_, _00316_, _42545_);
  or (_00318_, \oc8051_gm_cxrom_1.cell7.data [6], _42545_);
  and (_03578_, _00318_, _00317_);
  or (_00319_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_00320_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_00321_, _00320_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_00322_, _00321_, _00319_);
  nand (_00323_, _00322_, _42545_);
  or (_00324_, \oc8051_gm_cxrom_1.cell8.data [7], _42545_);
  and (_03600_, _00324_, _00323_);
  or (_00325_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00326_, \oc8051_gm_cxrom_1.cell8.data [0], _00320_);
  nand (_00327_, _00326_, _00325_);
  nand (_00328_, _00327_, _42545_);
  or (_00329_, \oc8051_gm_cxrom_1.cell8.data [0], _42545_);
  and (_03608_, _00329_, _00328_);
  or (_00330_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00331_, \oc8051_gm_cxrom_1.cell8.data [1], _00320_);
  nand (_00332_, _00331_, _00330_);
  nand (_00333_, _00332_, _42545_);
  or (_00334_, \oc8051_gm_cxrom_1.cell8.data [1], _42545_);
  and (_03612_, _00334_, _00333_);
  or (_00335_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00336_, \oc8051_gm_cxrom_1.cell8.data [2], _00320_);
  nand (_00337_, _00336_, _00335_);
  nand (_00338_, _00337_, _42545_);
  or (_00339_, \oc8051_gm_cxrom_1.cell8.data [2], _42545_);
  and (_03616_, _00339_, _00338_);
  or (_00340_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00341_, \oc8051_gm_cxrom_1.cell8.data [3], _00320_);
  nand (_00342_, _00341_, _00340_);
  nand (_00343_, _00342_, _42545_);
  or (_00344_, \oc8051_gm_cxrom_1.cell8.data [3], _42545_);
  and (_03620_, _00344_, _00343_);
  or (_00345_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00346_, \oc8051_gm_cxrom_1.cell8.data [4], _00320_);
  nand (_00347_, _00346_, _00345_);
  nand (_00348_, _00347_, _42545_);
  or (_00349_, \oc8051_gm_cxrom_1.cell8.data [4], _42545_);
  and (_03624_, _00349_, _00348_);
  or (_00350_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00351_, \oc8051_gm_cxrom_1.cell8.data [5], _00320_);
  nand (_00352_, _00351_, _00350_);
  nand (_00353_, _00352_, _42545_);
  or (_00354_, \oc8051_gm_cxrom_1.cell8.data [5], _42545_);
  and (_03628_, _00354_, _00353_);
  or (_00355_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00356_, \oc8051_gm_cxrom_1.cell8.data [6], _00320_);
  nand (_00357_, _00356_, _00355_);
  nand (_00358_, _00357_, _42545_);
  or (_00359_, \oc8051_gm_cxrom_1.cell8.data [6], _42545_);
  and (_03632_, _00359_, _00358_);
  or (_00360_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_00361_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_00362_, _00361_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_00363_, _00362_, _00360_);
  nand (_00364_, _00363_, _42545_);
  or (_00365_, \oc8051_gm_cxrom_1.cell9.data [7], _42545_);
  and (_03654_, _00365_, _00364_);
  or (_00366_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00367_, \oc8051_gm_cxrom_1.cell9.data [0], _00361_);
  nand (_00368_, _00367_, _00366_);
  nand (_00369_, _00368_, _42545_);
  or (_00370_, \oc8051_gm_cxrom_1.cell9.data [0], _42545_);
  and (_03661_, _00370_, _00369_);
  or (_00371_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00372_, \oc8051_gm_cxrom_1.cell9.data [1], _00361_);
  nand (_00373_, _00372_, _00371_);
  nand (_00374_, _00373_, _42545_);
  or (_00375_, \oc8051_gm_cxrom_1.cell9.data [1], _42545_);
  and (_03665_, _00375_, _00374_);
  or (_00376_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00377_, \oc8051_gm_cxrom_1.cell9.data [2], _00361_);
  nand (_00378_, _00377_, _00376_);
  nand (_00379_, _00378_, _42545_);
  or (_00380_, \oc8051_gm_cxrom_1.cell9.data [2], _42545_);
  and (_03669_, _00380_, _00379_);
  or (_00381_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00382_, \oc8051_gm_cxrom_1.cell9.data [3], _00361_);
  nand (_00383_, _00382_, _00381_);
  nand (_00384_, _00383_, _42545_);
  or (_00385_, \oc8051_gm_cxrom_1.cell9.data [3], _42545_);
  and (_03673_, _00385_, _00384_);
  or (_00386_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00387_, \oc8051_gm_cxrom_1.cell9.data [4], _00361_);
  nand (_00388_, _00387_, _00386_);
  nand (_00389_, _00388_, _42545_);
  or (_00390_, \oc8051_gm_cxrom_1.cell9.data [4], _42545_);
  and (_03677_, _00390_, _00389_);
  or (_00391_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00392_, \oc8051_gm_cxrom_1.cell9.data [5], _00361_);
  nand (_00393_, _00392_, _00391_);
  nand (_00394_, _00393_, _42545_);
  or (_00395_, \oc8051_gm_cxrom_1.cell9.data [5], _42545_);
  and (_03681_, _00395_, _00394_);
  or (_00396_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00397_, \oc8051_gm_cxrom_1.cell9.data [6], _00361_);
  nand (_00398_, _00397_, _00396_);
  nand (_00399_, _00398_, _42545_);
  or (_00400_, \oc8051_gm_cxrom_1.cell9.data [6], _42545_);
  and (_03685_, _00400_, _00399_);
  or (_00401_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_00402_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_00403_, _00402_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_00404_, _00403_, _00401_);
  nand (_00405_, _00404_, _42545_);
  or (_00406_, \oc8051_gm_cxrom_1.cell10.data [7], _42545_);
  and (_03707_, _00406_, _00405_);
  or (_00407_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00408_, \oc8051_gm_cxrom_1.cell10.data [0], _00402_);
  nand (_00409_, _00408_, _00407_);
  nand (_00410_, _00409_, _42545_);
  or (_00411_, \oc8051_gm_cxrom_1.cell10.data [0], _42545_);
  and (_03714_, _00411_, _00410_);
  or (_00412_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00413_, \oc8051_gm_cxrom_1.cell10.data [1], _00402_);
  nand (_00414_, _00413_, _00412_);
  nand (_00415_, _00414_, _42545_);
  or (_00416_, \oc8051_gm_cxrom_1.cell10.data [1], _42545_);
  and (_03718_, _00416_, _00415_);
  or (_00417_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00418_, \oc8051_gm_cxrom_1.cell10.data [2], _00402_);
  nand (_00419_, _00418_, _00417_);
  nand (_00420_, _00419_, _42545_);
  or (_00421_, \oc8051_gm_cxrom_1.cell10.data [2], _42545_);
  and (_03722_, _00421_, _00420_);
  or (_00422_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00423_, \oc8051_gm_cxrom_1.cell10.data [3], _00402_);
  nand (_00424_, _00423_, _00422_);
  nand (_00425_, _00424_, _42545_);
  or (_00426_, \oc8051_gm_cxrom_1.cell10.data [3], _42545_);
  and (_03726_, _00426_, _00425_);
  or (_00427_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00428_, \oc8051_gm_cxrom_1.cell10.data [4], _00402_);
  nand (_00429_, _00428_, _00427_);
  nand (_00430_, _00429_, _42545_);
  or (_00431_, \oc8051_gm_cxrom_1.cell10.data [4], _42545_);
  and (_03730_, _00431_, _00430_);
  or (_00432_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00433_, \oc8051_gm_cxrom_1.cell10.data [5], _00402_);
  nand (_00434_, _00433_, _00432_);
  nand (_00435_, _00434_, _42545_);
  or (_00436_, \oc8051_gm_cxrom_1.cell10.data [5], _42545_);
  and (_03734_, _00436_, _00435_);
  or (_00437_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00438_, \oc8051_gm_cxrom_1.cell10.data [6], _00402_);
  nand (_00439_, _00438_, _00437_);
  nand (_00440_, _00439_, _42545_);
  or (_00441_, \oc8051_gm_cxrom_1.cell10.data [6], _42545_);
  and (_03738_, _00441_, _00440_);
  or (_00442_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_00443_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_00444_, _00443_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_00445_, _00444_, _00442_);
  nand (_00446_, _00445_, _42545_);
  or (_00447_, \oc8051_gm_cxrom_1.cell11.data [7], _42545_);
  and (_03760_, _00447_, _00446_);
  or (_00448_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00449_, \oc8051_gm_cxrom_1.cell11.data [0], _00443_);
  nand (_00450_, _00449_, _00448_);
  nand (_00451_, _00450_, _42545_);
  or (_00452_, \oc8051_gm_cxrom_1.cell11.data [0], _42545_);
  and (_03767_, _00452_, _00451_);
  or (_00453_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00454_, \oc8051_gm_cxrom_1.cell11.data [1], _00443_);
  nand (_00455_, _00454_, _00453_);
  nand (_00456_, _00455_, _42545_);
  or (_00457_, \oc8051_gm_cxrom_1.cell11.data [1], _42545_);
  and (_03771_, _00457_, _00456_);
  or (_00458_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00459_, \oc8051_gm_cxrom_1.cell11.data [2], _00443_);
  nand (_00460_, _00459_, _00458_);
  nand (_00461_, _00460_, _42545_);
  or (_00462_, \oc8051_gm_cxrom_1.cell11.data [2], _42545_);
  and (_03775_, _00462_, _00461_);
  or (_00463_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00464_, \oc8051_gm_cxrom_1.cell11.data [3], _00443_);
  nand (_00465_, _00464_, _00463_);
  nand (_00466_, _00465_, _42545_);
  or (_00467_, \oc8051_gm_cxrom_1.cell11.data [3], _42545_);
  and (_03779_, _00467_, _00466_);
  or (_00468_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00469_, \oc8051_gm_cxrom_1.cell11.data [4], _00443_);
  nand (_00470_, _00469_, _00468_);
  nand (_00471_, _00470_, _42545_);
  or (_00472_, \oc8051_gm_cxrom_1.cell11.data [4], _42545_);
  and (_03783_, _00472_, _00471_);
  or (_00473_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00474_, \oc8051_gm_cxrom_1.cell11.data [5], _00443_);
  nand (_00475_, _00474_, _00473_);
  nand (_00476_, _00475_, _42545_);
  or (_00477_, \oc8051_gm_cxrom_1.cell11.data [5], _42545_);
  and (_03787_, _00477_, _00476_);
  or (_00478_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00479_, \oc8051_gm_cxrom_1.cell11.data [6], _00443_);
  nand (_00480_, _00479_, _00478_);
  nand (_00481_, _00480_, _42545_);
  or (_00482_, \oc8051_gm_cxrom_1.cell11.data [6], _42545_);
  and (_03791_, _00482_, _00481_);
  or (_00483_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_00484_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_00485_, _00484_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_00486_, _00485_, _00483_);
  nand (_00487_, _00486_, _42545_);
  or (_00488_, \oc8051_gm_cxrom_1.cell12.data [7], _42545_);
  and (_03813_, _00488_, _00487_);
  or (_00489_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00490_, \oc8051_gm_cxrom_1.cell12.data [0], _00484_);
  nand (_00491_, _00490_, _00489_);
  nand (_00492_, _00491_, _42545_);
  or (_00493_, \oc8051_gm_cxrom_1.cell12.data [0], _42545_);
  and (_03820_, _00493_, _00492_);
  or (_00494_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00495_, \oc8051_gm_cxrom_1.cell12.data [1], _00484_);
  nand (_00496_, _00495_, _00494_);
  nand (_00497_, _00496_, _42545_);
  or (_00498_, \oc8051_gm_cxrom_1.cell12.data [1], _42545_);
  and (_03824_, _00498_, _00497_);
  or (_00499_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00500_, \oc8051_gm_cxrom_1.cell12.data [2], _00484_);
  nand (_00501_, _00500_, _00499_);
  nand (_00502_, _00501_, _42545_);
  or (_00503_, \oc8051_gm_cxrom_1.cell12.data [2], _42545_);
  and (_03828_, _00503_, _00502_);
  or (_00504_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00505_, \oc8051_gm_cxrom_1.cell12.data [3], _00484_);
  nand (_00506_, _00505_, _00504_);
  nand (_00507_, _00506_, _42545_);
  or (_00508_, \oc8051_gm_cxrom_1.cell12.data [3], _42545_);
  and (_03832_, _00508_, _00507_);
  or (_00509_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00510_, \oc8051_gm_cxrom_1.cell12.data [4], _00484_);
  nand (_00511_, _00510_, _00509_);
  nand (_00512_, _00511_, _42545_);
  or (_00513_, \oc8051_gm_cxrom_1.cell12.data [4], _42545_);
  and (_03836_, _00513_, _00512_);
  or (_00514_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00515_, \oc8051_gm_cxrom_1.cell12.data [5], _00484_);
  nand (_00516_, _00515_, _00514_);
  nand (_00517_, _00516_, _42545_);
  or (_00518_, \oc8051_gm_cxrom_1.cell12.data [5], _42545_);
  and (_03840_, _00518_, _00517_);
  or (_00519_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00520_, \oc8051_gm_cxrom_1.cell12.data [6], _00484_);
  nand (_00521_, _00520_, _00519_);
  nand (_00522_, _00521_, _42545_);
  or (_00523_, \oc8051_gm_cxrom_1.cell12.data [6], _42545_);
  and (_03844_, _00523_, _00522_);
  or (_00524_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_00525_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_00526_, _00525_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_00527_, _00526_, _00524_);
  nand (_00528_, _00527_, _42545_);
  or (_00529_, \oc8051_gm_cxrom_1.cell13.data [7], _42545_);
  and (_03867_, _00529_, _00528_);
  or (_00530_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00531_, \oc8051_gm_cxrom_1.cell13.data [0], _00525_);
  nand (_00532_, _00531_, _00530_);
  nand (_00533_, _00532_, _42545_);
  or (_00534_, \oc8051_gm_cxrom_1.cell13.data [0], _42545_);
  and (_03874_, _00534_, _00533_);
  or (_00535_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00536_, \oc8051_gm_cxrom_1.cell13.data [1], _00525_);
  nand (_00537_, _00536_, _00535_);
  nand (_00538_, _00537_, _42545_);
  or (_00539_, \oc8051_gm_cxrom_1.cell13.data [1], _42545_);
  and (_03878_, _00539_, _00538_);
  or (_00540_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00541_, \oc8051_gm_cxrom_1.cell13.data [2], _00525_);
  nand (_00542_, _00541_, _00540_);
  nand (_00544_, _00542_, _42545_);
  or (_00545_, \oc8051_gm_cxrom_1.cell13.data [2], _42545_);
  and (_03882_, _00545_, _00544_);
  or (_00547_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00549_, \oc8051_gm_cxrom_1.cell13.data [3], _00525_);
  nand (_00550_, _00549_, _00547_);
  nand (_00552_, _00550_, _42545_);
  or (_00553_, \oc8051_gm_cxrom_1.cell13.data [3], _42545_);
  and (_03886_, _00553_, _00552_);
  or (_00555_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00557_, \oc8051_gm_cxrom_1.cell13.data [4], _00525_);
  nand (_00558_, _00557_, _00555_);
  nand (_00560_, _00558_, _42545_);
  or (_00561_, \oc8051_gm_cxrom_1.cell13.data [4], _42545_);
  and (_03890_, _00561_, _00560_);
  or (_00563_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00565_, \oc8051_gm_cxrom_1.cell13.data [5], _00525_);
  nand (_00566_, _00565_, _00563_);
  nand (_00568_, _00566_, _42545_);
  or (_00569_, \oc8051_gm_cxrom_1.cell13.data [5], _42545_);
  and (_03894_, _00569_, _00568_);
  or (_00571_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00573_, \oc8051_gm_cxrom_1.cell13.data [6], _00525_);
  nand (_00574_, _00573_, _00571_);
  nand (_00576_, _00574_, _42545_);
  or (_00577_, \oc8051_gm_cxrom_1.cell13.data [6], _42545_);
  and (_03898_, _00577_, _00576_);
  or (_00579_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_00581_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_00582_, _00581_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_00584_, _00582_, _00579_);
  nand (_00585_, _00584_, _42545_);
  or (_00587_, \oc8051_gm_cxrom_1.cell14.data [7], _42545_);
  and (_03920_, _00587_, _00585_);
  or (_00589_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00590_, \oc8051_gm_cxrom_1.cell14.data [0], _00581_);
  nand (_00592_, _00590_, _00589_);
  nand (_00593_, _00592_, _42545_);
  or (_00594_, \oc8051_gm_cxrom_1.cell14.data [0], _42545_);
  and (_03927_, _00594_, _00593_);
  or (_00595_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00596_, \oc8051_gm_cxrom_1.cell14.data [1], _00581_);
  nand (_00597_, _00596_, _00595_);
  nand (_00598_, _00597_, _42545_);
  or (_00599_, \oc8051_gm_cxrom_1.cell14.data [1], _42545_);
  and (_03931_, _00599_, _00598_);
  or (_00600_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00601_, \oc8051_gm_cxrom_1.cell14.data [2], _00581_);
  nand (_00602_, _00601_, _00600_);
  nand (_00603_, _00602_, _42545_);
  or (_00604_, \oc8051_gm_cxrom_1.cell14.data [2], _42545_);
  and (_03934_, _00604_, _00603_);
  or (_00605_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00606_, \oc8051_gm_cxrom_1.cell14.data [3], _00581_);
  nand (_00607_, _00606_, _00605_);
  nand (_00608_, _00607_, _42545_);
  or (_00609_, \oc8051_gm_cxrom_1.cell14.data [3], _42545_);
  and (_03938_, _00609_, _00608_);
  or (_00610_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00611_, \oc8051_gm_cxrom_1.cell14.data [4], _00581_);
  nand (_00612_, _00611_, _00610_);
  nand (_00613_, _00612_, _42545_);
  or (_00614_, \oc8051_gm_cxrom_1.cell14.data [4], _42545_);
  and (_03942_, _00614_, _00613_);
  or (_00615_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00616_, \oc8051_gm_cxrom_1.cell14.data [5], _00581_);
  nand (_00617_, _00616_, _00615_);
  nand (_00618_, _00617_, _42545_);
  or (_00619_, \oc8051_gm_cxrom_1.cell14.data [5], _42545_);
  and (_03946_, _00619_, _00618_);
  or (_00620_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00621_, \oc8051_gm_cxrom_1.cell14.data [6], _00581_);
  nand (_00622_, _00621_, _00620_);
  nand (_00623_, _00622_, _42545_);
  or (_00624_, \oc8051_gm_cxrom_1.cell14.data [6], _42545_);
  and (_03950_, _00624_, _00623_);
  or (_00625_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_00626_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_00627_, _00626_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_00628_, _00627_, _00625_);
  nand (_00629_, _00628_, _42545_);
  or (_00630_, \oc8051_gm_cxrom_1.cell15.data [7], _42545_);
  and (_03971_, _00630_, _00629_);
  or (_00631_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00632_, \oc8051_gm_cxrom_1.cell15.data [0], _00626_);
  nand (_00633_, _00632_, _00631_);
  nand (_00634_, _00633_, _42545_);
  or (_00635_, \oc8051_gm_cxrom_1.cell15.data [0], _42545_);
  and (_03978_, _00635_, _00634_);
  or (_00636_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00637_, \oc8051_gm_cxrom_1.cell15.data [1], _00626_);
  nand (_00638_, _00637_, _00636_);
  nand (_00639_, _00638_, _42545_);
  or (_00640_, \oc8051_gm_cxrom_1.cell15.data [1], _42545_);
  and (_03982_, _00640_, _00639_);
  or (_00641_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00642_, \oc8051_gm_cxrom_1.cell15.data [2], _00626_);
  nand (_00643_, _00642_, _00641_);
  nand (_00644_, _00643_, _42545_);
  or (_00645_, \oc8051_gm_cxrom_1.cell15.data [2], _42545_);
  and (_03986_, _00645_, _00644_);
  or (_00646_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00647_, \oc8051_gm_cxrom_1.cell15.data [3], _00626_);
  nand (_00648_, _00647_, _00646_);
  nand (_00649_, _00648_, _42545_);
  or (_00650_, \oc8051_gm_cxrom_1.cell15.data [3], _42545_);
  and (_03990_, _00650_, _00649_);
  or (_00651_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00652_, \oc8051_gm_cxrom_1.cell15.data [4], _00626_);
  nand (_00653_, _00652_, _00651_);
  nand (_00654_, _00653_, _42545_);
  or (_00655_, \oc8051_gm_cxrom_1.cell15.data [4], _42545_);
  and (_03994_, _00655_, _00654_);
  or (_00656_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00657_, \oc8051_gm_cxrom_1.cell15.data [5], _00626_);
  nand (_00658_, _00657_, _00656_);
  nand (_00659_, _00658_, _42545_);
  or (_00660_, \oc8051_gm_cxrom_1.cell15.data [5], _42545_);
  and (_03998_, _00660_, _00659_);
  or (_00661_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00662_, \oc8051_gm_cxrom_1.cell15.data [6], _00626_);
  nand (_00663_, _00662_, _00661_);
  nand (_00664_, _00663_, _42545_);
  or (_00665_, \oc8051_gm_cxrom_1.cell15.data [6], _42545_);
  and (_04002_, _00665_, _00664_);
  nor (_07729_, _37919_, rst);
  and (_00666_, _36955_, _42545_);
  nand (_00667_, _00666_, _37965_);
  nor (_00668_, _37908_, _37882_);
  or (_07732_, _00668_, _00667_);
  not (_00669_, _37779_);
  nor (_00670_, _00669_, _37600_);
  not (_00671_, _37327_);
  not (_00672_, _37875_);
  and (_00673_, _00672_, _37852_);
  not (_00674_, _37828_);
  and (_00675_, _00674_, _37804_);
  and (_00676_, _00675_, _00673_);
  and (_00677_, _00676_, _00671_);
  and (_00678_, _00677_, _00670_);
  not (_00679_, _37600_);
  not (_00680_, _37755_);
  and (_00681_, _37779_, _00680_);
  and (_00682_, _00681_, _00679_);
  and (_00683_, _00673_, _37828_);
  and (_00684_, _00683_, _37327_);
  and (_00685_, _00684_, _00682_);
  nor (_00686_, _00671_, _37852_);
  and (_00687_, _00686_, _00681_);
  and (_00688_, _00687_, _00679_);
  or (_00689_, _00688_, _00685_);
  and (_00690_, _00673_, _00674_);
  nor (_00691_, _37755_, _00671_);
  and (_00692_, _00691_, _00670_);
  and (_00693_, _00692_, _00690_);
  and (_00694_, _37875_, _37852_);
  and (_00695_, _00694_, _00675_);
  nor (_00696_, _37779_, _37600_);
  and (_00697_, _00696_, _00680_);
  and (_00698_, _00697_, _00695_);
  nor (_00699_, _00698_, _00693_);
  and (_00700_, _00696_, _37755_);
  and (_00701_, _00700_, _00686_);
  and (_00702_, _00669_, _37600_);
  and (_00703_, _00702_, _37327_);
  and (_00704_, _00703_, _00695_);
  nor (_00705_, _00704_, _00701_);
  nand (_00706_, _00705_, _00699_);
  or (_00707_, _00706_, _00689_);
  or (_00708_, _00707_, _00678_);
  not (_00709_, _37804_);
  nor (_00710_, _37755_, _37327_);
  and (_00711_, _00702_, _00710_);
  nor (_00712_, _00711_, _00709_);
  and (_00713_, _00694_, _00674_);
  not (_00714_, _00713_);
  nor (_00715_, _00714_, _00712_);
  not (_00716_, _00715_);
  and (_00717_, _37779_, _37600_);
  and (_00718_, _00717_, _00691_);
  and (_00719_, _00718_, _00695_);
  and (_00720_, _37755_, _00671_);
  and (_00721_, _00702_, _00720_);
  and (_00722_, _00721_, _00695_);
  nor (_00723_, _00722_, _00719_);
  and (_00724_, _00723_, _00716_);
  and (_00725_, _00702_, _00691_);
  and (_00726_, _00694_, _37828_);
  and (_00727_, _00726_, _00709_);
  and (_00728_, _00727_, _00725_);
  and (_00729_, _37755_, _37327_);
  or (_00730_, _00729_, _00710_);
  and (_00731_, _00717_, _00695_);
  and (_00732_, _00731_, _00730_);
  or (_00733_, _00732_, _00728_);
  and (_00734_, _00670_, _37755_);
  and (_00735_, _00727_, _00734_);
  and (_00736_, _00726_, _37804_);
  and (_00737_, _00717_, _37755_);
  and (_00738_, _00737_, _00736_);
  or (_00739_, _00738_, _00735_);
  or (_00740_, _00739_, _00733_);
  and (_00741_, _00729_, _00696_);
  and (_00742_, _00690_, _00709_);
  and (_00743_, _00742_, _00741_);
  and (_00744_, _00717_, _00680_);
  and (_00745_, _00736_, _00744_);
  or (_00746_, _00745_, _00743_);
  and (_00747_, _00720_, _00670_);
  and (_00748_, _00695_, _00747_);
  and (_00749_, _00726_, _00697_);
  or (_00750_, _00749_, _00748_);
  or (_00751_, _00750_, _00746_);
  nor (_00752_, _00751_, _00740_);
  nand (_00753_, _00752_, _00724_);
  or (_00754_, _00753_, _00708_);
  and (_00755_, _00754_, _36966_);
  not (_00756_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_00757_, _36944_, _18770_);
  and (_00758_, _00757_, _37909_);
  nor (_00759_, _00758_, _00756_);
  or (_00760_, _00759_, rst);
  or (_07735_, _00760_, _00755_);
  nand (_00761_, _37600_, _36890_);
  or (_00762_, _36890_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_00763_, _00762_, _42545_);
  and (_07738_, _00763_, _00761_);
  and (_00764_, \oc8051_top_1.oc8051_sfr1.wait_data , _42545_);
  and (_00765_, _00764_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00766_, _37908_, _37907_);
  or (_00767_, _00766_, _37985_);
  and (_00768_, _37883_, _37943_);
  and (_00769_, _37908_, _37896_);
  and (_00770_, _37974_, _37882_);
  or (_00771_, _00770_, _00769_);
  or (_00772_, _00771_, _00768_);
  or (_00773_, _00772_, _00767_);
  not (_00774_, _37962_);
  and (_00775_, _37900_, _37966_);
  and (_00776_, _37883_, _37887_);
  and (_00777_, _00776_, _37403_);
  or (_00778_, _00777_, _00775_);
  or (_00779_, _00778_, _00774_);
  or (_00780_, _00779_, _00773_);
  and (_00781_, _00780_, _00666_);
  or (_07741_, _00781_, _00765_);
  and (_00782_, _37908_, _37888_);
  or (_00783_, _00782_, _37884_);
  and (_00784_, _37403_, _37857_);
  and (_00785_, _00784_, _37942_);
  or (_00786_, _00785_, _38040_);
  and (_00787_, _37898_, _37926_);
  and (_00788_, _00787_, _37943_);
  or (_00789_, _00788_, _00786_);
  or (_00790_, _00789_, _00783_);
  and (_00791_, _00790_, _36955_);
  and (_00792_, _38011_, _00756_);
  not (_00793_, _37903_);
  and (_00794_, _00793_, _00792_);
  and (_00795_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00796_, _00795_, _00794_);
  or (_00797_, _00796_, _00791_);
  and (_07744_, _00797_, _42545_);
  and (_00798_, _00764_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nor (_00799_, _37974_, _37968_);
  nor (_00800_, _00799_, _37897_);
  and (_00801_, _37392_, _37857_);
  and (_00802_, _00801_, _37958_);
  or (_00803_, _00802_, _00800_);
  or (_00804_, _00803_, _38028_);
  and (_00805_, _37900_, _37968_);
  nor (_00806_, _00799_, _37996_);
  or (_00807_, _00806_, _00805_);
  and (_00808_, _00787_, _37959_);
  or (_00809_, _00808_, _00807_);
  not (_00810_, _37900_);
  nor (_00811_, _00810_, _37997_);
  and (_00812_, _37983_, _37857_);
  or (_00813_, _00812_, _00783_);
  or (_00814_, _00813_, _00811_);
  or (_00815_, _00814_, _00809_);
  or (_00816_, _00815_, _00804_);
  and (_00817_, _00816_, _00666_);
  or (_07747_, _00817_, _00798_);
  and (_00818_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00819_, _37929_, _36955_);
  or (_00820_, _00819_, _00818_);
  or (_00821_, _00820_, _00794_);
  and (_07750_, _00821_, _42545_);
  and (_00822_, _37959_, _37924_);
  and (_00823_, _37927_, _37881_);
  and (_00824_, _00823_, _37392_);
  or (_00825_, _00824_, _00822_);
  or (_00826_, _00825_, _00777_);
  and (_00827_, _00825_, _37911_);
  or (_00828_, _00827_, _36901_);
  and (_00829_, _00828_, _00826_);
  and (_00830_, _37966_, _37908_);
  and (_00831_, _37966_, _37882_);
  or (_00832_, _00831_, _00830_);
  or (_00833_, _00832_, _00776_);
  and (_00834_, _00833_, _00792_);
  or (_00835_, _00834_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00836_, _00835_, _00829_);
  or (_00837_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18770_);
  and (_00838_, _00837_, _42545_);
  and (_07753_, _00838_, _00836_);
  and (_00839_, _00764_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_00840_, _00770_, _38003_);
  and (_00841_, _38030_, _37942_);
  or (_00842_, _00808_, _00841_);
  or (_00843_, _00842_, _00840_);
  or (_00844_, _00785_, _37944_);
  and (_00845_, _38021_, _37958_);
  or (_00846_, _00845_, _37984_);
  or (_00847_, _00846_, _00844_);
  and (_00848_, _00801_, _37942_);
  or (_00849_, _00802_, _00848_);
  or (_00850_, _37884_, _37975_);
  or (_00851_, _00850_, _00849_);
  or (_00852_, _00851_, _00847_);
  or (_00853_, _00852_, _00843_);
  and (_00854_, _00853_, _00666_);
  or (_07756_, _00854_, _00839_);
  and (_00855_, _00764_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  not (_00856_, _37989_);
  and (_00857_, _37900_, _37979_);
  or (_00858_, _00857_, _00856_);
  or (_00859_, _38036_, _38032_);
  and (_00860_, _38040_, _37392_);
  or (_00861_, _00860_, _00859_);
  or (_00862_, _00861_, _00803_);
  or (_00863_, _00862_, _00858_);
  nor (_00864_, _38026_, _37992_);
  nand (_00865_, _00864_, _37981_);
  and (_00866_, _00787_, _37939_);
  or (_00867_, _00866_, _00788_);
  and (_00868_, _00784_, _37941_);
  and (_00869_, _00784_, _37891_);
  or (_00870_, _00869_, _00868_);
  and (_00871_, _37883_, _37931_);
  or (_00872_, _00871_, _00870_);
  or (_00873_, _00872_, _00867_);
  or (_00874_, _00873_, _00865_);
  or (_00875_, _00874_, _00809_);
  or (_00876_, _00875_, _00863_);
  and (_00877_, _00876_, _00666_);
  or (_07759_, _00877_, _00855_);
  and (_00878_, _00787_, _37932_);
  or (_00879_, _00878_, _38041_);
  and (_00880_, _00801_, _37886_);
  and (_00881_, _00880_, _37655_);
  or (_00882_, _00881_, _38023_);
  and (_00883_, _37932_, _37857_);
  or (_00884_, _00883_, _00882_);
  or (_00885_, _00884_, _00879_);
  and (_00886_, _00787_, _37888_);
  or (_00887_, _00886_, _00885_);
  and (_00888_, _00887_, _36955_);
  nand (_00889_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_00890_, _00889_, _37916_);
  or (_00891_, _00890_, _00888_);
  and (_07762_, _00891_, _42545_);
  or (_00892_, _38002_, _37944_);
  or (_00893_, _00806_, _37995_);
  or (_00894_, _00893_, _00892_);
  and (_00895_, _37890_, _37392_);
  and (_00896_, _00895_, _37928_);
  or (_00897_, _00896_, _37976_);
  or (_00898_, _00822_, _37988_);
  or (_00899_, _00898_, _00897_);
  nand (_00900_, _37986_, _37930_);
  or (_00901_, _00900_, _00899_);
  or (_00902_, _00901_, _00894_);
  and (_00903_, _00784_, _37887_);
  or (_00904_, _00903_, _00824_);
  and (_00905_, _38021_, _37890_);
  or (_00906_, _00905_, _38026_);
  or (_00907_, _00906_, _37936_);
  and (_00908_, _00801_, _37890_);
  or (_00909_, _00908_, _38035_);
  or (_00910_, _00909_, _00907_);
  or (_00911_, _00910_, _00904_);
  or (_00912_, _37963_, _37949_);
  or (_00913_, _00912_, _00786_);
  or (_00914_, _00913_, _00803_);
  or (_00915_, _00914_, _00911_);
  or (_00916_, _00915_, _00902_);
  and (_00917_, _00916_, _36955_);
  and (_00918_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00919_, _00827_, _00794_);
  and (_00920_, _37911_, _37960_);
  or (_00921_, _00920_, _00919_);
  or (_00922_, _00921_, _00918_);
  or (_00923_, _00922_, _00917_);
  and (_07765_, _00923_, _42545_);
  nor (_07824_, _38051_, rst);
  nor (_07826_, _38016_, rst);
  nand (_07829_, _00833_, _00666_);
  nand (_00924_, _00666_, _00776_);
  not (_00926_, _37908_);
  or (_00927_, _00667_, _00926_);
  and (_07832_, _00927_, _00924_);
  or (_00928_, _00735_, _00678_);
  or (_00929_, _00928_, _00745_);
  or (_00930_, _00929_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_00931_, _00930_, _00758_);
  nor (_00932_, _00757_, _37909_);
  or (_00933_, _00932_, rst);
  or (_07835_, _00933_, _00931_);
  nand (_00934_, _37804_, _36890_);
  or (_00935_, _36890_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_00936_, _00935_, _42545_);
  and (_07838_, _00936_, _00934_);
  not (_00937_, _36890_);
  or (_00938_, _37828_, _00937_);
  or (_00939_, _36890_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_00940_, _00939_, _42545_);
  and (_07841_, _00940_, _00938_);
  nand (_00941_, _37875_, _36890_);
  or (_00942_, _36890_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_00943_, _00942_, _42545_);
  and (_07844_, _00943_, _00941_);
  nand (_00944_, _37852_, _36890_);
  or (_00945_, _36890_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_00946_, _00945_, _42545_);
  and (_07847_, _00946_, _00944_);
  or (_00947_, _37327_, _00937_);
  or (_00948_, _36890_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_00949_, _00948_, _42545_);
  and (_07850_, _00949_, _00947_);
  nand (_00951_, _37755_, _36890_);
  or (_00952_, _36890_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_00953_, _00952_, _42545_);
  and (_07853_, _00953_, _00951_);
  nand (_00954_, _37779_, _36890_);
  or (_00955_, _36890_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_00956_, _00955_, _42545_);
  and (_07856_, _00956_, _00954_);
  or (_00957_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _18770_);
  and (_00958_, _00957_, _42545_);
  and (_00959_, _00958_, _00835_);
  and (_00960_, _37948_, _37857_);
  or (_00961_, _00960_, _00883_);
  or (_00962_, _00961_, _00882_);
  and (_00963_, _00787_, _37979_);
  or (_00964_, _00963_, _00782_);
  or (_00965_, _37974_, _37958_);
  and (_00966_, _00965_, _37900_);
  or (_00967_, _00966_, _00964_);
  or (_00969_, _00967_, _00962_);
  or (_00970_, _00879_, _37884_);
  or (_00971_, _38036_, _37967_);
  or (_00972_, _00971_, _00970_);
  and (_00973_, _00784_, _37965_);
  and (_00974_, _00784_, _37947_);
  or (_00975_, _00974_, _00869_);
  nor (_00976_, _00975_, _00973_);
  nand (_00977_, _00976_, _38034_);
  or (_00978_, _00977_, _00972_);
  and (_00979_, _37900_, _37892_);
  and (_00980_, _37948_, _37935_);
  or (_00981_, _00980_, _00979_);
  and (_00982_, _37965_, _37392_);
  and (_00983_, _00982_, _37900_);
  and (_00984_, _00787_, _37948_);
  or (_00985_, _00984_, _00983_);
  or (_00986_, _00985_, _00981_);
  or (_00987_, _00866_, _00775_);
  or (_00988_, _00886_, _00871_);
  or (_00989_, _00988_, _00987_);
  or (_00990_, _00989_, _00986_);
  or (_00991_, _00990_, _00978_);
  or (_00992_, _00991_, _00969_);
  and (_00993_, _00992_, _00666_);
  or (_07859_, _00993_, _00959_);
  and (_00994_, _00764_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor (_00995_, _00810_, _38000_);
  and (_00996_, _00801_, _37784_);
  and (_00997_, _00996_, _37655_);
  nor (_00998_, _00997_, _38025_);
  not (_00999_, _00998_);
  or (_01000_, _00999_, _00964_);
  or (_01001_, _01000_, _00995_);
  and (_01002_, _37900_, _37939_);
  and (_01003_, _37907_, _37403_);
  and (_01004_, _01003_, _37924_);
  or (_01005_, _01004_, _00870_);
  or (_01006_, _01005_, _01002_);
  not (_01007_, _37945_);
  or (_01008_, _00811_, _01007_);
  or (_01009_, _01008_, _01006_);
  or (_01010_, _00861_, _00778_);
  or (_01011_, _01010_, _01009_);
  or (_01012_, _01011_, _01001_);
  and (_01013_, _01012_, _00666_);
  or (_32090_, _01013_, _00994_);
  or (_01014_, _38035_, _37949_);
  or (_01015_, _01014_, _00904_);
  or (_01016_, _01015_, _00902_);
  and (_01017_, _01016_, _36955_);
  and (_01018_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01019_, _01018_, _00921_);
  or (_01020_, _01019_, _01017_);
  and (_32091_, _01020_, _42545_);
  and (_01021_, _37993_, _37403_);
  or (_01022_, _01021_, _38040_);
  or (_01023_, _01022_, _00907_);
  or (_01024_, _01023_, _00825_);
  and (_01025_, _01024_, _36955_);
  and (_01026_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01027_, _01026_, _00919_);
  or (_01028_, _01027_, _01025_);
  and (_32094_, _01028_, _42545_);
  or (_01029_, _00961_, _00871_);
  or (_01030_, _00882_, _38022_);
  or (_01031_, _37902_, _00776_);
  and (_01032_, _00878_, _37392_);
  or (_01033_, _01032_, _00984_);
  or (_01034_, _01033_, _01031_);
  or (_01035_, _01034_, _01030_);
  or (_01036_, _01035_, _01029_);
  or (_01037_, _00886_, _37901_);
  and (_01038_, _37900_, _37943_);
  or (_01039_, _00983_, _01038_);
  or (_01040_, _01039_, _01037_);
  and (_01041_, _00787_, _37983_);
  or (_01042_, _01041_, _00775_);
  or (_01043_, _01042_, _00966_);
  or (_01044_, _01043_, _01040_);
  or (_01045_, _00908_, _38041_);
  or (_01046_, _01045_, _00905_);
  or (_01047_, _00979_, _00857_);
  and (_01048_, _37883_, _37892_);
  or (_01049_, _01002_, _01048_);
  or (_01050_, _01049_, _01047_);
  or (_01051_, _01050_, _01046_);
  and (_01052_, _37948_, _37924_);
  and (_01053_, _00982_, _37928_);
  and (_01054_, _00878_, _37403_);
  or (_01055_, _01054_, _01053_);
  or (_01056_, _01055_, _01052_);
  or (_01057_, _01056_, _00825_);
  or (_01058_, _01057_, _01051_);
  or (_01059_, _01058_, _01044_);
  or (_01060_, _01059_, _01036_);
  and (_01061_, _01060_, _36955_);
  and (_01062_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_01063_, _37903_, _36901_);
  or (_01064_, _00834_, _01063_);
  or (_01065_, _01064_, _01062_);
  or (_01066_, _01065_, _01061_);
  and (_32096_, _01066_, _42545_);
  or (_01067_, _37902_, _37949_);
  and (_01068_, _37883_, _37939_);
  or (_01069_, _01068_, _00782_);
  or (_01070_, _01069_, _01067_);
  or (_01071_, _01070_, _01030_);
  or (_01072_, _01071_, _01029_);
  and (_01073_, _38021_, _37965_);
  and (_01074_, _00801_, _37965_);
  or (_01075_, _01074_, _01073_);
  or (_01076_, _00896_, _38041_);
  or (_01077_, _01076_, _01075_);
  or (_01078_, _01077_, _37894_);
  and (_01079_, _37988_, _37809_);
  or (_01080_, _01079_, _38001_);
  or (_01081_, _01080_, _01078_);
  or (_01082_, _01081_, _01044_);
  or (_01083_, _01082_, _01072_);
  and (_01084_, _01083_, _36955_);
  and (_01085_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01086_, _01085_, _01064_);
  or (_01087_, _01086_, _01084_);
  and (_32098_, _01087_, _42545_);
  and (_01088_, _00764_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_01089_, _42085_);
  or (_01090_, _00886_, _01089_);
  and (_01091_, _37883_, _37974_);
  and (_01092_, _37883_, _37958_);
  and (_01093_, _01092_, _37392_);
  or (_01094_, _01093_, _01091_);
  and (_01095_, _37883_, _37983_);
  and (_01096_, _00996_, _37889_);
  and (_01097_, _37883_, _37956_);
  or (_01098_, _01097_, _01096_);
  or (_01099_, _01098_, _01095_);
  or (_01100_, _01099_, _01094_);
  or (_01101_, _01100_, _01090_);
  or (_01102_, _00892_, _00849_);
  or (_01103_, _00881_, _00785_);
  and (_01104_, _37900_, _37974_);
  or (_01105_, _01104_, _00808_);
  or (_01106_, _01105_, _01103_);
  or (_01107_, _01106_, _01102_);
  and (_01108_, _38021_, _37931_);
  or (_01109_, _01108_, _38041_);
  or (_01110_, _01109_, _37925_);
  or (_01111_, _01032_, _00841_);
  or (_01112_, _01111_, _01110_);
  not (_01113_, _42083_);
  or (_01114_, _00850_, _01113_);
  or (_01115_, _01114_, _01112_);
  or (_01116_, _01115_, _01107_);
  or (_01117_, _01116_, _01101_);
  and (_01118_, _01117_, _00666_);
  or (_32100_, _01118_, _01088_);
  or (_01119_, _00860_, _01048_);
  or (_01120_, _01119_, _01054_);
  or (_01121_, _01120_, _00858_);
  or (_01122_, _01121_, _01034_);
  or (_01123_, _01097_, _01104_);
  or (_01124_, _01093_, _00961_);
  or (_01125_, _01124_, _01123_);
  not (_01126_, _38024_);
  nand (_01127_, _01126_, _37950_);
  or (_01128_, _00868_, _38032_);
  or (_01129_, _01128_, _37884_);
  or (_01130_, _00788_, _37980_);
  or (_01131_, _01130_, _01129_);
  or (_01132_, _01131_, _01127_);
  or (_01133_, _01132_, _01125_);
  or (_01134_, _01133_, _01122_);
  and (_01135_, _01134_, _00666_);
  and (_01136_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_01137_, _37902_, _36912_);
  or (_01138_, _01137_, _01136_);
  and (_01139_, _01138_, _42545_);
  or (_32102_, _01139_, _01135_);
  not (_01140_, _00984_);
  and (_01141_, _01140_, _37950_);
  and (_01142_, _37883_, _37932_);
  or (_01143_, _01142_, _00886_);
  or (_01144_, _00812_, _00788_);
  or (_01145_, _01144_, _01143_);
  not (_01146_, _38042_);
  or (_01147_, _01146_, _42082_);
  or (_01148_, _01147_, _01042_);
  nor (_01149_, _01148_, _01145_);
  nand (_01150_, _01149_, _01141_);
  and (_01151_, _37983_, _37882_);
  or (_01152_, _01151_, _00983_);
  or (_01153_, _00980_, _00960_);
  or (_01154_, _01153_, _01103_);
  or (_01155_, _01154_, _01152_);
  or (_01156_, _01155_, _00809_);
  or (_01157_, _01156_, _00804_);
  or (_01158_, _01157_, _01150_);
  and (_01159_, _01158_, _36955_);
  and (_01160_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01161_, _01160_, _37914_);
  or (_01162_, _01161_, _01159_);
  and (_32104_, _01162_, _42545_);
  or (_01163_, _01153_, _01105_);
  or (_01164_, _01163_, _01152_);
  or (_01165_, _38040_, _38026_);
  or (_01166_, _01165_, _37949_);
  or (_01167_, _01092_, _00984_);
  or (_01168_, _01167_, _01166_);
  or (_01169_, _00844_, _01089_);
  or (_01170_, _01169_, _01168_);
  or (_01171_, _00807_, _00803_);
  or (_01172_, _01171_, _01170_);
  or (_01173_, _01172_, _01164_);
  and (_01174_, _01173_, _36955_);
  and (_01175_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01176_, _01175_, _37915_);
  or (_01177_, _01176_, _01174_);
  and (_32106_, _01177_, _42545_);
  and (_01178_, _00764_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_01179_, _00768_, _38003_);
  not (_01180_, _37881_);
  and (_01181_, _37983_, _01180_);
  or (_01182_, _01181_, _01095_);
  or (_01183_, _01182_, _01179_);
  or (_01184_, _01123_, _01113_);
  or (_01185_, _01184_, _01183_);
  or (_01186_, _01094_, _00885_);
  or (_01187_, _01186_, _01090_);
  or (_01188_, _01187_, _01185_);
  and (_01189_, _01188_, _00666_);
  or (_32108_, _01189_, _01178_);
  nor (_38388_, _37600_, rst);
  nor (_38389_, _42076_, rst);
  and (_01190_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_01191_, _37120_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_01192_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01193_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_01194_, _01193_, _01192_);
  and (_01195_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_01196_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_01197_, _01196_, _01195_);
  and (_01198_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_01199_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_01200_, _01199_, _01198_);
  and (_01201_, _01200_, _01197_);
  and (_01202_, _01201_, _01194_);
  nor (_01203_, _01202_, _37120_);
  nor (_01204_, _01203_, _01191_);
  nor (_01205_, _01204_, _42060_);
  nor (_01206_, _01205_, _01190_);
  nor (_38391_, _01206_, rst);
  nor (_38401_, _37804_, rst);
  and (_38403_, _37828_, _42545_);
  nor (_38404_, _37875_, rst);
  nor (_38405_, _37852_, rst);
  and (_38406_, _37327_, _42545_);
  nor (_38407_, _37755_, rst);
  nor (_38408_, _37779_, rst);
  nor (_38409_, _42285_, rst);
  nor (_38410_, _42190_, rst);
  nor (_38412_, _42436_, rst);
  nor (_38413_, _42238_, rst);
  nor (_38414_, _42142_, rst);
  nor (_38415_, _42367_, rst);
  nor (_38416_, _42339_, rst);
  and (_01212_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_01214_, _37120_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_01216_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_01218_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_01220_, _01218_, _01216_);
  and (_01222_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_01224_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_01226_, _01224_, _01222_);
  and (_01228_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_01230_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_01232_, _01230_, _01228_);
  and (_01234_, _01232_, _01226_);
  and (_01236_, _01234_, _01220_);
  nor (_01238_, _01236_, _37120_);
  nor (_01240_, _01238_, _01214_);
  nor (_01242_, _01240_, _42060_);
  nor (_01244_, _01242_, _01212_);
  nor (_38418_, _01244_, rst);
  and (_01247_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_01249_, _37120_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_01251_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_01253_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_01255_, _01253_, _01251_);
  and (_01257_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_01259_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_01261_, _01259_, _01257_);
  and (_01263_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_01265_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_01267_, _01265_, _01263_);
  and (_01269_, _01267_, _01261_);
  and (_01271_, _01269_, _01255_);
  nor (_01273_, _01271_, _37120_);
  nor (_01275_, _01273_, _01249_);
  nor (_01277_, _01275_, _42060_);
  nor (_01279_, _01277_, _01247_);
  nor (_38419_, _01279_, rst);
  and (_01282_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_01284_, _37120_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_01286_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_01288_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_01290_, _01288_, _01286_);
  and (_01292_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_01294_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_01296_, _01294_, _01292_);
  and (_01298_, _01296_, _01290_);
  and (_01299_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_01300_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01301_, _01300_, _01299_);
  and (_01302_, _01301_, _01298_);
  nor (_01303_, _01302_, _37120_);
  nor (_01304_, _01303_, _01284_);
  nor (_01305_, _01304_, _42060_);
  nor (_01306_, _01305_, _01282_);
  nor (_38420_, _01306_, rst);
  and (_01307_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_01308_, _37120_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_01309_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_01310_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01311_, _01310_, _01309_);
  and (_01312_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_01313_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_01314_, _01313_, _01312_);
  and (_01315_, _01314_, _01311_);
  and (_01316_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_01317_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01318_, _01317_, _01316_);
  and (_01319_, _01318_, _01315_);
  nor (_01320_, _01319_, _37120_);
  nor (_01321_, _01320_, _01308_);
  nor (_01322_, _01321_, _42060_);
  nor (_01323_, _01322_, _01307_);
  nor (_38421_, _01323_, rst);
  and (_01324_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_01325_, _37120_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_01326_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_01327_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01328_, _01327_, _01326_);
  and (_01329_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_01330_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_01331_, _01330_, _01329_);
  and (_01332_, _01331_, _01328_);
  and (_01333_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_01334_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01335_, _01334_, _01333_);
  and (_01336_, _01335_, _01332_);
  nor (_01337_, _01336_, _37120_);
  nor (_01338_, _01337_, _01325_);
  nor (_01339_, _01338_, _42060_);
  nor (_01340_, _01339_, _01324_);
  nor (_38422_, _01340_, rst);
  and (_01341_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_01342_, _37120_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_01343_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_01344_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01345_, _01344_, _01343_);
  and (_01346_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_01347_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_01348_, _01347_, _01346_);
  and (_01349_, _01348_, _01345_);
  and (_01350_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_01351_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01352_, _01351_, _01350_);
  and (_01353_, _01352_, _01349_);
  nor (_01354_, _01353_, _37120_);
  nor (_01355_, _01354_, _01342_);
  nor (_01356_, _01355_, _42060_);
  nor (_01357_, _01356_, _01341_);
  nor (_38424_, _01357_, rst);
  and (_01358_, _42060_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_01359_, _37120_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_01360_, _37185_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_01361_, _37218_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01362_, _01361_, _01360_);
  and (_01363_, _37076_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_01364_, _37043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01365_, _01364_, _01363_);
  and (_01366_, _37010_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_01367_, _37153_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_01368_, _01367_, _01366_);
  and (_01369_, _01368_, _01365_);
  and (_01370_, _01369_, _01362_);
  nor (_01371_, _01370_, _37120_);
  nor (_01372_, _01371_, _01359_);
  nor (_01373_, _01372_, _42060_);
  nor (_01374_, _01373_, _01358_);
  nor (_38425_, _01374_, rst);
  and (_01375_, _36966_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_01376_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_01377_, _01375_, _38240_);
  and (_01378_, _01377_, _42545_);
  and (_38450_, _01378_, _01376_);
  not (_01379_, _01375_);
  or (_01380_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_01381_, _36966_, _42545_);
  and (_01382_, _01381_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_01383_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _42545_);
  or (_01384_, _01383_, _01382_);
  and (_38451_, _01384_, _01380_);
  nor (_38489_, _42081_, rst);
  nor (_38492_, _42054_, rst);
  nor (_01385_, _37962_, _38011_);
  nor (_01386_, _42147_, _28417_);
  and (_01387_, _42147_, _28417_);
  nor (_01388_, _01387_, _01386_);
  nor (_01389_, _42397_, _27935_);
  and (_01390_, _42397_, _27935_);
  nor (_01391_, _01390_, _01389_);
  nor (_01392_, _01391_, _01388_);
  nor (_01393_, _42344_, _38057_);
  and (_01394_, _42344_, _38057_);
  nor (_01395_, _01394_, _01393_);
  and (_01396_, _01395_, _42467_);
  nor (_01397_, _42248_, _28242_);
  and (_01398_, _42248_, _28242_);
  nor (_01399_, _01398_, _01397_);
  not (_01400_, _01399_);
  and (_01401_, _01400_, _01396_);
  and (_01402_, _01401_, _01392_);
  nor (_01403_, _31755_, _39547_);
  and (_01404_, _01403_, _01402_);
  and (_01405_, _01404_, _01385_);
  not (_01406_, _01405_);
  and (_01407_, _01392_, _01396_);
  nor (_01408_, _01399_, _39143_);
  and (_01409_, _42195_, _32994_);
  nor (_01410_, _42195_, _32994_);
  or (_01411_, _01410_, _01409_);
  or (_01412_, _42294_, _27573_);
  nand (_01413_, _42294_, _27573_);
  and (_01414_, _01413_, _01412_);
  or (_01415_, _42443_, _27332_);
  nand (_01416_, _42443_, _27332_);
  and (_01417_, _01416_, _01415_);
  or (_01418_, _01417_, _01414_);
  nor (_01419_, _01418_, _01411_);
  and (_01420_, _01419_, _01408_);
  and (_01421_, _01420_, _01407_);
  nor (_01422_, _28088_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_01423_, _01422_, _01421_);
  not (_01424_, _37933_);
  nor (_01425_, _00769_, _01048_);
  not (_01426_, _00848_);
  nor (_01427_, _01041_, _37975_);
  and (_01428_, _01427_, _01426_);
  and (_01429_, _01428_, _00998_);
  nor (_01430_, _01385_, _37913_);
  nor (_01431_, _31906_, _30006_);
  and (_01432_, _01431_, _33266_);
  and (_01433_, _01432_, _33886_);
  not (_01434_, _01433_);
  nor (_01435_, _01434_, _34616_);
  and (_01436_, _01435_, _35465_);
  and (_01437_, _01436_, _36238_);
  and (_01438_, _01437_, _01430_);
  and (_01439_, _01438_, _30203_);
  and (_01440_, _01385_, _29152_);
  not (_01441_, _37913_);
  and (_01442_, _37912_, _37947_);
  nor (_01443_, _01442_, _01385_);
  nor (_01444_, _01443_, _01441_);
  and (_01445_, _01444_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_01446_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_01447_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01448_, _01447_, _01446_);
  nor (_01449_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_01450_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01451_, _01450_, _01449_);
  and (_01452_, _01451_, _01448_);
  and (_01453_, _01452_, _38049_);
  or (_01454_, _01453_, _01445_);
  or (_01455_, _01454_, _01440_);
  nor (_01456_, _01455_, _01439_);
  or (_01457_, _37892_, _37956_);
  nor (_01458_, _01457_, _37948_);
  nor (_01459_, _01458_, _00926_);
  not (_01460_, _01459_);
  and (_01461_, _01460_, _01456_);
  and (_01462_, _01461_, _01429_);
  and (_01463_, _00766_, _37403_);
  or (_01464_, _01463_, _37960_);
  nor (_01465_, _01464_, _01456_);
  and (_01466_, _01465_, _37955_);
  or (_01467_, _01466_, _01462_);
  and (_01468_, _01467_, _01425_);
  and (_01469_, _01468_, _01424_);
  nor (_01470_, _01469_, _42093_);
  and (_01471_, _37958_, _37924_);
  nor (_01472_, _01471_, _00823_);
  nor (_01473_, _01472_, _36912_);
  nor (_01474_, _01473_, _38013_);
  not (_01475_, _01474_);
  nor (_01476_, _01475_, _01470_);
  nor (_01477_, _38636_, _38627_);
  and (_01478_, _01477_, _38678_);
  not (_01479_, _01478_);
  and (_01480_, _01479_, _01444_);
  not (_01481_, _39004_);
  and (_01482_, _01481_, _38049_);
  nor (_01483_, _01482_, _01480_);
  not (_01484_, _01483_);
  nor (_01485_, _01484_, _01476_);
  not (_01486_, _01485_);
  nor (_01487_, _01486_, _01423_);
  and (_01488_, _01487_, _01406_);
  nor (_01489_, _38013_, rst);
  and (_38496_, _01489_, _01488_);
  and (_38497_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _42545_);
  and (_38498_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _42545_);
  and (_01490_, _38013_, _31111_);
  and (_01491_, _01048_, _37911_);
  and (_01492_, _01491_, _38288_);
  and (_01493_, _00998_, _37962_);
  and (_01494_, _01493_, _01427_);
  nor (_01495_, _01494_, _42093_);
  and (_01496_, _01471_, _36901_);
  nor (_01497_, _01496_, _38013_);
  not (_01498_, _01497_);
  nor (_01499_, _01498_, _01495_);
  and (_01500_, _01499_, _01473_);
  and (_01501_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01502_, _01501_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01503_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01504_, _01503_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01505_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01506_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01507_, _01506_, _01505_);
  and (_01508_, _01507_, _01504_);
  and (_01509_, _01508_, _01502_);
  and (_01510_, _01509_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01511_, _01510_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01512_, _01511_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_01513_, _01512_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01514_, _01513_, _38240_);
  or (_01515_, _01513_, _38240_);
  and (_01516_, _01515_, _01514_);
  and (_01517_, _01516_, _01500_);
  nor (_01518_, _01491_, _01473_);
  nand (_01519_, _01518_, _01499_);
  not (_01520_, _00766_);
  and (_01521_, _01425_, _01520_);
  and (_01522_, _01521_, _01428_);
  and (_01523_, _01522_, _01493_);
  nor (_01524_, _01523_, _42093_);
  and (_01525_, _37932_, _36901_);
  and (_01526_, _01525_, _37908_);
  or (_01527_, _01526_, _01524_);
  nor (_01528_, _01527_, _01519_);
  and (_01529_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01530_, _01496_, _42077_);
  or (_01531_, _01530_, _01529_);
  or (_01532_, _01531_, _01517_);
  nor (_01533_, _01532_, _01492_);
  nand (_01534_, _01533_, _01488_);
  or (_01535_, _01534_, _01490_);
  not (_01536_, _01526_);
  and (_01537_, _01536_, _01499_);
  and (_01538_, _01537_, _42076_);
  not (_01539_, _01206_);
  nor (_01540_, _01537_, _01539_);
  nor (_01541_, _01540_, _01538_);
  and (_01542_, _01541_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_01543_, _01541_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01544_, _01537_, _42339_);
  not (_01545_, _01374_);
  nor (_01546_, _01537_, _01545_);
  nor (_01547_, _01546_, _01544_);
  and (_01548_, _01547_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_01549_, _01547_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_01550_, _01549_, _01548_);
  and (_01551_, _01537_, _42367_);
  not (_01552_, _01357_);
  nor (_01553_, _01537_, _01552_);
  nor (_01554_, _01553_, _01551_);
  and (_01555_, _01554_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_01556_, _01554_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_01557_, _01537_, _42142_);
  not (_01558_, _01340_);
  nor (_01559_, _01537_, _01558_);
  nor (_01560_, _01559_, _01557_);
  nand (_01561_, _01560_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01562_, _01537_, _42238_);
  not (_01563_, _01323_);
  nor (_01564_, _01537_, _01563_);
  nor (_01565_, _01564_, _01562_);
  and (_01566_, _01565_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_01567_, _01565_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01568_, _01537_, _42436_);
  not (_01569_, _01306_);
  nor (_01570_, _01537_, _01569_);
  nor (_01571_, _01570_, _01568_);
  and (_01572_, _01571_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01573_, _01537_, _42190_);
  not (_01574_, _01279_);
  nor (_01575_, _01537_, _01574_);
  nor (_01576_, _01575_, _01573_);
  and (_01577_, _01576_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01578_, _01537_, _42285_);
  not (_01579_, _01244_);
  nor (_01580_, _01537_, _01579_);
  nor (_01581_, _01580_, _01578_);
  and (_01582_, _01581_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_01583_, _01576_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_01584_, _01583_, _01577_);
  and (_01585_, _01584_, _01582_);
  nor (_01586_, _01585_, _01577_);
  not (_01587_, _01586_);
  nor (_01588_, _01571_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_01589_, _01588_, _01572_);
  and (_01590_, _01589_, _01587_);
  nor (_01591_, _01590_, _01572_);
  nor (_01592_, _01591_, _01567_);
  or (_01593_, _01592_, _01566_);
  or (_01594_, _01560_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01595_, _01594_, _01561_);
  nand (_01596_, _01595_, _01593_);
  and (_01597_, _01596_, _01561_);
  nor (_01598_, _01597_, _01556_);
  or (_01599_, _01598_, _01555_);
  and (_01600_, _01599_, _01550_);
  nor (_01601_, _01600_, _01548_);
  nor (_01602_, _01601_, _01543_);
  or (_01603_, _01602_, _01542_);
  and (_01604_, _01603_, _01502_);
  and (_01605_, _01604_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01606_, _01605_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01607_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_01608_, _01607_, _01541_);
  not (_01609_, _01541_);
  nor (_01610_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01611_, _01610_, _38214_);
  and (_01612_, _01611_, _38219_);
  and (_01613_, _01612_, _38204_);
  nor (_01614_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01615_, _01614_, _01613_);
  nor (_01616_, _01615_, _01609_);
  nor (_01617_, _01616_, _01608_);
  or (_01618_, _01541_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01619_, _01541_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01620_, _01619_, _01618_);
  and (_01621_, _01620_, _01617_);
  or (_01623_, _01621_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_01624_, _01621_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_01626_, _01624_, _01623_);
  not (_01627_, _01518_);
  and (_01629_, _01627_, _01537_);
  and (_01630_, _37908_, _36901_);
  and (_01632_, _01630_, _37932_);
  nor (_01633_, _01632_, _01524_);
  nor (_01635_, _01633_, _01629_);
  and (_01636_, _01635_, _01626_);
  or (_01638_, _01636_, _01535_);
  and (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01641_, _37065_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01642_, _01641_, _42060_);
  nor (_01644_, _01642_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_01645_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_01647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_01648_, _01647_, _01645_);
  not (_01650_, _01648_);
  nor (_01651_, _01650_, _01644_);
  and (_01653_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_01654_, _01653_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01655_, _01654_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01656_, _01655_, _01651_);
  and (_01657_, _01656_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01658_, _01657_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01659_, _01658_, _01639_);
  and (_01660_, _01659_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01661_, _01660_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_01662_, _01660_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01663_, _01662_, _01661_);
  or (_01664_, _01663_, _01488_);
  and (_01665_, _01664_, _42545_);
  and (_38499_, _01665_, _01638_);
  and (_01666_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _42545_);
  and (_01667_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01668_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_01669_, _36955_, _01668_);
  not (_01670_, _01669_);
  not (_01671_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01672_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01673_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01674_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_01675_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_01676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_01677_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_01678_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_01679_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_01680_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_01681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01682_, _01681_, _01680_);
  and (_01683_, _01682_, _01679_);
  and (_01684_, _01683_, _01678_);
  and (_01685_, _01684_, _01677_);
  and (_01686_, _01685_, _01676_);
  and (_01687_, _01686_, _01675_);
  and (_01688_, _01687_, _01674_);
  and (_01689_, _01688_, _01673_);
  and (_01690_, _01689_, _01672_);
  nor (_01691_, _01690_, _01671_);
  and (_01692_, _01690_, _01671_);
  nor (_01693_, _01692_, _01691_);
  nor (_01694_, _01689_, _01672_);
  nor (_01695_, _01694_, _01690_);
  not (_01696_, _01695_);
  not (_01697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01698_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01700_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01701_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01702_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_01703_, _01702_, _01700_);
  and (_01704_, _01703_, _01701_);
  nor (_01705_, _01704_, _01700_);
  nor (_01706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01707_, _01706_, _01699_);
  not (_01708_, _01707_);
  nor (_01709_, _01708_, _01705_);
  nor (_01710_, _01709_, _01699_);
  not (_01711_, _01710_);
  and (_01712_, _01711_, _01688_);
  and (_01713_, _01712_, _01698_);
  and (_01714_, _01713_, _01697_);
  and (_01715_, _01714_, _01696_);
  nor (_01716_, _01714_, _01696_);
  or (_01717_, _01716_, _01715_);
  not (_01718_, _01717_);
  and (_01719_, _01710_, _01689_);
  and (_01720_, _01710_, _01688_);
  and (_01721_, _01720_, _01698_);
  nor (_01722_, _01721_, _01697_);
  or (_01723_, _01722_, _01719_);
  nor (_01724_, _01720_, _01698_);
  nor (_01725_, _01724_, _01721_);
  not (_01726_, _01725_);
  and (_01727_, _01710_, _01687_);
  nor (_01728_, _01727_, _01674_);
  nor (_01729_, _01728_, _01720_);
  not (_01730_, _01729_);
  and (_01731_, _01710_, _01685_);
  and (_01732_, _01731_, _01676_);
  nor (_01733_, _01732_, _01675_);
  nor (_01734_, _01733_, _01727_);
  not (_01735_, _01734_);
  nor (_01736_, _01731_, _01676_);
  nor (_01737_, _01736_, _01732_);
  and (_01738_, _01710_, _01683_);
  and (_01739_, _01738_, _01678_);
  nor (_01740_, _01738_, _01678_);
  nor (_01741_, _01740_, _01739_);
  not (_01742_, _01741_);
  and (_01743_, _01710_, _01682_);
  nor (_01744_, _01743_, _01679_);
  or (_01745_, _01744_, _01738_);
  nand (_01746_, _01710_, _01681_);
  and (_01747_, _01746_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_01748_, _01747_, _01743_);
  not (_01749_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01750_, _01710_, _01749_);
  nor (_01751_, _01710_, _01749_);
  nor (_01752_, _01751_, _01750_);
  not (_01753_, _01752_);
  and (_01754_, _00692_, _00676_);
  or (_01755_, _01754_, _00732_);
  nor (_01756_, _01755_, _00743_);
  and (_01757_, _01756_, _00724_);
  not (_01758_, _00742_);
  nor (_01759_, _00725_, _00747_);
  nor (_01760_, _01759_, _01758_);
  and (_01761_, _00742_, _00692_);
  and (_01762_, _00702_, _00729_);
  and (_01763_, _00727_, _01762_);
  or (_01764_, _01763_, _01761_);
  nor (_01765_, _01764_, _01760_);
  not (_01766_, _01765_);
  not (_01767_, _00721_);
  not (_01768_, _00727_);
  nor (_01769_, _00736_, _00676_);
  and (_01770_, _01769_, _01768_);
  nor (_01771_, _01770_, _01767_);
  nor (_01772_, _01771_, _01766_);
  and (_01773_, _01772_, _01757_);
  not (_01774_, _00689_);
  and (_01775_, _00729_, _00670_);
  and (_01776_, _01775_, _00695_);
  and (_01777_, _00695_, _00692_);
  nor (_01778_, _01777_, _01776_);
  and (_01779_, _01778_, _00705_);
  and (_01780_, _01779_, _01774_);
  and (_01781_, _00744_, _00677_);
  and (_01782_, _00726_, _00711_);
  nor (_01783_, _01782_, _00690_);
  and (_01784_, _00725_, _37804_);
  not (_01785_, _01784_);
  nor (_01786_, _01775_, _00711_);
  and (_01787_, _01786_, _01785_);
  nor (_01788_, _01787_, _01783_);
  nor (_01789_, _01788_, _01781_);
  and (_01790_, _01789_, _01780_);
  not (_01791_, _00683_);
  and (_01792_, _00670_, _00671_);
  nor (_01793_, _01792_, _00725_);
  nor (_01794_, _01793_, _01791_);
  not (_01795_, _01794_);
  and (_01796_, _00718_, _00676_);
  not (_01797_, _00695_);
  and (_01798_, _00710_, _00670_);
  nor (_01799_, _00700_, _01798_);
  nor (_01800_, _01799_, _01797_);
  nor (_01801_, _01800_, _01796_);
  and (_01802_, _01801_, _01795_);
  nor (_01803_, _00748_, _00738_);
  nor (_01804_, _01793_, _37852_);
  and (_01805_, _00742_, _00717_);
  nor (_01806_, _01805_, _01804_);
  and (_01807_, _01806_, _01803_);
  and (_01808_, _01807_, _01802_);
  and (_01809_, _01808_, _01790_);
  not (_01810_, _00736_);
  and (_01811_, _00730_, _00670_);
  not (_01812_, _01811_);
  and (_01813_, _00696_, _00720_);
  not (_01814_, _01813_);
  nor (_01815_, _00741_, _00692_);
  and (_01816_, _01815_, _01814_);
  and (_01817_, _01816_, _01812_);
  and (_01818_, _01817_, _01759_);
  nor (_01819_, _01818_, _01810_);
  not (_01820_, _01819_);
  and (_01821_, _00696_, _00710_);
  nor (_01822_, _01813_, _01821_);
  nor (_01823_, _01822_, _01758_);
  not (_01824_, _01823_);
  and (_01825_, _00696_, _00691_);
  nor (_01826_, _00721_, _01825_);
  nor (_01827_, _01826_, _01758_);
  not (_01828_, _01762_);
  nor (_01829_, _00736_, _00690_);
  nor (_01830_, _01829_, _01828_);
  nor (_01831_, _01830_, _01827_);
  and (_01832_, _01831_, _01824_);
  and (_01833_, _01832_, _01820_);
  and (_01834_, _01833_, _01809_);
  and (_01835_, _01834_, _01773_);
  not (_01836_, _01835_);
  nor (_01837_, _01703_, _01701_);
  nor (_01838_, _01837_, _01704_);
  nand (_01839_, _01838_, _01836_);
  or (_01840_, _01776_, _00719_);
  and (_01841_, _00702_, _00671_);
  and (_01842_, _00727_, _01841_);
  or (_01843_, _01842_, _00738_);
  or (_01844_, _01843_, _01840_);
  or (_01845_, _01844_, _00689_);
  nand (_01846_, _01765_, _01756_);
  or (_01847_, _01846_, _01845_);
  or (_01848_, _01847_, _01835_);
  nor (_01849_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01850_, _01849_, _01701_);
  and (_01851_, _01850_, _01848_);
  or (_01852_, _01838_, _01836_);
  and (_01853_, _01852_, _01839_);
  nand (_01854_, _01853_, _01851_);
  and (_01855_, _01854_, _01839_);
  not (_01856_, _01855_);
  and (_01857_, _01708_, _01705_);
  nor (_01858_, _01857_, _01709_);
  and (_01859_, _01858_, _01856_);
  and (_01860_, _01859_, _01753_);
  not (_01861_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_01862_, _01750_, _01861_);
  nand (_01863_, _01862_, _01746_);
  and (_01864_, _01863_, _01860_);
  and (_01865_, _01864_, _01748_);
  and (_01866_, _01865_, _01745_);
  and (_01867_, _01866_, _01742_);
  nor (_01868_, _01739_, _01677_);
  or (_01869_, _01868_, _01731_);
  nand (_01870_, _01869_, _01867_);
  nor (_01871_, _01870_, _01737_);
  and (_01872_, _01871_, _01735_);
  and (_01873_, _01872_, _01730_);
  and (_01874_, _01873_, _01726_);
  and (_01875_, _01874_, _01723_);
  and (_01876_, _01875_, _01718_);
  nor (_01877_, _01876_, _01715_);
  not (_01878_, _01877_);
  nor (_01879_, _01878_, _01693_);
  and (_01880_, _01878_, _01693_);
  or (_01881_, _01880_, _01879_);
  or (_01882_, _01881_, _01670_);
  or (_01883_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_01884_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_01885_, _01884_, _01883_);
  and (_01886_, _01885_, _01882_);
  or (_38501_, _01886_, _01667_);
  nor (_01887_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_38502_, _01887_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_38503_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _42545_);
  nor (_01888_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_01889_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01890_, _01889_, _01888_);
  nor (_01891_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_01892_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_01893_, _01892_, _01891_);
  and (_01894_, _01893_, _01890_);
  nor (_01895_, _01894_, rst);
  and (_01896_, \oc8051_top_1.oc8051_rom1.ea_int , _36922_);
  nand (_01897_, _01896_, _36955_);
  and (_01898_, _01897_, _38503_);
  or (_38504_, _01898_, _01895_);
  and (_01899_, _01894_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_01900_, _01899_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_38506_, _01900_, _42545_);
  nor (_01901_, _01644_, _42060_);
  or (_01902_, _01835_, _37131_);
  and (_01903_, _01848_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_01904_, _01835_, _37131_);
  and (_01905_, _01904_, _01902_);
  nand (_01906_, _01905_, _01903_);
  and (_01907_, _01906_, _01902_);
  nor (_01908_, _01907_, _42060_);
  and (_01909_, _01908_, _37032_);
  nor (_01910_, _01908_, _37032_);
  nor (_01911_, _01910_, _01909_);
  nor (_01912_, _01911_, _01901_);
  and (_01913_, _37207_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01914_, _01913_, _01901_);
  and (_01915_, _01914_, _01847_);
  or (_01916_, _01915_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01917_, _01916_, _01912_);
  and (_38507_, _01917_, _42545_);
  or (_01918_, _37556_, _37800_);
  nor (_01919_, _01918_, _37848_);
  not (_01920_, _37822_);
  and (_01921_, _37775_, _01920_);
  and (_01922_, _01921_, _37870_);
  not (_01923_, _01381_);
  nor (_01924_, _01923_, _37262_);
  and (_01925_, _01924_, _37751_);
  and (_01926_, _01925_, _01922_);
  and (_38510_, _01926_, _01919_);
  nor (_01927_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_01928_, _01927_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_01929_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_38513_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _42545_);
  and (_01930_, _38513_, _01929_);
  or (_38511_, _01930_, _01928_);
  not (_01931_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01932_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01933_, _01932_, _01931_);
  and (_01934_, _01932_, _01931_);
  nor (_01935_, _01934_, _01933_);
  not (_01936_, _01935_);
  and (_01937_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01938_, _01937_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01939_, _01937_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01940_, _01939_, _01938_);
  or (_01941_, _01940_, _01932_);
  and (_01942_, _01941_, _01936_);
  nor (_01943_, _01933_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01944_, _01933_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_01945_, _01944_, _01943_);
  or (_01946_, _01938_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_38515_, _01946_, _42545_);
  and (_01947_, _38515_, _01945_);
  and (_38514_, _01947_, _01942_);
  not (_01948_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_01949_, _01644_, _01948_);
  and (_01950_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_01951_, _01949_);
  and (_01952_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_01953_, _01952_, _01950_);
  and (_38516_, _01953_, _42545_);
  and (_01954_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01955_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_01956_, _01955_, _01954_);
  and (_38517_, _01956_, _42545_);
  and (_01957_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_01958_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01959_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _01958_);
  and (_01960_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01961_, _01960_, _01957_);
  and (_38518_, _01961_, _42545_);
  and (_01962_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01963_, _01962_, _01959_);
  and (_38519_, _01963_, _42545_);
  or (_01964_, _01958_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_38521_, _01964_, _42545_);
  not (_01965_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_01966_, _01965_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01967_, _01966_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01968_, _01958_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_01969_, _01968_, _42545_);
  and (_38522_, _01969_, _01967_);
  or (_01970_, _01958_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_38523_, _01970_, _42545_);
  nor (_01971_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_01972_, _01971_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01973_, _01972_, _42545_);
  and (_01974_, _38513_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_38524_, _01974_, _01973_);
  and (_01975_, _01948_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_01976_, _01975_, _01972_);
  and (_38525_, _01976_, _42545_);
  not (_01977_, _01972_);
  or (_01978_, _01977_, _38288_);
  or (_01979_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_01980_, _01979_, _42545_);
  and (_38526_, _01980_, _01978_);
  nand (_01981_, _37921_, _42545_);
  nor (_38527_, _01981_, _38053_);
  or (_01982_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_01983_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_01984_, _01375_, _01983_);
  and (_01985_, _01984_, _42545_);
  and (_38565_, _01985_, _01982_);
  or (_01986_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_01987_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_01988_, _01375_, _01987_);
  and (_01989_, _01988_, _42545_);
  and (_38566_, _01989_, _01986_);
  or (_01990_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_01991_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_01992_, _01375_, _01991_);
  and (_01993_, _01992_, _42545_);
  and (_38567_, _01993_, _01990_);
  or (_01994_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_01995_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_01996_, _01375_, _01995_);
  and (_01997_, _01996_, _42545_);
  and (_38568_, _01997_, _01994_);
  or (_01998_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_01999_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_02000_, _01999_, _42545_);
  and (_38569_, _02000_, _01998_);
  or (_02001_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_02002_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_02003_, _01375_, _02002_);
  and (_02004_, _02003_, _42545_);
  and (_38571_, _02004_, _02001_);
  or (_02005_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_02006_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_02007_, _02006_, _42545_);
  and (_38572_, _02007_, _02005_);
  or (_02008_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_02009_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_02010_, _01375_, _02009_);
  and (_02011_, _02010_, _42545_);
  and (_38573_, _02011_, _02008_);
  or (_02012_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_02013_, _01375_, _38208_);
  and (_02014_, _02013_, _42545_);
  and (_38574_, _02014_, _02012_);
  or (_02015_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_02016_, _01375_, _38214_);
  and (_02017_, _02016_, _42545_);
  and (_38575_, _02017_, _02015_);
  or (_02018_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_02019_, _01375_, _38219_);
  and (_02020_, _02019_, _42545_);
  and (_38576_, _02020_, _02018_);
  or (_02021_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_02022_, _01375_, _38204_);
  and (_02023_, _02022_, _42545_);
  and (_38577_, _02023_, _02021_);
  or (_02024_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_02025_, _01375_, _38225_);
  and (_02026_, _02025_, _42545_);
  and (_38578_, _02026_, _02024_);
  or (_02027_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_02028_, _01375_, _38230_);
  and (_02029_, _02028_, _42545_);
  and (_38579_, _02029_, _02027_);
  or (_02030_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_02031_, _01375_, _38235_);
  and (_02032_, _02031_, _42545_);
  and (_38580_, _02032_, _02030_);
  and (_02033_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_02034_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_02035_, _02034_, _02033_);
  and (_38584_, _02035_, _42545_);
  and (_02036_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_02037_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_02038_, _02037_, _02036_);
  and (_38585_, _02038_, _42545_);
  and (_02039_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_02040_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_02041_, _02040_, _02039_);
  and (_38586_, _02041_, _42545_);
  and (_02042_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_02043_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_02044_, _02043_, _02042_);
  and (_38587_, _02044_, _42545_);
  and (_02045_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_02046_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or (_02047_, _02046_, _02045_);
  and (_38588_, _02047_, _42545_);
  and (_02048_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_02049_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or (_02050_, _02049_, _02048_);
  and (_38589_, _02050_, _42545_);
  and (_02051_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_02052_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or (_02053_, _02052_, _02051_);
  and (_38590_, _02053_, _42545_);
  and (_02054_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_02055_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or (_02056_, _02055_, _02054_);
  and (_38591_, _02056_, _42545_);
  and (_02057_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_02058_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or (_02059_, _02058_, _02057_);
  and (_38592_, _02059_, _42545_);
  and (_02060_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_02061_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02062_, _02061_, _02060_);
  and (_38593_, _02062_, _42545_);
  and (_02063_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_02064_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or (_02065_, _02064_, _02063_);
  and (_38594_, _02065_, _42545_);
  and (_02066_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_02067_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or (_02068_, _02067_, _02066_);
  and (_38595_, _02068_, _42545_);
  and (_02069_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_02070_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or (_02071_, _02070_, _02069_);
  and (_38596_, _02071_, _42545_);
  and (_02072_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_02073_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or (_02074_, _02073_, _02072_);
  and (_38597_, _02074_, _42545_);
  and (_02075_, _01375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_02076_, _01379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or (_02077_, _02076_, _02075_);
  and (_38598_, _02077_, _42545_);
  and (_38772_, _37809_, _42545_);
  and (_38773_, _37833_, _42545_);
  and (_38774_, _37880_, _42545_);
  nor (_38775_, _41981_, rst);
  and (_02078_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_02079_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_02080_, _02079_, _02078_);
  and (_38776_, _02080_, _42545_);
  and (_02081_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02082_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_02083_, _02082_, _01949_);
  or (_02084_, _02083_, _02081_);
  and (_38777_, _02084_, _42545_);
  and (_02085_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02086_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_02087_, _02086_, _02085_);
  and (_38778_, _02087_, _42545_);
  and (_02088_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02089_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_02090_, _02089_, _02088_);
  and (_38779_, _02090_, _42545_);
  and (_02091_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02092_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_02093_, _02092_, _02091_);
  and (_38781_, _02093_, _42545_);
  and (_02094_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02095_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_02096_, _02095_, _01949_);
  or (_02097_, _02096_, _02094_);
  and (_38782_, _02097_, _42545_);
  and (_02098_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02099_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_02100_, _02099_, _02098_);
  and (_38783_, _02100_, _42545_);
  and (_02101_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02102_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_02103_, _02102_, _02101_);
  and (_38784_, _02103_, _42545_);
  and (_02104_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_02105_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_02106_, _02105_, _02104_);
  and (_38785_, _02106_, _42545_);
  and (_02107_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_02108_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_02109_, _02108_, _02107_);
  and (_38786_, _02109_, _42545_);
  and (_02110_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_02111_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_02112_, _02111_, _02110_);
  and (_38787_, _02112_, _42545_);
  and (_02113_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_02114_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_02116_, _02114_, _02113_);
  and (_38788_, _02116_, _42545_);
  and (_02119_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_02121_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_02123_, _02121_, _02119_);
  and (_38789_, _02123_, _42545_);
  and (_02126_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_02128_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_02130_, _02128_, _02126_);
  and (_38790_, _02130_, _42545_);
  and (_02133_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_02135_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_02137_, _02135_, _02133_);
  and (_38792_, _02137_, _42545_);
  and (_02140_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_02142_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_02144_, _02142_, _02140_);
  and (_38793_, _02144_, _42545_);
  and (_02147_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_02149_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_02151_, _02149_, _02147_);
  and (_38794_, _02151_, _42545_);
  and (_02154_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_02156_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_02158_, _02156_, _02154_);
  and (_38795_, _02158_, _42545_);
  and (_02161_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_02163_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_02165_, _02163_, _02161_);
  and (_38796_, _02165_, _42545_);
  and (_02168_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_02170_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_02172_, _02170_, _02168_);
  and (_38797_, _02172_, _42545_);
  and (_02175_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_02176_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_02177_, _02176_, _02175_);
  and (_38798_, _02177_, _42545_);
  and (_02178_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_02179_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_02180_, _02179_, _02178_);
  and (_38799_, _02180_, _42545_);
  and (_02181_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_02182_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_02183_, _02182_, _02181_);
  and (_38800_, _02183_, _42545_);
  and (_02184_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_02185_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_02186_, _02185_, _02184_);
  and (_38801_, _02186_, _42545_);
  and (_02187_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_02188_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_02189_, _02188_, _02187_);
  and (_38803_, _02189_, _42545_);
  and (_02190_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_02191_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_02192_, _02191_, _02190_);
  and (_38804_, _02192_, _42545_);
  and (_02193_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_02194_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_02195_, _02194_, _02193_);
  and (_38805_, _02195_, _42545_);
  and (_02196_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_02197_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_02198_, _02197_, _02196_);
  and (_38806_, _02198_, _42545_);
  and (_02199_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_02200_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_02201_, _02200_, _02199_);
  and (_38807_, _02201_, _42545_);
  and (_02202_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_02203_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_02204_, _02203_, _02202_);
  and (_38808_, _02204_, _42545_);
  and (_02205_, _01949_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_02206_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_02207_, _02206_, _02205_);
  and (_38809_, _02207_, _42545_);
  nor (_38810_, _42268_, rst);
  nor (_38812_, _42168_, rst);
  nor (_38813_, _42418_, rst);
  nor (_38814_, _42221_, rst);
  nor (_38815_, _42117_, rst);
  nor (_38816_, _42388_, rst);
  nor (_38818_, _42321_, rst);
  and (_38833_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _42545_);
  and (_38834_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _42545_);
  and (_38835_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _42545_);
  and (_38836_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _42545_);
  and (_38837_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _42545_);
  and (_38839_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _42545_);
  and (_38840_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _42545_);
  or (_02208_, _01528_, _01491_);
  and (_02209_, _02208_, _32276_);
  and (_02210_, _01500_, _42286_);
  and (_02211_, _01496_, _01579_);
  and (_02212_, _38013_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_02213_, _02212_, _02211_);
  or (_02214_, _02213_, _02210_);
  nor (_02215_, _01581_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_02216_, _02215_, _01582_);
  and (_02217_, _02216_, _01635_);
  nor (_02218_, _02217_, _02214_);
  nand (_02219_, _02218_, _01488_);
  or (_02220_, _02219_, _02209_);
  or (_02221_, _01488_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_02222_, _02221_, _42545_);
  and (_38841_, _02222_, _02220_);
  and (_02223_, _02208_, _32918_);
  and (_02224_, _01500_, _42191_);
  and (_02225_, _01496_, _01574_);
  and (_02226_, _38013_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_02227_, _02226_, _02225_);
  or (_02228_, _02227_, _02224_);
  or (_02229_, _02228_, _02223_);
  nor (_02230_, _01584_, _01582_);
  nor (_02231_, _02230_, _01585_);
  nand (_02232_, _02231_, _01635_);
  nand (_02233_, _02232_, _01488_);
  or (_02234_, _02233_, _02229_);
  or (_02235_, _01488_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_02236_, _02235_, _42545_);
  and (_38842_, _02236_, _02234_);
  and (_02237_, _02208_, _33593_);
  and (_02238_, _01500_, _42437_);
  and (_02239_, _01496_, _01569_);
  and (_02240_, _38013_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_02241_, _02240_, _02239_);
  or (_02242_, _02241_, _02238_);
  or (_02243_, _02242_, _02237_);
  nor (_02244_, _01589_, _01587_);
  nor (_02245_, _02244_, _01590_);
  nand (_02246_, _02245_, _01635_);
  nand (_02247_, _02246_, _01488_);
  or (_02248_, _02247_, _02243_);
  not (_02249_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02250_, _01644_, _02249_);
  and (_02251_, _01644_, _02249_);
  nor (_02252_, _02251_, _02250_);
  or (_02253_, _02252_, _01488_);
  and (_02254_, _02253_, _42545_);
  and (_38843_, _02254_, _02248_);
  and (_02255_, _02208_, _34344_);
  and (_02256_, _01500_, _42239_);
  and (_02257_, _01496_, _01563_);
  and (_02258_, _38013_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_02259_, _02258_, _02257_);
  or (_02260_, _02259_, _02256_);
  or (_02261_, _01567_, _01566_);
  nand (_02262_, _02261_, _01591_);
  not (_02263_, _01629_);
  and (_02264_, _01527_, _02263_);
  or (_02265_, _02261_, _01591_);
  and (_02266_, _02265_, _02264_);
  and (_02267_, _02266_, _02262_);
  nor (_02268_, _02267_, _02260_);
  nand (_02269_, _02268_, _01488_);
  or (_02270_, _02269_, _02255_);
  and (_02271_, _02250_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02272_, _02250_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02273_, _02272_, _02271_);
  or (_02274_, _02273_, _01488_);
  and (_02275_, _02274_, _42545_);
  and (_38844_, _02275_, _02270_);
  and (_02276_, _02208_, _35139_);
  or (_02277_, _01595_, _01593_);
  and (_02278_, _02264_, _01596_);
  and (_02279_, _02278_, _02277_);
  and (_02280_, _01500_, _42143_);
  and (_02281_, _01496_, _01558_);
  and (_02282_, _38013_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_02283_, _02282_, _02281_);
  or (_02284_, _02283_, _02280_);
  nor (_02285_, _02284_, _02279_);
  nand (_02286_, _02285_, _01488_);
  or (_02287_, _02286_, _02276_);
  and (_02288_, _02271_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02289_, _02271_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02290_, _02289_, _02288_);
  or (_02291_, _02290_, _01488_);
  and (_02292_, _02291_, _42545_);
  and (_38845_, _02292_, _02287_);
  and (_02293_, _02208_, _35967_);
  and (_02294_, _01500_, _42368_);
  and (_02295_, _01496_, _01552_);
  and (_02296_, _38013_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_02297_, _02296_, _02295_);
  or (_02298_, _02297_, _02294_);
  or (_02299_, _01556_, _01555_);
  nand (_02300_, _02299_, _01597_);
  or (_02301_, _02299_, _01597_);
  and (_02302_, _02301_, _02264_);
  and (_02303_, _02302_, _02300_);
  nor (_02304_, _02303_, _02298_);
  nand (_02305_, _02304_, _01488_);
  or (_02306_, _02305_, _02293_);
  nor (_02307_, _02288_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02308_, _02307_, _01651_);
  or (_02309_, _02308_, _01488_);
  and (_02310_, _02309_, _42545_);
  and (_38846_, _02310_, _02306_);
  nor (_02311_, _01651_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02312_, _01651_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_02313_, _02312_, _02311_);
  or (_02314_, _02313_, _01488_);
  and (_02315_, _02314_, _42545_);
  not (_02316_, _01488_);
  and (_02317_, _38013_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02318_, _02208_, _36695_);
  and (_02319_, _01500_, _42340_);
  and (_02320_, _01496_, _01545_);
  or (_02321_, _02320_, _02319_);
  or (_02322_, _01599_, _01550_);
  not (_02323_, _01635_);
  nor (_02324_, _02323_, _01600_);
  and (_02325_, _02324_, _02322_);
  or (_02326_, _02325_, _02321_);
  or (_02327_, _02326_, _02318_);
  or (_02328_, _02327_, _02317_);
  or (_02329_, _02328_, _02316_);
  and (_38847_, _02329_, _02315_);
  or (_02330_, _01542_, _01543_);
  nor (_02331_, _02330_, _01601_);
  and (_02332_, _02330_, _01601_);
  or (_02333_, _02332_, _02331_);
  or (_02334_, _02333_, _02323_);
  and (_02335_, _02208_, _31111_);
  and (_02336_, _01500_, _42077_);
  and (_02337_, _01496_, _01539_);
  and (_02338_, _38013_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_02339_, _02338_, _02337_);
  or (_02340_, _02339_, _02336_);
  nor (_02341_, _02340_, _02335_);
  and (_02342_, _02341_, _02334_);
  nand (_02343_, _02342_, _01488_);
  nor (_02344_, _02312_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02345_, _02312_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_02346_, _02345_, _02344_);
  or (_02347_, _02346_, _01488_);
  and (_02348_, _02347_, _42545_);
  and (_38848_, _02348_, _02343_);
  not (_02349_, _38013_);
  nor (_02350_, _02349_, _32265_);
  not (_02352_, _38325_);
  and (_02353_, _01491_, _02352_);
  and (_02354_, _01603_, _38208_);
  nor (_02355_, _01603_, _38208_);
  nor (_02356_, _02355_, _02354_);
  nand (_02357_, _02356_, _01609_);
  or (_02358_, _02356_, _01609_);
  and (_02359_, _02358_, _02264_);
  and (_02360_, _02359_, _02357_);
  and (_02361_, _01500_, _00680_);
  and (_02362_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_02363_, _01496_, _42286_);
  or (_02364_, _02363_, _02362_);
  nor (_02365_, _02364_, _02361_);
  nand (_02366_, _02365_, _01488_);
  or (_02367_, _02366_, _02360_);
  or (_02368_, _02367_, _02353_);
  or (_02369_, _02368_, _02350_);
  or (_02370_, _02345_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_02371_, _01654_, _01651_);
  and (_02372_, _02371_, _02370_);
  or (_02373_, _02372_, _01488_);
  and (_02374_, _02373_, _42545_);
  and (_38850_, _02374_, _02369_);
  nor (_02375_, _02349_, _32907_);
  and (_02376_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02377_, _02376_, _01609_);
  and (_02378_, _01610_, _01541_);
  nor (_02379_, _02378_, _02377_);
  nand (_02380_, _02379_, _38214_);
  or (_02381_, _02379_, _38214_);
  and (_02382_, _02381_, _02264_);
  and (_02383_, _02382_, _02380_);
  not (_02384_, _38356_);
  and (_02385_, _01491_, _02384_);
  and (_02386_, _01500_, _00669_);
  and (_02387_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_02388_, _01496_, _42191_);
  or (_02389_, _02388_, _02387_);
  or (_02390_, _02389_, _02386_);
  nor (_02391_, _02390_, _02385_);
  nand (_02392_, _02391_, _01488_);
  or (_02393_, _02392_, _02383_);
  or (_02394_, _02393_, _02375_);
  nand (_02395_, _02371_, _01676_);
  or (_02396_, _02371_, _01676_);
  and (_02397_, _02396_, _02395_);
  or (_02398_, _02397_, _01488_);
  and (_02399_, _02398_, _42545_);
  and (_38851_, _02399_, _02394_);
  and (_02400_, _01611_, _01541_);
  and (_02401_, _02377_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_02402_, _02401_, _02400_);
  nand (_02403_, _02402_, _38219_);
  or (_02404_, _02402_, _38219_);
  and (_02405_, _02404_, _02264_);
  and (_02406_, _02405_, _02403_);
  nor (_02407_, _02349_, _33582_);
  not (_02408_, _38386_);
  and (_02409_, _01491_, _02408_);
  and (_02410_, _01500_, _00679_);
  and (_02411_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_02412_, _01496_, _42437_);
  or (_02413_, _02412_, _02411_);
  or (_02414_, _02413_, _02410_);
  nor (_02415_, _02414_, _02409_);
  nand (_02416_, _02415_, _01488_);
  or (_02417_, _02416_, _02407_);
  or (_02418_, _02417_, _02406_);
  nor (_02419_, _01656_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_02420_, _02419_, _01657_);
  or (_02421_, _02420_, _01488_);
  and (_02422_, _02421_, _42545_);
  and (_38852_, _02422_, _02418_);
  nor (_02423_, _02349_, _34333_);
  and (_02424_, _01604_, _01609_);
  and (_02425_, _01612_, _01541_);
  nor (_02426_, _02425_, _02424_);
  nand (_02427_, _02426_, _38204_);
  or (_02428_, _02426_, _38204_);
  and (_02429_, _02428_, _02264_);
  and (_02430_, _02429_, _02427_);
  not (_02431_, _38439_);
  and (_02432_, _01491_, _02431_);
  nor (_02433_, _01509_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_02434_, _02433_, _01510_);
  and (_02435_, _02434_, _01500_);
  and (_02436_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_02437_, _01496_, _42239_);
  or (_02438_, _02437_, _02436_);
  or (_02439_, _02438_, _02435_);
  nor (_02440_, _02439_, _02432_);
  nand (_02441_, _02440_, _01488_);
  or (_02442_, _02441_, _02430_);
  or (_02443_, _02442_, _02423_);
  nor (_02444_, _01657_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02445_, _02444_, _01658_);
  or (_02446_, _02445_, _01488_);
  and (_02447_, _02446_, _42545_);
  and (_38853_, _02447_, _02443_);
  and (_02448_, _01605_, _01609_);
  and (_02449_, _01613_, _01541_);
  nor (_02450_, _02449_, _02448_);
  nand (_02451_, _02450_, _38225_);
  or (_02452_, _02450_, _38225_);
  and (_02453_, _02452_, _02264_);
  and (_02454_, _02453_, _02451_);
  nor (_02455_, _02349_, _35128_);
  not (_02456_, _38472_);
  and (_02457_, _01491_, _02456_);
  nor (_02458_, _01510_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02459_, _02458_, _01511_);
  and (_02460_, _02459_, _01500_);
  and (_02461_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_02462_, _01496_, _42143_);
  or (_02463_, _02462_, _02461_);
  or (_02464_, _02463_, _02460_);
  nor (_02465_, _02464_, _02457_);
  nand (_02466_, _02465_, _01488_);
  or (_02467_, _02466_, _02455_);
  or (_02468_, _02467_, _02454_);
  nor (_02469_, _01658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_02470_, _01658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02471_, _02470_, _02469_);
  or (_02472_, _02471_, _01488_);
  and (_02473_, _02472_, _42545_);
  and (_38854_, _02473_, _02468_);
  and (_02474_, _01606_, _01609_);
  and (_02475_, _02449_, _38225_);
  nor (_02476_, _02475_, _02474_);
  nand (_02477_, _02476_, _38230_);
  or (_02478_, _02476_, _38230_);
  and (_02479_, _02478_, _02264_);
  and (_02480_, _02479_, _02477_);
  nor (_02481_, _02349_, _35956_);
  not (_02482_, _38537_);
  and (_02483_, _01491_, _02482_);
  nor (_02484_, _01511_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_02485_, _02484_, _01512_);
  and (_02486_, _02485_, _01500_);
  and (_02487_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_02488_, _01496_, _42368_);
  or (_02489_, _02488_, _02487_);
  or (_02490_, _02489_, _02486_);
  nor (_02491_, _02490_, _02483_);
  nand (_02492_, _02491_, _01488_);
  or (_02493_, _02492_, _02481_);
  or (_02494_, _02493_, _02480_);
  or (_02495_, _02470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_02496_, _02470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_02497_, _02496_, _02495_);
  or (_02498_, _02497_, _01488_);
  and (_02499_, _02498_, _42545_);
  and (_38855_, _02499_, _02494_);
  or (_02500_, _01617_, _38235_);
  nand (_02501_, _01617_, _38235_);
  nand (_02502_, _02501_, _02500_);
  and (_02503_, _02502_, _02264_);
  or (_02504_, _02349_, _36684_);
  nand (_02505_, _01491_, _38563_);
  or (_02506_, _01512_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02507_, _02506_, _01513_);
  nand (_02508_, _02507_, _01500_);
  nand (_02509_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_02510_, _01496_, _42340_);
  and (_02511_, _02510_, _02509_);
  and (_02512_, _02511_, _02508_);
  and (_02513_, _02512_, _02505_);
  and (_02514_, _02513_, _01488_);
  nand (_02515_, _02514_, _02504_);
  or (_02516_, _02515_, _02503_);
  nor (_02517_, _01659_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_02518_, _02517_, _01660_);
  or (_02519_, _02518_, _01488_);
  and (_02520_, _02519_, _42545_);
  and (_38856_, _02520_, _02516_);
  and (_02521_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_02522_, _01850_, _01848_);
  nor (_02523_, _02522_, _01851_);
  or (_02524_, _02523_, _01670_);
  or (_02525_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_02526_, _02525_, _01884_);
  and (_02527_, _02526_, _02524_);
  or (_38857_, _02527_, _02521_);
  or (_02528_, _01853_, _01851_);
  and (_02529_, _02528_, _01854_);
  or (_02530_, _02529_, _01670_);
  or (_02531_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_02532_, _02531_, _01884_);
  and (_02533_, _02532_, _02530_);
  and (_02534_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_38858_, _02534_, _02533_);
  and (_02535_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02536_, _01858_, _01856_);
  nor (_02537_, _02536_, _01859_);
  or (_02538_, _02537_, _01670_);
  or (_02539_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_02540_, _02539_, _01884_);
  and (_02541_, _02540_, _02538_);
  or (_38859_, _02541_, _02535_);
  and (_02543_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02544_, _01859_, _01753_);
  nor (_02545_, _02544_, _01860_);
  or (_02546_, _02545_, _01670_);
  or (_02547_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_02548_, _02547_, _01884_);
  and (_02549_, _02548_, _02546_);
  or (_38861_, _02549_, _02543_);
  and (_02550_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02551_, _01863_, _01860_);
  nor (_02552_, _02551_, _01864_);
  or (_02553_, _02552_, _01670_);
  or (_02554_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_02555_, _02554_, _01884_);
  and (_02556_, _02555_, _02553_);
  or (_38862_, _02556_, _02550_);
  or (_02557_, _01864_, _01748_);
  nor (_02558_, _01670_, _01865_);
  and (_02559_, _02558_, _02557_);
  nor (_02560_, _01669_, _02002_);
  or (_02561_, _02560_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02562_, _02561_, _02559_);
  or (_02563_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _36922_);
  and (_02564_, _02563_, _42545_);
  and (_38863_, _02564_, _02562_);
  nor (_02566_, _01865_, _01745_);
  nor (_02567_, _02566_, _01866_);
  or (_02568_, _02567_, _01670_);
  or (_02569_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_02570_, _02569_, _01884_);
  and (_02571_, _02570_, _02568_);
  and (_02572_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_38864_, _02572_, _02571_);
  nor (_02574_, _01866_, _01742_);
  nor (_02575_, _02574_, _01867_);
  or (_02576_, _02575_, _01670_);
  or (_02577_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_02578_, _02577_, _01884_);
  and (_02579_, _02578_, _02576_);
  and (_02580_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_38865_, _02580_, _02579_);
  or (_02581_, _01869_, _01867_);
  and (_02582_, _02581_, _01870_);
  or (_02583_, _02582_, _01670_);
  or (_02584_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02585_, _02584_, _01884_);
  and (_02586_, _02585_, _02583_);
  and (_02587_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_38866_, _02587_, _02586_);
  and (_02588_, _01870_, _01737_);
  nor (_02589_, _02588_, _01871_);
  or (_02590_, _02589_, _01670_);
  or (_02591_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_02592_, _02591_, _01884_);
  and (_02593_, _02592_, _02590_);
  and (_02594_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_38867_, _02594_, _02593_);
  nor (_02595_, _01871_, _01735_);
  nor (_02596_, _02595_, _01872_);
  or (_02597_, _02596_, _01670_);
  or (_02598_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_02599_, _02598_, _01884_);
  and (_02600_, _02599_, _02597_);
  and (_02601_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_38868_, _02601_, _02600_);
  and (_02602_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02603_, _01872_, _01730_);
  nor (_02604_, _02603_, _01873_);
  or (_02605_, _02604_, _01670_);
  or (_02606_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_02607_, _02606_, _01884_);
  and (_02608_, _02607_, _02605_);
  or (_38869_, _02608_, _02602_);
  nor (_02609_, _01873_, _01726_);
  nor (_02610_, _02609_, _01874_);
  or (_02611_, _02610_, _01670_);
  or (_02612_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02613_, _02612_, _01884_);
  and (_02614_, _02613_, _02611_);
  and (_02615_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_38870_, _02615_, _02614_);
  nor (_02616_, _01874_, _01723_);
  nor (_02618_, _02616_, _01875_);
  or (_02619_, _02618_, _01670_);
  or (_02620_, _01669_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_02621_, _02620_, _01884_);
  and (_02622_, _02621_, _02619_);
  and (_02624_, _01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_38872_, _02624_, _02622_);
  or (_02625_, _01875_, _01718_);
  nor (_02626_, _01670_, _01876_);
  and (_02627_, _02626_, _02625_);
  nor (_02629_, _01669_, _38235_);
  or (_02630_, _02629_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02631_, _02630_, _02627_);
  or (_02632_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _36922_);
  and (_02633_, _02632_, _42545_);
  and (_38873_, _02633_, _02631_);
  and (_02635_, _01894_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_02636_, _02635_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_38874_, _02636_, _42545_);
  and (_02637_, _01894_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_02639_, _02637_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_38875_, _02639_, _42545_);
  and (_02640_, _01894_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_02641_, _02640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_38876_, _02641_, _42545_);
  and (_02643_, _01894_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_02644_, _02643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_38877_, _02644_, _42545_);
  and (_02645_, _01894_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_02646_, _02645_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_38878_, _02646_, _42545_);
  and (_02648_, _01894_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_02650_, _02648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_38879_, _02650_, _42545_);
  and (_02651_, _01894_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_02652_, _02651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_38880_, _02652_, _42545_);
  and (_02653_, _01848_, _36955_);
  nand (_02654_, _02653_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_02656_, _02653_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_02657_, _02656_, _01884_);
  and (_38881_, _02657_, _02654_);
  or (_02659_, _01905_, _01903_);
  and (_02660_, _02659_, _01906_);
  or (_02661_, _02660_, _42060_);
  or (_02663_, _36955_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_02664_, _02663_, _01884_);
  and (_38883_, _02664_, _02661_);
  and (_02666_, _01927_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_02667_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_02668_, _02667_, _38513_);
  or (_38899_, _02668_, _02666_);
  and (_02670_, _01927_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_02671_, _02082_, _38513_);
  or (_38900_, _02671_, _02670_);
  and (_02673_, _01927_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_02674_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_02676_, _02674_, _38513_);
  or (_38901_, _02676_, _02673_);
  and (_02678_, _01927_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_02679_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_02680_, _02679_, _38513_);
  or (_38902_, _02680_, _02678_);
  and (_02681_, _01927_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_02682_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_02683_, _02682_, _38513_);
  or (_38903_, _02683_, _02681_);
  and (_02685_, _01927_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_02686_, _02095_, _38513_);
  or (_38905_, _02686_, _02685_);
  and (_02688_, _01927_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_02689_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_02691_, _02689_, _38513_);
  or (_38906_, _02691_, _02688_);
  and (_38907_, _01935_, _42545_);
  nor (_38908_, _01945_, rst);
  and (_38909_, _01941_, _42545_);
  and (_02693_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02695_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_02696_, _02695_, _02693_);
  and (_38910_, _02696_, _42545_);
  and (_02698_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02699_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_02700_, _02699_, _02698_);
  and (_38911_, _02700_, _42545_);
  and (_02702_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02704_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_02705_, _02704_, _02702_);
  and (_38912_, _02705_, _42545_);
  and (_02706_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02707_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_02709_, _02707_, _02706_);
  and (_38913_, _02709_, _42545_);
  and (_02710_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02712_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_02713_, _02712_, _02710_);
  and (_38914_, _02713_, _42545_);
  and (_02715_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02716_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_02717_, _02716_, _02715_);
  and (_38916_, _02717_, _42545_);
  and (_02719_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02720_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_02722_, _02720_, _02719_);
  and (_38917_, _02722_, _42545_);
  and (_02723_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02725_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_02726_, _02725_, _02723_);
  and (_38918_, _02726_, _42545_);
  and (_02728_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_02729_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_02731_, _02729_, _02728_);
  and (_38919_, _02731_, _42545_);
  and (_02732_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_02733_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_02734_, _02733_, _02732_);
  and (_38920_, _02734_, _42545_);
  and (_02735_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_02738_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_02739_, _02738_, _02735_);
  and (_38921_, _02739_, _42545_);
  and (_02741_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_02742_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_02743_, _02742_, _02741_);
  and (_38922_, _02743_, _42545_);
  and (_02745_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_02746_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_02748_, _02746_, _02745_);
  and (_38923_, _02748_, _42545_);
  and (_02749_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_02751_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_02752_, _02751_, _02749_);
  and (_38924_, _02752_, _42545_);
  and (_02754_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_02755_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_02756_, _02755_, _02754_);
  and (_38925_, _02756_, _42545_);
  and (_02758_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_02760_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_02761_, _02760_, _02758_);
  and (_38927_, _02761_, _42545_);
  and (_02762_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_02764_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_02765_, _02764_, _02762_);
  and (_38928_, _02765_, _42545_);
  and (_02767_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_02768_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_02769_, _02768_, _02767_);
  and (_38929_, _02769_, _42545_);
  and (_02771_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_02772_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_02774_, _02772_, _02771_);
  and (_38930_, _02774_, _42545_);
  and (_02775_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_02777_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_02778_, _02777_, _02775_);
  and (_38931_, _02778_, _42545_);
  and (_02780_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_02781_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_02782_, _02781_, _02780_);
  and (_38932_, _02782_, _42545_);
  and (_02784_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_02786_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_02787_, _02786_, _02784_);
  and (_38933_, _02787_, _42545_);
  and (_02788_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_02790_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_02791_, _02790_, _02788_);
  and (_38934_, _02791_, _42545_);
  and (_02793_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_02794_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_02795_, _02794_, _02793_);
  and (_38935_, _02795_, _42545_);
  and (_02797_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_02798_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_02800_, _02798_, _02797_);
  and (_38936_, _02800_, _42545_);
  and (_02801_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_02803_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_02804_, _02803_, _02801_);
  and (_38938_, _02804_, _42545_);
  and (_02806_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_02807_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_02808_, _02807_, _02806_);
  and (_38939_, _02808_, _42545_);
  and (_02810_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_02812_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_02813_, _02812_, _02810_);
  and (_38940_, _02813_, _42545_);
  and (_02814_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_02816_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_02817_, _02816_, _02814_);
  and (_38941_, _02817_, _42545_);
  and (_02819_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_02820_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_02821_, _02820_, _02819_);
  and (_38942_, _02821_, _42545_);
  and (_02823_, _01949_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_02824_, _01951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_02826_, _02824_, _02823_);
  and (_38943_, _02826_, _42545_);
  and (_02827_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02829_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_02830_, _02829_, _02827_);
  and (_38944_, _02830_, _42545_);
  and (_02832_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02833_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_02834_, _02833_, _02832_);
  and (_38945_, _02834_, _42545_);
  and (_02836_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02838_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_02839_, _02838_, _02836_);
  and (_38946_, _02839_, _42545_);
  and (_02840_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02841_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_02842_, _02841_, _02840_);
  and (_38947_, _02842_, _42545_);
  and (_02844_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02845_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_02846_, _02845_, _02844_);
  and (_38949_, _02846_, _42545_);
  and (_02848_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02849_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_02851_, _02849_, _02848_);
  and (_38950_, _02851_, _42545_);
  and (_02852_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02854_, _01959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_02855_, _02854_, _02852_);
  and (_38951_, _02855_, _42545_);
  and (_02857_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02858_, _42268_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02859_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_02861_, _02859_, _01958_);
  and (_02862_, _02861_, _02858_);
  or (_02863_, _02862_, _02857_);
  and (_38952_, _02863_, _42545_);
  and (_02865_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02867_, _42168_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02868_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_02869_, _02868_, _01958_);
  and (_02870_, _02869_, _02867_);
  or (_02872_, _02870_, _02865_);
  and (_38953_, _02872_, _42545_);
  and (_02873_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02875_, _42418_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02876_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_02877_, _02876_, _01958_);
  and (_02879_, _02877_, _02875_);
  or (_02880_, _02879_, _02873_);
  and (_38954_, _02880_, _42545_);
  and (_02882_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02883_, _42221_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02884_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_02886_, _02884_, _01958_);
  and (_02887_, _02886_, _02883_);
  or (_02888_, _02887_, _02882_);
  and (_38955_, _02888_, _42545_);
  and (_02890_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02891_, _42117_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02893_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_02894_, _02893_, _01958_);
  and (_02896_, _02894_, _02891_);
  or (_02897_, _02896_, _02890_);
  and (_38956_, _02897_, _42545_);
  and (_02898_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02900_, _42388_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02901_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_02902_, _02901_, _01958_);
  and (_02904_, _02902_, _02900_);
  or (_02905_, _02904_, _02898_);
  and (_38957_, _02905_, _42545_);
  and (_02907_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02908_, _42321_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02909_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_02911_, _02909_, _01958_);
  and (_02912_, _02911_, _02908_);
  or (_02913_, _02912_, _02907_);
  and (_38958_, _02913_, _42545_);
  and (_02916_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02917_, _42054_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02919_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_02920_, _02919_, _01958_);
  and (_02921_, _02920_, _02917_);
  or (_02923_, _02921_, _02916_);
  and (_38960_, _02923_, _42545_);
  and (_02925_, _01965_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_02926_, _02925_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02927_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _01958_);
  and (_02929_, _02927_, _42545_);
  and (_38961_, _02929_, _02926_);
  and (_02931_, _01965_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_02932_, _02931_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02934_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _01958_);
  and (_02935_, _02934_, _42545_);
  and (_38962_, _02935_, _02932_);
  and (_02937_, _01965_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_02938_, _02937_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02939_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _01958_);
  and (_02941_, _02939_, _42545_);
  and (_38963_, _02941_, _02938_);
  and (_02942_, _01965_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_02944_, _02942_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02945_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _01958_);
  and (_02946_, _02945_, _42545_);
  and (_38964_, _02946_, _02944_);
  and (_02948_, _01965_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_02949_, _02948_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02951_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _01958_);
  and (_02953_, _02951_, _42545_);
  and (_38965_, _02953_, _02949_);
  and (_02955_, _01965_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_02956_, _02955_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02957_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _01958_);
  and (_02958_, _02957_, _42545_);
  and (_38966_, _02958_, _02956_);
  and (_02960_, _01965_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_02961_, _02960_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02963_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _01958_);
  and (_02965_, _02963_, _42545_);
  and (_38967_, _02965_, _02961_);
  nand (_02967_, _01972_, _32265_);
  or (_02968_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_02969_, _02968_, _42545_);
  and (_38968_, _02969_, _02967_);
  nand (_02971_, _01972_, _32907_);
  or (_02972_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_02974_, _02972_, _42545_);
  and (_38969_, _02974_, _02971_);
  nand (_02976_, _01972_, _33582_);
  or (_02978_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_02979_, _02978_, _42545_);
  and (_38971_, _02979_, _02976_);
  nand (_02981_, _01972_, _34333_);
  or (_02982_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_02984_, _02982_, _42545_);
  and (_38972_, _02984_, _02981_);
  nand (_02985_, _01972_, _35128_);
  or (_02986_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_02988_, _02986_, _42545_);
  and (_38973_, _02988_, _02985_);
  nand (_02989_, _01972_, _35956_);
  or (_02991_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_02992_, _02991_, _42545_);
  and (_38974_, _02992_, _02989_);
  nand (_02994_, _01972_, _36684_);
  or (_02995_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_02996_, _02995_, _42545_);
  and (_38975_, _02996_, _02994_);
  or (_02999_, _01977_, _31111_);
  or (_03000_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_03002_, _03000_, _42545_);
  and (_38976_, _03002_, _02999_);
  nand (_03003_, _01972_, _38325_);
  or (_03005_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_03006_, _03005_, _42545_);
  and (_38977_, _03006_, _03003_);
  nand (_03008_, _01972_, _38356_);
  or (_03009_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_03012_, _03009_, _42545_);
  and (_38978_, _03012_, _03008_);
  nand (_03013_, _01972_, _38386_);
  or (_03014_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_03016_, _03014_, _42545_);
  and (_38979_, _03016_, _03013_);
  nand (_03017_, _01972_, _38439_);
  or (_03019_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_03020_, _03019_, _42545_);
  and (_38980_, _03020_, _03017_);
  nand (_03023_, _01972_, _38472_);
  or (_03024_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_03025_, _03024_, _42545_);
  and (_38982_, _03025_, _03023_);
  nand (_03027_, _01972_, _38537_);
  or (_03028_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_03030_, _03028_, _42545_);
  and (_38983_, _03030_, _03027_);
  or (_03031_, _01977_, _38563_);
  or (_03033_, _01972_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_03035_, _03033_, _42545_);
  and (_38984_, _03035_, _03031_);
  nor (_39204_, _42095_, rst);
  and (_03037_, _41996_, _41990_);
  nand (_03039_, _03037_, _38146_);
  or (_03040_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_03041_, _03040_, _42545_);
  and (_39205_, _03041_, _03039_);
  not (_03043_, _41997_);
  nor (_03044_, _03043_, _38146_);
  and (_03046_, _03043_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03048_, _03046_, _41991_);
  or (_03049_, _03048_, _03044_);
  or (_03050_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03052_, _03050_, _42545_);
  and (_39206_, _03052_, _03049_);
  and (_03053_, _42000_, _41990_);
  not (_03055_, _03053_);
  nor (_03056_, _03055_, _38146_);
  nand (_03057_, _41998_, _41990_);
  or (_03060_, _03057_, _42002_);
  and (_03061_, _03060_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_03062_, _03061_, _03056_);
  and (_39207_, _03062_, _42545_);
  and (_03064_, _41994_, _41990_);
  not (_03065_, _03064_);
  and (_03067_, _03065_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_03068_, _03065_, _38146_);
  or (_03069_, _03068_, _03067_);
  and (_39209_, _03069_, _42545_);
  or (_03071_, _41994_, _42000_);
  or (_03072_, _03071_, _41997_);
  nor (_03073_, _42007_, _42004_);
  or (_03074_, _41996_, _41991_);
  or (_03075_, _03074_, _03073_);
  or (_03076_, _03075_, _03072_);
  and (_03077_, _03076_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_03078_, _42007_, _41990_);
  not (_03079_, _03078_);
  nor (_03080_, _03079_, _38146_);
  or (_03082_, _03080_, _03077_);
  and (_39210_, _03082_, _42545_);
  and (_03083_, _42009_, _41995_);
  and (_03084_, _03083_, _42002_);
  or (_03085_, _03057_, _03084_);
  or (_03086_, _42007_, _03071_);
  and (_03087_, _03086_, _41990_);
  or (_03088_, _03087_, _03085_);
  and (_03089_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_03090_, _42008_, _41990_);
  and (_03092_, _03090_, _41533_);
  or (_03093_, _03092_, _03089_);
  and (_39211_, _03093_, _42545_);
  nand (_03094_, _42013_, _03084_);
  and (_03095_, _03094_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_03096_, _42006_, _41990_);
  and (_03097_, _03096_, _41533_);
  or (_03098_, _03097_, _03095_);
  and (_39212_, _03098_, _42545_);
  or (_03099_, _42016_, _42004_);
  and (_03100_, _03099_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_03101_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_03102_, _03101_, _42011_);
  and (_03103_, _41990_, _41052_);
  and (_03104_, _03103_, _42005_);
  not (_03105_, _03104_);
  nor (_03106_, _03105_, _38146_);
  or (_03107_, _03106_, _03102_);
  or (_03108_, _03107_, _03100_);
  and (_39213_, _03108_, _42545_);
  nand (_03109_, _03037_, _38123_);
  or (_03110_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03111_, _03110_, _03109_);
  and (_39304_, _03111_, _42545_);
  nand (_03112_, _03037_, _38115_);
  or (_03113_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_03114_, _03113_, _42545_);
  and (_39305_, _03114_, _03112_);
  nand (_03115_, _03037_, _38108_);
  or (_03116_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_03117_, _03116_, _42545_);
  and (_39306_, _03117_, _03115_);
  nand (_03118_, _03037_, _38100_);
  or (_03119_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_03120_, _03119_, _42545_);
  and (_39307_, _03120_, _03118_);
  nand (_03121_, _03037_, _38092_);
  or (_03122_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_03123_, _03122_, _42545_);
  and (_39308_, _03123_, _03121_);
  nand (_03124_, _03037_, _38085_);
  or (_03125_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_03126_, _03125_, _42545_);
  and (_39309_, _03126_, _03124_);
  nand (_03127_, _03037_, _38078_);
  or (_03128_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_03129_, _03128_, _42545_);
  and (_39310_, _03129_, _03127_);
  nor (_03130_, _41991_, _38123_);
  and (_03131_, _03130_, _41997_);
  nand (_03132_, _41997_, _41990_);
  and (_03133_, _03132_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_03134_, _03133_, _03131_);
  and (_39311_, _03134_, _42545_);
  nor (_03135_, _03043_, _38115_);
  and (_03136_, _03043_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_03137_, _03136_, _41991_);
  or (_03138_, _03137_, _03135_);
  or (_03139_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03140_, _03139_, _42545_);
  and (_39312_, _03140_, _03138_);
  nor (_03141_, _03043_, _38108_);
  and (_03142_, _03043_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_03143_, _03142_, _41991_);
  or (_03144_, _03143_, _03141_);
  or (_03145_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_03146_, _03145_, _42545_);
  and (_39313_, _03146_, _03144_);
  nor (_03147_, _03043_, _38100_);
  and (_03148_, _03043_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03149_, _03148_, _41991_);
  or (_03150_, _03149_, _03147_);
  or (_03151_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03152_, _03151_, _42545_);
  and (_39315_, _03152_, _03150_);
  nor (_03153_, _03043_, _38092_);
  and (_03154_, _03043_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_03155_, _03154_, _41991_);
  or (_03156_, _03155_, _03153_);
  or (_03157_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_03158_, _03157_, _42545_);
  and (_39316_, _03158_, _03156_);
  nor (_03159_, _03043_, _38085_);
  and (_03160_, _03043_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_03161_, _03160_, _41991_);
  or (_03162_, _03161_, _03159_);
  or (_03163_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_03164_, _03163_, _42545_);
  and (_39317_, _03164_, _03162_);
  nor (_03165_, _03043_, _38078_);
  and (_03167_, _03043_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03168_, _03167_, _41991_);
  or (_03169_, _03168_, _03165_);
  or (_03170_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03171_, _03170_, _42545_);
  and (_39318_, _03171_, _03169_);
  and (_03172_, _03055_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_03173_, _03130_, _42000_);
  or (_03174_, _03173_, _03172_);
  and (_39319_, _03174_, _42545_);
  nor (_03175_, _03055_, _38115_);
  and (_03176_, _03060_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_03177_, _03176_, _03175_);
  and (_39320_, _03177_, _42545_);
  nor (_03178_, _03055_, _38108_);
  and (_03179_, _03060_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_03180_, _03179_, _03178_);
  and (_39321_, _03180_, _42545_);
  nor (_03181_, _03055_, _38100_);
  and (_03182_, _03060_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_03183_, _03182_, _03181_);
  and (_39322_, _03183_, _42545_);
  and (_03184_, _03055_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_03185_, _03055_, _38092_);
  or (_03186_, _03185_, _03184_);
  and (_39323_, _03186_, _42545_);
  nor (_03187_, _03055_, _38085_);
  and (_03188_, _03060_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_03189_, _03188_, _03187_);
  and (_39324_, _03189_, _42545_);
  nor (_03190_, _03055_, _38078_);
  and (_03191_, _03060_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_03192_, _03191_, _03190_);
  and (_39326_, _03192_, _42545_);
  and (_03195_, _03065_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_03197_, _03130_, _41994_);
  or (_03199_, _03197_, _03195_);
  and (_39327_, _03199_, _42545_);
  and (_03202_, _03065_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_03204_, _03065_, _38115_);
  or (_03205_, _03204_, _03202_);
  and (_39328_, _03205_, _42545_);
  and (_03206_, _03065_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_03207_, _03065_, _38108_);
  or (_03208_, _03207_, _03206_);
  and (_39329_, _03208_, _42545_);
  nor (_03210_, _03065_, _38100_);
  and (_03211_, _03065_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_03213_, _03211_, _03210_);
  and (_39330_, _03213_, _42545_);
  and (_03214_, _03065_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_03216_, _03065_, _38092_);
  or (_03217_, _03216_, _03214_);
  and (_39331_, _03217_, _42545_);
  nor (_03219_, _03065_, _38085_);
  and (_03220_, _03065_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_03221_, _03220_, _03219_);
  and (_39332_, _03221_, _42545_);
  nor (_03223_, _03065_, _38078_);
  and (_03224_, _03065_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_03226_, _03224_, _03223_);
  and (_39333_, _03226_, _42545_);
  and (_03227_, _03075_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_03229_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_03230_, _03229_, _03072_);
  and (_03231_, _03078_, _38124_);
  or (_03233_, _03231_, _03230_);
  or (_03234_, _03233_, _03227_);
  and (_39334_, _03234_, _42545_);
  and (_03236_, _03075_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_03237_, _03079_, _38115_);
  and (_03238_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_03239_, _03238_, _03072_);
  or (_03240_, _03239_, _03237_);
  or (_03241_, _03240_, _03236_);
  and (_39335_, _03241_, _42545_);
  and (_03242_, _03076_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_03243_, _03079_, _38108_);
  or (_03244_, _03243_, _03242_);
  and (_39337_, _03244_, _42545_);
  and (_03245_, _03075_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_03246_, _03079_, _38100_);
  and (_03247_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03248_, _03247_, _03072_);
  or (_03249_, _03248_, _03246_);
  or (_03250_, _03249_, _03245_);
  and (_39338_, _03250_, _42545_);
  and (_03251_, _03075_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_03252_, _03079_, _38092_);
  and (_03253_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03255_, _03253_, _03072_);
  or (_03256_, _03255_, _03252_);
  or (_03258_, _03256_, _03251_);
  and (_39339_, _03258_, _42545_);
  nor (_03259_, _03079_, _38085_);
  and (_03261_, _03079_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_03262_, _03261_, _03259_);
  and (_39340_, _03262_, _42545_);
  nor (_03264_, _03079_, _38078_);
  and (_03265_, _03076_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or (_03266_, _03265_, _03264_);
  and (_39341_, _03266_, _42545_);
  and (_03268_, _03085_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_03269_, _03130_, _42008_);
  and (_03271_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_03272_, _03271_, _03086_);
  or (_03273_, _03272_, _03269_);
  or (_03275_, _03273_, _03268_);
  and (_39342_, _03275_, _42545_);
  and (_03276_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_03278_, _03090_, _42166_);
  or (_03279_, _03278_, _03276_);
  and (_39343_, _03279_, _42545_);
  and (_03281_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_03282_, _03090_, _42416_);
  or (_03283_, _03282_, _03281_);
  and (_39344_, _03283_, _42545_);
  and (_03284_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_03285_, _03090_, _42219_);
  or (_03286_, _03285_, _03284_);
  and (_39345_, _03286_, _42545_);
  and (_03287_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_03288_, _03090_, _42115_);
  or (_03289_, _03288_, _03287_);
  and (_39346_, _03289_, _42545_);
  and (_03290_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_03291_, _03090_, _42386_);
  or (_03292_, _03291_, _03290_);
  and (_39348_, _03292_, _42545_);
  and (_03293_, _03088_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_03294_, _03090_, _40183_);
  or (_03295_, _03294_, _03293_);
  and (_39349_, _03295_, _42545_);
  nand (_03296_, _42013_, _42002_);
  and (_03298_, _03296_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nand (_03299_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor (_03301_, _03299_, _03083_);
  and (_03302_, _03096_, _38124_);
  or (_03303_, _03302_, _03301_);
  or (_03305_, _03303_, _03298_);
  and (_39350_, _03305_, _42545_);
  and (_03306_, _03296_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_03308_, _03096_, _42166_);
  nand (_03309_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_03310_, _03309_, _03083_);
  or (_03312_, _03310_, _03308_);
  or (_03313_, _03312_, _03306_);
  and (_39351_, _03313_, _42545_);
  and (_03315_, _03094_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_03316_, _03096_, _42416_);
  or (_03317_, _03316_, _03315_);
  and (_39352_, _03317_, _42545_);
  and (_03319_, _03296_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_03320_, _03096_, _42219_);
  nand (_03322_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_03323_, _03322_, _03083_);
  or (_03324_, _03323_, _03320_);
  or (_03326_, _03324_, _03319_);
  and (_39353_, _03326_, _42545_);
  and (_03327_, _03096_, _42115_);
  nand (_03328_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_03329_, _03328_, _03084_);
  not (_03330_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_03331_, _42013_, _03330_);
  or (_03332_, _03331_, _03329_);
  or (_03333_, _03332_, _03327_);
  and (_39354_, _03333_, _42545_);
  and (_03334_, _03296_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_03335_, _03096_, _42386_);
  nand (_03336_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_03337_, _03336_, _03083_);
  or (_03338_, _03337_, _03335_);
  or (_03339_, _03338_, _03334_);
  and (_39355_, _03339_, _42545_);
  and (_03340_, _03096_, _40183_);
  and (_03341_, _03296_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nand (_03342_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor (_03343_, _03342_, _03083_);
  or (_03345_, _03343_, _03341_);
  or (_03346_, _03345_, _03340_);
  and (_39356_, _03346_, _42545_);
  and (_03348_, _03099_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03349_, _03104_, _38124_);
  and (_03351_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03352_, _03351_, _42011_);
  or (_03353_, _03352_, _03349_);
  or (_03355_, _03353_, _03348_);
  and (_39357_, _03355_, _42545_);
  and (_03356_, _03099_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_03358_, _03105_, _38115_);
  and (_03359_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_03360_, _03359_, _42011_);
  or (_03362_, _03360_, _03358_);
  or (_03363_, _03362_, _03356_);
  and (_39358_, _03363_, _42545_);
  and (_03365_, _03099_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_03366_, _03105_, _38108_);
  and (_03367_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_03369_, _03367_, _42011_);
  or (_03370_, _03369_, _03366_);
  or (_03372_, _03370_, _03365_);
  and (_39359_, _03372_, _42545_);
  and (_03374_, _03099_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_03375_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_03376_, _03375_, _42011_);
  nor (_03377_, _03105_, _38100_);
  or (_03378_, _03377_, _03376_);
  or (_03379_, _03378_, _03374_);
  and (_39360_, _03379_, _42545_);
  and (_03380_, _03105_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_03381_, _03105_, _38092_);
  or (_03382_, _03381_, _03380_);
  and (_39361_, _03382_, _42545_);
  and (_03383_, _03099_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_03384_, _03105_, _38085_);
  and (_03385_, _41990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_03386_, _03385_, _42011_);
  or (_03387_, _03386_, _03384_);
  or (_03388_, _03387_, _03383_);
  and (_39362_, _03388_, _42545_);
  nor (_03389_, _03105_, _38078_);
  or (_03390_, _03105_, _42013_);
  and (_03392_, _03390_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_03393_, _03392_, _03389_);
  and (_39363_, _03393_, _42545_);
  not (_03395_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03396_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_03398_, _03396_, _03395_);
  and (_03399_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _42545_);
  and (_39423_, _03399_, _03398_);
  nor (_03401_, _03398_, rst);
  nand (_03402_, _03396_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03403_, _03396_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03405_, _03403_, _03402_);
  and (_39425_, _03405_, _03401_);
  not (_03406_, _42081_);
  and (_03408_, _42147_, _03406_);
  and (_03409_, _03408_, _42248_);
  nor (_03410_, _42344_, _42397_);
  and (_03412_, _03410_, _03409_);
  and (_03413_, _03412_, _38735_);
  nor (_03414_, _03413_, _01404_);
  not (_03416_, _42294_);
  nor (_03417_, _03416_, _42195_);
  and (_03418_, _03417_, _40183_);
  or (_03420_, _03418_, _42443_);
  nor (_03421_, _42294_, _42195_);
  and (_03422_, _03421_, _41533_);
  and (_03423_, _42294_, _42195_);
  and (_03424_, _03423_, _42115_);
  and (_03425_, _03416_, _42195_);
  and (_03426_, _03425_, _42386_);
  or (_03427_, _03426_, _03424_);
  or (_03428_, _03427_, _03422_);
  or (_03429_, _03428_, _03420_);
  not (_03430_, _42443_);
  and (_03431_, _03417_, _42416_);
  or (_03432_, _03431_, _03430_);
  and (_03433_, _03421_, _42219_);
  and (_03434_, _03423_, _38124_);
  and (_03435_, _03425_, _42166_);
  or (_03436_, _03435_, _03434_);
  or (_03437_, _03436_, _03433_);
  or (_03438_, _03437_, _03432_);
  nand (_03439_, _03438_, _03429_);
  nor (_03440_, _03439_, _03414_);
  not (_03442_, _42344_);
  and (_03443_, _03442_, _42397_);
  and (_03445_, _42248_, _42148_);
  and (_03446_, _03445_, _03406_);
  and (_03447_, _03446_, _03443_);
  nor (_03449_, _39015_, _39001_);
  and (_03450_, _39015_, _39001_);
  nor (_03451_, _03450_, _03449_);
  and (_03453_, _38987_, _38817_);
  nor (_03454_, _38987_, _38817_);
  or (_03455_, _03454_, _03453_);
  nor (_03457_, _03455_, _03451_);
  and (_03458_, _03455_, _03451_);
  nor (_03459_, _03458_, _03457_);
  nor (_03461_, _39039_, _39027_);
  and (_03462_, _39039_, _39027_);
  nor (_03463_, _03462_, _03461_);
  not (_03465_, _39052_);
  and (_03466_, _03465_, _38758_);
  nor (_03467_, _03465_, _38758_);
  nor (_03469_, _03467_, _03466_);
  nor (_03470_, _03469_, _03463_);
  and (_03471_, _03469_, _03463_);
  or (_03473_, _03471_, _03470_);
  nor (_03474_, _03473_, _03459_);
  and (_03475_, _03473_, _03459_);
  nor (_03476_, _03475_, _03474_);
  nand (_03477_, _03476_, _42443_);
  or (_03478_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03479_, _03478_, _03423_);
  and (_03480_, _03479_, _03477_);
  and (_03481_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_03482_, _42443_, _38622_);
  or (_03483_, _03482_, _03481_);
  and (_03484_, _03483_, _03421_);
  or (_03485_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_03486_, _03430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03487_, _03486_, _03425_);
  and (_03488_, _03487_, _03485_);
  or (_03489_, _03488_, _03484_);
  or (_03490_, _03430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03491_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_03492_, _03491_, _03417_);
  and (_03493_, _03492_, _03490_);
  or (_03495_, _03493_, _03489_);
  or (_03496_, _03495_, _03480_);
  and (_03498_, _03496_, _03447_);
  and (_03499_, _42344_, _42398_);
  nor (_03500_, _00800_, _37969_);
  and (_03502_, _03500_, _00864_);
  and (_03503_, _38030_, _37907_);
  or (_03504_, _03503_, _37940_);
  nor (_03506_, _03504_, _38022_);
  and (_03507_, _37947_, _37857_);
  or (_03508_, _03507_, _00802_);
  or (_03510_, _03508_, _00869_);
  nor (_03511_, _03510_, _38002_);
  and (_03512_, _03511_, _03506_);
  and (_03514_, _03512_, _01141_);
  and (_03515_, _03514_, _03502_);
  and (_03516_, _03515_, _37991_);
  nor (_03518_, _03516_, _36912_);
  nor (_03519_, _03518_, p3_in[0]);
  and (_03520_, _03518_, _39461_);
  nor (_03522_, _03520_, _03519_);
  or (_03523_, _03522_, _03430_);
  or (_03524_, _03518_, p3_in[4]);
  not (_03526_, _03518_);
  or (_03527_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03528_, _03527_, _03524_);
  or (_03529_, _03528_, _42443_);
  and (_03530_, _03529_, _03423_);
  and (_03531_, _03530_, _03523_);
  or (_03532_, _03518_, p3_in[5]);
  or (_03533_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03534_, _03533_, _03532_);
  and (_03535_, _03534_, _03430_);
  or (_03536_, _03518_, p3_in[1]);
  or (_03537_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03538_, _03537_, _03536_);
  and (_03539_, _03538_, _42443_);
  or (_03540_, _03539_, _03535_);
  and (_03541_, _03540_, _03425_);
  or (_03542_, _03541_, _03531_);
  or (_03543_, _03518_, p3_in[3]);
  or (_03544_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03545_, _03544_, _03543_);
  or (_03546_, _03545_, _03430_);
  nor (_03548_, _03518_, p3_in[7]);
  and (_03549_, _03518_, _39106_);
  nor (_03551_, _03549_, _03548_);
  or (_03552_, _03551_, _42443_);
  and (_03553_, _03552_, _03421_);
  and (_03555_, _03553_, _03546_);
  or (_03556_, _03518_, p3_in[6]);
  or (_03557_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03559_, _03557_, _03556_);
  and (_03560_, _03559_, _03430_);
  or (_03561_, _03518_, p3_in[2]);
  or (_03563_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03564_, _03563_, _03561_);
  and (_03565_, _03564_, _42443_);
  or (_03567_, _03565_, _03560_);
  and (_03568_, _03567_, _03417_);
  or (_03569_, _03568_, _03555_);
  or (_03571_, _03569_, _03542_);
  nand (_03572_, _03571_, _03499_);
  nand (_03573_, _03572_, _03446_);
  and (_03575_, _03408_, _42249_);
  and (_03576_, _03575_, _03443_);
  not (_03577_, _03443_);
  nand (_03579_, _03577_, _03409_);
  nor (_03580_, _42248_, _42081_);
  and (_03581_, _03580_, _42344_);
  nor (_03582_, _03581_, _28834_);
  nand (_03583_, _03582_, _03579_);
  nor (_03584_, _03583_, _03576_);
  or (_03585_, _03584_, _03446_);
  and (_03586_, _03585_, _03573_);
  and (_03587_, _42344_, _42397_);
  and (_03588_, _03580_, _42148_);
  and (_03589_, _03588_, _03587_);
  and (_03590_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_03591_, _42443_, _40942_);
  or (_03592_, _03591_, _03590_);
  and (_03593_, _03592_, _03421_);
  and (_03594_, _03430_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_03595_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03596_, _03595_, _03594_);
  and (_03597_, _03596_, _03417_);
  or (_03598_, _03597_, _03593_);
  and (_03599_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_03601_, _42443_, _40967_);
  or (_03602_, _03601_, _03599_);
  and (_03605_, _03602_, _03423_);
  and (_03606_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor (_03607_, _42443_, _41368_);
  or (_03609_, _03607_, _03606_);
  and (_03610_, _03609_, _03425_);
  or (_03611_, _03610_, _03605_);
  or (_03613_, _03611_, _03598_);
  and (_03614_, _03613_, _03589_);
  nor (_03615_, _42397_, _42147_);
  and (_03617_, _03615_, _03581_);
  or (_03618_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand (_03619_, _42443_, _40543_);
  and (_03621_, _03619_, _03421_);
  and (_03622_, _03621_, _03618_);
  and (_03623_, _03430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03625_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03626_, _03625_, _03623_);
  and (_03627_, _03626_, _03417_);
  or (_03629_, _03627_, _03622_);
  and (_03630_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_03631_, _42443_, _40530_);
  or (_03633_, _03631_, _03630_);
  and (_03634_, _03633_, _03423_);
  and (_03635_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_03636_, _42443_, _40534_);
  or (_03637_, _03636_, _03635_);
  and (_03638_, _03637_, _03425_);
  or (_03639_, _03638_, _03634_);
  or (_03640_, _03639_, _03629_);
  and (_03641_, _03640_, _03617_);
  and (_03642_, _03446_, _03410_);
  and (_03643_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_03644_, _42443_, _35161_);
  or (_03645_, _03644_, _03643_);
  and (_03646_, _03645_, _03423_);
  and (_03647_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_03648_, _42443_, _35988_);
  or (_03649_, _03648_, _03647_);
  and (_03650_, _03649_, _03425_);
  or (_03651_, _03650_, _03646_);
  and (_03652_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_03653_, _42443_, _31188_);
  or (_03655_, _03653_, _03652_);
  and (_03656_, _03655_, _03421_);
  nor (_03658_, _42443_, _36716_);
  and (_03659_, _42443_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03660_, _03659_, _03658_);
  and (_03662_, _03660_, _03417_);
  or (_03663_, _03662_, _03656_);
  or (_03664_, _03663_, _03651_);
  and (_03666_, _03664_, _03642_);
  or (_03667_, _03666_, _03641_);
  or (_03668_, _03667_, _03614_);
  and (_03670_, _01421_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_03671_, _03417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03672_, _03671_, _42443_);
  and (_03674_, _03421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03675_, _03423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03676_, _03425_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_03678_, _03676_, _03675_);
  or (_03679_, _03678_, _03674_);
  or (_03680_, _03679_, _03672_);
  and (_03682_, _03417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03683_, _03682_, _03430_);
  and (_03684_, _03421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_03686_, _03423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03687_, _03425_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03688_, _03687_, _03686_);
  or (_03689_, _03688_, _03684_);
  or (_03690_, _03689_, _03683_);
  and (_03691_, _03690_, _03576_);
  and (_03692_, _03691_, _03680_);
  or (_03693_, _03692_, _03670_);
  or (_03694_, _03693_, _03668_);
  or (_03695_, _03694_, _03586_);
  and (_03696_, _03423_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03697_, _03417_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03698_, _03697_, _03696_);
  and (_03699_, _03421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03700_, _03425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03701_, _03700_, _03699_);
  or (_03702_, _03701_, _03698_);
  and (_03703_, _03702_, _03430_);
  and (_03704_, _03423_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_03705_, _03417_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03706_, _03705_, _03704_);
  and (_03708_, _03421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_03709_, _03425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03711_, _03709_, _03708_);
  or (_03712_, _03711_, _03706_);
  and (_03713_, _03712_, _42443_);
  or (_03715_, _03713_, _03703_);
  and (_03716_, _03715_, _03410_);
  nor (_03717_, _03518_, p2_in[0]);
  and (_03719_, _03518_, _39371_);
  nor (_03720_, _03719_, _03717_);
  or (_03721_, _03720_, _03430_);
  or (_03723_, _03518_, p2_in[4]);
  or (_03724_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03725_, _03724_, _03723_);
  or (_03727_, _03725_, _42443_);
  and (_03728_, _03727_, _03423_);
  and (_03729_, _03728_, _03721_);
  or (_03731_, _03518_, p2_in[5]);
  or (_03732_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03733_, _03732_, _03731_);
  and (_03735_, _03733_, _03430_);
  or (_03736_, _03518_, p2_in[1]);
  or (_03737_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03739_, _03737_, _03736_);
  and (_03740_, _03739_, _42443_);
  or (_03741_, _03740_, _03735_);
  and (_03742_, _03741_, _03425_);
  or (_03743_, _03742_, _03729_);
  or (_03744_, _03518_, p2_in[3]);
  or (_03745_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03746_, _03745_, _03744_);
  or (_03747_, _03746_, _03430_);
  nor (_03748_, _03518_, p2_in[7]);
  and (_03749_, _03518_, _39096_);
  nor (_03750_, _03749_, _03748_);
  or (_03751_, _03750_, _42443_);
  and (_03752_, _03751_, _03421_);
  and (_03753_, _03752_, _03747_);
  or (_03754_, _03518_, p2_in[6]);
  or (_03755_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03756_, _03755_, _03754_);
  and (_03757_, _03756_, _03430_);
  or (_03758_, _03518_, p2_in[2]);
  or (_03759_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03761_, _03759_, _03758_);
  and (_03762_, _03761_, _42443_);
  or (_03764_, _03762_, _03757_);
  and (_03765_, _03764_, _03417_);
  or (_03766_, _03765_, _03753_);
  or (_03768_, _03766_, _03743_);
  and (_03769_, _03768_, _03499_);
  or (_03770_, _03769_, _03716_);
  and (_03772_, _03770_, _03409_);
  and (_03773_, _03421_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03774_, _03425_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03776_, _03774_, _03773_);
  and (_03777_, _03417_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_03778_, _03423_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_03780_, _03778_, _03777_);
  or (_03781_, _03780_, _03776_);
  and (_03782_, _03781_, _03587_);
  and (_03784_, _03417_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_03785_, _03423_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_03786_, _03785_, _03784_);
  and (_03788_, _03421_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03789_, _03425_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_03790_, _03789_, _03788_);
  or (_03792_, _03790_, _03786_);
  and (_03793_, _03792_, _03499_);
  or (_03794_, _03793_, _03430_);
  or (_03795_, _03794_, _03782_);
  and (_03796_, _03417_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03797_, _03423_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_03798_, _03797_, _03796_);
  and (_03799_, _03421_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03800_, _03425_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_03801_, _03800_, _03799_);
  or (_03802_, _03801_, _03798_);
  and (_03803_, _03802_, _03499_);
  and (_03804_, _03417_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03805_, _03423_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_03806_, _03805_, _03804_);
  and (_03807_, _03421_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03808_, _03425_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03809_, _03808_, _03807_);
  or (_03810_, _03809_, _03806_);
  and (_03811_, _03810_, _03587_);
  or (_03812_, _03811_, _42443_);
  or (_03814_, _03812_, _03803_);
  and (_03815_, _03814_, _03575_);
  and (_03817_, _03815_, _03795_);
  or (_03818_, _03518_, p0_in[2]);
  or (_03819_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03821_, _03819_, _03818_);
  and (_03822_, _03821_, _03417_);
  nor (_03823_, _03518_, p0_in[0]);
  and (_03825_, _03518_, _39129_);
  nor (_03826_, _03825_, _03823_);
  and (_03827_, _03826_, _03423_);
  or (_03829_, _03827_, _03822_);
  or (_03830_, _03518_, p0_in[3]);
  or (_03831_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03833_, _03831_, _03830_);
  and (_03834_, _03833_, _03421_);
  or (_03835_, _03518_, p0_in[1]);
  or (_03837_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03838_, _03837_, _03835_);
  and (_03839_, _03838_, _03425_);
  or (_03841_, _03839_, _03834_);
  or (_03842_, _03841_, _03829_);
  and (_03843_, _03842_, _03409_);
  or (_03845_, _03518_, p1_in[3]);
  or (_03846_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03847_, _03846_, _03845_);
  and (_03849_, _03847_, _03421_);
  or (_03850_, _03518_, p1_in[1]);
  or (_03851_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03852_, _03851_, _03850_);
  and (_03853_, _03852_, _03425_);
  or (_03854_, _03853_, _03849_);
  or (_03855_, _03518_, p1_in[2]);
  or (_03856_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03857_, _03856_, _03855_);
  and (_03858_, _03857_, _03417_);
  nor (_03859_, _03518_, p1_in[0]);
  and (_03860_, _03518_, _39232_);
  nor (_03861_, _03860_, _03859_);
  and (_03862_, _03861_, _03423_);
  or (_03863_, _03862_, _03858_);
  or (_03864_, _03863_, _03854_);
  and (_03865_, _03864_, _03446_);
  or (_03866_, _03865_, _03843_);
  and (_03868_, _03866_, _42443_);
  or (_03869_, _03518_, p1_in[6]);
  or (_03871_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03872_, _03871_, _03869_);
  and (_03873_, _03872_, _03417_);
  or (_03875_, _03518_, p1_in[4]);
  or (_03876_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03877_, _03876_, _03875_);
  and (_03879_, _03877_, _03423_);
  or (_03880_, _03879_, _03873_);
  nor (_03881_, _03518_, p1_in[7]);
  and (_03883_, _03518_, _39081_);
  nor (_03884_, _03883_, _03881_);
  and (_03885_, _03884_, _03421_);
  or (_03887_, _03518_, p1_in[5]);
  or (_03888_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03889_, _03888_, _03887_);
  and (_03891_, _03889_, _03425_);
  or (_03892_, _03891_, _03885_);
  or (_03893_, _03892_, _03880_);
  and (_03895_, _03893_, _03446_);
  or (_03896_, _03518_, p0_in[6]);
  or (_03897_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03899_, _03897_, _03896_);
  and (_03900_, _03899_, _03417_);
  or (_03901_, _03518_, p0_in[4]);
  or (_03902_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03903_, _03902_, _03901_);
  and (_03904_, _03903_, _03423_);
  or (_03905_, _03904_, _03900_);
  nor (_03906_, _03518_, p0_in[7]);
  and (_03907_, _03518_, _39065_);
  nor (_03908_, _03907_, _03906_);
  and (_03909_, _03908_, _03421_);
  or (_03910_, _03518_, p0_in[5]);
  or (_03911_, _03526_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03912_, _03911_, _03910_);
  and (_03913_, _03912_, _03425_);
  or (_03914_, _03913_, _03909_);
  or (_03915_, _03914_, _03905_);
  and (_03916_, _03915_, _03409_);
  or (_03917_, _03916_, _03895_);
  and (_03918_, _03917_, _03430_);
  or (_03919_, _03918_, _03868_);
  and (_03921_, _03919_, _03587_);
  or (_03922_, _03921_, _03817_);
  or (_03924_, _03922_, _03772_);
  or (_03925_, _03924_, _03695_);
  or (_03926_, _03925_, _03498_);
  nand (_03928_, _03670_, _31732_);
  and (_03929_, _03928_, _03414_);
  and (_03930_, _03929_, _03926_);
  or (_03932_, _03930_, _03440_);
  and (_39426_, _03932_, _42545_);
  and (_03933_, _03587_, _03408_);
  and (_03935_, _42248_, _42443_);
  and (_03936_, _03935_, _03421_);
  and (_03937_, _03936_, _03933_);
  and (_03939_, _03937_, _38194_);
  and (_03940_, _42397_, _42148_);
  and (_03941_, _03935_, _03423_);
  and (_03943_, _03941_, _03406_);
  and (_03944_, _03943_, _03442_);
  and (_03945_, _03944_, _03940_);
  and (_03947_, _03945_, _38627_);
  and (_03948_, _03410_, _03408_);
  and (_03949_, _03948_, _03941_);
  and (_03951_, _03949_, _38731_);
  or (_03952_, _03951_, _03947_);
  nor (_03953_, _03952_, _03939_);
  nor (_03954_, _03953_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_03955_, _03421_, _03430_);
  not (_03956_, _03955_);
  and (_03957_, _03956_, _38748_);
  and (_03958_, _03957_, _01402_);
  and (_03959_, _03949_, _38735_);
  or (_03960_, _03959_, _01423_);
  or (_03961_, _03960_, _03958_);
  nor (_03962_, _03961_, _03954_);
  and (_03963_, _03933_, _03417_);
  and (_03964_, _03963_, _03935_);
  and (_03965_, _03964_, _38194_);
  or (_03966_, _03965_, rst);
  nor (_39427_, _03966_, _03962_);
  not (_03967_, _03962_);
  nand (_03968_, _03943_, _03577_);
  and (_03969_, _03955_, _42248_);
  and (_03970_, _42344_, _03406_);
  and (_03972_, _03615_, _03970_);
  and (_03973_, _03972_, _03969_);
  and (_03975_, _03443_, _03408_);
  nor (_03976_, _42248_, _42443_);
  and (_03977_, _03976_, _03423_);
  and (_03979_, _03977_, _03975_);
  nor (_03980_, _03979_, _03973_);
  and (_03981_, _03980_, _03968_);
  and (_03983_, _42249_, _42443_);
  and (_03984_, _03983_, _03417_);
  and (_03985_, _03984_, _03975_);
  and (_03987_, _03976_, _03425_);
  and (_03988_, _03987_, _03975_);
  nor (_03989_, _03988_, _03985_);
  and (_03991_, _03983_, _03421_);
  and (_03992_, _03991_, _03975_);
  and (_03993_, _03983_, _03423_);
  and (_03995_, _03499_, _03408_);
  and (_03996_, _03995_, _03993_);
  nor (_03997_, _03996_, _03992_);
  and (_03999_, _03997_, _03989_);
  and (_04000_, _03991_, _03933_);
  and (_04001_, _03983_, _03425_);
  and (_04003_, _03940_, _03970_);
  and (_04004_, _04003_, _04001_);
  nor (_04005_, _04004_, _04000_);
  and (_04006_, _03993_, _03975_);
  and (_04007_, _04003_, _03993_);
  nor (_04008_, _04007_, _04006_);
  and (_04009_, _04008_, _04005_);
  and (_04010_, _04009_, _03999_);
  and (_04011_, _04010_, _03981_);
  and (_04012_, _04001_, _03933_);
  and (_04013_, _03933_, _03425_);
  and (_04014_, _04013_, _03976_);
  nor (_04015_, _04014_, _04012_);
  nand (_04016_, _03983_, _03963_);
  nand (_04017_, _04013_, _03935_);
  and (_04018_, _04017_, _04016_);
  and (_04019_, _04018_, _04015_);
  and (_04020_, _03977_, _03933_);
  nor (_04021_, _04020_, _03937_);
  and (_04022_, _03993_, _03933_);
  and (_04023_, _03969_, _03933_);
  nor (_04024_, _04023_, _04022_);
  and (_04025_, _04024_, _04021_);
  nor (_04026_, _03964_, _03945_);
  and (_04027_, _04026_, _04025_);
  and (_04028_, _04027_, _04019_);
  and (_04029_, _04028_, _04011_);
  nor (_04030_, _04029_, _03967_);
  or (_04031_, _04030_, _20620_);
  nand (_04032_, _03992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_04033_, _04022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_04034_, _04033_, _04032_);
  nand (_04035_, _03973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand (_04036_, _03996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_04037_, _04036_, _04035_);
  and (_04038_, _04037_, _04034_);
  nand (_04039_, _03979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_04040_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_04041_, _04040_, _04039_);
  nand (_04042_, _03985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand (_04043_, _03988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_04044_, _04043_, _04042_);
  and (_04045_, _04044_, _04041_);
  and (_04046_, _04045_, _04038_);
  nand (_04047_, _04012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nand (_04048_, _04000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_04049_, _04048_, _04047_);
  and (_04050_, _03987_, _03933_);
  nand (_04051_, _04050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_04052_, _03984_, _03933_);
  nand (_04053_, _04052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_04054_, _04053_, _04051_);
  and (_04055_, _04054_, _04049_);
  nand (_04056_, _04004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_04057_, _04007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_04058_, _04057_, _04056_);
  nand (_04059_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_04060_, _04023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_04061_, _04060_, _04059_);
  and (_04062_, _04061_, _04058_);
  and (_04063_, _04062_, _04055_);
  and (_04064_, _04063_, _04046_);
  nand (_04065_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand (_04066_, _03964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_04067_, _04066_, _04065_);
  and (_04068_, _03944_, _03615_);
  nand (_04069_, _04068_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_04070_, _03935_, _03425_);
  and (_04071_, _04070_, _03933_);
  nand (_04072_, _04071_, _38148_);
  and (_04073_, _04072_, _04069_);
  and (_04075_, _04073_, _04067_);
  and (_04076_, _03972_, _03941_);
  nand (_04077_, _04076_, _03551_);
  and (_04078_, _03995_, _03941_);
  nand (_04079_, _04078_, _03750_);
  and (_04080_, _04079_, _04077_);
  and (_04081_, _03933_, _03941_);
  nand (_04082_, _04081_, _03908_);
  and (_04083_, _04003_, _03941_);
  nand (_04084_, _04083_, _03884_);
  and (_04085_, _04084_, _04082_);
  and (_04086_, _04085_, _04080_);
  and (_04087_, _04086_, _04075_);
  nand (_04088_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_04089_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_04090_, _04089_, _04088_);
  and (_04091_, _04090_, _04087_);
  nand (_04092_, _04091_, _04064_);
  nand (_04093_, _04092_, _03962_);
  and (_04094_, _04093_, _04031_);
  nor (_04095_, _04094_, _03965_);
  and (_04096_, _03965_, _31111_);
  or (_04097_, _04096_, _04095_);
  and (_39428_, _04097_, _42545_);
  nor (_39505_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_04098_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_04099_, _03396_, rst);
  and (_39506_, _04099_, _04098_);
  nor (_04100_, _03396_, _03395_);
  or (_04101_, _04100_, _03398_);
  and (_04102_, _03402_, _42545_);
  and (_39507_, _04102_, _04101_);
  nand (_04103_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_04104_, _03979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_04105_, _04104_, _04103_);
  nand (_04106_, _03985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_04107_, _03988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_04108_, _04107_, _04106_);
  and (_04109_, _04108_, _04105_);
  nand (_04110_, _04022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_04111_, _03992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_04112_, _04111_, _04110_);
  nand (_04113_, _03973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand (_04114_, _03996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_04115_, _04114_, _04113_);
  and (_04116_, _04115_, _04112_);
  and (_04117_, _04116_, _04109_);
  nand (_04118_, _04000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_04119_, _04012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_04120_, _04119_, _04118_);
  nand (_04121_, _04050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_04122_, _04052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_04123_, _04122_, _04121_);
  and (_04124_, _04123_, _04120_);
  nand (_04125_, _04023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand (_04126_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_04127_, _04126_, _04125_);
  nand (_04128_, _04004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand (_04129_, _04007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_04130_, _04129_, _04128_);
  and (_04131_, _04130_, _04127_);
  and (_04132_, _04131_, _04124_);
  and (_04133_, _04132_, _04117_);
  nand (_04134_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand (_04135_, _03964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_04136_, _04135_, _04134_);
  nand (_04137_, _04068_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_04138_, _04071_, _42289_);
  and (_04139_, _04138_, _04137_);
  and (_04140_, _04139_, _04136_);
  nand (_04141_, _04076_, _03522_);
  nand (_04142_, _04078_, _03720_);
  and (_04143_, _04142_, _04141_);
  nand (_04144_, _04083_, _03861_);
  nand (_04145_, _04081_, _03826_);
  and (_04146_, _04145_, _04144_);
  and (_04147_, _04146_, _04143_);
  and (_04148_, _04147_, _04140_);
  not (_04149_, _03945_);
  or (_04150_, _04149_, _03476_);
  nand (_04151_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_04152_, _04151_, _04150_);
  and (_04153_, _04152_, _04148_);
  and (_04154_, _04153_, _04133_);
  nor (_04155_, _04154_, _03967_);
  nor (_04156_, _04030_, _19460_);
  or (_04157_, _04156_, _03965_);
  or (_04158_, _04157_, _04155_);
  nand (_04159_, _03965_, _32265_);
  and (_04160_, _04159_, _42545_);
  and (_39509_, _04160_, _04158_);
  nand (_04161_, _03965_, _32907_);
  nor (_04162_, _04030_, _20446_);
  and (_04163_, _03979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_04164_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_04165_, _04164_, _04163_);
  and (_04166_, _03985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_04167_, _03988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_04168_, _04167_, _04166_);
  or (_04169_, _04168_, _04165_);
  and (_04171_, _04022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_04172_, _03992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_04173_, _04172_, _04171_);
  and (_04174_, _03996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_04175_, _03973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_04176_, _04175_, _04174_);
  or (_04177_, _04176_, _04173_);
  or (_04178_, _04177_, _04169_);
  and (_04179_, _04000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_04180_, _04012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_04181_, _04180_, _04179_);
  and (_04182_, _04050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_04183_, _04052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_04184_, _04183_, _04182_);
  or (_04185_, _04184_, _04181_);
  and (_04186_, _04004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_04187_, _04007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_04188_, _04187_, _04186_);
  and (_04189_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_04190_, _04023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_04191_, _04190_, _04189_);
  or (_04192_, _04191_, _04188_);
  or (_04193_, _04192_, _04185_);
  or (_04194_, _04193_, _04178_);
  and (_04195_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_04196_, _03964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_04197_, _04196_, _04195_);
  and (_04198_, _04068_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_04199_, _04071_, _42173_);
  or (_04200_, _04199_, _04198_);
  or (_04201_, _04200_, _04197_);
  and (_04202_, _04076_, _03538_);
  and (_04203_, _04078_, _03739_);
  or (_04204_, _04203_, _04202_);
  and (_04205_, _04083_, _03852_);
  and (_04206_, _04081_, _03838_);
  or (_04207_, _04206_, _04205_);
  or (_04208_, _04207_, _04204_);
  or (_04209_, _04208_, _04201_);
  and (_04210_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_04211_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_04212_, _04211_, _04210_);
  or (_04213_, _04212_, _04209_);
  or (_04214_, _04213_, _04194_);
  and (_04215_, _04214_, _03962_);
  or (_04216_, _04215_, _04162_);
  or (_04217_, _04216_, _03965_);
  and (_04218_, _04217_, _42545_);
  and (_39510_, _04218_, _04161_);
  nand (_04219_, _03965_, _33582_);
  nor (_04220_, _04030_, _19099_);
  and (_04221_, _04004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_04222_, _04007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_04223_, _04222_, _04221_);
  and (_04224_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_04225_, _04023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_04226_, _04225_, _04224_);
  or (_04227_, _04226_, _04223_);
  and (_04228_, _04012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_04229_, _04000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_04230_, _04229_, _04228_);
  and (_04231_, _04050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_04232_, _04052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_04233_, _04232_, _04231_);
  or (_04234_, _04233_, _04230_);
  or (_04235_, _04234_, _04227_);
  and (_04236_, _03979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_04237_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_04238_, _04237_, _04236_);
  and (_04239_, _03988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_04240_, _03985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_04241_, _04240_, _04239_);
  or (_04242_, _04241_, _04238_);
  and (_04243_, _03992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_04244_, _04022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_04245_, _04244_, _04243_);
  and (_04246_, _03996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_04247_, _03973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_04248_, _04247_, _04246_);
  or (_04249_, _04248_, _04245_);
  or (_04250_, _04249_, _04242_);
  or (_04251_, _04250_, _04235_);
  and (_04252_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_04253_, _03964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or (_04254_, _04253_, _04252_);
  and (_04255_, _04068_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_04256_, _04071_, _42439_);
  or (_04257_, _04256_, _04255_);
  or (_04258_, _04257_, _04254_);
  and (_04259_, _04078_, _03761_);
  and (_04260_, _04076_, _03564_);
  or (_04261_, _04260_, _04259_);
  and (_04262_, _04081_, _03821_);
  and (_04263_, _04083_, _03857_);
  or (_04264_, _04263_, _04262_);
  or (_04265_, _04264_, _04261_);
  or (_04266_, _04265_, _04258_);
  and (_04267_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_04268_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_04269_, _04268_, _04267_);
  or (_04271_, _04269_, _04266_);
  or (_04272_, _04271_, _04251_);
  and (_04273_, _04272_, _03962_);
  or (_04274_, _04273_, _04220_);
  or (_04275_, _04274_, _03965_);
  and (_04276_, _04275_, _42545_);
  and (_39511_, _04276_, _04219_);
  nand (_04277_, _03965_, _34333_);
  nor (_04278_, _04030_, _20130_);
  and (_04279_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_04280_, _03979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_04281_, _04280_, _04279_);
  and (_04282_, _03985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_04283_, _03988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_04284_, _04283_, _04282_);
  or (_04285_, _04284_, _04281_);
  and (_04286_, _03992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_04287_, _04022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_04288_, _04287_, _04286_);
  and (_04289_, _03996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_04290_, _03973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_04291_, _04290_, _04289_);
  or (_04292_, _04291_, _04288_);
  or (_04293_, _04292_, _04285_);
  and (_04294_, _04004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_04295_, _04007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_04296_, _04295_, _04294_);
  and (_04297_, _04023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_04298_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_04299_, _04298_, _04297_);
  or (_04300_, _04299_, _04296_);
  and (_04301_, _04012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_04302_, _04000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_04303_, _04302_, _04301_);
  and (_04304_, _04050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_04305_, _04052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_04306_, _04305_, _04304_);
  or (_04307_, _04306_, _04303_);
  or (_04308_, _04307_, _04300_);
  or (_04309_, _04308_, _04293_);
  and (_04310_, _03964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_04311_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_04312_, _04311_, _04310_);
  and (_04313_, _04068_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_04314_, _04071_, _42242_);
  or (_04315_, _04314_, _04313_);
  or (_04316_, _04315_, _04312_);
  and (_04317_, _04078_, _03746_);
  and (_04318_, _04076_, _03545_);
  or (_04319_, _04318_, _04317_);
  and (_04320_, _04081_, _03833_);
  and (_04321_, _04083_, _03847_);
  or (_04322_, _04321_, _04320_);
  or (_04323_, _04322_, _04319_);
  or (_04324_, _04323_, _04316_);
  and (_04325_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_04326_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_04327_, _04326_, _04325_);
  or (_04328_, _04327_, _04324_);
  or (_04329_, _04328_, _04309_);
  and (_04330_, _04329_, _03962_);
  or (_04331_, _04330_, _04278_);
  or (_04332_, _04331_, _03965_);
  and (_04333_, _04332_, _42545_);
  and (_39512_, _04333_, _04277_);
  nand (_04334_, _03965_, _35128_);
  nor (_04335_, _04030_, _19297_);
  and (_04336_, _03979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_04337_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_04338_, _04337_, _04336_);
  and (_04339_, _03988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_04340_, _03985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_04341_, _04340_, _04339_);
  or (_04342_, _04341_, _04338_);
  and (_04343_, _03992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_04344_, _04022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_04345_, _04344_, _04343_);
  and (_04346_, _03973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_04347_, _03996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_04348_, _04347_, _04346_);
  or (_04349_, _04348_, _04345_);
  or (_04350_, _04349_, _04342_);
  and (_04351_, _04012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_04352_, _04000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_04353_, _04352_, _04351_);
  and (_04354_, _04050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_04355_, _04052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_04356_, _04355_, _04354_);
  or (_04357_, _04356_, _04353_);
  and (_04358_, _04007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_04359_, _04004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_04360_, _04359_, _04358_);
  and (_04361_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_04362_, _04023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_04363_, _04362_, _04361_);
  or (_04364_, _04363_, _04360_);
  or (_04365_, _04364_, _04357_);
  or (_04366_, _04365_, _04350_);
  and (_04367_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_04368_, _03964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or (_04370_, _04368_, _04367_);
  and (_04371_, _04068_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_04372_, _04071_, _42122_);
  or (_04373_, _04372_, _04371_);
  or (_04374_, _04373_, _04370_);
  and (_04375_, _04081_, _03903_);
  and (_04376_, _04083_, _03877_);
  or (_04377_, _04376_, _04375_);
  and (_04378_, _04076_, _03528_);
  and (_04379_, _04078_, _03725_);
  or (_04380_, _04379_, _04378_);
  or (_04381_, _04380_, _04377_);
  or (_04382_, _04381_, _04374_);
  and (_04383_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_04384_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_04385_, _04384_, _04383_);
  or (_04386_, _04385_, _04382_);
  or (_04387_, _04386_, _04366_);
  and (_04388_, _04387_, _03962_);
  or (_04389_, _04388_, _04335_);
  or (_04390_, _04389_, _03965_);
  and (_04391_, _04390_, _42545_);
  and (_39513_, _04391_, _04334_);
  nand (_04392_, _03965_, _35956_);
  nor (_04393_, _04030_, _20283_);
  and (_04394_, _03992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04395_, _04022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_04396_, _04395_, _04394_);
  and (_04397_, _03996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_04398_, _03973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_04399_, _04398_, _04397_);
  or (_04400_, _04399_, _04396_);
  and (_04401_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04402_, _03979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_04403_, _04402_, _04401_);
  and (_04404_, _03985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_04405_, _03988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_04406_, _04405_, _04404_);
  or (_04407_, _04406_, _04403_);
  or (_04408_, _04407_, _04400_);
  and (_04409_, _04004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_04410_, _04007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_04411_, _04410_, _04409_);
  and (_04412_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_04413_, _04023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_04414_, _04413_, _04412_);
  or (_04415_, _04414_, _04411_);
  and (_04416_, _04000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_04417_, _04012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_04418_, _04417_, _04416_);
  and (_04419_, _04050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_04420_, _04052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_04421_, _04420_, _04419_);
  or (_04422_, _04421_, _04418_);
  or (_04423_, _04422_, _04415_);
  or (_04424_, _04423_, _04408_);
  and (_04425_, _04078_, _03733_);
  and (_04426_, _04083_, _03889_);
  or (_04427_, _04426_, _04425_);
  and (_04428_, _04076_, _03534_);
  and (_04429_, _04081_, _03912_);
  or (_04430_, _04429_, _04428_);
  or (_04431_, _04430_, _04427_);
  and (_04432_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_04433_, _03964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_04434_, _04433_, _04432_);
  and (_04435_, _04068_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_04436_, _04071_, _42393_);
  or (_04437_, _04436_, _04435_);
  or (_04438_, _04437_, _04434_);
  or (_04439_, _04438_, _04431_);
  and (_04440_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_04441_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_04442_, _04441_, _04440_);
  or (_04443_, _04442_, _04439_);
  or (_04444_, _04443_, _04424_);
  and (_04445_, _04444_, _03962_);
  or (_04446_, _04445_, _04393_);
  or (_04447_, _04446_, _03965_);
  and (_04448_, _04447_, _42545_);
  and (_39514_, _04448_, _04392_);
  nand (_04449_, _03965_, _36684_);
  nor (_04450_, _04030_, _19634_);
  and (_04451_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_04452_, _03979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_04453_, _04452_, _04451_);
  and (_04454_, _03988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_04455_, _03985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_04456_, _04455_, _04454_);
  or (_04457_, _04456_, _04453_);
  and (_04458_, _03992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_04459_, _04022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_04460_, _04459_, _04458_);
  and (_04461_, _03996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_04462_, _03973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_04463_, _04462_, _04461_);
  or (_04464_, _04463_, _04460_);
  or (_04465_, _04464_, _04457_);
  and (_04466_, _04000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_04467_, _04012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or (_04469_, _04467_, _04466_);
  and (_04470_, _04050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_04471_, _04052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_04472_, _04471_, _04470_);
  or (_04473_, _04472_, _04469_);
  and (_04474_, _04004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_04475_, _04007_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_04476_, _04475_, _04474_);
  and (_04477_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_04478_, _04023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_04479_, _04478_, _04477_);
  or (_04480_, _04479_, _04476_);
  or (_04481_, _04480_, _04473_);
  or (_04482_, _04481_, _04465_);
  and (_04483_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_04484_, _03964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_04485_, _04484_, _04483_);
  and (_04486_, _04068_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_04487_, _04071_, _42301_);
  or (_04488_, _04487_, _04486_);
  or (_04489_, _04488_, _04485_);
  and (_04490_, _04076_, _03559_);
  and (_04491_, _04078_, _03756_);
  or (_04492_, _04491_, _04490_);
  and (_04493_, _04081_, _03899_);
  and (_04494_, _04083_, _03872_);
  or (_04495_, _04494_, _04493_);
  or (_04496_, _04495_, _04492_);
  or (_04497_, _04496_, _04489_);
  and (_04498_, _03949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_04499_, _03945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_04500_, _04499_, _04498_);
  or (_04501_, _04500_, _04497_);
  or (_04502_, _04501_, _04482_);
  and (_04503_, _04502_, _03962_);
  or (_04504_, _04503_, _04450_);
  or (_04505_, _04504_, _03965_);
  and (_04506_, _04505_, _42545_);
  and (_39515_, _04506_, _04449_);
  and (_39584_, _42476_, _42545_);
  nor (_39587_, _42443_, rst);
  nor (_39611_, _42294_, rst);
  nor (_39613_, _42195_, rst);
  not (_04507_, _00628_);
  nor (_04508_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_04509_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04510_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04509_);
  nor (_04511_, _04510_, _04508_);
  nor (_04512_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04513_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04509_);
  nor (_04514_, _04513_, _04512_);
  nor (_04515_, _04514_, _04511_);
  nor (_04516_, _02273_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04517_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04509_);
  or (_04518_, _04517_, _04516_);
  and (_04519_, _04514_, _04511_);
  nor (_04520_, _02252_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04521_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04509_);
  nor (_04522_, _04521_, _04520_);
  and (_04523_, _04522_, _04519_);
  nor (_04524_, _04522_, _04519_);
  nor (_04525_, _04524_, _04523_);
  not (_04526_, _04525_);
  nor (_04527_, _04526_, _04518_);
  and (_04528_, _04527_, _04515_);
  not (_04529_, _04511_);
  nor (_04530_, _04514_, _04529_);
  and (_04531_, _04527_, _04530_);
  nor (_04532_, _04531_, _04528_);
  and (_04533_, _04527_, _04519_);
  and (_04534_, _04525_, _04518_);
  not (_04535_, _04523_);
  not (_04536_, _04524_);
  or (_04537_, _04536_, _04518_);
  nand (_04538_, _04537_, _04535_);
  or (_04539_, _04538_, _04534_);
  nor (_04540_, _04539_, _04533_);
  and (_04541_, _04540_, _04532_);
  and (_04542_, _04523_, _04518_);
  nor (_04543_, _04523_, _04518_);
  or (_04544_, _04543_, _04542_);
  nor (_04545_, _04544_, _04525_);
  and (_04546_, _04545_, _04515_);
  and (_04547_, _04545_, _04530_);
  and (_04548_, _04514_, _04529_);
  and (_04549_, _04545_, _04548_);
  or (_04550_, _04549_, _04547_);
  nor (_04551_, _04550_, _04546_);
  and (_04552_, _04551_, _04541_);
  and (_04553_, _04552_, _04507_);
  not (_04554_, _00527_);
  and (_04555_, _04528_, _04554_);
  not (_04556_, _00584_);
  and (_04557_, _04531_, _04556_);
  or (_04558_, _04557_, _04555_);
  not (_04559_, _00486_);
  and (_04560_, _04533_, _04559_);
  not (_04561_, _00445_);
  and (_04562_, _04544_, _04526_);
  and (_04564_, _04562_, _04548_);
  and (_04565_, _04564_, _04561_);
  or (_04566_, _04565_, _04560_);
  or (_04567_, _04566_, _04558_);
  not (_04568_, _00404_);
  and (_04569_, _04562_, _04530_);
  and (_04570_, _04569_, _04568_);
  not (_04571_, _00363_);
  and (_04572_, _04562_, _04515_);
  and (_04573_, _04572_, _04571_);
  or (_04574_, _04573_, _04570_);
  not (_04575_, _00281_);
  and (_04576_, _04534_, _04548_);
  and (_04577_, _04576_, _04575_);
  not (_04578_, _00322_);
  and (_04579_, _04542_, _04578_);
  or (_04580_, _04579_, _04577_);
  or (_04581_, _04580_, _04574_);
  or (_04582_, _04581_, _04567_);
  not (_04583_, _00004_);
  and (_04584_, _04546_, _04583_);
  not (_04585_, _00045_);
  and (_04586_, _04547_, _04585_);
  not (_04587_, _43422_);
  nor (_04588_, _04535_, _04518_);
  and (_04589_, _04588_, _04587_);
  or (_04590_, _04589_, _04586_);
  or (_04591_, _04590_, _04584_);
  not (_04592_, _00240_);
  and (_04593_, _04534_, _04530_);
  and (_04594_, _04593_, _04592_);
  not (_04595_, _00199_);
  and (_04596_, _04534_, _04515_);
  and (_04597_, _04596_, _04595_);
  or (_04598_, _04597_, _04594_);
  not (_04599_, _00127_);
  and (_04600_, _04534_, _04519_);
  and (_04601_, _04600_, _04599_);
  not (_04602_, _00086_);
  and (_04603_, _04549_, _04602_);
  or (_04604_, _04603_, _04601_);
  or (_04605_, _04604_, _04598_);
  or (_04606_, _04605_, _04591_);
  or (_04607_, _04606_, _04582_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04607_, _04553_);
  and (_04608_, _04547_, _04602_);
  and (_04609_, _04588_, _04583_);
  or (_04610_, _04609_, _04608_);
  and (_04611_, _04572_, _04568_);
  and (_04612_, _04569_, _04561_);
  and (_04613_, _04564_, _04559_);
  or (_04614_, _04613_, _04612_);
  or (_04615_, _04614_, _04611_);
  or (_04616_, _04615_, _04610_);
  and (_04617_, _04552_, _04587_);
  and (_04618_, _04528_, _04556_);
  and (_04619_, _04531_, _04507_);
  and (_04620_, _04542_, _04571_);
  or (_04621_, _04620_, _04619_);
  or (_04622_, _04621_, _04618_);
  and (_04623_, _04576_, _04578_);
  and (_04624_, _04533_, _04554_);
  or (_04625_, _04624_, _04623_);
  or (_04626_, _04625_, _04622_);
  and (_04627_, _04600_, _04595_);
  and (_04628_, _04596_, _04592_);
  and (_04629_, _04593_, _04575_);
  or (_04630_, _04629_, _04628_);
  or (_04631_, _04630_, _04627_);
  and (_04632_, _04546_, _04585_);
  and (_04633_, _04549_, _04599_);
  or (_04634_, _04633_, _04632_);
  or (_04635_, _04634_, _04631_);
  or (_04636_, _04635_, _04626_);
  or (_04637_, _04636_, _04617_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04637_, _04616_);
  and (_04638_, _04552_, _04583_);
  and (_04639_, _04569_, _04559_);
  and (_04640_, _04547_, _04599_);
  or (_04641_, _04640_, _04639_);
  and (_04642_, _04549_, _04595_);
  and (_04643_, _04546_, _04602_);
  or (_04644_, _04643_, _04642_);
  or (_04645_, _04644_, _04641_);
  and (_04646_, _04596_, _04575_);
  and (_04647_, _04600_, _04592_);
  or (_04648_, _04647_, _04646_);
  and (_04649_, _04528_, _04507_);
  and (_04650_, _04533_, _04556_);
  or (_04651_, _04650_, _04649_);
  or (_04652_, _04651_, _04648_);
  and (_04653_, _04576_, _04571_);
  and (_04654_, _04542_, _04568_);
  and (_04655_, _04588_, _04585_);
  or (_04656_, _04655_, _04654_);
  or (_04657_, _04656_, _04653_);
  and (_04658_, _04593_, _04578_);
  and (_04659_, _04531_, _04587_);
  or (_04660_, _04659_, _04658_);
  or (_04661_, _04660_, _04657_);
  and (_04663_, _04564_, _04554_);
  and (_04664_, _04572_, _04561_);
  or (_04665_, _04664_, _04663_);
  or (_04666_, _04665_, _04661_);
  or (_04667_, _04666_, _04652_);
  or (_04668_, _04667_, _04645_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04668_, _04638_);
  and (_04669_, _04552_, _04556_);
  and (_04670_, _04564_, _04568_);
  and (_04671_, _04549_, _04585_);
  or (_04672_, _04671_, _04670_);
  and (_04673_, _04546_, _04587_);
  and (_04674_, _04547_, _04583_);
  or (_04675_, _04674_, _04673_);
  or (_04676_, _04675_, _04672_);
  and (_04677_, _04533_, _04561_);
  and (_04678_, _04596_, _04599_);
  or (_04679_, _04678_, _04677_);
  and (_04680_, _04531_, _04554_);
  and (_04681_, _04528_, _04559_);
  or (_04682_, _04681_, _04680_);
  or (_04683_, _04682_, _04679_);
  and (_04684_, _04593_, _04595_);
  and (_04685_, _04576_, _04592_);
  or (_04686_, _04685_, _04684_);
  and (_04687_, _04600_, _04602_);
  and (_04688_, _04588_, _04507_);
  and (_04689_, _04542_, _04575_);
  or (_04690_, _04689_, _04688_);
  or (_04691_, _04690_, _04687_);
  or (_04692_, _04691_, _04686_);
  and (_04693_, _04569_, _04571_);
  and (_04694_, _04572_, _04578_);
  or (_04695_, _04694_, _04693_);
  or (_04696_, _04695_, _04692_);
  or (_04697_, _04696_, _04683_);
  or (_04698_, _04697_, _04676_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04698_, _04669_);
  not (_04699_, _00204_);
  and (_04700_, _04593_, _04699_);
  not (_04701_, _00245_);
  and (_04702_, _04576_, _04701_);
  or (_04703_, _04702_, _04700_);
  not (_04704_, _00135_);
  and (_04705_, _04596_, _04704_);
  not (_04706_, _00091_);
  and (_04707_, _04600_, _04706_);
  or (_04708_, _04707_, _04705_);
  or (_04709_, _04708_, _04703_);
  not (_04710_, _00327_);
  and (_04711_, _04572_, _04710_);
  not (_04712_, _00409_);
  and (_04713_, _04564_, _04712_);
  not (_04714_, _00450_);
  and (_04715_, _04533_, _04714_);
  or (_04716_, _04715_, _04713_);
  or (_04717_, _04716_, _04711_);
  or (_04718_, _04717_, _04709_);
  not (_04719_, _00592_);
  and (_04720_, _04552_, _04719_);
  not (_04721_, _00050_);
  and (_04722_, _04549_, _04721_);
  not (_04723_, _43427_);
  and (_04724_, _04546_, _04723_);
  not (_04725_, _00009_);
  and (_04726_, _04547_, _04725_);
  or (_04727_, _04726_, _04724_);
  or (_04728_, _04727_, _04722_);
  not (_04729_, _00368_);
  and (_04730_, _04569_, _04729_);
  not (_04731_, _00491_);
  and (_04732_, _04528_, _04731_);
  not (_04733_, _00532_);
  and (_04734_, _04531_, _04733_);
  not (_04735_, _00633_);
  and (_04736_, _04588_, _04735_);
  not (_04737_, _00286_);
  and (_04738_, _04542_, _04737_);
  or (_04739_, _04738_, _04736_);
  or (_04740_, _04739_, _04734_);
  or (_04741_, _04740_, _04732_);
  or (_04742_, _04741_, _04730_);
  or (_04743_, _04742_, _04728_);
  or (_04744_, _04743_, _04720_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _04744_, _04718_);
  not (_04745_, _00597_);
  and (_04746_, _04552_, _04745_);
  not (_04747_, _00414_);
  and (_04748_, _04564_, _04747_);
  not (_04749_, _00055_);
  and (_04750_, _04549_, _04749_);
  or (_04751_, _04750_, _04748_);
  not (_04752_, _43432_);
  and (_04753_, _04546_, _04752_);
  not (_04754_, _00014_);
  and (_04755_, _04547_, _04754_);
  or (_04756_, _04755_, _04753_);
  or (_04757_, _04756_, _04751_);
  not (_04758_, _00455_);
  and (_04759_, _04533_, _04758_);
  not (_04761_, _00146_);
  and (_04762_, _04596_, _04761_);
  or (_04763_, _04762_, _04759_);
  not (_04764_, _00537_);
  and (_04765_, _04531_, _04764_);
  not (_04766_, _00496_);
  and (_04767_, _04528_, _04766_);
  or (_04768_, _04767_, _04765_);
  or (_04769_, _04768_, _04763_);
  not (_04770_, _00209_);
  and (_04771_, _04593_, _04770_);
  not (_04772_, _00250_);
  and (_04773_, _04576_, _04772_);
  or (_04774_, _04773_, _04771_);
  not (_04775_, _00096_);
  and (_04776_, _04600_, _04775_);
  not (_04777_, _00638_);
  and (_04778_, _04588_, _04777_);
  not (_04779_, _00291_);
  and (_04780_, _04542_, _04779_);
  or (_04781_, _04780_, _04778_);
  or (_04782_, _04781_, _04776_);
  or (_04783_, _04782_, _04774_);
  not (_04784_, _00373_);
  and (_04785_, _04569_, _04784_);
  not (_04786_, _00332_);
  and (_04787_, _04572_, _04786_);
  or (_04788_, _04787_, _04785_);
  or (_04789_, _04788_, _04783_);
  or (_04790_, _04789_, _04769_);
  or (_04791_, _04790_, _04757_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _04791_, _04746_);
  not (_04792_, _00060_);
  and (_04793_, _04549_, _04792_);
  not (_04794_, _43437_);
  and (_04795_, _04546_, _04794_);
  or (_04796_, _04795_, _04793_);
  not (_04797_, _00255_);
  and (_04798_, _04576_, _04797_);
  not (_04799_, _00101_);
  and (_04800_, _04600_, _04799_);
  or (_04801_, _04800_, _04798_);
  not (_04802_, _00214_);
  and (_04803_, _04593_, _04802_);
  not (_04804_, _00157_);
  and (_04805_, _04596_, _04804_);
  or (_04806_, _04805_, _04803_);
  or (_04807_, _04806_, _04801_);
  not (_04808_, _00019_);
  and (_04809_, _04547_, _04808_);
  or (_04810_, _04809_, _04807_);
  or (_04811_, _04810_, _04796_);
  not (_04812_, _00602_);
  and (_04813_, _04552_, _04812_);
  not (_04814_, _00378_);
  and (_04815_, _04569_, _04814_);
  not (_04816_, _00460_);
  and (_04817_, _04533_, _04816_);
  not (_04818_, _00419_);
  and (_04819_, _04564_, _04818_);
  or (_04820_, _04819_, _04817_);
  or (_04821_, _04820_, _04815_);
  not (_04822_, _00337_);
  and (_04823_, _04572_, _04822_);
  not (_04824_, _00501_);
  and (_04825_, _04528_, _04824_);
  not (_04826_, _00542_);
  and (_04827_, _04531_, _04826_);
  not (_04828_, _00643_);
  and (_04829_, _04588_, _04828_);
  not (_04830_, _00296_);
  and (_04831_, _04542_, _04830_);
  or (_04832_, _04831_, _04829_);
  or (_04833_, _04832_, _04827_);
  or (_04834_, _04833_, _04825_);
  or (_04835_, _04834_, _04823_);
  or (_04836_, _04835_, _04821_);
  or (_04837_, _04836_, _04813_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _04837_, _04811_);
  not (_04838_, _00607_);
  and (_04839_, _04552_, _04838_);
  not (_04840_, _00424_);
  and (_04841_, _04564_, _04840_);
  not (_04842_, _00065_);
  and (_04843_, _04549_, _04842_);
  or (_04844_, _04843_, _04841_);
  not (_04845_, _43442_);
  and (_04846_, _04546_, _04845_);
  not (_04847_, _00024_);
  and (_04848_, _04547_, _04847_);
  or (_04849_, _04848_, _04846_);
  or (_04850_, _04849_, _04844_);
  not (_04851_, _00465_);
  and (_04852_, _04533_, _04851_);
  not (_04853_, _00106_);
  and (_04854_, _04600_, _04853_);
  or (_04855_, _04854_, _04852_);
  not (_04856_, _00550_);
  and (_04857_, _04531_, _04856_);
  not (_04858_, _00506_);
  and (_04859_, _04528_, _04858_);
  or (_04860_, _04859_, _04857_);
  or (_04861_, _04860_, _04855_);
  not (_04862_, _00219_);
  and (_04863_, _04593_, _04862_);
  not (_04864_, _00260_);
  and (_04865_, _04576_, _04864_);
  or (_04866_, _04865_, _04863_);
  not (_04867_, _00168_);
  and (_04868_, _04596_, _04867_);
  not (_04869_, _00648_);
  and (_04870_, _04588_, _04869_);
  not (_04871_, _00301_);
  and (_04872_, _04542_, _04871_);
  or (_04873_, _04872_, _04870_);
  or (_04874_, _04873_, _04868_);
  or (_04875_, _04874_, _04866_);
  not (_04876_, _00383_);
  and (_04877_, _04569_, _04876_);
  not (_04878_, _00342_);
  and (_04879_, _04572_, _04878_);
  or (_04880_, _04879_, _04877_);
  or (_04881_, _04880_, _04875_);
  or (_04882_, _04881_, _04861_);
  or (_04883_, _04882_, _04850_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _04883_, _04839_);
  not (_04884_, _00612_);
  and (_04885_, _04552_, _04884_);
  not (_04886_, _00429_);
  and (_04887_, _04564_, _04886_);
  not (_04888_, _00070_);
  and (_04889_, _04549_, _04888_);
  or (_04890_, _04889_, _04887_);
  not (_04891_, _43447_);
  and (_04892_, _04546_, _04891_);
  not (_04893_, _00029_);
  and (_04894_, _04547_, _04893_);
  or (_04895_, _04894_, _04892_);
  or (_04896_, _04895_, _04890_);
  not (_04897_, _00470_);
  and (_04898_, _04533_, _04897_);
  not (_04899_, _00111_);
  and (_04900_, _04600_, _04899_);
  or (_04901_, _04900_, _04898_);
  not (_04902_, _00558_);
  and (_04903_, _04531_, _04902_);
  not (_04904_, _00511_);
  and (_04905_, _04528_, _04904_);
  or (_04906_, _04905_, _04903_);
  or (_04907_, _04906_, _04901_);
  not (_04908_, _00224_);
  and (_04909_, _04593_, _04908_);
  not (_04910_, _00265_);
  and (_04911_, _04576_, _04910_);
  or (_04912_, _04911_, _04909_);
  not (_04913_, _00179_);
  and (_04914_, _04596_, _04913_);
  not (_04915_, _00653_);
  and (_04916_, _04588_, _04915_);
  not (_04917_, _00306_);
  and (_04918_, _04542_, _04917_);
  or (_04919_, _04918_, _04916_);
  or (_04920_, _04919_, _04914_);
  or (_04921_, _04920_, _04912_);
  not (_04922_, _00388_);
  and (_04923_, _04569_, _04922_);
  not (_04924_, _00347_);
  and (_04925_, _04572_, _04924_);
  or (_04926_, _04925_, _04923_);
  or (_04927_, _04926_, _04921_);
  or (_04928_, _04927_, _04907_);
  or (_04929_, _04928_, _04896_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _04929_, _04885_);
  not (_04930_, _00075_);
  and (_04931_, _04549_, _04930_);
  not (_04932_, _43452_);
  and (_04933_, _04546_, _04932_);
  or (_04934_, _04933_, _04931_);
  not (_04935_, _00270_);
  and (_04936_, _04576_, _04935_);
  not (_04937_, _00116_);
  and (_04938_, _04600_, _04937_);
  or (_04939_, _04938_, _04936_);
  not (_04940_, _00229_);
  and (_04941_, _04593_, _04940_);
  not (_04942_, _00188_);
  and (_04943_, _04596_, _04942_);
  or (_04944_, _04943_, _04941_);
  or (_04945_, _04944_, _04939_);
  not (_04946_, _00034_);
  and (_04947_, _04547_, _04946_);
  or (_04948_, _04947_, _04945_);
  or (_04949_, _04948_, _04934_);
  not (_04950_, _00617_);
  and (_04951_, _04552_, _04950_);
  not (_04952_, _00352_);
  and (_04953_, _04572_, _04952_);
  not (_04954_, _00475_);
  and (_04955_, _04533_, _04954_);
  not (_04956_, _00434_);
  and (_04957_, _04564_, _04956_);
  or (_04958_, _04957_, _04955_);
  or (_04959_, _04958_, _04953_);
  not (_04960_, _00393_);
  and (_04961_, _04569_, _04960_);
  not (_04962_, _00516_);
  and (_04963_, _04528_, _04962_);
  not (_04964_, _00566_);
  and (_04965_, _04531_, _04964_);
  not (_04966_, _00658_);
  and (_04967_, _04588_, _04966_);
  not (_04968_, _00311_);
  and (_04969_, _04542_, _04968_);
  or (_04970_, _04969_, _04967_);
  or (_04971_, _04970_, _04965_);
  or (_04972_, _04971_, _04963_);
  or (_04973_, _04972_, _04961_);
  or (_04974_, _04973_, _04959_);
  or (_04975_, _04974_, _04951_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _04975_, _04949_);
  not (_04976_, _00234_);
  and (_04977_, _04593_, _04976_);
  not (_04978_, _00275_);
  and (_04979_, _04576_, _04978_);
  or (_04980_, _04979_, _04977_);
  not (_04981_, _00193_);
  and (_04982_, _04596_, _04981_);
  not (_04983_, _00121_);
  and (_04984_, _04600_, _04983_);
  or (_04985_, _04984_, _04982_);
  or (_04986_, _04985_, _04980_);
  not (_04987_, _00357_);
  and (_04988_, _04572_, _04987_);
  not (_04989_, _00439_);
  and (_04990_, _04564_, _04989_);
  not (_04991_, _00480_);
  and (_04992_, _04533_, _04991_);
  or (_04993_, _04992_, _04990_);
  or (_04994_, _04993_, _04988_);
  or (_04995_, _04994_, _04986_);
  not (_04996_, _00622_);
  and (_04997_, _04552_, _04996_);
  not (_04998_, _00080_);
  and (_04999_, _04549_, _04998_);
  not (_05000_, _43457_);
  and (_05001_, _04546_, _05000_);
  not (_05002_, _00039_);
  and (_05003_, _04547_, _05002_);
  or (_05004_, _05003_, _05001_);
  or (_05005_, _05004_, _04999_);
  not (_05006_, _00398_);
  and (_05007_, _04569_, _05006_);
  not (_05008_, _00521_);
  and (_05009_, _04528_, _05008_);
  not (_05010_, _00574_);
  and (_05011_, _04531_, _05010_);
  not (_05012_, _00663_);
  and (_05013_, _04588_, _05012_);
  not (_05014_, _00316_);
  and (_05015_, _04542_, _05014_);
  or (_05016_, _05015_, _05013_);
  or (_05017_, _05016_, _05011_);
  or (_05018_, _05017_, _05009_);
  or (_05019_, _05018_, _05007_);
  or (_05020_, _05019_, _05005_);
  or (_05021_, _05020_, _04997_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _05021_, _04995_);
  and (_05022_, _04564_, _04733_);
  and (_05023_, _04533_, _04719_);
  and (_05024_, _04528_, _04735_);
  and (_05025_, _04542_, _04712_);
  or (_05026_, _05025_, _05024_);
  or (_05027_, _05026_, _05023_);
  or (_05028_, _05027_, _05022_);
  and (_05029_, _04549_, _04699_);
  and (_05030_, _04600_, _04701_);
  and (_05031_, _04596_, _04737_);
  or (_05032_, _05031_, _05030_);
  or (_05033_, _05032_, _05029_);
  or (_05034_, _05033_, _05028_);
  and (_05035_, _04552_, _04725_);
  and (_05036_, _04576_, _04729_);
  and (_05037_, _04593_, _04710_);
  or (_05038_, _05037_, _05036_);
  and (_05039_, _04572_, _04714_);
  and (_05040_, _04569_, _04731_);
  or (_05041_, _05040_, _05039_);
  or (_05042_, _05041_, _05038_);
  and (_05043_, _04547_, _04704_);
  and (_05044_, _04546_, _04706_);
  and (_05045_, _04531_, _04723_);
  and (_05046_, _04588_, _04721_);
  or (_05047_, _05046_, _05045_);
  or (_05048_, _05047_, _05044_);
  or (_05049_, _05048_, _05043_);
  or (_05050_, _05049_, _05042_);
  or (_05051_, _05050_, _05035_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _05051_, _05034_);
  and (_05052_, _04552_, _04754_);
  and (_05053_, _04569_, _04766_);
  and (_05054_, _04547_, _04761_);
  or (_05055_, _05054_, _05053_);
  and (_05056_, _04549_, _04770_);
  and (_05057_, _04546_, _04775_);
  or (_05058_, _05057_, _05056_);
  or (_05059_, _05058_, _05055_);
  and (_05060_, _04596_, _04779_);
  and (_05061_, _04600_, _04772_);
  or (_05062_, _05061_, _05060_);
  and (_05063_, _04528_, _04777_);
  and (_05064_, _04533_, _04745_);
  or (_05065_, _05064_, _05063_);
  or (_05066_, _05065_, _05062_);
  and (_05067_, _04576_, _04784_);
  and (_05068_, _04542_, _04747_);
  and (_05069_, _04588_, _04749_);
  or (_05070_, _05069_, _05068_);
  or (_05071_, _05070_, _05067_);
  and (_05072_, _04593_, _04786_);
  and (_05073_, _04531_, _04752_);
  or (_05074_, _05073_, _05072_);
  or (_05075_, _05074_, _05071_);
  and (_05076_, _04564_, _04764_);
  and (_05077_, _04572_, _04758_);
  or (_05078_, _05077_, _05076_);
  or (_05079_, _05078_, _05075_);
  or (_05080_, _05079_, _05066_);
  or (_05081_, _05080_, _05059_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _05081_, _05052_);
  and (_05082_, _04552_, _04808_);
  and (_05083_, _04572_, _04816_);
  and (_05084_, _04547_, _04804_);
  or (_05085_, _05084_, _05083_);
  and (_05086_, _04549_, _04802_);
  and (_05087_, _04546_, _04799_);
  or (_05088_, _05087_, _05086_);
  or (_05089_, _05088_, _05085_);
  and (_05090_, _04528_, _04828_);
  and (_05091_, _04531_, _04794_);
  or (_05092_, _05091_, _05090_);
  and (_05093_, _04533_, _04812_);
  and (_05094_, _04596_, _04830_);
  or (_05095_, _05094_, _05093_);
  or (_05096_, _05095_, _05092_);
  and (_05097_, _04593_, _04822_);
  and (_05098_, _04542_, _04818_);
  and (_05099_, _04588_, _04792_);
  or (_05100_, _05099_, _05098_);
  or (_05101_, _05100_, _05097_);
  and (_05102_, _04576_, _04814_);
  and (_05103_, _04600_, _04797_);
  or (_05104_, _05103_, _05102_);
  or (_05105_, _05104_, _05101_);
  and (_05106_, _04569_, _04824_);
  and (_05107_, _04564_, _04826_);
  or (_05108_, _05107_, _05106_);
  or (_05109_, _05108_, _05105_);
  or (_05110_, _05109_, _05096_);
  or (_05111_, _05110_, _05089_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _05111_, _05082_);
  and (_05112_, _04564_, _04856_);
  and (_05113_, _04533_, _04838_);
  and (_05114_, _04528_, _04869_);
  and (_05115_, _04542_, _04840_);
  or (_05116_, _05115_, _05114_);
  or (_05117_, _05116_, _05113_);
  or (_05118_, _05117_, _05112_);
  and (_05119_, _04549_, _04862_);
  and (_05120_, _04600_, _04864_);
  and (_05121_, _04596_, _04871_);
  or (_05122_, _05121_, _05120_);
  or (_05123_, _05122_, _05119_);
  or (_05124_, _05123_, _05118_);
  and (_05125_, _04552_, _04847_);
  and (_05126_, _04576_, _04876_);
  and (_05127_, _04593_, _04878_);
  or (_05128_, _05127_, _05126_);
  and (_05129_, _04572_, _04851_);
  and (_05130_, _04569_, _04858_);
  or (_05131_, _05130_, _05129_);
  or (_05132_, _05131_, _05128_);
  and (_05133_, _04547_, _04867_);
  and (_05134_, _04546_, _04853_);
  and (_05135_, _04531_, _04845_);
  and (_05136_, _04588_, _04842_);
  or (_05137_, _05136_, _05135_);
  or (_05138_, _05137_, _05134_);
  or (_05139_, _05138_, _05133_);
  or (_05140_, _05139_, _05132_);
  or (_05141_, _05140_, _05125_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _05141_, _05124_);
  and (_05142_, _04552_, _04893_);
  and (_05143_, _04569_, _04904_);
  and (_05144_, _04547_, _04913_);
  or (_05145_, _05144_, _05143_);
  and (_05146_, _04572_, _04897_);
  and (_05147_, _04546_, _04899_);
  or (_05148_, _05147_, _05146_);
  or (_05149_, _05148_, _05145_);
  and (_05150_, _04596_, _04917_);
  and (_05151_, _04600_, _04910_);
  or (_05152_, _05151_, _05150_);
  and (_05153_, _04528_, _04915_);
  and (_05154_, _04533_, _04884_);
  or (_05155_, _05154_, _05153_);
  or (_05156_, _05155_, _05152_);
  and (_05157_, _04576_, _04922_);
  and (_05158_, _04542_, _04886_);
  and (_05159_, _04588_, _04888_);
  or (_05160_, _05159_, _05158_);
  or (_05161_, _05160_, _05157_);
  and (_05162_, _04593_, _04924_);
  and (_05163_, _04531_, _04891_);
  or (_05164_, _05163_, _05162_);
  or (_05165_, _05164_, _05161_);
  and (_05166_, _04564_, _04902_);
  and (_05167_, _04549_, _04908_);
  or (_05168_, _05167_, _05166_);
  or (_05169_, _05168_, _05165_);
  or (_05170_, _05169_, _05156_);
  or (_05171_, _05170_, _05149_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _05171_, _05142_);
  and (_05172_, _04552_, _04946_);
  and (_05173_, _04569_, _04962_);
  and (_05174_, _04547_, _04942_);
  or (_05175_, _05174_, _05173_);
  and (_05176_, _04572_, _04954_);
  and (_05177_, _04546_, _04937_);
  or (_05178_, _05177_, _05176_);
  or (_05179_, _05178_, _05175_);
  and (_05180_, _04596_, _04968_);
  and (_05181_, _04600_, _04935_);
  or (_05182_, _05181_, _05180_);
  and (_05183_, _04528_, _04966_);
  and (_05184_, _04533_, _04950_);
  or (_05185_, _05184_, _05183_);
  or (_05186_, _05185_, _05182_);
  and (_05187_, _04593_, _04952_);
  and (_05188_, _04542_, _04956_);
  and (_05189_, _04588_, _04930_);
  or (_05190_, _05189_, _05188_);
  or (_05191_, _05190_, _05187_);
  and (_05192_, _04576_, _04960_);
  and (_05193_, _04531_, _04932_);
  or (_05194_, _05193_, _05192_);
  or (_05195_, _05194_, _05191_);
  and (_05196_, _04564_, _04964_);
  and (_05197_, _04549_, _04940_);
  or (_05198_, _05197_, _05196_);
  or (_05199_, _05198_, _05195_);
  or (_05200_, _05199_, _05186_);
  or (_05201_, _05200_, _05179_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _05201_, _05172_);
  and (_05202_, _04564_, _05010_);
  and (_05203_, _04533_, _04996_);
  and (_05204_, _04528_, _05012_);
  and (_05205_, _04542_, _04989_);
  or (_05206_, _05205_, _05204_);
  or (_05207_, _05206_, _05203_);
  or (_05208_, _05207_, _05202_);
  and (_05209_, _04549_, _04976_);
  and (_05210_, _04600_, _04978_);
  and (_05211_, _04596_, _05014_);
  or (_05212_, _05211_, _05210_);
  or (_05213_, _05212_, _05209_);
  or (_05214_, _05213_, _05208_);
  and (_05215_, _04552_, _05002_);
  and (_05216_, _04576_, _05006_);
  and (_05217_, _04593_, _04987_);
  or (_05218_, _05217_, _05216_);
  and (_05219_, _04572_, _04991_);
  and (_05220_, _04569_, _05008_);
  or (_05221_, _05220_, _05219_);
  or (_05222_, _05221_, _05218_);
  and (_05223_, _04547_, _04981_);
  and (_05224_, _04546_, _04983_);
  and (_05225_, _04531_, _05000_);
  and (_05226_, _04588_, _04998_);
  or (_05227_, _05226_, _05225_);
  or (_05228_, _05227_, _05224_);
  or (_05229_, _05228_, _05223_);
  or (_05230_, _05229_, _05222_);
  or (_05231_, _05230_, _05215_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _05231_, _05214_);
  and (_05232_, _04552_, _04735_);
  and (_05233_, _04531_, _04719_);
  and (_05234_, _04528_, _04733_);
  or (_05235_, _05234_, _05233_);
  and (_05236_, _04564_, _04714_);
  and (_05237_, _04533_, _04731_);
  or (_05238_, _05237_, _05236_);
  or (_05239_, _05238_, _05235_);
  and (_05240_, _04572_, _04729_);
  and (_05241_, _04569_, _04712_);
  or (_05242_, _05241_, _05240_);
  and (_05243_, _04576_, _04737_);
  and (_05244_, _04542_, _04710_);
  or (_05245_, _05244_, _05243_);
  or (_05246_, _05245_, _05242_);
  or (_05247_, _05246_, _05239_);
  and (_05248_, _04546_, _04725_);
  and (_05249_, _04547_, _04721_);
  and (_05250_, _04588_, _04723_);
  or (_05251_, _05250_, _05249_);
  or (_05252_, _05251_, _05248_);
  and (_05253_, _04593_, _04701_);
  and (_05254_, _04596_, _04699_);
  or (_05255_, _05254_, _05253_);
  and (_05256_, _04549_, _04706_);
  and (_05257_, _04600_, _04704_);
  or (_05258_, _05257_, _05256_);
  or (_05259_, _05258_, _05255_);
  or (_05260_, _05259_, _05252_);
  or (_05261_, _05260_, _05247_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _05261_, _05232_);
  and (_05262_, _04552_, _04777_);
  and (_05263_, _04531_, _04745_);
  and (_05264_, _04528_, _04764_);
  or (_05265_, _05264_, _05263_);
  and (_05266_, _04533_, _04766_);
  and (_05267_, _04564_, _04758_);
  or (_05268_, _05267_, _05266_);
  or (_05269_, _05268_, _05265_);
  and (_05270_, _04569_, _04747_);
  and (_05271_, _04572_, _04784_);
  or (_05272_, _05271_, _05270_);
  and (_05273_, _04576_, _04779_);
  and (_05274_, _04542_, _04786_);
  or (_05275_, _05274_, _05273_);
  or (_05276_, _05275_, _05272_);
  or (_05277_, _05276_, _05269_);
  and (_05278_, _04596_, _04770_);
  and (_05279_, _04593_, _04772_);
  or (_05280_, _05279_, _05278_);
  and (_05281_, _04549_, _04775_);
  and (_05282_, _04600_, _04761_);
  or (_05283_, _05282_, _05281_);
  or (_05284_, _05283_, _05280_);
  and (_05285_, _04588_, _04752_);
  and (_05286_, _04547_, _04749_);
  and (_05287_, _04546_, _04754_);
  or (_05288_, _05287_, _05286_);
  or (_05289_, _05288_, _05285_);
  or (_05290_, _05289_, _05284_);
  or (_05291_, _05290_, _05277_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _05291_, _05262_);
  and (_05292_, _04552_, _04828_);
  and (_05293_, _04528_, _04826_);
  and (_05294_, _04531_, _04812_);
  or (_05295_, _05294_, _05293_);
  and (_05296_, _04564_, _04816_);
  and (_05297_, _04533_, _04824_);
  or (_05298_, _05297_, _05296_);
  or (_05299_, _05298_, _05295_);
  and (_05300_, _04572_, _04814_);
  and (_05301_, _04569_, _04818_);
  or (_05302_, _05301_, _05300_);
  and (_05303_, _04542_, _04822_);
  and (_05304_, _04576_, _04830_);
  or (_05305_, _05304_, _05303_);
  or (_05306_, _05305_, _05302_);
  or (_05307_, _05306_, _05299_);
  and (_05308_, _04596_, _04802_);
  and (_05309_, _04593_, _04797_);
  or (_05310_, _05309_, _05308_);
  and (_05311_, _04549_, _04799_);
  and (_05312_, _04600_, _04804_);
  or (_05313_, _05312_, _05311_);
  or (_05314_, _05313_, _05310_);
  and (_05315_, _04588_, _04794_);
  and (_05316_, _04546_, _04808_);
  and (_05317_, _04547_, _04792_);
  or (_05318_, _05317_, _05316_);
  or (_05319_, _05318_, _05315_);
  or (_05320_, _05319_, _05314_);
  or (_05321_, _05320_, _05307_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05321_, _05292_);
  and (_05322_, _04552_, _04869_);
  and (_05323_, _04531_, _04838_);
  and (_05324_, _04528_, _04856_);
  or (_05325_, _05324_, _05323_);
  and (_05326_, _04533_, _04858_);
  and (_05327_, _04564_, _04851_);
  or (_05328_, _05327_, _05326_);
  or (_05329_, _05328_, _05325_);
  and (_05330_, _04569_, _04840_);
  and (_05331_, _04572_, _04876_);
  or (_05332_, _05331_, _05330_);
  and (_05333_, _04576_, _04871_);
  and (_05334_, _04542_, _04878_);
  or (_05335_, _05334_, _05333_);
  or (_05336_, _05335_, _05332_);
  or (_05337_, _05336_, _05329_);
  and (_05338_, _04596_, _04862_);
  and (_05339_, _04593_, _04864_);
  or (_05340_, _05339_, _05338_);
  and (_05341_, _04549_, _04853_);
  and (_05342_, _04600_, _04867_);
  or (_05343_, _05342_, _05341_);
  or (_05344_, _05343_, _05340_);
  and (_05345_, _04588_, _04845_);
  and (_05346_, _04547_, _04842_);
  and (_05347_, _04546_, _04847_);
  or (_05348_, _05347_, _05346_);
  or (_05349_, _05348_, _05345_);
  or (_05350_, _05349_, _05344_);
  or (_05351_, _05350_, _05337_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05351_, _05322_);
  and (_05352_, _04552_, _04915_);
  and (_05353_, _04531_, _04884_);
  and (_05354_, _04528_, _04902_);
  or (_05355_, _05354_, _05353_);
  and (_05356_, _04533_, _04904_);
  and (_05357_, _04564_, _04897_);
  or (_05358_, _05357_, _05356_);
  or (_05359_, _05358_, _05355_);
  and (_05360_, _04569_, _04886_);
  and (_05361_, _04572_, _04922_);
  or (_05362_, _05361_, _05360_);
  and (_05363_, _04576_, _04917_);
  and (_05364_, _04542_, _04924_);
  or (_05365_, _05364_, _05363_);
  or (_05366_, _05365_, _05362_);
  or (_05367_, _05366_, _05359_);
  and (_05368_, _04596_, _04908_);
  and (_05369_, _04593_, _04910_);
  or (_05370_, _05369_, _05368_);
  and (_05371_, _04600_, _04913_);
  and (_05372_, _04549_, _04899_);
  or (_05373_, _05372_, _05371_);
  or (_05374_, _05373_, _05370_);
  and (_05375_, _04588_, _04891_);
  and (_05376_, _04547_, _04888_);
  and (_05377_, _04546_, _04893_);
  or (_05378_, _05377_, _05376_);
  or (_05379_, _05378_, _05375_);
  or (_05380_, _05379_, _05374_);
  or (_05381_, _05380_, _05367_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05381_, _05352_);
  and (_05382_, _04552_, _04966_);
  and (_05383_, _04531_, _04950_);
  and (_05384_, _04528_, _04964_);
  or (_05385_, _05384_, _05383_);
  and (_05386_, _04564_, _04954_);
  and (_05387_, _04533_, _04962_);
  or (_05388_, _05387_, _05386_);
  or (_05389_, _05388_, _05385_);
  and (_05390_, _04572_, _04960_);
  and (_05391_, _04569_, _04956_);
  or (_05392_, _05391_, _05390_);
  and (_05393_, _04576_, _04968_);
  and (_05394_, _04542_, _04952_);
  or (_05395_, _05394_, _05393_);
  or (_05396_, _05395_, _05392_);
  or (_05397_, _05396_, _05389_);
  and (_05398_, _04546_, _04946_);
  and (_05399_, _04547_, _04930_);
  and (_05400_, _04588_, _04932_);
  or (_05401_, _05400_, _05399_);
  or (_05402_, _05401_, _05398_);
  and (_05403_, _04593_, _04935_);
  and (_05404_, _04596_, _04940_);
  or (_05405_, _05404_, _05403_);
  and (_05406_, _04549_, _04937_);
  and (_05407_, _04600_, _04942_);
  or (_05408_, _05407_, _05406_);
  or (_05409_, _05408_, _05405_);
  or (_05410_, _05409_, _05402_);
  or (_05411_, _05410_, _05397_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05411_, _05382_);
  and (_05412_, _04552_, _05012_);
  and (_05413_, _04528_, _05010_);
  and (_05414_, _04531_, _04996_);
  or (_05415_, _05414_, _05413_);
  and (_05416_, _04564_, _04991_);
  and (_05417_, _04533_, _05008_);
  or (_05418_, _05417_, _05416_);
  or (_05419_, _05418_, _05415_);
  and (_05420_, _04572_, _05006_);
  and (_05421_, _04569_, _04989_);
  or (_05422_, _05421_, _05420_);
  and (_05423_, _04576_, _05014_);
  and (_05424_, _04542_, _04987_);
  or (_05425_, _05424_, _05423_);
  or (_05426_, _05425_, _05422_);
  or (_05427_, _05426_, _05419_);
  and (_05428_, _04596_, _04976_);
  and (_05429_, _04593_, _04978_);
  or (_05430_, _05429_, _05428_);
  and (_05431_, _04549_, _04983_);
  and (_05432_, _04600_, _04981_);
  or (_05433_, _05432_, _05431_);
  or (_05434_, _05433_, _05430_);
  and (_05435_, _04588_, _05000_);
  and (_05436_, _04547_, _04998_);
  and (_05437_, _04546_, _05002_);
  or (_05438_, _05437_, _05436_);
  or (_05439_, _05438_, _05435_);
  or (_05440_, _05439_, _05434_);
  or (_05441_, _05440_, _05427_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05441_, _05412_);
  and (_05442_, _04552_, _04723_);
  and (_05443_, _04547_, _04706_);
  and (_05444_, _04549_, _04704_);
  or (_05445_, _05444_, _05443_);
  and (_05446_, _04564_, _04731_);
  and (_05447_, _04546_, _04721_);
  or (_05448_, _05447_, _05446_);
  or (_05449_, _05448_, _05445_);
  and (_05450_, _04593_, _04737_);
  and (_05451_, _04576_, _04710_);
  or (_05452_, _05451_, _05450_);
  and (_05453_, _04531_, _04735_);
  and (_05454_, _04533_, _04733_);
  or (_05455_, _05454_, _05453_);
  or (_05456_, _05455_, _05452_);
  and (_05457_, _04600_, _04699_);
  and (_05458_, _04542_, _04729_);
  and (_05459_, _04588_, _04725_);
  or (_05460_, _05459_, _05458_);
  or (_05461_, _05460_, _05457_);
  and (_05462_, _04528_, _04719_);
  and (_05463_, _04596_, _04701_);
  or (_05464_, _05463_, _05462_);
  or (_05465_, _05464_, _05461_);
  and (_05466_, _04569_, _04714_);
  and (_05467_, _04572_, _04712_);
  or (_05468_, _05467_, _05466_);
  or (_05469_, _05468_, _05465_);
  or (_05470_, _05469_, _05456_);
  or (_05471_, _05470_, _05449_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _05471_, _05442_);
  and (_05472_, _04552_, _04752_);
  and (_05473_, _04547_, _04775_);
  and (_05474_, _04549_, _04761_);
  or (_05475_, _05474_, _05473_);
  and (_05476_, _04564_, _04766_);
  and (_05477_, _04546_, _04749_);
  or (_05478_, _05477_, _05476_);
  or (_05479_, _05478_, _05475_);
  and (_05480_, _04593_, _04779_);
  and (_05481_, _04576_, _04786_);
  or (_05482_, _05481_, _05480_);
  and (_05483_, _04531_, _04777_);
  and (_05484_, _04533_, _04764_);
  or (_05485_, _05484_, _05483_);
  or (_05486_, _05485_, _05482_);
  and (_05487_, _04600_, _04770_);
  and (_05488_, _04542_, _04784_);
  and (_05489_, _04588_, _04754_);
  or (_05490_, _05489_, _05488_);
  or (_05491_, _05490_, _05487_);
  and (_05492_, _04528_, _04745_);
  and (_05493_, _04596_, _04772_);
  or (_05494_, _05493_, _05492_);
  or (_05495_, _05494_, _05491_);
  and (_05496_, _04569_, _04758_);
  and (_05497_, _04572_, _04747_);
  or (_05498_, _05497_, _05496_);
  or (_05499_, _05498_, _05495_);
  or (_05500_, _05499_, _05486_);
  or (_05501_, _05500_, _05479_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _05501_, _05472_);
  and (_05502_, _04552_, _04794_);
  and (_05503_, _04547_, _04799_);
  and (_05504_, _04549_, _04804_);
  or (_05505_, _05504_, _05503_);
  and (_05506_, _04564_, _04824_);
  and (_05507_, _04546_, _04792_);
  or (_05508_, _05507_, _05506_);
  or (_05509_, _05508_, _05505_);
  and (_05510_, _04593_, _04830_);
  and (_05511_, _04576_, _04822_);
  or (_05512_, _05511_, _05510_);
  and (_05513_, _04531_, _04828_);
  and (_05514_, _04533_, _04826_);
  or (_05515_, _05514_, _05513_);
  or (_05516_, _05515_, _05512_);
  and (_05517_, _04596_, _04797_);
  and (_05518_, _04542_, _04814_);
  and (_05519_, _04588_, _04808_);
  or (_05520_, _05519_, _05518_);
  or (_05521_, _05520_, _05517_);
  and (_05522_, _04528_, _04812_);
  and (_05523_, _04600_, _04802_);
  or (_05524_, _05523_, _05522_);
  or (_05525_, _05524_, _05521_);
  and (_05526_, _04569_, _04816_);
  and (_05527_, _04572_, _04818_);
  or (_05528_, _05527_, _05526_);
  or (_05529_, _05528_, _05525_);
  or (_05530_, _05529_, _05516_);
  or (_05531_, _05530_, _05509_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _05531_, _05502_);
  and (_05532_, _04547_, _04853_);
  and (_05533_, _04588_, _04847_);
  or (_05534_, _05533_, _05532_);
  and (_05535_, _04572_, _04840_);
  and (_05536_, _04569_, _04851_);
  and (_05537_, _04564_, _04858_);
  or (_05538_, _05537_, _05536_);
  or (_05539_, _05538_, _05535_);
  or (_05540_, _05539_, _05534_);
  and (_05541_, _04552_, _04845_);
  and (_05542_, _04528_, _04838_);
  and (_05543_, _04531_, _04869_);
  and (_05544_, _04542_, _04876_);
  or (_05545_, _05544_, _05543_);
  or (_05546_, _05545_, _05542_);
  and (_05547_, _04576_, _04878_);
  and (_05548_, _04533_, _04856_);
  or (_05549_, _05548_, _05547_);
  or (_05550_, _05549_, _05546_);
  and (_05551_, _04600_, _04862_);
  and (_05552_, _04596_, _04864_);
  and (_05553_, _04593_, _04871_);
  or (_05554_, _05553_, _05552_);
  or (_05555_, _05554_, _05551_);
  and (_05556_, _04549_, _04867_);
  and (_05557_, _04546_, _04842_);
  or (_05558_, _05557_, _05556_);
  or (_05559_, _05558_, _05555_);
  or (_05560_, _05559_, _05550_);
  or (_05561_, _05560_, _05541_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _05561_, _05540_);
  and (_05562_, _04546_, _04888_);
  and (_05563_, _04547_, _04899_);
  and (_05564_, _04588_, _04893_);
  or (_05565_, _05564_, _05563_);
  or (_05566_, _05565_, _05562_);
  and (_05567_, _04533_, _04902_);
  and (_05568_, _04528_, _04884_);
  and (_05569_, _04531_, _04915_);
  and (_05570_, _04542_, _04922_);
  or (_05571_, _05570_, _05569_);
  or (_05572_, _05571_, _05568_);
  or (_05573_, _05572_, _05567_);
  or (_05574_, _05573_, _05566_);
  and (_05575_, _04552_, _04891_);
  and (_05576_, _04569_, _04897_);
  and (_05577_, _04564_, _04904_);
  or (_05578_, _05577_, _05576_);
  and (_05579_, _04572_, _04886_);
  and (_05580_, _04576_, _04924_);
  or (_05581_, _05580_, _05579_);
  or (_05582_, _05581_, _05578_);
  and (_05583_, _04593_, _04917_);
  and (_05584_, _04596_, _04910_);
  or (_05585_, _05584_, _05583_);
  and (_05586_, _04600_, _04908_);
  and (_05587_, _04549_, _04913_);
  or (_05588_, _05587_, _05586_);
  or (_05589_, _05588_, _05585_);
  or (_05590_, _05589_, _05582_);
  or (_05591_, _05590_, _05575_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _05591_, _05574_);
  and (_05592_, _04547_, _04937_);
  and (_05593_, _04588_, _04946_);
  or (_05594_, _05593_, _05592_);
  and (_05595_, _04572_, _04956_);
  and (_05596_, _04569_, _04954_);
  and (_05597_, _04564_, _04962_);
  or (_05598_, _05597_, _05596_);
  or (_05599_, _05598_, _05595_);
  or (_05600_, _05599_, _05594_);
  and (_05601_, _04552_, _04932_);
  and (_05602_, _04528_, _04950_);
  and (_05603_, _04531_, _04966_);
  and (_05604_, _04542_, _04960_);
  or (_05605_, _05604_, _05603_);
  or (_05606_, _05605_, _05602_);
  and (_05607_, _04576_, _04952_);
  and (_05608_, _04533_, _04964_);
  or (_05609_, _05608_, _05607_);
  or (_05610_, _05609_, _05606_);
  and (_05611_, _04600_, _04940_);
  and (_05612_, _04596_, _04935_);
  and (_05613_, _04593_, _04968_);
  or (_05614_, _05613_, _05612_);
  or (_05615_, _05614_, _05611_);
  and (_05616_, _04546_, _04930_);
  and (_05617_, _04549_, _04942_);
  or (_05618_, _05617_, _05616_);
  or (_05619_, _05618_, _05615_);
  or (_05620_, _05619_, _05610_);
  or (_05621_, _05620_, _05601_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _05621_, _05600_);
  and (_05622_, _04546_, _04998_);
  and (_05623_, _04547_, _04983_);
  and (_05624_, _04588_, _05002_);
  or (_05625_, _05624_, _05623_);
  or (_05626_, _05625_, _05622_);
  and (_05627_, _04533_, _05010_);
  and (_05628_, _04528_, _04996_);
  and (_05629_, _04531_, _05012_);
  and (_05630_, _04542_, _05006_);
  or (_05631_, _05630_, _05629_);
  or (_05632_, _05631_, _05628_);
  or (_05633_, _05632_, _05627_);
  or (_05634_, _05633_, _05626_);
  and (_05635_, _04552_, _05000_);
  and (_05636_, _04569_, _04991_);
  and (_05637_, _04564_, _05008_);
  or (_05638_, _05637_, _05636_);
  and (_05639_, _04576_, _04987_);
  and (_05640_, _04572_, _04989_);
  or (_05641_, _05640_, _05639_);
  or (_05642_, _05641_, _05638_);
  and (_05643_, _04593_, _05014_);
  and (_05644_, _04596_, _04978_);
  or (_05645_, _05644_, _05643_);
  and (_05646_, _04549_, _04981_);
  and (_05647_, _04600_, _04976_);
  or (_05648_, _05647_, _05646_);
  or (_05649_, _05648_, _05645_);
  or (_05650_, _05649_, _05642_);
  or (_05651_, _05650_, _05635_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _05651_, _05634_);
  not (_05652_, \uc8051golden_1.IRAM[15] [7]);
  not (_05653_, \uc8051golden_1.PC [1]);
  nand (_05654_, \uc8051golden_1.PC [1], \uc8051golden_1.PC [0]);
  not (_05655_, \uc8051golden_1.PC [3]);
  or (_05656_, \uc8051golden_1.PC [2], _05655_);
  or (_05657_, _05656_, _05654_);
  or (_05658_, _05657_, _00450_);
  or (_05659_, _05653_, \uc8051golden_1.PC [0]);
  or (_05660_, _05659_, _05656_);
  or (_05661_, _05660_, _00409_);
  and (_05662_, _05661_, _05658_);
  not (_05663_, \uc8051golden_1.PC [2]);
  or (_05664_, _05663_, \uc8051golden_1.PC [3]);
  or (_05665_, _05664_, _05654_);
  or (_05666_, _05665_, _00286_);
  or (_05667_, _05664_, _05659_);
  or (_05668_, _05667_, _00245_);
  and (_05669_, _05668_, _05666_);
  and (_05670_, _05669_, _05662_);
  nand (_05671_, \uc8051golden_1.PC [2], \uc8051golden_1.PC [3]);
  or (_05672_, _05671_, _05654_);
  or (_05673_, _05672_, _00633_);
  or (_05674_, _05671_, _05659_);
  or (_05675_, _05674_, _00592_);
  and (_05676_, _05675_, _05673_);
  or (_05677_, \uc8051golden_1.PC [2], \uc8051golden_1.PC [3]);
  or (_05678_, _05677_, _05654_);
  or (_05679_, _05678_, _00091_);
  or (_05680_, _05677_, _05659_);
  or (_05681_, _05680_, _00050_);
  and (_05682_, _05681_, _05679_);
  and (_05683_, _05682_, _05676_);
  and (_05684_, _05683_, _05670_);
  not (_05685_, \uc8051golden_1.PC [0]);
  or (_05686_, \uc8051golden_1.PC [1], _05685_);
  or (_05687_, _05686_, _05671_);
  or (_05688_, _05687_, _00532_);
  or (_05689_, \uc8051golden_1.PC [1], \uc8051golden_1.PC [0]);
  or (_05690_, _05689_, _05671_);
  or (_05691_, _05690_, _00491_);
  and (_05692_, _05691_, _05688_);
  or (_05693_, _05677_, _05689_);
  or (_05694_, _05693_, _43427_);
  or (_05695_, _05677_, _05686_);
  or (_05696_, _05695_, _00009_);
  and (_05697_, _05696_, _05694_);
  and (_05698_, _05697_, _05692_);
  or (_05699_, _05686_, _05656_);
  or (_05700_, _05699_, _00368_);
  or (_05701_, _05689_, _05656_);
  or (_05702_, _05701_, _00327_);
  and (_05703_, _05702_, _05700_);
  or (_05704_, _05686_, _05664_);
  or (_05705_, _05704_, _00204_);
  or (_05706_, _05689_, _05664_);
  or (_05707_, _05706_, _00135_);
  and (_05708_, _05707_, _05705_);
  and (_05709_, _05708_, _05703_);
  and (_05710_, _05709_, _05698_);
  and (_05711_, _05710_, _05684_);
  or (_05712_, _05657_, _00455_);
  or (_05713_, _05660_, _00414_);
  and (_05714_, _05713_, _05712_);
  or (_05715_, _05665_, _00291_);
  or (_05716_, _05667_, _00250_);
  and (_05717_, _05716_, _05715_);
  and (_05718_, _05717_, _05714_);
  or (_05719_, _05672_, _00638_);
  or (_05720_, _05674_, _00597_);
  and (_05721_, _05720_, _05719_);
  or (_05722_, _05678_, _00096_);
  or (_05723_, _05680_, _00055_);
  and (_05724_, _05723_, _05722_);
  and (_05725_, _05724_, _05721_);
  and (_05726_, _05725_, _05718_);
  or (_05727_, _05687_, _00537_);
  or (_05728_, _05690_, _00496_);
  and (_05729_, _05728_, _05727_);
  or (_05730_, _05693_, _43432_);
  or (_05731_, _05695_, _00014_);
  and (_05732_, _05731_, _05730_);
  and (_05733_, _05732_, _05729_);
  or (_05734_, _05699_, _00373_);
  or (_05735_, _05701_, _00332_);
  and (_05736_, _05735_, _05734_);
  or (_05737_, _05704_, _00209_);
  or (_05738_, _05706_, _00146_);
  and (_05739_, _05738_, _05737_);
  and (_05740_, _05739_, _05736_);
  and (_05741_, _05740_, _05733_);
  nand (_05742_, _05741_, _05726_);
  or (_05743_, _05742_, _05711_);
  or (_05744_, _05657_, _00460_);
  or (_05745_, _05660_, _00419_);
  and (_05746_, _05745_, _05744_);
  or (_05747_, _05665_, _00296_);
  or (_05748_, _05667_, _00255_);
  and (_05749_, _05748_, _05747_);
  and (_05750_, _05749_, _05746_);
  or (_05751_, _05672_, _00643_);
  or (_05752_, _05674_, _00602_);
  and (_05753_, _05752_, _05751_);
  or (_05754_, _05678_, _00101_);
  or (_05755_, _05680_, _00060_);
  and (_05756_, _05755_, _05754_);
  and (_05757_, _05756_, _05753_);
  and (_05758_, _05757_, _05750_);
  or (_05759_, _05687_, _00542_);
  or (_05760_, _05690_, _00501_);
  and (_05761_, _05760_, _05759_);
  or (_05762_, _05693_, _43437_);
  or (_05763_, _05695_, _00019_);
  and (_05764_, _05763_, _05762_);
  and (_05765_, _05764_, _05761_);
  or (_05766_, _05699_, _00378_);
  or (_05767_, _05701_, _00337_);
  and (_05768_, _05767_, _05766_);
  or (_05769_, _05704_, _00214_);
  or (_05770_, _05706_, _00157_);
  and (_05771_, _05770_, _05769_);
  and (_05772_, _05771_, _05768_);
  and (_05773_, _05772_, _05765_);
  nand (_05774_, _05773_, _05758_);
  or (_05775_, _05657_, _00465_);
  or (_05776_, _05660_, _00424_);
  and (_05777_, _05776_, _05775_);
  or (_05778_, _05665_, _00301_);
  or (_05779_, _05667_, _00260_);
  and (_05780_, _05779_, _05778_);
  and (_05781_, _05780_, _05777_);
  or (_05782_, _05672_, _00648_);
  or (_05783_, _05674_, _00607_);
  and (_05784_, _05783_, _05782_);
  or (_05785_, _05678_, _00106_);
  or (_05786_, _05680_, _00065_);
  and (_05787_, _05786_, _05785_);
  and (_05788_, _05787_, _05784_);
  and (_05789_, _05788_, _05781_);
  or (_05790_, _05687_, _00550_);
  or (_05791_, _05690_, _00506_);
  and (_05792_, _05791_, _05790_);
  or (_05793_, _05693_, _43442_);
  or (_05794_, _05695_, _00024_);
  and (_05795_, _05794_, _05793_);
  and (_05796_, _05795_, _05792_);
  or (_05797_, _05699_, _00383_);
  or (_05798_, _05701_, _00342_);
  and (_05799_, _05798_, _05797_);
  or (_05800_, _05704_, _00219_);
  or (_05801_, _05706_, _00168_);
  and (_05802_, _05801_, _05800_);
  and (_05803_, _05802_, _05799_);
  and (_05804_, _05803_, _05796_);
  nand (_05805_, _05804_, _05789_);
  or (_05806_, _05805_, _05774_);
  or (_05807_, _05806_, _05743_);
  not (_05808_, _05807_);
  or (_05809_, _05657_, _00470_);
  or (_05810_, _05660_, _00429_);
  and (_05811_, _05810_, _05809_);
  or (_05812_, _05665_, _00306_);
  or (_05813_, _05667_, _00265_);
  and (_05814_, _05813_, _05812_);
  and (_05815_, _05814_, _05811_);
  or (_05816_, _05672_, _00653_);
  or (_05817_, _05674_, _00612_);
  and (_05818_, _05817_, _05816_);
  or (_05819_, _05678_, _00111_);
  or (_05820_, _05680_, _00070_);
  and (_05821_, _05820_, _05819_);
  and (_05822_, _05821_, _05818_);
  and (_05823_, _05822_, _05815_);
  or (_05824_, _05687_, _00558_);
  or (_05825_, _05690_, _00511_);
  and (_05826_, _05825_, _05824_);
  or (_05827_, _05693_, _43447_);
  or (_05828_, _05695_, _00029_);
  and (_05829_, _05828_, _05827_);
  and (_05830_, _05829_, _05826_);
  or (_05831_, _05699_, _00388_);
  or (_05832_, _05701_, _00347_);
  and (_05833_, _05832_, _05831_);
  or (_05834_, _05704_, _00224_);
  or (_05835_, _05706_, _00179_);
  and (_05836_, _05835_, _05834_);
  and (_05837_, _05836_, _05833_);
  and (_05838_, _05837_, _05830_);
  nand (_05839_, _05838_, _05823_);
  or (_05840_, _05657_, _00475_);
  or (_05841_, _05660_, _00434_);
  and (_05842_, _05841_, _05840_);
  or (_05843_, _05665_, _00311_);
  or (_05844_, _05667_, _00270_);
  and (_05845_, _05844_, _05843_);
  and (_05846_, _05845_, _05842_);
  or (_05847_, _05672_, _00658_);
  or (_05848_, _05674_, _00617_);
  and (_05849_, _05848_, _05847_);
  or (_05850_, _05678_, _00116_);
  or (_05851_, _05680_, _00075_);
  and (_05852_, _05851_, _05850_);
  and (_05853_, _05852_, _05849_);
  and (_05854_, _05853_, _05846_);
  or (_05855_, _05687_, _00566_);
  or (_05856_, _05690_, _00516_);
  and (_05857_, _05856_, _05855_);
  or (_05858_, _05693_, _43452_);
  or (_05859_, _05695_, _00034_);
  and (_05860_, _05859_, _05858_);
  and (_05861_, _05860_, _05857_);
  or (_05862_, _05699_, _00393_);
  or (_05863_, _05701_, _00352_);
  and (_05864_, _05863_, _05862_);
  or (_05865_, _05704_, _00229_);
  or (_05866_, _05706_, _00188_);
  and (_05867_, _05866_, _05865_);
  and (_05868_, _05867_, _05864_);
  and (_05869_, _05868_, _05861_);
  nand (_05870_, _05869_, _05854_);
  or (_05871_, _05870_, _05839_);
  or (_05872_, _05657_, _00480_);
  or (_05873_, _05660_, _00439_);
  and (_05874_, _05873_, _05872_);
  or (_05875_, _05665_, _00316_);
  or (_05876_, _05667_, _00275_);
  and (_05877_, _05876_, _05875_);
  and (_05878_, _05877_, _05874_);
  or (_05879_, _05672_, _00663_);
  or (_05880_, _05674_, _00622_);
  and (_05881_, _05880_, _05879_);
  or (_05882_, _05678_, _00121_);
  or (_05883_, _05680_, _00080_);
  and (_05884_, _05883_, _05882_);
  and (_05885_, _05884_, _05881_);
  and (_05886_, _05885_, _05878_);
  or (_05887_, _05687_, _00574_);
  or (_05888_, _05690_, _00521_);
  and (_05889_, _05888_, _05887_);
  or (_05890_, _05693_, _43457_);
  or (_05891_, _05695_, _00039_);
  and (_05892_, _05891_, _05890_);
  and (_05893_, _05892_, _05889_);
  or (_05894_, _05699_, _00398_);
  or (_05895_, _05701_, _00357_);
  and (_05896_, _05895_, _05894_);
  or (_05897_, _05704_, _00234_);
  or (_05898_, _05706_, _00193_);
  and (_05899_, _05898_, _05897_);
  and (_05900_, _05899_, _05896_);
  and (_05901_, _05900_, _05893_);
  nand (_05902_, _05901_, _05886_);
  or (_05903_, _05657_, _00445_);
  or (_05904_, _05660_, _00404_);
  and (_05905_, _05904_, _05903_);
  or (_05906_, _05665_, _00281_);
  or (_05907_, _05667_, _00240_);
  and (_05908_, _05907_, _05906_);
  and (_05909_, _05908_, _05905_);
  or (_05910_, _05672_, _00628_);
  or (_05911_, _05674_, _00584_);
  and (_05912_, _05911_, _05910_);
  or (_05913_, _05678_, _00086_);
  or (_05914_, _05680_, _00045_);
  and (_05915_, _05914_, _05913_);
  and (_05916_, _05915_, _05912_);
  and (_05917_, _05916_, _05909_);
  or (_05918_, _05687_, _00527_);
  or (_05919_, _05690_, _00486_);
  and (_05920_, _05919_, _05918_);
  or (_05921_, _05693_, _43422_);
  or (_05922_, _05695_, _00004_);
  and (_05923_, _05922_, _05921_);
  and (_05924_, _05923_, _05920_);
  or (_05925_, _05699_, _00363_);
  or (_05926_, _05701_, _00322_);
  and (_05927_, _05926_, _05925_);
  or (_05928_, _05704_, _00199_);
  or (_05929_, _05706_, _00127_);
  and (_05930_, _05929_, _05928_);
  and (_05931_, _05930_, _05927_);
  and (_05932_, _05931_, _05924_);
  and (_05933_, _05932_, _05917_);
  or (_05934_, _05933_, _05902_);
  nor (_05935_, _05934_, _05871_);
  and (_05936_, _05935_, _05808_);
  and (_05937_, _05933_, _05902_);
  and (_05938_, _05838_, _05823_);
  and (_05939_, _05869_, _05854_);
  or (_05940_, _05939_, _05938_);
  not (_05941_, _05940_);
  and (_05942_, _05941_, _05937_);
  and (_05943_, _05942_, _05808_);
  nor (_05944_, _05943_, _05936_);
  not (_05945_, _05871_);
  and (_05946_, _05937_, _05945_);
  and (_05947_, _05946_, _05808_);
  not (_05948_, _05947_);
  or (_05949_, _05939_, _05839_);
  not (_05950_, _05949_);
  and (_05951_, _05950_, _05937_);
  and (_05952_, _05951_, _05808_);
  or (_05953_, _05870_, _05938_);
  not (_05954_, _05953_);
  and (_05955_, _05954_, _05937_);
  and (_05956_, _05955_, _05808_);
  nor (_05957_, _05956_, _05952_);
  and (_05958_, _05957_, _05948_);
  and (_05959_, _05958_, _05944_);
  and (_05960_, _05901_, _05886_);
  and (_05961_, _05933_, _05960_);
  and (_05962_, _05961_, _05945_);
  and (_05963_, _05962_, _05808_);
  not (_05964_, _05963_);
  and (_05965_, _05961_, _05941_);
  and (_05966_, _05965_, _05808_);
  not (_05967_, _05966_);
  and (_05968_, _05954_, _05961_);
  and (_05969_, _05968_, _05808_);
  and (_05970_, _05961_, _05950_);
  and (_05971_, _05970_, _05808_);
  nor (_05972_, _05971_, _05969_);
  and (_05973_, _05972_, _05967_);
  and (_05974_, _05973_, _05964_);
  and (_05975_, _05974_, _05959_);
  nor (_05976_, _05975_, _05653_);
  not (_05977_, _05976_);
  not (_05978_, _05806_);
  not (_05979_, _05711_);
  and (_05980_, _05742_, _05979_);
  and (_05981_, _05980_, _05978_);
  and (_05982_, _05981_, _05935_);
  and (_05983_, \uc8051golden_1.ACC [0], _05685_);
  not (_05984_, \uc8051golden_1.ACC [1]);
  and (_05985_, _05686_, _05659_);
  nor (_05986_, _05985_, _05984_);
  and (_05987_, _05985_, _05984_);
  nor (_05988_, _05987_, _05986_);
  and (_05989_, _05988_, _05983_);
  nor (_05990_, _05988_, _05983_);
  nor (_05991_, _05990_, _05989_);
  and (_05992_, _05991_, _05982_);
  or (_05993_, _05940_, _05934_);
  or (_05994_, _05993_, _05807_);
  or (_05995_, _05933_, _05960_);
  or (_05996_, _05995_, _05953_);
  or (_05997_, _05996_, _05807_);
  and (_05998_, _05997_, _05994_);
  or (_05999_, _05995_, _05871_);
  or (_06000_, _05999_, _05807_);
  or (_06001_, _05995_, _05949_);
  or (_06002_, _06001_, _05807_);
  and (_06003_, _06002_, _06000_);
  or (_06004_, _05995_, _05940_);
  or (_06005_, _06004_, _05807_);
  or (_06006_, _05934_, _05949_);
  or (_06007_, _06006_, _05807_);
  and (_06008_, _06007_, _06005_);
  and (_06009_, _06008_, _06003_);
  and (_06010_, _06009_, _05998_);
  not (_06011_, _05743_);
  not (_06012_, _05805_);
  and (_06013_, _06012_, _05774_);
  and (_06014_, _06013_, _06011_);
  and (_06015_, _06014_, _05935_);
  nor (_06016_, _05953_, _05934_);
  and (_06017_, _06016_, _05808_);
  nor (_06018_, _06017_, _06015_);
  and (_06019_, _06018_, _06010_);
  or (_06020_, _06019_, _05653_);
  not (_06021_, _05982_);
  and (_06022_, _06016_, _05981_);
  not (_06023_, _06022_);
  not (_06024_, _05985_);
  nand (_06025_, _06009_, _05998_);
  or (_06026_, _06025_, _06024_);
  nand (_06027_, _06026_, _06023_);
  and (_06028_, \uc8051golden_1.DPL [0], \uc8051golden_1.ACC [0]);
  and (_06029_, \uc8051golden_1.DPL [1], \uc8051golden_1.ACC [1]);
  nor (_06030_, \uc8051golden_1.DPL [1], \uc8051golden_1.ACC [1]);
  nor (_06031_, _06030_, _06029_);
  and (_06032_, _06031_, _06028_);
  nor (_06033_, _06031_, _06028_);
  nor (_06034_, _06033_, _06032_);
  nand (_06035_, _06034_, _06022_);
  and (_06036_, _06035_, _06018_);
  nand (_06037_, _06036_, _06027_);
  nand (_06038_, _06037_, _06021_);
  nand (_06039_, _06038_, _05975_);
  and (_06040_, _06039_, _06020_);
  or (_06041_, _06040_, _05992_);
  nand (_06042_, _06041_, _05977_);
  nor (_06043_, _05975_, \uc8051golden_1.PC [0]);
  not (_06044_, _06043_);
  not (_06045_, \uc8051golden_1.ACC [0]);
  and (_06046_, _06045_, \uc8051golden_1.PC [0]);
  nor (_06047_, _06046_, _05983_);
  and (_06048_, _06047_, _05982_);
  or (_06049_, _06019_, \uc8051golden_1.PC [0]);
  or (_06050_, _06025_, _05685_);
  nand (_06051_, _06050_, _06023_);
  nor (_06052_, \uc8051golden_1.DPL [0], \uc8051golden_1.ACC [0]);
  nor (_06053_, _06052_, _06028_);
  nand (_06054_, _06053_, _06022_);
  and (_06055_, _06054_, _06018_);
  nand (_06056_, _06055_, _06051_);
  nand (_06057_, _06056_, _06021_);
  nand (_06058_, _06057_, _05975_);
  and (_06059_, _06058_, _06049_);
  or (_06060_, _06059_, _06048_);
  nand (_06061_, _06060_, _06044_);
  or (_06062_, _06061_, _06042_);
  and (_06063_, \uc8051golden_1.PC [2], \uc8051golden_1.PC [1]);
  nor (_06064_, \uc8051golden_1.PC [2], \uc8051golden_1.PC [1]);
  nor (_06065_, _06064_, _06063_);
  nor (_06066_, _06065_, _05975_);
  not (_06067_, _06066_);
  nor (_06068_, _05989_, _05986_);
  nor (_06069_, _05654_, _05663_);
  and (_06070_, _05654_, _05663_);
  nor (_06071_, _06070_, _06069_);
  and (_06072_, _06071_, \uc8051golden_1.ACC [2]);
  nor (_06073_, _06071_, \uc8051golden_1.ACC [2]);
  nor (_06074_, _06073_, _06072_);
  not (_06075_, _06074_);
  nor (_06076_, _06075_, _06068_);
  and (_06077_, _06075_, _06068_);
  nor (_06078_, _06077_, _06076_);
  and (_06079_, _06078_, _05982_);
  or (_06080_, _06065_, _06019_);
  nor (_06081_, _06032_, _06029_);
  and (_06082_, \uc8051golden_1.DPL [2], \uc8051golden_1.ACC [2]);
  nor (_06083_, \uc8051golden_1.DPL [2], \uc8051golden_1.ACC [2]);
  nor (_06084_, _06083_, _06082_);
  not (_06085_, _06084_);
  nor (_06086_, _06085_, _06081_);
  and (_06087_, _06085_, _06081_);
  nor (_06088_, _06087_, _06086_);
  nand (_06089_, _06088_, _06022_);
  and (_06090_, _06089_, _06018_);
  or (_06091_, _06071_, _06025_);
  nand (_06092_, _06091_, _06023_);
  nand (_06093_, _06092_, _06090_);
  nand (_06094_, _06093_, _06021_);
  nand (_06095_, _06094_, _05975_);
  and (_06096_, _06095_, _06080_);
  or (_06097_, _06096_, _06079_);
  and (_06098_, _06097_, _06067_);
  nor (_06099_, _06076_, _06072_);
  not (_06100_, _05665_);
  nor (_06101_, _06069_, _05655_);
  nor (_06102_, _06101_, _06100_);
  nor (_06103_, _06102_, \uc8051golden_1.ACC [3]);
  and (_06104_, _06102_, \uc8051golden_1.ACC [3]);
  nor (_06105_, _06104_, _06103_);
  and (_06106_, _06105_, _06099_);
  nor (_06107_, _06105_, _06099_);
  nor (_06108_, _06107_, _06106_);
  and (_06109_, _06108_, _05982_);
  nor (_06110_, _06086_, _06082_);
  and (_06111_, \uc8051golden_1.DPL [3], \uc8051golden_1.ACC [3]);
  nor (_06112_, \uc8051golden_1.DPL [3], \uc8051golden_1.ACC [3]);
  nor (_06113_, _06112_, _06111_);
  not (_06114_, _06113_);
  nor (_06115_, _06114_, _06110_);
  and (_06116_, _06114_, _06110_);
  nor (_06117_, _06116_, _06115_);
  nand (_06118_, _06117_, _06022_);
  and (_06119_, _06118_, _06018_);
  not (_06120_, _06102_);
  or (_06121_, _06025_, _06120_);
  nor (_06122_, _05671_, _05653_);
  nor (_06123_, _06063_, \uc8051golden_1.PC [3]);
  nor (_06124_, _06123_, _06122_);
  or (_06125_, _06124_, _06010_);
  and (_06126_, _06125_, _06121_);
  nand (_06127_, _06126_, _06023_);
  nand (_06128_, _06127_, _06119_);
  or (_06129_, _06124_, _06018_);
  and (_06130_, _06129_, _06021_);
  and (_06131_, _06130_, _06128_);
  or (_06132_, _06131_, _06109_);
  and (_06133_, _06132_, _05975_);
  not (_06134_, _06124_);
  nor (_06135_, _06134_, _05975_);
  nor (_06136_, _06135_, _06133_);
  or (_06137_, _06136_, _06098_);
  or (_06138_, _06137_, _06062_);
  or (_06139_, _06138_, _00445_);
  nand (_06140_, _06097_, _06067_);
  or (_06141_, _06135_, _06133_);
  or (_06142_, _06141_, _06140_);
  or (_06143_, _06142_, _06062_);
  or (_06144_, _06143_, _00281_);
  and (_06145_, _06144_, _06139_);
  and (_06146_, _06041_, _05977_);
  or (_06147_, _06061_, _06146_);
  or (_06148_, _06147_, _06142_);
  or (_06149_, _06148_, _00199_);
  and (_06150_, _06060_, _06044_);
  or (_06151_, _06150_, _06146_);
  or (_06152_, _06141_, _06098_);
  or (_06153_, _06152_, _06151_);
  or (_06154_, _06153_, _43422_);
  and (_06155_, _06154_, _06149_);
  and (_06156_, _06155_, _06145_);
  or (_06157_, _06136_, _06140_);
  or (_06158_, _06157_, _06062_);
  or (_06159_, _06158_, _00628_);
  or (_06160_, _06152_, _06062_);
  or (_06161_, _06160_, _00086_);
  and (_06162_, _06161_, _06159_);
  or (_06163_, _06150_, _06042_);
  or (_06164_, _06163_, _06157_);
  or (_06165_, _06164_, _00584_);
  or (_06166_, _06147_, _06137_);
  or (_06167_, _06166_, _00363_);
  and (_06168_, _06167_, _06165_);
  and (_06169_, _06168_, _06162_);
  and (_06170_, _06169_, _06156_);
  or (_06171_, _06163_, _06142_);
  or (_06172_, _06171_, _00240_);
  or (_06173_, _06151_, _06142_);
  or (_06174_, _06173_, _00127_);
  and (_06175_, _06174_, _06172_);
  or (_06176_, _06163_, _06137_);
  or (_06177_, _06176_, _00404_);
  or (_06178_, _06152_, _06147_);
  or (_06179_, _06178_, _00004_);
  and (_06180_, _06179_, _06177_);
  and (_06181_, _06180_, _06175_);
  or (_06182_, _06157_, _06151_);
  or (_06183_, _06182_, _00486_);
  or (_06184_, _06163_, _06152_);
  or (_06185_, _06184_, _00045_);
  and (_06186_, _06185_, _06183_);
  or (_06187_, _06157_, _06147_);
  or (_06188_, _06187_, _00527_);
  or (_06189_, _06151_, _06137_);
  or (_06190_, _06189_, _00322_);
  and (_06191_, _06190_, _06188_);
  and (_06192_, _06191_, _06186_);
  and (_06193_, _06192_, _06181_);
  nand (_06194_, _06193_, _06170_);
  and (_06195_, _06014_, _05962_);
  not (_06196_, _06195_);
  nor (_06197_, _06196_, _06194_);
  nor (_06198_, _06158_, _00638_);
  nor (_06199_, _06138_, _00455_);
  nor (_06200_, _06199_, _06198_);
  nor (_06201_, _06173_, _00146_);
  nor (_06202_, _06153_, _43432_);
  nor (_06203_, _06202_, _06201_);
  and (_06204_, _06203_, _06200_);
  nor (_06205_, _06176_, _00414_);
  nor (_06206_, _06166_, _00373_);
  nor (_06207_, _06206_, _06205_);
  nor (_06208_, _06164_, _00597_);
  nor (_06209_, _06182_, _00496_);
  nor (_06210_, _06209_, _06208_);
  and (_06211_, _06210_, _06207_);
  and (_06212_, _06211_, _06204_);
  nor (_06213_, _06143_, _00291_);
  nor (_06214_, _06171_, _00250_);
  nor (_06215_, _06214_, _06213_);
  nor (_06216_, _06148_, _00209_);
  nor (_06217_, _06160_, _00096_);
  nor (_06218_, _06217_, _06216_);
  and (_06219_, _06218_, _06215_);
  nor (_06220_, _06184_, _00055_);
  nor (_06221_, _06178_, _00014_);
  nor (_06222_, _06221_, _06220_);
  nor (_06223_, _06187_, _00537_);
  nor (_06224_, _06189_, _00332_);
  nor (_06225_, _06224_, _06223_);
  and (_06226_, _06225_, _06222_);
  and (_06227_, _06226_, _06219_);
  and (_06228_, _06227_, _06212_);
  not (_06229_, _06228_);
  and (_06230_, _06229_, _06197_);
  not (_06231_, _05742_);
  and (_06232_, _06231_, _05711_);
  and (_06233_, _06232_, _05978_);
  and (_06234_, _06233_, _05968_);
  nor (_06235_, _06178_, _00029_);
  nor (_06236_, _06184_, _00070_);
  nor (_06237_, _06236_, _06235_);
  nor (_06238_, _06187_, _00558_);
  nor (_06239_, _06143_, _00306_);
  nor (_06240_, _06239_, _06238_);
  and (_06241_, _06240_, _06237_);
  nor (_06242_, _06138_, _00470_);
  nor (_06243_, _06166_, _00388_);
  nor (_06244_, _06243_, _06242_);
  nor (_06245_, _06173_, _00179_);
  nor (_06246_, _06153_, _43447_);
  nor (_06247_, _06246_, _06245_);
  and (_06248_, _06247_, _06244_);
  and (_06249_, _06248_, _06241_);
  nor (_06250_, _06158_, _00653_);
  nor (_06251_, _06164_, _00612_);
  nor (_06252_, _06251_, _06250_);
  nor (_06253_, _06182_, _00511_);
  nor (_06254_, _06189_, _00347_);
  nor (_06255_, _06254_, _06253_);
  and (_06256_, _06255_, _06252_);
  nor (_06257_, _06148_, _00224_);
  nor (_06258_, _06171_, _00265_);
  nor (_06259_, _06258_, _06257_);
  nor (_06260_, _06176_, _00429_);
  nor (_06261_, _06160_, _00111_);
  nor (_06262_, _06261_, _06260_);
  and (_06263_, _06262_, _06259_);
  and (_06264_, _06263_, _06256_);
  and (_06265_, _06264_, _06249_);
  nor (_06266_, _06265_, _06194_);
  and (_06267_, _06266_, _06234_);
  not (_06268_, \uc8051golden_1.SP [1]);
  and (_06269_, _06268_, \uc8051golden_1.SP [0]);
  not (_06270_, \uc8051golden_1.SP [0]);
  and (_06271_, \uc8051golden_1.SP [1], _06270_);
  nor (_06272_, _06271_, _06269_);
  not (_06273_, _06272_);
  and (_06274_, _06273_, _05966_);
  and (_06275_, _06014_, _05942_);
  not (_06276_, _06275_);
  nor (_06277_, _06276_, _06194_);
  and (_06278_, _06277_, _06229_);
  not (_06279_, _06015_);
  and (_06280_, _06013_, _05742_);
  and (_06281_, _06280_, _05935_);
  not (_06282_, _06281_);
  not (_06283_, _05774_);
  and (_06284_, _05805_, _06231_);
  and (_06285_, _06284_, _06283_);
  and (_06286_, _06285_, _05935_);
  not (_06287_, _05935_);
  and (_06288_, _05805_, _06283_);
  and (_06289_, _06288_, _05742_);
  and (_06290_, _05805_, _05774_);
  nor (_06291_, _06290_, _06289_);
  nor (_06292_, _06291_, _06287_);
  nor (_06293_, _06292_, _06286_);
  and (_06294_, _06293_, _06282_);
  and (_06295_, _06294_, _06279_);
  or (_06296_, _06295_, _06194_);
  nor (_06297_, _06296_, _06229_);
  and (_06298_, _05742_, _05711_);
  and (_06299_, _06298_, _05978_);
  and (_06300_, _06299_, _06016_);
  and (_06301_, _06300_, _06266_);
  not (_06302_, _06004_);
  and (_06303_, _06280_, _06302_);
  not (_06304_, _06005_);
  and (_06305_, _06299_, _05970_);
  not (_06306_, _06305_);
  and (_06307_, _06014_, _05970_);
  not (_06308_, _06307_);
  not (_06309_, _06194_);
  nor (_06310_, _06143_, _00316_);
  nor (_06311_, _06160_, _00121_);
  nor (_06312_, _06311_, _06310_);
  nor (_06313_, _06176_, _00439_);
  nor (_06314_, _06189_, _00357_);
  nor (_06315_, _06314_, _06313_);
  and (_06316_, _06315_, _06312_);
  nor (_06317_, _06171_, _00275_);
  nor (_06318_, _06148_, _00234_);
  nor (_06319_, _06318_, _06317_);
  nor (_06320_, _06184_, _00080_);
  nor (_06321_, _06178_, _00039_);
  nor (_06322_, _06321_, _06320_);
  and (_06323_, _06322_, _06319_);
  and (_06324_, _06323_, _06316_);
  nor (_06325_, _06164_, _00622_);
  nor (_06326_, _06166_, _00398_);
  nor (_06327_, _06326_, _06325_);
  nor (_06328_, _06187_, _00574_);
  nor (_06329_, _06138_, _00480_);
  nor (_06330_, _06329_, _06328_);
  and (_06331_, _06330_, _06327_);
  nor (_06332_, _06173_, _00193_);
  nor (_06333_, _06153_, _43457_);
  nor (_06334_, _06333_, _06332_);
  nor (_06335_, _06158_, _00663_);
  nor (_06336_, _06182_, _00521_);
  nor (_06337_, _06336_, _06335_);
  and (_06338_, _06337_, _06334_);
  and (_06339_, _06338_, _06331_);
  and (_06340_, _06339_, _06324_);
  and (_06341_, _06340_, _06309_);
  or (_06342_, _06171_, _00260_);
  or (_06343_, _06148_, _00219_);
  and (_06344_, _06343_, _06342_);
  or (_06345_, _06158_, _00648_);
  or (_06346_, _06138_, _00465_);
  and (_06347_, _06346_, _06345_);
  and (_06348_, _06347_, _06344_);
  or (_06349_, _06176_, _00424_);
  or (_06350_, _06166_, _00383_);
  and (_06351_, _06350_, _06349_);
  or (_06352_, _06164_, _00607_);
  or (_06353_, _06182_, _00506_);
  and (_06354_, _06353_, _06352_);
  and (_06355_, _06354_, _06351_);
  and (_06356_, _06355_, _06348_);
  or (_06357_, _06153_, _43442_);
  or (_06358_, _06184_, _00065_);
  and (_06359_, _06358_, _06357_);
  or (_06360_, _06143_, _00301_);
  or (_06361_, _06173_, _00168_);
  and (_06362_, _06361_, _06360_);
  and (_06363_, _06362_, _06359_);
  or (_06364_, _06187_, _00550_);
  or (_06365_, _06189_, _00342_);
  and (_06366_, _06365_, _06364_);
  or (_06367_, _06160_, _00106_);
  or (_06368_, _06178_, _00024_);
  and (_06369_, _06368_, _06367_);
  and (_06370_, _06369_, _06366_);
  and (_06371_, _06370_, _06363_);
  and (_06372_, _06371_, _06356_);
  and (_06373_, _06372_, _06194_);
  nor (_06374_, _06373_, _06341_);
  and (_06375_, _06299_, _05942_);
  and (_06376_, _06299_, _05935_);
  nor (_06377_, _06376_, _06375_);
  nor (_06378_, _06377_, _06374_);
  not (_06379_, _06290_);
  nor (_06380_, _06379_, _06006_);
  not (_06381_, _06006_);
  and (_06382_, _06288_, _06381_);
  nor (_06383_, _06382_, _06380_);
  not (_06384_, _06383_);
  and (_06385_, _06384_, _06372_);
  not (_06386_, _05993_);
  and (_06387_, _06299_, _06386_);
  and (_06388_, _06233_, _06386_);
  nor (_06389_, _06388_, _06387_);
  not (_06390_, _06389_);
  and (_06391_, _06390_, _06374_);
  not (_06392_, _05999_);
  and (_06393_, _06299_, _06392_);
  not (_06394_, _05996_);
  and (_06395_, _06299_, _06394_);
  not (_06396_, _06395_);
  nor (_06397_, _06396_, _06374_);
  not (_06398_, \uc8051golden_1.SP [3]);
  and (_06399_, _06233_, _06394_);
  and (_06400_, _06399_, _06398_);
  and (_06401_, _06014_, _06394_);
  not (_06402_, _06001_);
  and (_06403_, _06014_, _06402_);
  nor (_06404_, _06403_, _06401_);
  or (_06405_, _06404_, _06372_);
  and (_06406_, _06014_, _06392_);
  nor (_06407_, _06399_, _06395_);
  nand (_06408_, _06404_, \uc8051golden_1.PSW [3]);
  and (_06409_, _06408_, _06407_);
  or (_06410_, _06409_, _06406_);
  and (_06411_, _06410_, _06405_);
  or (_06412_, _06411_, _06400_);
  nor (_06413_, _06412_, _06397_);
  not (_06414_, _06406_);
  nor (_06415_, _06414_, _06372_);
  nor (_06416_, _06415_, _06413_);
  nor (_06417_, _06416_, _06393_);
  and (_06418_, _06393_, _06374_);
  and (_06419_, _06233_, _06392_);
  and (_06420_, _06014_, _06386_);
  nor (_06421_, _06420_, _06419_);
  not (_06422_, _06421_);
  nor (_06423_, _06422_, _06418_);
  not (_06424_, _06423_);
  nor (_06425_, _06424_, _06417_);
  and (_06426_, _06422_, _06372_);
  or (_06427_, _06390_, _06426_);
  nor (_06428_, _06427_, _06425_);
  or (_06429_, _06428_, _06384_);
  nor (_06430_, _06429_, _06391_);
  nor (_06431_, _06430_, _06385_);
  and (_06432_, _06233_, _06381_);
  and (_06433_, _06299_, _06381_);
  nor (_06434_, _06433_, _06432_);
  not (_06435_, _06434_);
  nor (_06436_, _06435_, _06431_);
  and (_06437_, _06016_, _06014_);
  nor (_06438_, _06434_, _06374_);
  nor (_06439_, _06438_, _06437_);
  not (_06440_, _06439_);
  or (_06441_, _06440_, _06436_);
  not (_06442_, _06437_);
  nor (_06443_, _06442_, _06372_);
  nor (_06444_, _06443_, _06300_);
  nand (_06445_, _06444_, _06441_);
  not (_06446_, _06300_);
  nor (_06447_, _06374_, _06446_);
  nor (_06448_, _06447_, _06015_);
  nand (_06449_, _06448_, _06445_);
  not (_06450_, _06377_);
  and (_06451_, _06290_, _05980_);
  and (_06452_, _06288_, _06232_);
  and (_06453_, _06290_, _06011_);
  or (_06454_, _06453_, _06452_);
  nor (_06455_, _06454_, _06451_);
  or (_06456_, _06455_, _05993_);
  and (_06457_, _06280_, _06386_);
  nor (_06458_, _06457_, _06401_);
  and (_06459_, _06458_, _06456_);
  and (_06460_, _06233_, _05965_);
  nor (_06461_, _06460_, _06234_);
  and (_06462_, _06290_, _06232_);
  nor (_06463_, _06462_, _06289_);
  or (_06464_, _06463_, _05993_);
  and (_06465_, _06299_, _05968_);
  and (_06466_, _06288_, _06011_);
  and (_06467_, _06466_, _06386_);
  nor (_06468_, _06467_, _06465_);
  and (_06469_, _06468_, _06464_);
  and (_06470_, _06469_, _06461_);
  and (_06471_, _06470_, _06459_);
  and (_06472_, _06233_, _06016_);
  not (_06473_, _06472_);
  and (_06474_, _05981_, _05951_);
  and (_06475_, _06299_, _05962_);
  nor (_06476_, _06475_, _06474_);
  and (_06477_, _06476_, _06473_);
  and (_06478_, _05981_, _05955_);
  and (_06479_, _05981_, _05946_);
  nor (_06480_, _06479_, _06478_);
  and (_06481_, _06232_, _06013_);
  and (_06482_, _06481_, _06386_);
  and (_06483_, _06290_, _06298_);
  and (_06484_, _06483_, _06386_);
  nor (_06485_, _06484_, _06482_);
  and (_06486_, _06485_, _06480_);
  and (_06487_, _06233_, _05970_);
  nor (_06488_, _06487_, _06420_);
  and (_06489_, _06488_, _06276_);
  and (_06490_, _06489_, _06486_);
  and (_06491_, _06490_, _06477_);
  and (_06492_, _06491_, _06471_);
  and (_06493_, _06492_, _05685_);
  nor (_06494_, _06493_, _05653_);
  and (_06495_, _06493_, _05653_);
  nor (_06496_, _06495_, _06494_);
  nor (_06497_, _06492_, _05685_);
  or (_06498_, _06497_, _06493_);
  nor (_06499_, _06498_, _06496_);
  not (_06500_, _06065_);
  nor (_06501_, _06492_, _06500_);
  and (_06502_, _06492_, _06071_);
  nor (_06503_, _06502_, _06501_);
  nor (_06504_, _06492_, _06134_);
  and (_06505_, _06492_, _06120_);
  nor (_06506_, _06505_, _06504_);
  and (_06507_, _06506_, _06503_);
  and (_06508_, _06507_, _06499_);
  and (_06509_, _06508_, _04845_);
  not (_06510_, _06496_);
  nor (_06511_, _06498_, _06510_);
  and (_06512_, _06511_, _06507_);
  and (_06513_, _06512_, _04842_);
  nor (_06514_, _06513_, _06509_);
  nor (_06515_, _06506_, _06503_);
  and (_06516_, _06515_, _06499_);
  and (_06517_, _06516_, _04858_);
  not (_06518_, _06506_);
  nor (_06519_, _06518_, _06503_);
  and (_06520_, _06519_, _06511_);
  and (_06521_, _06520_, _04864_);
  nor (_06522_, _06521_, _06517_);
  and (_06523_, _06522_, _06514_);
  and (_06524_, _06518_, _06503_);
  and (_06525_, _06498_, _06496_);
  and (_06526_, _06525_, _06524_);
  and (_06527_, _06526_, _04851_);
  and (_06528_, _06524_, _06499_);
  and (_06529_, _06528_, _04878_);
  nor (_06530_, _06529_, _06527_);
  and (_06531_, _06498_, _06510_);
  and (_06532_, _06531_, _06519_);
  and (_06533_, _06532_, _04862_);
  and (_06534_, _06531_, _06507_);
  and (_06535_, _06534_, _04847_);
  nor (_06536_, _06535_, _06533_);
  and (_06537_, _06536_, _06530_);
  and (_06538_, _06537_, _06523_);
  and (_06539_, _06525_, _06515_);
  and (_06540_, _06539_, _04869_);
  and (_06541_, _06515_, _06511_);
  and (_06542_, _06541_, _04838_);
  nor (_06543_, _06542_, _06540_);
  and (_06544_, _06531_, _06515_);
  and (_06545_, _06544_, _04856_);
  and (_06546_, _06531_, _06524_);
  and (_06547_, _06546_, _04876_);
  nor (_06548_, _06547_, _06545_);
  and (_06549_, _06548_, _06543_);
  and (_06550_, _06524_, _06511_);
  and (_06551_, _06550_, _04840_);
  and (_06552_, _06525_, _06507_);
  and (_06553_, _06552_, _04853_);
  nor (_06554_, _06553_, _06551_);
  and (_06555_, _06525_, _06519_);
  and (_06556_, _06555_, _04871_);
  and (_06557_, _06519_, _06499_);
  and (_06558_, _06557_, _04867_);
  nor (_06559_, _06558_, _06556_);
  and (_06560_, _06559_, _06554_);
  and (_06561_, _06560_, _06549_);
  and (_06562_, _06561_, _06538_);
  nor (_06563_, _06562_, _06279_);
  nor (_06564_, _06563_, _06450_);
  and (_06565_, _06564_, _06449_);
  or (_06566_, _06565_, _06378_);
  and (_06567_, _06014_, _05955_);
  not (_06568_, _06567_);
  and (_06569_, _06299_, _05955_);
  nor (_06570_, _06569_, _06478_);
  and (_06571_, _06570_, _06568_);
  and (_06572_, _06299_, _05946_);
  nor (_06573_, _06572_, _06479_);
  and (_06574_, _06014_, _05946_);
  not (_06575_, _06574_);
  and (_06576_, _06575_, _06573_);
  and (_06577_, _06576_, _06571_);
  and (_06578_, _06014_, _05965_);
  not (_06579_, _06578_);
  and (_06580_, _06014_, _05951_);
  not (_06581_, _06580_);
  and (_06582_, _06299_, _05951_);
  nor (_06583_, _06582_, _06474_);
  and (_06584_, _06583_, _06581_);
  and (_06585_, _06584_, _06579_);
  and (_06586_, _06585_, _06577_);
  nand (_06587_, _06586_, _06566_);
  and (_06588_, _06299_, _05965_);
  not (_06589_, _06372_);
  nor (_06590_, _06586_, _06589_);
  nor (_06591_, _06590_, _06588_);
  and (_06592_, _06591_, _06587_);
  and (_06593_, _06588_, \uc8051golden_1.SP [3]);
  or (_06594_, _06593_, _06460_);
  nor (_06595_, _06594_, _06592_);
  not (_06596_, _06460_);
  nor (_06597_, _06374_, _06596_);
  or (_06598_, _06597_, _06595_);
  and (_06599_, _06598_, _06308_);
  and (_06600_, _06307_, _06372_);
  or (_06601_, _06600_, _06599_);
  nand (_06602_, _06601_, _06306_);
  and (_06603_, _06305_, _06398_);
  nor (_06604_, _06603_, _06487_);
  nand (_06605_, _06604_, _06602_);
  and (_06606_, _06014_, _05968_);
  and (_06607_, _06487_, _06374_);
  nor (_06608_, _06607_, _06606_);
  nand (_06609_, _06608_, _06605_);
  and (_06610_, _06606_, _06372_);
  nor (_06611_, _06610_, _06234_);
  and (_06612_, _06611_, _06609_);
  and (_06613_, _06374_, _06234_);
  or (_06614_, _06613_, _06612_);
  nand (_06615_, _06614_, _06196_);
  nor (_06616_, _06372_, _06196_);
  not (_06617_, _06616_);
  and (_06618_, _06617_, _06615_);
  nor (_06619_, _06143_, _00311_);
  nor (_06620_, _06160_, _00116_);
  nor (_06621_, _06620_, _06619_);
  nor (_06622_, _06182_, _00516_);
  nor (_06623_, _06189_, _00352_);
  nor (_06625_, _06623_, _06622_);
  and (_06626_, _06625_, _06621_);
  nor (_06627_, _06184_, _00075_);
  nor (_06628_, _06178_, _00034_);
  nor (_06629_, _06628_, _06627_);
  nor (_06630_, _06171_, _00270_);
  nor (_06631_, _06173_, _00188_);
  nor (_06632_, _06631_, _06630_);
  and (_06633_, _06632_, _06629_);
  and (_06634_, _06633_, _06626_);
  nor (_06635_, _06138_, _00475_);
  nor (_06636_, _06176_, _00434_);
  nor (_06637_, _06636_, _06635_);
  nor (_06638_, _06158_, _00658_);
  nor (_06639_, _06166_, _00393_);
  nor (_06640_, _06639_, _06638_);
  and (_06641_, _06640_, _06637_);
  nor (_06642_, _06164_, _00617_);
  nor (_06643_, _06187_, _00566_);
  nor (_06644_, _06643_, _06642_);
  nor (_06645_, _06148_, _00229_);
  nor (_06646_, _06153_, _43452_);
  nor (_06647_, _06646_, _06645_);
  and (_06648_, _06647_, _06644_);
  and (_06649_, _06648_, _06641_);
  and (_06650_, _06649_, _06634_);
  nor (_06651_, _06650_, _06194_);
  nor (_06652_, _06487_, _06393_);
  and (_06653_, _06652_, _06461_);
  and (_06654_, _06396_, _06377_);
  and (_06655_, _06434_, _06389_);
  and (_06656_, _06655_, _06654_);
  and (_06657_, _06656_, _06653_);
  not (_06658_, _06657_);
  and (_06659_, _06658_, _06651_);
  not (_06660_, _06659_);
  and (_06661_, _06651_, _06300_);
  not (_06662_, _06661_);
  nor (_06663_, _06153_, _43437_);
  nor (_06664_, _06184_, _00060_);
  nor (_06665_, _06664_, _06663_);
  nor (_06666_, _06182_, _00501_);
  nor (_06667_, _06143_, _00296_);
  nor (_06668_, _06667_, _06666_);
  and (_06669_, _06668_, _06665_);
  nor (_06670_, _06138_, _00460_);
  nor (_06671_, _06189_, _00337_);
  nor (_06672_, _06671_, _06670_);
  nor (_06673_, _06148_, _00214_);
  nor (_06674_, _06178_, _00019_);
  nor (_06675_, _06674_, _06673_);
  and (_06676_, _06675_, _06672_);
  and (_06677_, _06676_, _06669_);
  nor (_06678_, _06158_, _00643_);
  nor (_06679_, _06164_, _00602_);
  nor (_06680_, _06679_, _06678_);
  nor (_06681_, _06187_, _00542_);
  nor (_06682_, _06166_, _00378_);
  nor (_06683_, _06682_, _06681_);
  and (_06684_, _06683_, _06680_);
  nor (_06685_, _06176_, _00419_);
  nor (_06686_, _06160_, _00101_);
  nor (_06687_, _06686_, _06685_);
  nor (_06688_, _06171_, _00255_);
  nor (_06689_, _06173_, _00157_);
  nor (_06690_, _06689_, _06688_);
  and (_06691_, _06690_, _06687_);
  and (_06692_, _06691_, _06684_);
  and (_06693_, _06692_, _06677_);
  nor (_06694_, _06437_, _06406_);
  and (_06695_, _06694_, _06421_);
  and (_06696_, _06695_, _06404_);
  and (_06697_, _06696_, _06584_);
  and (_06698_, _06697_, _06577_);
  and (_06699_, _06698_, _06383_);
  nor (_06700_, _06606_, _06195_);
  and (_06701_, _06700_, _06579_);
  and (_06702_, _06701_, _06308_);
  and (_06703_, _06702_, _06699_);
  nor (_06704_, _06703_, _06693_);
  not (_06705_, _06704_);
  and (_06706_, _06539_, _04828_);
  and (_06707_, _06526_, _04816_);
  nor (_06708_, _06707_, _06706_);
  and (_06709_, _06557_, _04804_);
  and (_06710_, _06508_, _04794_);
  nor (_06711_, _06710_, _06709_);
  and (_06712_, _06711_, _06708_);
  and (_06713_, _06541_, _04812_);
  and (_06714_, _06544_, _04826_);
  nor (_06715_, _06714_, _06713_);
  and (_06716_, _06516_, _04824_);
  and (_06717_, _06528_, _04822_);
  nor (_06718_, _06717_, _06716_);
  and (_06719_, _06718_, _06715_);
  and (_06720_, _06719_, _06712_);
  and (_06721_, _06555_, _04830_);
  and (_06722_, _06520_, _04797_);
  nor (_06723_, _06722_, _06721_);
  and (_06724_, _06532_, _04802_);
  and (_06725_, _06552_, _04799_);
  nor (_06726_, _06725_, _06724_);
  and (_06727_, _06726_, _06723_);
  and (_06728_, _06550_, _04818_);
  and (_06729_, _06546_, _04814_);
  nor (_06730_, _06729_, _06728_);
  and (_06731_, _06512_, _04792_);
  and (_06732_, _06534_, _04808_);
  nor (_06733_, _06732_, _06731_);
  and (_06734_, _06733_, _06730_);
  and (_06735_, _06734_, _06727_);
  and (_06736_, _06735_, _06720_);
  nor (_06737_, _06736_, _06279_);
  not (_06738_, \uc8051golden_1.SP [2]);
  nor (_06739_, _06399_, _06588_);
  nor (_06740_, _06739_, _06738_);
  not (_06741_, _06740_);
  and (_06742_, _06290_, _05742_);
  not (_06743_, _06742_);
  nor (_06744_, _05953_, _05933_);
  not (_06745_, _06744_);
  nor (_06746_, _05965_, _05951_);
  and (_06747_, _06746_, _06745_);
  nor (_06748_, _06747_, _06743_);
  not (_06749_, _06748_);
  and (_06750_, _06742_, _06392_);
  and (_06751_, _06290_, _06231_);
  and (_06752_, _06751_, _05951_);
  nor (_06753_, _06752_, _06750_);
  and (_06754_, _06462_, _05965_);
  and (_06755_, _06462_, _06402_);
  nor (_06756_, _06755_, _06754_);
  and (_06757_, _06756_, _06753_);
  and (_06758_, _06757_, _06749_);
  and (_06759_, _06758_, _06741_);
  and (_06760_, _06001_, _05993_);
  nor (_06761_, _06760_, _06743_);
  not (_06762_, _06761_);
  and (_06763_, _06742_, _05970_);
  and (_06764_, _06742_, _05962_);
  nor (_06765_, _06764_, _06763_);
  not (_06766_, _06765_);
  not (_06767_, _06751_);
  and (_06768_, _05993_, _06287_);
  nor (_06769_, _06768_, _06767_);
  nor (_06770_, _06769_, _06766_);
  and (_06771_, _06770_, _06762_);
  and (_06772_, _06751_, _05968_);
  and (_06773_, _06751_, _06392_);
  nor (_06774_, _06773_, _06772_);
  not (_06775_, _06774_);
  or (_06776_, _05970_, _05955_);
  and (_06777_, _06776_, _06751_);
  nor (_06778_, _06777_, _06775_);
  and (_06779_, _06305_, \uc8051golden_1.SP [2]);
  and (_06780_, _06751_, _06016_);
  nor (_06781_, _06780_, _06779_);
  and (_06782_, _06781_, _06778_);
  and (_06783_, _06742_, _05968_);
  and (_06784_, _06290_, _05946_);
  nor (_06785_, _06784_, _06783_);
  and (_06786_, _06751_, _05962_);
  and (_06787_, _06751_, _06394_);
  nor (_06788_, _06787_, _06786_);
  and (_06789_, _06788_, _06785_);
  and (_06790_, _06453_, _06402_);
  and (_06791_, _06742_, _05935_);
  nor (_06792_, _06791_, _06790_);
  and (_06793_, _06453_, _05965_);
  and (_06794_, _06742_, _05955_);
  nor (_06795_, _06794_, _06793_);
  and (_06796_, _06795_, _06792_);
  and (_06797_, _06796_, _06789_);
  and (_06798_, _06797_, _06782_);
  and (_06799_, _06798_, _06771_);
  and (_06800_, _06799_, _06759_);
  not (_06801_, _06800_);
  nor (_06802_, _06801_, _06737_);
  and (_06803_, _06802_, _06705_);
  and (_06804_, _06803_, _06662_);
  and (_06805_, _06804_, _06660_);
  not (_06806_, \uc8051golden_1.IRAM[1] [1]);
  not (_06807_, _06234_);
  or (_06808_, _06372_, _06194_);
  nor (_06809_, _06808_, _06446_);
  or (_06810_, _06164_, _00592_);
  or (_06811_, _06187_, _00532_);
  and (_06812_, _06811_, _06810_);
  or (_06813_, _06138_, _00450_);
  or (_06814_, _06176_, _00409_);
  and (_06815_, _06814_, _06813_);
  and (_06816_, _06815_, _06812_);
  or (_06817_, _06153_, _43427_);
  or (_06818_, _06178_, _00009_);
  and (_06819_, _06818_, _06817_);
  or (_06820_, _06148_, _00204_);
  or (_06821_, _06173_, _00135_);
  and (_06822_, _06821_, _06820_);
  and (_06823_, _06822_, _06819_);
  and (_06824_, _06823_, _06816_);
  or (_06825_, _06166_, _00368_);
  or (_06826_, _06189_, _00327_);
  and (_06827_, _06826_, _06825_);
  or (_06828_, _06158_, _00633_);
  or (_06829_, _06182_, _00491_);
  and (_06830_, _06829_, _06828_);
  and (_06831_, _06830_, _06827_);
  or (_06832_, _06143_, _00286_);
  or (_06833_, _06171_, _00245_);
  and (_06834_, _06833_, _06832_);
  or (_06835_, _06160_, _00091_);
  or (_06836_, _06184_, _00050_);
  and (_06837_, _06836_, _06835_);
  and (_06838_, _06837_, _06834_);
  and (_06839_, _06838_, _06831_);
  and (_06840_, _06839_, _06824_);
  nor (_06841_, _06840_, _06442_);
  not (_06842_, _06420_);
  nor (_06843_, _06840_, _06842_);
  not (_06844_, _06393_);
  or (_06845_, _06840_, _06414_);
  nor (_06846_, _06840_, _06404_);
  and (_06847_, _06288_, _05711_);
  not (_06848_, _06847_);
  and (_06849_, _06298_, _06013_);
  nor (_06850_, _06849_, _06014_);
  and (_06851_, _06850_, _06848_);
  nor (_06852_, _06851_, _06001_);
  not (_06853_, _06852_);
  and (_06854_, _06483_, _06402_);
  not (_06855_, _06854_);
  and (_06856_, _06849_, _06302_);
  nor (_06857_, _06755_, _06856_);
  and (_06858_, _06857_, _06855_);
  not (_06859_, _06858_);
  and (_06860_, _06290_, _05711_);
  not (_06861_, _06860_);
  and (_06862_, _06861_, _06851_);
  nor (_06863_, _06862_, _05996_);
  nor (_06864_, _06863_, _06859_);
  and (_06865_, _06864_, _06853_);
  or (_06866_, _06865_, _06846_);
  nand (_06867_, _06866_, _06396_);
  or (_06868_, _06808_, _06396_);
  nand (_06869_, _06868_, _06867_);
  and (_06870_, _06399_, _06270_);
  nor (_06871_, _06870_, _06406_);
  and (_06872_, _06462_, _06392_);
  and (_06873_, _06483_, _06392_);
  or (_06874_, _06873_, _06872_);
  not (_06875_, _06874_);
  nor (_06876_, _06452_, _06849_);
  nor (_06877_, _06876_, _05999_);
  and (_06878_, _06289_, _06392_);
  and (_06879_, _06878_, _05711_);
  nor (_06880_, _06879_, _06877_);
  and (_06881_, _06880_, _06875_);
  and (_06882_, _06881_, _06871_);
  nand (_06883_, _06882_, _06869_);
  nand (_06884_, _06883_, _06845_);
  and (_06885_, _06884_, _06844_);
  nor (_06886_, _06808_, _06844_);
  or (_06887_, _06886_, _06885_);
  and (_06888_, _06840_, _06419_);
  nor (_06889_, _06862_, _05993_);
  nor (_06890_, _06889_, _06888_);
  and (_06891_, _06890_, _06887_);
  or (_06892_, _06891_, _06843_);
  nand (_06893_, _06892_, _06389_);
  nor (_06894_, _06808_, _06389_);
  nor (_06895_, _06894_, _06384_);
  nand (_06896_, _06895_, _06893_);
  and (_06897_, _06840_, _06384_);
  and (_06898_, _06849_, _06381_);
  nor (_06899_, _06898_, _06435_);
  not (_06900_, _06899_);
  nor (_06901_, _06900_, _06897_);
  and (_06902_, _06901_, _06896_);
  nor (_06903_, _06808_, _06434_);
  nor (_06904_, _06903_, _06902_);
  not (_06905_, _06016_);
  nor (_06906_, _06862_, _06905_);
  nor (_06907_, _06906_, _06904_);
  or (_06908_, _06907_, _06841_);
  and (_06909_, _06908_, _06446_);
  nor (_06910_, _06909_, _06809_);
  nor (_06911_, _06862_, _06287_);
  nor (_06912_, _06911_, _06910_);
  and (_06913_, _06555_, _04737_);
  and (_06914_, _06552_, _04706_);
  nor (_06915_, _06914_, _06913_);
  and (_06916_, _06544_, _04733_);
  and (_06917_, _06516_, _04731_);
  nor (_06918_, _06917_, _06916_);
  and (_06919_, _06918_, _06915_);
  and (_06920_, _06512_, _04721_);
  and (_06921_, _06534_, _04725_);
  nor (_06922_, _06921_, _06920_);
  and (_06923_, _06532_, _04699_);
  and (_06924_, _06557_, _04704_);
  nor (_06925_, _06924_, _06923_);
  and (_06926_, _06925_, _06922_);
  and (_06927_, _06926_, _06919_);
  and (_06928_, _06526_, _04714_);
  and (_06929_, _06550_, _04712_);
  nor (_06930_, _06929_, _06928_);
  and (_06931_, _06539_, _04735_);
  and (_06932_, _06546_, _04729_);
  nor (_06933_, _06932_, _06931_);
  and (_06934_, _06933_, _06930_);
  and (_06935_, _06520_, _04701_);
  and (_06936_, _06508_, _04723_);
  nor (_06937_, _06936_, _06935_);
  and (_06938_, _06541_, _04719_);
  and (_06939_, _06528_, _04710_);
  nor (_06940_, _06939_, _06938_);
  and (_06941_, _06940_, _06937_);
  and (_06942_, _06941_, _06934_);
  and (_06943_, _06942_, _06927_);
  nor (_06944_, _06943_, _06279_);
  or (_06945_, _06944_, _06912_);
  and (_06946_, _06808_, _06376_);
  and (_06947_, _06849_, _05942_);
  nor (_06948_, _06947_, _06375_);
  not (_06949_, _06948_);
  nor (_06950_, _06949_, _06946_);
  and (_06951_, _06950_, _06945_);
  not (_06952_, _06375_);
  nor (_06953_, _06808_, _06952_);
  or (_06954_, _06953_, _06951_);
  and (_06955_, _06288_, _06298_);
  and (_06956_, _06955_, _05951_);
  not (_06957_, _06956_);
  and (_06958_, _06462_, _05951_);
  and (_06959_, _06452_, _05951_);
  nor (_06960_, _06959_, _06958_);
  and (_06961_, _06483_, _05951_);
  and (_06962_, _06849_, _05951_);
  nor (_06963_, _06962_, _06961_);
  and (_06964_, _06963_, _06960_);
  and (_06965_, _06964_, _06957_);
  and (_06966_, _06965_, _06954_);
  not (_06967_, _06840_);
  nor (_06968_, _06967_, _06584_);
  and (_06969_, _06849_, _05955_);
  and (_06970_, _06452_, _05955_);
  nor (_06971_, _06970_, _06969_);
  and (_06972_, _06955_, _05955_);
  and (_06973_, _06462_, _05955_);
  and (_06974_, _06483_, _05955_);
  or (_06975_, _06974_, _06973_);
  nor (_06976_, _06975_, _06972_);
  and (_06977_, _06976_, _06971_);
  not (_06978_, _06977_);
  nor (_06979_, _06978_, _06968_);
  and (_06980_, _06979_, _06966_);
  nor (_06981_, _06967_, _06577_);
  and (_06982_, _06452_, _05965_);
  not (_06983_, _06982_);
  and (_06984_, _06849_, _05965_);
  nor (_06985_, _06984_, _06754_);
  and (_06986_, _06985_, _06983_);
  and (_06987_, _06955_, _05965_);
  not (_06988_, _05965_);
  nor (_06989_, _06483_, _06014_);
  nor (_06990_, _06989_, _06988_);
  nor (_06991_, _06990_, _06987_);
  and (_06992_, _06991_, _06986_);
  not (_06993_, _06992_);
  not (_06994_, _06955_);
  and (_06995_, _06876_, _06994_);
  and (_06996_, _06861_, _06995_);
  not (_06997_, _06996_);
  and (_06998_, _06576_, _05946_);
  and (_06999_, _06998_, _06997_);
  nor (_07000_, _06999_, _06993_);
  not (_07001_, _07000_);
  nor (_07002_, _07001_, _06981_);
  and (_07003_, _07002_, _06980_);
  nor (_07004_, _06840_, _06579_);
  nor (_07005_, _07004_, _07003_);
  and (_07006_, _06588_, _06270_);
  nor (_07007_, _07006_, _07005_);
  and (_07008_, _06808_, _06460_);
  not (_07009_, _05970_);
  nor (_07010_, _06462_, _06014_);
  and (_07011_, _07010_, _06994_);
  or (_07012_, _07011_, _07009_);
  and (_07013_, _06849_, _05970_);
  and (_07014_, _06452_, _05970_);
  nor (_07015_, _07014_, _07013_);
  nand (_07016_, _06763_, _05711_);
  and (_07017_, _07016_, _07015_);
  and (_07018_, _07017_, _07012_);
  not (_07019_, _07018_);
  nor (_07020_, _07019_, _07008_);
  and (_07021_, _07020_, _07007_);
  nor (_07022_, _06840_, _06308_);
  nor (_07023_, _07022_, _07021_);
  and (_07024_, _06305_, _06270_);
  nor (_07025_, _07024_, _07023_);
  and (_07026_, _06808_, _06487_);
  nand (_07027_, _05805_, _05711_);
  not (_07028_, _07027_);
  and (_07029_, _07028_, _05968_);
  not (_07030_, _07029_);
  and (_07031_, _06849_, _05968_);
  nor (_07032_, _07031_, _06606_);
  and (_07033_, _07032_, _07030_);
  not (_07034_, _07033_);
  nor (_07035_, _07034_, _07026_);
  and (_07036_, _07035_, _07025_);
  not (_07037_, _06606_);
  nor (_07038_, _06840_, _07037_);
  or (_07039_, _07038_, _07036_);
  and (_07040_, _07039_, _06807_);
  nor (_07041_, _06808_, _06807_);
  or (_07042_, _07041_, _07040_);
  or (_07043_, _06462_, _06955_);
  and (_07044_, _07043_, _05962_);
  and (_07045_, _06849_, _05962_);
  nor (_07046_, _07045_, _07044_);
  and (_07047_, _06483_, _05962_);
  and (_07048_, _06452_, _05962_);
  nor (_07049_, _07048_, _07047_);
  and (_07050_, _07049_, _07046_);
  nand (_07051_, _07050_, _07042_);
  and (_07052_, _06840_, _06195_);
  or (_07053_, _07052_, _07051_);
  or (_07054_, _07053_, _06806_);
  not (_07055_, _06301_);
  and (_07056_, _06658_, _06266_);
  not (_07057_, _07056_);
  nor (_07058_, _06703_, _06228_);
  not (_07059_, _07058_);
  and (_07060_, _06544_, _04764_);
  and (_07061_, _06555_, _04779_);
  nor (_07062_, _07061_, _07060_);
  and (_07063_, _06520_, _04772_);
  and (_07064_, _06508_, _04752_);
  nor (_07065_, _07064_, _07063_);
  and (_07066_, _07065_, _07062_);
  and (_07067_, _06526_, _04758_);
  and (_07068_, _06552_, _04775_);
  nor (_07069_, _07068_, _07067_);
  and (_07070_, _06550_, _04747_);
  and (_07071_, _06528_, _04786_);
  nor (_07072_, _07071_, _07070_);
  and (_07073_, _07072_, _07069_);
  and (_07074_, _07073_, _07066_);
  and (_07075_, _06532_, _04770_);
  and (_07076_, _06557_, _04761_);
  nor (_07077_, _07076_, _07075_);
  and (_07078_, _06541_, _04745_);
  and (_07079_, _06534_, _04754_);
  nor (_07080_, _07079_, _07078_);
  and (_07081_, _07080_, _07077_);
  and (_07082_, _06539_, _04777_);
  and (_07083_, _06512_, _04749_);
  nor (_07084_, _07083_, _07082_);
  and (_07085_, _06516_, _04766_);
  and (_07086_, _06546_, _04784_);
  nor (_07087_, _07086_, _07085_);
  and (_07088_, _07087_, _07084_);
  and (_07089_, _07088_, _07081_);
  and (_07090_, _07089_, _07074_);
  nor (_07091_, _07090_, _06279_);
  nor (_07092_, _06399_, _06305_);
  nor (_07093_, _07092_, _06268_);
  not (_07094_, _07093_);
  and (_07095_, _06289_, _05946_);
  and (_07096_, _06289_, _05962_);
  nor (_07097_, _07096_, _07095_);
  and (_07098_, _06289_, _06016_);
  nor (_07099_, _07098_, _06878_);
  and (_07100_, _07099_, _07097_);
  and (_07101_, _07100_, _06749_);
  and (_07102_, _07101_, _07094_);
  and (_07103_, _06288_, _05980_);
  and (_07104_, _07103_, _05951_);
  nor (_07105_, _07104_, _06987_);
  and (_07106_, _06784_, _05742_);
  not (_07107_, _06289_);
  nor (_07108_, _05970_, _05935_);
  nor (_07109_, _07108_, _07107_);
  nor (_07110_, _07109_, _07106_);
  and (_07111_, _07110_, _07105_);
  and (_07112_, _06289_, _06386_);
  nor (_07113_, _06791_, _07112_);
  and (_07114_, _06289_, _05955_);
  nor (_07115_, _07114_, _06794_);
  and (_07116_, _07115_, _07113_);
  and (_07117_, _06765_, _06762_);
  and (_07118_, _07117_, _07116_);
  and (_07119_, _07118_, _07111_);
  and (_07120_, _06588_, \uc8051golden_1.SP [1]);
  not (_07121_, _07120_);
  and (_07122_, _06955_, _06402_);
  and (_07123_, _07103_, _06402_);
  nor (_07124_, _07123_, _07122_);
  and (_07125_, _07124_, _07121_);
  nor (_07126_, _06783_, _06750_);
  and (_07127_, _07103_, _05965_);
  not (_07128_, _07127_);
  and (_07129_, _07128_, _07126_);
  nor (_07130_, _06394_, _05968_);
  nor (_07131_, _07130_, _07107_);
  nor (_07132_, _07131_, _06956_);
  and (_07133_, _07132_, _07129_);
  and (_07134_, _07133_, _07125_);
  and (_07135_, _07134_, _07119_);
  and (_07136_, _07135_, _07102_);
  not (_07137_, _07136_);
  nor (_07138_, _07137_, _07091_);
  and (_07139_, _07138_, _07059_);
  and (_07140_, _07139_, _07057_);
  and (_07141_, _07140_, _07055_);
  nand (_07142_, _07053_, \uc8051golden_1.IRAM[0] [1]);
  and (_07143_, _07142_, _07141_);
  nand (_07144_, _07143_, _07054_);
  not (_07145_, \uc8051golden_1.IRAM[2] [1]);
  nor (_07146_, _07052_, _07051_);
  or (_07147_, _07146_, _07145_);
  not (_07148_, _07141_);
  not (_07149_, \uc8051golden_1.IRAM[3] [1]);
  or (_07150_, _07053_, _07149_);
  and (_07151_, _07150_, _07148_);
  nand (_07152_, _07151_, _07147_);
  nand (_07153_, _07152_, _07144_);
  nand (_07154_, _07153_, _06805_);
  not (_07155_, _06805_);
  not (_07156_, \uc8051golden_1.IRAM[6] [1]);
  or (_07157_, _07146_, _07156_);
  not (_07158_, \uc8051golden_1.IRAM[7] [1]);
  or (_07159_, _07053_, _07158_);
  and (_07160_, _07159_, _07148_);
  nand (_07161_, _07160_, _07157_);
  not (_07162_, \uc8051golden_1.IRAM[5] [1]);
  or (_07163_, _07053_, _07162_);
  not (_07164_, \uc8051golden_1.IRAM[4] [1]);
  or (_07165_, _07146_, _07164_);
  and (_07166_, _07165_, _07141_);
  nand (_07167_, _07166_, _07163_);
  nand (_07168_, _07167_, _07161_);
  nand (_07169_, _07168_, _07155_);
  nand (_07170_, _07169_, _07154_);
  nand (_07171_, _07170_, _06618_);
  not (_07172_, _06618_);
  nand (_07173_, _07053_, \uc8051golden_1.IRAM[10] [1]);
  nand (_07174_, _07146_, \uc8051golden_1.IRAM[11] [1]);
  and (_07175_, _07174_, _07148_);
  nand (_07176_, _07175_, _07173_);
  nand (_07177_, _07146_, \uc8051golden_1.IRAM[9] [1]);
  nand (_07178_, _07053_, \uc8051golden_1.IRAM[8] [1]);
  and (_07179_, _07178_, _07141_);
  nand (_07180_, _07179_, _07177_);
  nand (_07181_, _07180_, _07176_);
  nand (_07182_, _07181_, _06805_);
  nand (_07183_, _07053_, \uc8051golden_1.IRAM[14] [1]);
  nand (_07184_, _07146_, \uc8051golden_1.IRAM[15] [1]);
  and (_07185_, _07184_, _07148_);
  nand (_07186_, _07185_, _07183_);
  not (_07187_, \uc8051golden_1.IRAM[13] [1]);
  or (_07188_, _07053_, _07187_);
  nand (_07189_, _07053_, \uc8051golden_1.IRAM[12] [1]);
  and (_07190_, _07189_, _07141_);
  nand (_07191_, _07190_, _07188_);
  nand (_07192_, _07191_, _07186_);
  nand (_07193_, _07192_, _07155_);
  nand (_07194_, _07193_, _07182_);
  nand (_07195_, _07194_, _07172_);
  nand (_07196_, _07195_, _07171_);
  and (_07197_, _07196_, _06304_);
  or (_07198_, _07197_, _06303_);
  and (_07199_, _06451_, _06402_);
  not (_07200_, _07199_);
  nor (_07201_, _07200_, _06194_);
  and (_07202_, _07201_, _06228_);
  nor (_07203_, _07202_, _07198_);
  and (_07204_, _06790_, _06272_);
  not (_07205_, _07204_);
  and (_07206_, _06285_, _06394_);
  nor (_07207_, _07206_, _06787_);
  and (_07208_, _07207_, _07205_);
  and (_07209_, _07208_, _07203_);
  not (_07210_, _06401_);
  nor (_07211_, _07210_, _06194_);
  and (_07212_, _06280_, _06394_);
  and (_07213_, _07212_, _07196_);
  nor (_07214_, _07213_, _07211_);
  and (_07215_, _07214_, _07209_);
  and (_07216_, _07211_, _06229_);
  nor (_07217_, _07216_, _07215_);
  nor (_07218_, _06396_, _06194_);
  and (_07219_, _07218_, _06265_);
  nor (_07220_, _07219_, _07217_);
  not (_07221_, _06399_);
  nor (_07222_, _07221_, _06194_);
  nor (_07223_, _06273_, _05997_);
  nor (_07224_, _07223_, _07222_);
  and (_07225_, _07224_, _07220_);
  and (_07226_, _07222_, _06229_);
  nor (_07227_, _07226_, _07225_);
  and (_07228_, _06285_, _06392_);
  nor (_07229_, _07228_, _06773_);
  not (_07230_, _07229_);
  nor (_07231_, _07230_, _07227_);
  nor (_07232_, _06414_, _06194_);
  and (_07233_, _06280_, _06392_);
  and (_07234_, _07233_, _07196_);
  nor (_07235_, _07234_, _07232_);
  and (_07236_, _07235_, _07231_);
  and (_07237_, _07232_, _06229_);
  nor (_07238_, _07237_, _07236_);
  nor (_07239_, _06844_, _06194_);
  and (_07240_, _07239_, _06265_);
  or (_07241_, _07240_, _06419_);
  nor (_07242_, _07241_, _07238_);
  and (_07243_, _06419_, _06273_);
  nor (_07244_, _07243_, _07242_);
  not (_07245_, _06387_);
  nor (_07246_, _07245_, _06194_);
  and (_07247_, _07246_, _06265_);
  nor (_07248_, _07247_, _07244_);
  nor (_07249_, _06273_, _05994_);
  not (_07250_, _07249_);
  and (_07251_, _06285_, _06381_);
  and (_07252_, _06751_, _06381_);
  nor (_07253_, _07252_, _07251_);
  and (_07254_, _07253_, _07250_);
  and (_07255_, _07254_, _07248_);
  nor (_07256_, _06446_, _06194_);
  and (_07257_, _06280_, _06381_);
  and (_07258_, _07257_, _07196_);
  nor (_07259_, _07258_, _07256_);
  and (_07260_, _07259_, _07255_);
  nor (_07261_, _07260_, _06301_);
  nor (_07262_, _07261_, _06017_);
  and (_07263_, _06273_, _06017_);
  nor (_07264_, _07263_, _07262_);
  and (_07265_, _06284_, _05942_);
  or (_07266_, _07265_, _07264_);
  nor (_07267_, _07266_, _06297_);
  and (_07268_, _06280_, _05942_);
  and (_07269_, _07268_, _07196_);
  nor (_07270_, _07269_, _06277_);
  and (_07271_, _07270_, _07267_);
  nor (_07272_, _07271_, _06278_);
  nor (_07273_, _07272_, _05943_);
  and (_07274_, _06273_, _05943_);
  nor (_07275_, _07274_, _07273_);
  not (_07276_, _06569_);
  nor (_07277_, _07276_, _06194_);
  not (_07278_, _07277_);
  not (_07279_, _06478_);
  nor (_07280_, _07279_, _06194_);
  not (_07281_, _07280_);
  not (_07282_, _06474_);
  nor (_07283_, _07282_, _06194_);
  not (_07284_, _06582_);
  nor (_07285_, _07284_, _06194_);
  nor (_07286_, _07285_, _07283_);
  and (_07287_, _07286_, _07281_);
  and (_07288_, _07287_, _07278_);
  nor (_07289_, _07288_, _06229_);
  nor (_07290_, _07289_, _05956_);
  not (_07291_, _07290_);
  nor (_07292_, _07291_, _07275_);
  and (_07293_, _06273_, _05956_);
  nor (_07294_, _07293_, _07292_);
  nor (_07295_, _06573_, _06194_);
  and (_07296_, _07295_, _06228_);
  or (_07297_, _07296_, _05966_);
  nor (_07298_, _07297_, _07294_);
  nor (_07299_, _07298_, _06274_);
  and (_07300_, _06285_, _05968_);
  nor (_07301_, _07300_, _06772_);
  not (_07302_, _07301_);
  nor (_07303_, _07302_, _07299_);
  nor (_07304_, _07037_, _06194_);
  and (_07305_, _06280_, _05968_);
  and (_07306_, _07305_, _07196_);
  nor (_07307_, _07306_, _07304_);
  and (_07308_, _07307_, _07303_);
  and (_07309_, _07304_, _06229_);
  nor (_07310_, _07309_, _07308_);
  nor (_07311_, _06807_, _06194_);
  nor (_07312_, _06465_, _05969_);
  nor (_07313_, _07312_, _06273_);
  nor (_07314_, _07313_, _07311_);
  not (_07315_, _07314_);
  nor (_07316_, _07315_, _07310_);
  nor (_07317_, _07316_, _06267_);
  and (_07318_, _06284_, _05962_);
  nor (_07319_, _07318_, _07317_);
  and (_07320_, _06280_, _05962_);
  and (_07321_, _07320_, _07196_);
  nor (_07322_, _07321_, _06197_);
  and (_07323_, _07322_, _07319_);
  nor (_07324_, _07323_, _06230_);
  not (_07325_, _01382_);
  nor (_07326_, _06285_, _06280_);
  nor (_07327_, _07326_, _06004_);
  not (_07328_, _06014_);
  nor (_07329_, _06481_, _05808_);
  and (_07330_, _07329_, _07328_);
  nor (_07331_, _07330_, _06004_);
  or (_07332_, _07331_, _07327_);
  not (_07333_, _07332_);
  and (_07334_, _06290_, _05942_);
  nor (_07335_, _07334_, _07300_);
  and (_07336_, _06288_, _05942_);
  not (_07337_, _07336_);
  nor (_07338_, _07337_, _06232_);
  nor (_07339_, _07338_, _07206_);
  and (_07340_, _07339_, _07335_);
  not (_07341_, _07131_);
  and (_07342_, _07341_, _07126_);
  and (_07343_, _06013_, _05980_);
  and (_07344_, _07343_, _05962_);
  nor (_07345_, _07344_, _07251_);
  and (_07346_, _07345_, _07342_);
  and (_07347_, _07346_, _07340_);
  and (_07348_, _07347_, _07333_);
  not (_07349_, _05994_);
  nor (_07350_, _06017_, _07349_);
  not (_07351_, _05997_);
  nor (_07352_, _07351_, _05943_);
  and (_07353_, _07352_, _07350_);
  and (_07354_, _06466_, _06392_);
  nor (_07355_, _06379_, _05996_);
  nor (_07356_, _07355_, _07354_);
  and (_07357_, _06452_, _05942_);
  and (_07358_, _06289_, _06381_);
  nor (_07359_, _07358_, _07357_);
  and (_07360_, _07359_, _07356_);
  and (_07361_, _07360_, _07353_);
  and (_07362_, _06466_, _05962_);
  not (_07363_, _05962_);
  nor (_07364_, _06463_, _07363_);
  nor (_07365_, _07364_, _07362_);
  not (_07366_, _06790_);
  and (_07367_, _07312_, _07366_);
  and (_07368_, _07367_, _07365_);
  and (_07369_, _07368_, _07361_);
  nor (_07370_, _07305_, _07268_);
  nor (_07371_, _07257_, _06419_);
  and (_07372_, _07371_, _07370_);
  nor (_07373_, _05956_, _05966_);
  and (_07374_, _06774_, _07373_);
  and (_07375_, _07374_, _07372_);
  nor (_07376_, _07212_, _07045_);
  and (_07377_, _06452_, _06392_);
  or (_07378_, _06742_, _06453_);
  and (_07379_, _07378_, _05962_);
  nor (_07380_, _07379_, _07377_);
  and (_07381_, _07380_, _07376_);
  nor (_07382_, _07233_, _06380_);
  nor (_07383_, _07048_, _06878_);
  and (_07384_, _07383_, _07382_);
  and (_07385_, _07384_, _07381_);
  and (_07386_, _07385_, _07375_);
  and (_07387_, _07386_, _07369_);
  and (_07388_, _07387_, _07348_);
  and (_07389_, _07388_, _07278_);
  nor (_07390_, _07239_, _06277_);
  nor (_07391_, _07232_, _07218_);
  and (_07392_, _07391_, _07390_);
  and (_07393_, _07392_, _07389_);
  nor (_07394_, _07311_, _06197_);
  nor (_07395_, _06463_, _06287_);
  not (_07396_, _07395_);
  nor (_07397_, _06401_, _06399_);
  nor (_07398_, _06281_, _06387_);
  and (_07399_, _07398_, _07397_);
  and (_07400_, _07399_, _07396_);
  nor (_07401_, _07400_, _06194_);
  and (_07402_, _07378_, _05935_);
  not (_07403_, _07402_);
  nor (_07404_, _06286_, _06015_);
  and (_07405_, _07404_, _07403_);
  nor (_07406_, _07405_, _06194_);
  nor (_07407_, _07406_, _07401_);
  and (_07408_, _07407_, _07394_);
  nor (_07409_, _07201_, _07256_);
  nor (_07410_, _07304_, _07295_);
  and (_07411_, _07410_, _07409_);
  and (_07412_, _07411_, _07408_);
  and (_07413_, _07412_, _07287_);
  and (_07414_, _07413_, _07393_);
  nor (_07415_, _07414_, _07325_);
  not (_07416_, _07415_);
  nor (_07417_, _07416_, _07324_);
  not (_07418_, _07311_);
  and (_07419_, _05966_, _06270_);
  and (_07420_, _06967_, _06277_);
  nor (_07421_, _05994_, _06270_);
  nor (_07422_, _06808_, _07245_);
  not (_07423_, _07246_);
  not (_07424_, \uc8051golden_1.IRAM[1] [0]);
  or (_07425_, _07053_, _07424_);
  nand (_07426_, _07053_, \uc8051golden_1.IRAM[0] [0]);
  and (_07427_, _07426_, _07141_);
  nand (_07428_, _07427_, _07425_);
  not (_07429_, \uc8051golden_1.IRAM[2] [0]);
  or (_07430_, _07146_, _07429_);
  nand (_07431_, _07146_, \uc8051golden_1.IRAM[3] [0]);
  and (_07432_, _07431_, _07148_);
  nand (_07433_, _07432_, _07430_);
  nand (_07434_, _07433_, _07428_);
  nand (_07435_, _07434_, _06805_);
  nand (_07436_, _07053_, \uc8051golden_1.IRAM[6] [0]);
  nand (_07437_, _07146_, \uc8051golden_1.IRAM[7] [0]);
  and (_07438_, _07437_, _07148_);
  nand (_07439_, _07438_, _07436_);
  nand (_07440_, _07146_, \uc8051golden_1.IRAM[5] [0]);
  not (_07441_, \uc8051golden_1.IRAM[4] [0]);
  or (_07442_, _07146_, _07441_);
  and (_07443_, _07442_, _07141_);
  nand (_07444_, _07443_, _07440_);
  nand (_07445_, _07444_, _07439_);
  nand (_07446_, _07445_, _07155_);
  nand (_07447_, _07446_, _07435_);
  nand (_07448_, _07447_, _06618_);
  nand (_07449_, _07053_, \uc8051golden_1.IRAM[10] [0]);
  nand (_07450_, _07146_, \uc8051golden_1.IRAM[11] [0]);
  and (_07451_, _07450_, _07148_);
  nand (_07452_, _07451_, _07449_);
  nand (_07453_, _07146_, \uc8051golden_1.IRAM[9] [0]);
  nand (_07454_, _07053_, \uc8051golden_1.IRAM[8] [0]);
  and (_07455_, _07454_, _07141_);
  nand (_07456_, _07455_, _07453_);
  nand (_07457_, _07456_, _07452_);
  nand (_07458_, _07457_, _06805_);
  nand (_07459_, _07053_, \uc8051golden_1.IRAM[14] [0]);
  not (_07460_, \uc8051golden_1.IRAM[15] [0]);
  or (_07461_, _07053_, _07460_);
  and (_07462_, _07461_, _07148_);
  nand (_07463_, _07462_, _07459_);
  not (_07464_, \uc8051golden_1.IRAM[13] [0]);
  or (_07465_, _07053_, _07464_);
  nand (_07466_, _07053_, \uc8051golden_1.IRAM[12] [0]);
  and (_07467_, _07466_, _07141_);
  nand (_07468_, _07467_, _07465_);
  nand (_07469_, _07468_, _07463_);
  nand (_07470_, _07469_, _07155_);
  nand (_07471_, _07470_, _07458_);
  nand (_07472_, _07471_, _07172_);
  and (_07473_, _07472_, _07448_);
  and (_07474_, _07473_, _06304_);
  and (_07475_, _07329_, _06876_);
  nor (_07476_, _07475_, _06004_);
  not (_07477_, _07476_);
  nor (_07478_, _07477_, _07474_);
  and (_07479_, _07201_, _06840_);
  nor (_07480_, _07479_, _07478_);
  and (_07481_, _06790_, \uc8051golden_1.SP [0]);
  nor (_07482_, _07027_, _05996_);
  nor (_07483_, _07482_, _07481_);
  and (_07484_, _07483_, _07480_);
  nand (_07485_, _07472_, _07448_);
  and (_07486_, _07485_, _07212_);
  not (_07487_, _07486_);
  and (_07488_, _07487_, _07484_);
  and (_07489_, _07211_, _06840_);
  nor (_07490_, _07489_, _07218_);
  and (_07491_, _07490_, _07488_);
  not (_07492_, _07491_);
  and (_07493_, _07492_, _06868_);
  nor (_07494_, _05997_, _06270_);
  nor (_07495_, _07494_, _07493_);
  and (_07496_, _07222_, _06840_);
  nor (_07497_, _07377_, _06879_);
  and (_07498_, _07497_, _06875_);
  not (_07499_, _07498_);
  nor (_07500_, _07499_, _07496_);
  and (_07501_, _07500_, _07495_);
  and (_07502_, _07485_, _07233_);
  not (_07503_, _07502_);
  and (_07504_, _07503_, _07501_);
  and (_07505_, _07232_, _06840_);
  nor (_07506_, _07505_, _07239_);
  and (_07507_, _07506_, _07504_);
  nor (_07508_, _07507_, _06886_);
  or (_07509_, _07508_, _06419_);
  nand (_07510_, _06419_, _06270_);
  nand (_07511_, _07510_, _07509_);
  and (_07512_, _07511_, _07423_);
  nor (_07513_, _07512_, _07422_);
  and (_07514_, _06847_, _06381_);
  and (_07515_, _06380_, _05711_);
  or (_07516_, _07515_, _07514_);
  or (_07517_, _07516_, _07513_);
  nor (_07518_, _07517_, _07421_);
  and (_07519_, _07485_, _07257_);
  nor (_07520_, _07519_, _07256_);
  and (_07521_, _07520_, _07518_);
  nor (_07522_, _07521_, _06809_);
  nor (_07523_, _07522_, _06017_);
  and (_07524_, _06017_, _06270_);
  nor (_07525_, _07524_, _07523_);
  nor (_07526_, _06296_, _06967_);
  and (_07527_, _07028_, _05942_);
  nor (_07528_, _07527_, _07526_);
  not (_07529_, _07528_);
  nor (_07530_, _07529_, _07525_);
  and (_07531_, _07485_, _07268_);
  nor (_07532_, _07531_, _06277_);
  and (_07533_, _07532_, _07530_);
  nor (_07534_, _07533_, _07420_);
  nor (_07535_, _07534_, _05943_);
  and (_07536_, _05943_, _06270_);
  nor (_07537_, _07536_, _07535_);
  nor (_07538_, _07288_, _06967_);
  nor (_07539_, _07538_, _05956_);
  not (_07540_, _07539_);
  nor (_07541_, _07540_, _07537_);
  and (_07542_, _05956_, _06270_);
  nor (_07543_, _07542_, _07541_);
  and (_07544_, _07295_, _06840_);
  or (_07545_, _07544_, _05966_);
  nor (_07546_, _07545_, _07543_);
  nor (_07547_, _07546_, _07419_);
  nor (_07548_, _07547_, _07029_);
  and (_07549_, _07485_, _07305_);
  nor (_07550_, _07549_, _07304_);
  and (_07551_, _07550_, _07548_);
  and (_07552_, _07304_, _06967_);
  nor (_07553_, _07552_, _07551_);
  nor (_07554_, _07312_, _06270_);
  nor (_07555_, _07554_, _07553_);
  and (_07556_, _07555_, _07418_);
  nor (_07557_, _07556_, _07041_);
  and (_07558_, _07028_, _05962_);
  nor (_07559_, _07558_, _07557_);
  and (_07560_, _07485_, _07320_);
  nor (_07561_, _07560_, _06197_);
  and (_07562_, _07561_, _07559_);
  and (_07563_, _06967_, _06197_);
  nor (_07564_, _07563_, _07562_);
  nor (_07565_, _07564_, _07416_);
  and (_07566_, _07565_, _07417_);
  and (_07567_, _06651_, _06234_);
  and (_07568_, \uc8051golden_1.SP [1], \uc8051golden_1.SP [0]);
  and (_07569_, _07568_, \uc8051golden_1.SP [2]);
  nor (_07570_, _07568_, \uc8051golden_1.SP [2]);
  nor (_07571_, _07570_, _07569_);
  and (_07572_, _07571_, _05966_);
  not (_07573_, _06693_);
  and (_07574_, _07573_, _06277_);
  nand (_07575_, _07146_, \uc8051golden_1.IRAM[1] [2]);
  nand (_07576_, _07053_, \uc8051golden_1.IRAM[0] [2]);
  and (_07577_, _07576_, _07141_);
  nand (_07578_, _07577_, _07575_);
  nand (_07579_, _07053_, \uc8051golden_1.IRAM[2] [2]);
  not (_07580_, \uc8051golden_1.IRAM[3] [2]);
  or (_07581_, _07053_, _07580_);
  and (_07582_, _07581_, _07148_);
  nand (_07583_, _07582_, _07579_);
  nand (_07584_, _07583_, _07578_);
  nand (_07585_, _07584_, _06805_);
  nand (_07586_, _07053_, \uc8051golden_1.IRAM[6] [2]);
  nand (_07587_, _07146_, \uc8051golden_1.IRAM[7] [2]);
  and (_07588_, _07587_, _07148_);
  nand (_07589_, _07588_, _07586_);
  nand (_07590_, _07146_, \uc8051golden_1.IRAM[5] [2]);
  not (_07591_, \uc8051golden_1.IRAM[4] [2]);
  or (_07592_, _07146_, _07591_);
  and (_07593_, _07592_, _07141_);
  nand (_07594_, _07593_, _07590_);
  nand (_07595_, _07594_, _07589_);
  nand (_07596_, _07595_, _07155_);
  nand (_07597_, _07596_, _07585_);
  nand (_07598_, _07597_, _06618_);
  nand (_07599_, _07053_, \uc8051golden_1.IRAM[10] [2]);
  nand (_07600_, _07146_, \uc8051golden_1.IRAM[11] [2]);
  and (_07601_, _07600_, _07148_);
  nand (_07602_, _07601_, _07599_);
  nand (_07603_, _07146_, \uc8051golden_1.IRAM[9] [2]);
  nand (_07604_, _07053_, \uc8051golden_1.IRAM[8] [2]);
  and (_07605_, _07604_, _07141_);
  nand (_07606_, _07605_, _07603_);
  nand (_07607_, _07606_, _07602_);
  nand (_07608_, _07607_, _06805_);
  not (_07609_, \uc8051golden_1.IRAM[14] [2]);
  or (_07610_, _07146_, _07609_);
  not (_07611_, \uc8051golden_1.IRAM[15] [2]);
  or (_07612_, _07053_, _07611_);
  and (_07613_, _07612_, _07148_);
  nand (_07614_, _07613_, _07610_);
  nand (_07615_, _07146_, \uc8051golden_1.IRAM[13] [2]);
  nand (_07616_, _07053_, \uc8051golden_1.IRAM[12] [2]);
  and (_07617_, _07616_, _07141_);
  nand (_07618_, _07617_, _07615_);
  nand (_07619_, _07618_, _07614_);
  nand (_07620_, _07619_, _07155_);
  nand (_07621_, _07620_, _07608_);
  nand (_07622_, _07621_, _07172_);
  nand (_07623_, _07622_, _07598_);
  or (_07624_, _07623_, _05807_);
  and (_07625_, _07624_, _07331_);
  and (_07626_, _07201_, _06693_);
  nor (_07627_, _07626_, _07625_);
  not (_07628_, _07571_);
  and (_07629_, _07628_, _06790_);
  not (_07630_, _07629_);
  and (_07631_, _07103_, _06394_);
  or (_07632_, _06285_, _06955_);
  and (_07633_, _07632_, _06394_);
  nor (_07634_, _07633_, _07631_);
  and (_07635_, _07634_, _07630_);
  and (_07636_, _07635_, _07627_);
  and (_07637_, _07623_, _07212_);
  nor (_07638_, _07637_, _07211_);
  and (_07639_, _07638_, _07636_);
  and (_07640_, _07211_, _07573_);
  nor (_07641_, _07640_, _07639_);
  and (_07642_, _07218_, _06650_);
  nor (_07643_, _07642_, _07641_);
  or (_07644_, _07571_, _05997_);
  nand (_07645_, _07644_, _07643_);
  and (_07646_, _07222_, _06693_);
  and (_07647_, _06288_, _06392_);
  nor (_07648_, _07647_, _07646_);
  not (_07649_, _07648_);
  nor (_07650_, _07649_, _07645_);
  and (_07651_, _07623_, _07233_);
  nor (_07652_, _07651_, _07232_);
  and (_07653_, _07652_, _07650_);
  and (_07654_, _07232_, _07573_);
  nor (_07655_, _07654_, _07653_);
  and (_07656_, _07239_, _06650_);
  or (_07657_, _07656_, _06419_);
  nor (_07658_, _07657_, _07655_);
  and (_07659_, _07571_, _06419_);
  nor (_07660_, _07659_, _07658_);
  and (_07661_, _06650_, _05994_);
  and (_07662_, _07661_, _07246_);
  nor (_07663_, _07571_, _05994_);
  or (_07664_, _07663_, _06382_);
  or (_07665_, _07664_, _07662_);
  nor (_07666_, _07665_, _07660_);
  and (_07667_, _07623_, _07257_);
  nor (_07668_, _07667_, _07256_);
  and (_07669_, _07668_, _07666_);
  nor (_07670_, _07669_, _06661_);
  nor (_07671_, _07670_, _06017_);
  and (_07672_, _07571_, _06017_);
  nor (_07673_, _07672_, _07671_);
  nor (_07674_, _06296_, _07573_);
  or (_07675_, _07674_, _07336_);
  nor (_07676_, _07675_, _07673_);
  and (_07677_, _07623_, _07268_);
  nor (_07678_, _07677_, _06277_);
  and (_07679_, _07678_, _07676_);
  nor (_07680_, _07679_, _07574_);
  nor (_07681_, _07680_, _05943_);
  and (_07682_, _07571_, _05943_);
  nor (_07683_, _07682_, _07681_);
  nor (_07684_, _07288_, _07573_);
  nor (_07685_, _07684_, _05956_);
  not (_07686_, _07685_);
  nor (_07687_, _07686_, _07683_);
  and (_07688_, _07571_, _05956_);
  nor (_07689_, _07688_, _07687_);
  and (_07690_, _07295_, _06693_);
  or (_07691_, _07690_, _05966_);
  nor (_07692_, _07691_, _07689_);
  nor (_07693_, _07692_, _07572_);
  and (_07694_, _06288_, _05968_);
  nor (_07695_, _07694_, _07693_);
  and (_07696_, _07623_, _07305_);
  nor (_07697_, _07696_, _07304_);
  and (_07698_, _07697_, _07695_);
  and (_07699_, _07304_, _07573_);
  nor (_07700_, _07699_, _07698_);
  nor (_07701_, _07571_, _07312_);
  nor (_07702_, _07701_, _07311_);
  not (_07703_, _07702_);
  nor (_07704_, _07703_, _07700_);
  nor (_07705_, _07704_, _07567_);
  and (_07706_, _06288_, _05962_);
  nor (_07707_, _07706_, _07705_);
  and (_07708_, _07623_, _07320_);
  nor (_07709_, _07708_, _06197_);
  and (_07710_, _07709_, _07707_);
  and (_07711_, _07573_, _06197_);
  nor (_07712_, _07711_, _07710_);
  nor (_07713_, _07712_, _07416_);
  not (_07714_, _07713_);
  nand (_07715_, _07146_, \uc8051golden_1.IRAM[1] [3]);
  nand (_07716_, _07053_, \uc8051golden_1.IRAM[0] [3]);
  and (_07717_, _07716_, _07141_);
  nand (_07718_, _07717_, _07715_);
  nand (_07719_, _07053_, \uc8051golden_1.IRAM[2] [3]);
  nand (_07720_, _07146_, \uc8051golden_1.IRAM[3] [3]);
  and (_07721_, _07720_, _07148_);
  nand (_07722_, _07721_, _07719_);
  nand (_07723_, _07722_, _07718_);
  nand (_07724_, _07723_, _06805_);
  nand (_07725_, _07053_, \uc8051golden_1.IRAM[6] [3]);
  nand (_07726_, _07146_, \uc8051golden_1.IRAM[7] [3]);
  and (_07727_, _07726_, _07148_);
  nand (_07728_, _07727_, _07725_);
  nand (_07730_, _07146_, \uc8051golden_1.IRAM[5] [3]);
  nand (_07731_, _07053_, \uc8051golden_1.IRAM[4] [3]);
  and (_07733_, _07731_, _07141_);
  nand (_07734_, _07733_, _07730_);
  nand (_07736_, _07734_, _07728_);
  nand (_07737_, _07736_, _07155_);
  nand (_07739_, _07737_, _07724_);
  nand (_07740_, _07739_, _06618_);
  nand (_07742_, _07053_, \uc8051golden_1.IRAM[10] [3]);
  nand (_07743_, _07146_, \uc8051golden_1.IRAM[11] [3]);
  and (_07745_, _07743_, _07148_);
  nand (_07746_, _07745_, _07742_);
  nand (_07748_, _07146_, \uc8051golden_1.IRAM[9] [3]);
  nand (_07749_, _07053_, \uc8051golden_1.IRAM[8] [3]);
  and (_07751_, _07749_, _07141_);
  nand (_07752_, _07751_, _07748_);
  nand (_07754_, _07752_, _07746_);
  nand (_07755_, _07754_, _06805_);
  not (_07757_, \uc8051golden_1.IRAM[14] [3]);
  or (_07758_, _07146_, _07757_);
  not (_07760_, \uc8051golden_1.IRAM[15] [3]);
  or (_07761_, _07053_, _07760_);
  and (_07763_, _07761_, _07148_);
  nand (_07764_, _07763_, _07758_);
  nand (_07766_, _07146_, \uc8051golden_1.IRAM[13] [3]);
  not (_07767_, \uc8051golden_1.IRAM[12] [3]);
  or (_07768_, _07146_, _07767_);
  and (_07769_, _07768_, _07141_);
  nand (_07770_, _07769_, _07766_);
  nand (_07771_, _07770_, _07764_);
  nand (_07772_, _07771_, _07155_);
  nand (_07773_, _07772_, _07755_);
  nand (_07774_, _07773_, _07172_);
  nand (_07775_, _07774_, _07740_);
  and (_07776_, _07775_, _07305_);
  not (_07777_, _07256_);
  nor (_07778_, _06341_, _07777_);
  nor (_07779_, _07569_, \uc8051golden_1.SP [3]);
  and (_07780_, \uc8051golden_1.SP [2], \uc8051golden_1.SP [1]);
  and (_07781_, _07780_, \uc8051golden_1.SP [3]);
  and (_07782_, _07781_, \uc8051golden_1.SP [0]);
  nor (_07783_, _07782_, _07779_);
  and (_07784_, _07783_, _07349_);
  not (_07785_, _06419_);
  and (_07786_, _07775_, _07212_);
  and (_07787_, _07783_, _06790_);
  and (_07788_, _07775_, _06304_);
  not (_07789_, \uc8051golden_1.PSW [3]);
  and (_07790_, _06005_, _07789_);
  nor (_07791_, _07790_, _07788_);
  nor (_07792_, _07791_, _07201_);
  and (_07793_, _07201_, _06372_);
  nor (_07794_, _07793_, _06790_);
  not (_07795_, _07794_);
  nor (_07796_, _07795_, _07792_);
  or (_07797_, _07796_, _07212_);
  nor (_07798_, _07797_, _07787_);
  or (_07799_, _07798_, _07211_);
  nor (_07800_, _07799_, _07786_);
  and (_07801_, _07211_, _06589_);
  or (_07802_, _07801_, _07218_);
  nor (_07803_, _07802_, _07800_);
  and (_07804_, _06395_, _06341_);
  nor (_07805_, _07804_, _07803_);
  nor (_07806_, _07805_, _07351_);
  nor (_07807_, _07783_, _05997_);
  nor (_07808_, _07807_, _07222_);
  not (_07809_, _07808_);
  nor (_07810_, _07809_, _07806_);
  and (_07811_, _07222_, _06589_);
  nor (_07812_, _07811_, _07233_);
  not (_07813_, _07812_);
  nor (_07814_, _07813_, _07810_);
  and (_07815_, _07775_, _07233_);
  nor (_07816_, _07815_, _07232_);
  not (_07817_, _07816_);
  nor (_07818_, _07817_, _07814_);
  and (_07819_, _07232_, _06589_);
  or (_07820_, _07819_, _07239_);
  nor (_07821_, _07820_, _07818_);
  and (_07822_, _07239_, _06340_);
  nor (_07823_, _07822_, _07821_);
  and (_07825_, _07823_, _07785_);
  and (_07827_, _07783_, _06419_);
  nor (_07828_, _07827_, _07825_);
  nor (_07830_, _07828_, _07246_);
  and (_07831_, _07246_, _06374_);
  or (_07833_, _07831_, _07830_);
  and (_07834_, _07833_, _05994_);
  or (_07836_, _07834_, _07257_);
  nor (_07837_, _07836_, _07784_);
  and (_07839_, _07775_, _07257_);
  or (_07840_, _07839_, _07256_);
  nor (_07842_, _07840_, _07837_);
  or (_07843_, _07842_, _07778_);
  or (_07845_, _07843_, _06017_);
  not (_07846_, _06017_);
  or (_07848_, _07783_, _07846_);
  and (_07849_, _07848_, _06296_);
  and (_07851_, _07849_, _07845_);
  nor (_07852_, _06296_, _06372_);
  nor (_07854_, _07852_, _07268_);
  not (_07855_, _07854_);
  nor (_07857_, _07855_, _07851_);
  and (_07858_, _07775_, _07268_);
  nor (_07860_, _07858_, _06277_);
  not (_07861_, _07860_);
  nor (_07862_, _07861_, _07857_);
  nor (_07863_, _06808_, _06276_);
  nor (_07864_, _07863_, _07862_);
  nor (_07865_, _07864_, _05943_);
  and (_07866_, _07783_, _05943_);
  not (_07867_, _07866_);
  and (_07868_, _07867_, _07288_);
  not (_07869_, _07868_);
  nor (_07870_, _07869_, _07865_);
  nor (_07871_, _07288_, _06589_);
  nor (_07872_, _07871_, _05956_);
  not (_07873_, _07872_);
  nor (_07874_, _07873_, _07870_);
  and (_07875_, _07783_, _05956_);
  or (_07876_, _07875_, _07295_);
  nor (_07877_, _07876_, _07874_);
  and (_07878_, _07295_, _06372_);
  or (_07879_, _07878_, _05966_);
  nor (_07880_, _07879_, _07877_);
  and (_07881_, _07783_, _05966_);
  nor (_07882_, _07881_, _07305_);
  not (_07883_, _07882_);
  nor (_07884_, _07883_, _07880_);
  or (_07885_, _07884_, _07304_);
  nor (_07886_, _07885_, _07776_);
  not (_07887_, _07312_);
  and (_07888_, _07304_, _06589_);
  nor (_07889_, _07888_, _07887_);
  not (_07890_, _07889_);
  nor (_07891_, _07890_, _07886_);
  nor (_07892_, _07783_, _07312_);
  nor (_07893_, _07892_, _07311_);
  not (_07894_, _07893_);
  nor (_07895_, _07894_, _07891_);
  not (_07896_, _06340_);
  and (_07897_, _07311_, _07896_);
  nor (_07898_, _07897_, _07320_);
  not (_07899_, _07898_);
  nor (_07900_, _07899_, _07895_);
  and (_07901_, _07775_, _07320_);
  nor (_07902_, _07901_, _06197_);
  not (_07903_, _07902_);
  nor (_07904_, _07903_, _07900_);
  and (_07905_, _06589_, _06197_);
  nor (_07906_, _07905_, _07904_);
  nor (_07907_, _07906_, _07714_);
  nand (_07908_, _07907_, _07566_);
  nand (_07909_, _07908_, _05652_);
  and (_07910_, _07780_, _06270_);
  nor (_07911_, _07571_, _06271_);
  nor (_07912_, _07911_, _07910_);
  and (_07913_, _07781_, _06270_);
  nor (_07914_, _07910_, _07783_);
  nor (_07915_, _07914_, _07913_);
  and (_07916_, _07353_, _07373_);
  and (_07917_, _07916_, _07367_);
  nor (_07918_, _07917_, _07325_);
  and (_07919_, _07918_, _07915_);
  and (_07920_, _07919_, _07912_);
  and (_07921_, _07920_, _06269_);
  not (_07922_, _07921_);
  and (_07923_, _07922_, _07909_);
  and (_07924_, _06840_, _06228_);
  and (_07925_, _06693_, _06372_);
  and (_07926_, _07925_, _07924_);
  and (_07927_, _06340_, _06194_);
  not (_07928_, _06650_);
  and (_07929_, _07928_, _06265_);
  and (_07930_, _07929_, _07927_);
  and (_07931_, _07930_, _07926_);
  and (_07932_, _07931_, \uc8051golden_1.P2 [7]);
  not (_07933_, _07932_);
  not (_07934_, _06265_);
  and (_07935_, _06650_, _07934_);
  and (_07936_, _07935_, _07927_);
  and (_07937_, _06693_, _06589_);
  and (_07938_, _06967_, _06228_);
  and (_07939_, _07938_, _07937_);
  and (_07940_, _07939_, _07936_);
  and (_07941_, _07940_, \uc8051golden_1.SBUF [7]);
  not (_07942_, _07941_);
  nor (_07943_, _06650_, _06265_);
  and (_07944_, _07943_, _07927_);
  and (_07945_, _07926_, _07944_);
  and (_07946_, _07945_, \uc8051golden_1.P3 [7]);
  and (_07947_, _07937_, _07924_);
  and (_07948_, _07930_, _07947_);
  and (_07949_, _07948_, \uc8051golden_1.IE [7]);
  nor (_07950_, _07949_, _07946_);
  and (_07951_, _07950_, _07942_);
  and (_07952_, _07951_, _07933_);
  and (_07953_, _06650_, _06265_);
  and (_07954_, _07953_, _07927_);
  and (_07955_, _07938_, _07925_);
  and (_07956_, _07955_, _07954_);
  and (_07957_, _07956_, \uc8051golden_1.SP [7]);
  not (_07958_, _07957_);
  and (_07959_, _07954_, _06372_);
  nor (_07960_, _06967_, _06228_);
  and (_07961_, _07960_, _06693_);
  and (_07962_, _07961_, _07959_);
  and (_07963_, _07962_, \uc8051golden_1.DPL [7]);
  nor (_07964_, _06840_, _06228_);
  and (_07965_, _07964_, _07925_);
  and (_07966_, _07965_, _07954_);
  and (_07967_, _07966_, \uc8051golden_1.DPH [7]);
  nor (_07968_, _07967_, _07963_);
  and (_07969_, _07968_, _07958_);
  and (_07970_, _07936_, _07926_);
  and (_07971_, _07970_, \uc8051golden_1.P1 [7]);
  and (_07972_, _07936_, _07947_);
  and (_07973_, _07972_, \uc8051golden_1.SCON [7]);
  nor (_07974_, _07973_, _07971_);
  and (_07975_, _07964_, _07937_);
  and (_07976_, _07975_, _07954_);
  and (_07977_, _07976_, \uc8051golden_1.TL1 [7]);
  nor (_07978_, _06693_, _06372_);
  and (_07979_, _07978_, _07938_);
  and (_07980_, _07979_, _07954_);
  and (_07981_, _07980_, \uc8051golden_1.TH1 [7]);
  nor (_07982_, _07981_, _07977_);
  and (_07983_, _07982_, _07974_);
  and (_07984_, _07983_, _07969_);
  and (_07985_, _07984_, _07952_);
  nor (_07986_, _06340_, _06309_);
  and (_07987_, _07986_, _07935_);
  and (_07988_, _07987_, _07926_);
  and (_07989_, _07988_, \uc8051golden_1.PSW [7]);
  not (_07990_, _07989_);
  and (_07991_, _07986_, _07943_);
  and (_07992_, _07991_, _07926_);
  and (_07993_, _07992_, \uc8051golden_1.B [7]);
  and (_07994_, _07929_, _07986_);
  and (_07995_, _07994_, _07926_);
  and (_07996_, _07995_, \uc8051golden_1.ACC [7]);
  nor (_07997_, _07996_, _07993_);
  and (_07998_, _07997_, _07990_);
  and (_07999_, _07944_, _07947_);
  and (_08000_, _07999_, \uc8051golden_1.IP [7]);
  and (_08001_, _07964_, _07573_);
  and (_08002_, _08001_, _07959_);
  and (_08003_, _08002_, \uc8051golden_1.PCON [7]);
  nor (_08004_, _08003_, _08000_);
  and (_08005_, _08004_, _07998_);
  and (_08006_, _07939_, _07954_);
  and (_08007_, _08006_, \uc8051golden_1.TMOD [7]);
  not (_08008_, _08007_);
  and (_08009_, _07960_, _07937_);
  and (_08010_, _08009_, _07954_);
  and (_08011_, _08010_, \uc8051golden_1.TL0 [7]);
  and (_08012_, _07978_, _07924_);
  and (_08013_, _08012_, _07954_);
  and (_08014_, _08013_, \uc8051golden_1.TH0 [7]);
  nor (_08015_, _08014_, _08011_);
  and (_08016_, _08015_, _08008_);
  and (_08017_, _07947_, _07954_);
  and (_08018_, _08017_, \uc8051golden_1.TCON [7]);
  and (_08019_, _07926_, _07954_);
  and (_08020_, _08019_, \uc8051golden_1.P0 [7]);
  nor (_08021_, _08020_, _08018_);
  and (_08022_, _08021_, _08016_);
  and (_08023_, _08022_, _08005_);
  and (_08024_, _08023_, _07985_);
  not (_08025_, \uc8051golden_1.IRAM[1] [7]);
  or (_08026_, _07053_, _08025_);
  nand (_08027_, _07053_, \uc8051golden_1.IRAM[0] [7]);
  and (_08028_, _08027_, _07141_);
  nand (_08029_, _08028_, _08026_);
  nand (_08030_, _07053_, \uc8051golden_1.IRAM[2] [7]);
  nand (_08031_, _07146_, \uc8051golden_1.IRAM[3] [7]);
  and (_08032_, _08031_, _07148_);
  nand (_08033_, _08032_, _08030_);
  nand (_08034_, _08033_, _08029_);
  nand (_08035_, _08034_, _06805_);
  nand (_08036_, _07053_, \uc8051golden_1.IRAM[6] [7]);
  nand (_08037_, _07146_, \uc8051golden_1.IRAM[7] [7]);
  and (_08038_, _08037_, _07148_);
  nand (_08039_, _08038_, _08036_);
  nand (_08040_, _07146_, \uc8051golden_1.IRAM[5] [7]);
  nand (_08041_, _07053_, \uc8051golden_1.IRAM[4] [7]);
  and (_08042_, _08041_, _07141_);
  nand (_08043_, _08042_, _08040_);
  nand (_08044_, _08043_, _08039_);
  nand (_08045_, _08044_, _07155_);
  nand (_08046_, _08045_, _08035_);
  nand (_08047_, _08046_, _06618_);
  nand (_08048_, _07053_, \uc8051golden_1.IRAM[10] [7]);
  nand (_08049_, _07146_, \uc8051golden_1.IRAM[11] [7]);
  and (_08050_, _08049_, _07148_);
  nand (_08051_, _08050_, _08048_);
  nand (_08052_, _07146_, \uc8051golden_1.IRAM[9] [7]);
  nand (_08053_, _07053_, \uc8051golden_1.IRAM[8] [7]);
  and (_08054_, _08053_, _07141_);
  nand (_08055_, _08054_, _08052_);
  nand (_08056_, _08055_, _08051_);
  nand (_08057_, _08056_, _06805_);
  nand (_08058_, _07053_, \uc8051golden_1.IRAM[14] [7]);
  or (_08059_, _07053_, _05652_);
  and (_08060_, _08059_, _07148_);
  nand (_08061_, _08060_, _08058_);
  nand (_08062_, _07146_, \uc8051golden_1.IRAM[13] [7]);
  nand (_08063_, _07053_, \uc8051golden_1.IRAM[12] [7]);
  and (_08064_, _08063_, _07141_);
  nand (_08065_, _08064_, _08062_);
  nand (_08066_, _08065_, _08061_);
  nand (_08067_, _08066_, _07155_);
  nand (_08068_, _08067_, _08057_);
  nand (_08069_, _08068_, _07172_);
  nand (_08070_, _08069_, _08047_);
  or (_08071_, _08070_, _06194_);
  and (_08072_, _08071_, _08024_);
  not (_08073_, _08072_);
  nand (_08074_, _07146_, \uc8051golden_1.IRAM[1] [6]);
  nand (_08075_, _07053_, \uc8051golden_1.IRAM[0] [6]);
  and (_08076_, _08075_, _07141_);
  nand (_08077_, _08076_, _08074_);
  nand (_08078_, _07053_, \uc8051golden_1.IRAM[2] [6]);
  nand (_08079_, _07146_, \uc8051golden_1.IRAM[3] [6]);
  and (_08080_, _08079_, _07148_);
  nand (_08081_, _08080_, _08078_);
  nand (_08082_, _08081_, _08077_);
  nand (_08083_, _08082_, _06805_);
  nand (_08084_, _07053_, \uc8051golden_1.IRAM[6] [6]);
  nand (_08085_, _07146_, \uc8051golden_1.IRAM[7] [6]);
  and (_08086_, _08085_, _07148_);
  nand (_08087_, _08086_, _08084_);
  nand (_08088_, _07146_, \uc8051golden_1.IRAM[5] [6]);
  nand (_08089_, _07053_, \uc8051golden_1.IRAM[4] [6]);
  and (_08090_, _08089_, _07141_);
  nand (_08091_, _08090_, _08088_);
  nand (_08092_, _08091_, _08087_);
  nand (_08093_, _08092_, _07155_);
  nand (_08094_, _08093_, _08083_);
  nand (_08095_, _08094_, _06618_);
  nand (_08096_, _07053_, \uc8051golden_1.IRAM[10] [6]);
  nand (_08097_, _07146_, \uc8051golden_1.IRAM[11] [6]);
  and (_08098_, _08097_, _07148_);
  nand (_08099_, _08098_, _08096_);
  nand (_08100_, _07146_, \uc8051golden_1.IRAM[9] [6]);
  nand (_08101_, _07053_, \uc8051golden_1.IRAM[8] [6]);
  and (_08102_, _08101_, _07141_);
  nand (_08103_, _08102_, _08100_);
  nand (_08104_, _08103_, _08099_);
  nand (_08105_, _08104_, _06805_);
  nand (_08106_, _07053_, \uc8051golden_1.IRAM[14] [6]);
  nand (_08107_, _07146_, \uc8051golden_1.IRAM[15] [6]);
  and (_08108_, _08107_, _07148_);
  nand (_08109_, _08108_, _08106_);
  nand (_08110_, _07146_, \uc8051golden_1.IRAM[13] [6]);
  nand (_08111_, _07053_, \uc8051golden_1.IRAM[12] [6]);
  and (_08112_, _08111_, _07141_);
  nand (_08113_, _08112_, _08110_);
  nand (_08114_, _08113_, _08109_);
  nand (_08115_, _08114_, _07155_);
  nand (_08116_, _08115_, _08105_);
  nand (_08117_, _08116_, _07172_);
  nand (_08118_, _08117_, _08095_);
  or (_08119_, _08118_, _06194_);
  and (_08120_, _07940_, \uc8051golden_1.SBUF [6]);
  and (_08121_, _07931_, \uc8051golden_1.P2 [6]);
  and (_08122_, _07948_, \uc8051golden_1.IE [6]);
  and (_08123_, _07945_, \uc8051golden_1.P3 [6]);
  or (_08124_, _08123_, _08122_);
  or (_08125_, _08124_, _08121_);
  nor (_08126_, _08125_, _08120_);
  and (_08127_, _07970_, \uc8051golden_1.P1 [6]);
  and (_08128_, _07972_, \uc8051golden_1.SCON [6]);
  nor (_08129_, _08128_, _08127_);
  and (_08130_, _07976_, \uc8051golden_1.TL1 [6]);
  and (_08131_, _07980_, \uc8051golden_1.TH1 [6]);
  nor (_08132_, _08131_, _08130_);
  and (_08133_, _08132_, _08129_);
  and (_08134_, _08133_, _08126_);
  and (_08135_, _07988_, \uc8051golden_1.PSW [6]);
  and (_08136_, _07992_, \uc8051golden_1.B [6]);
  and (_08137_, _07995_, \uc8051golden_1.ACC [6]);
  or (_08138_, _08137_, _08136_);
  nor (_08139_, _08138_, _08135_);
  and (_08140_, _08002_, \uc8051golden_1.PCON [6]);
  and (_08141_, _07999_, \uc8051golden_1.IP [6]);
  nor (_08142_, _08141_, _08140_);
  and (_08143_, _08142_, _08139_);
  and (_08144_, _08017_, \uc8051golden_1.TCON [6]);
  and (_08145_, _08010_, \uc8051golden_1.TL0 [6]);
  and (_08146_, _08013_, \uc8051golden_1.TH0 [6]);
  or (_08147_, _08146_, _08145_);
  nor (_08148_, _08147_, _08144_);
  and (_08149_, _08006_, \uc8051golden_1.TMOD [6]);
  and (_08150_, _07962_, \uc8051golden_1.DPL [6]);
  and (_08151_, _07966_, \uc8051golden_1.DPH [6]);
  or (_08152_, _08151_, _08150_);
  and (_08153_, _08019_, \uc8051golden_1.P0 [6]);
  and (_08154_, _07956_, \uc8051golden_1.SP [6]);
  or (_08155_, _08154_, _08153_);
  or (_08156_, _08155_, _08152_);
  nor (_08157_, _08156_, _08149_);
  and (_08158_, _08157_, _08148_);
  and (_08159_, _08158_, _08143_);
  and (_08160_, _08159_, _08134_);
  and (_08161_, _08160_, _08119_);
  not (_08162_, _08161_);
  nand (_08163_, _07146_, \uc8051golden_1.IRAM[1] [5]);
  nand (_08164_, _07053_, \uc8051golden_1.IRAM[0] [5]);
  and (_08165_, _08164_, _07141_);
  nand (_08166_, _08165_, _08163_);
  nand (_08167_, _07053_, \uc8051golden_1.IRAM[2] [5]);
  nand (_08168_, _07146_, \uc8051golden_1.IRAM[3] [5]);
  and (_08169_, _08168_, _07148_);
  nand (_08170_, _08169_, _08167_);
  nand (_08171_, _08170_, _08166_);
  nand (_08172_, _08171_, _06805_);
  nand (_08173_, _07053_, \uc8051golden_1.IRAM[6] [5]);
  nand (_08174_, _07146_, \uc8051golden_1.IRAM[7] [5]);
  and (_08175_, _08174_, _07148_);
  nand (_08176_, _08175_, _08173_);
  nand (_08177_, _07146_, \uc8051golden_1.IRAM[5] [5]);
  nand (_08178_, _07053_, \uc8051golden_1.IRAM[4] [5]);
  and (_08179_, _08178_, _07141_);
  nand (_08180_, _08179_, _08177_);
  nand (_08181_, _08180_, _08176_);
  nand (_08182_, _08181_, _07155_);
  nand (_08183_, _08182_, _08172_);
  nand (_08184_, _08183_, _06618_);
  nand (_08185_, _07053_, \uc8051golden_1.IRAM[10] [5]);
  nand (_08186_, _07146_, \uc8051golden_1.IRAM[11] [5]);
  and (_08187_, _08186_, _07148_);
  nand (_08188_, _08187_, _08185_);
  nand (_08189_, _07146_, \uc8051golden_1.IRAM[9] [5]);
  nand (_08190_, _07053_, \uc8051golden_1.IRAM[8] [5]);
  and (_08191_, _08190_, _07141_);
  nand (_08192_, _08191_, _08189_);
  nand (_08193_, _08192_, _08188_);
  nand (_08194_, _08193_, _06805_);
  nand (_08195_, _07053_, \uc8051golden_1.IRAM[14] [5]);
  nand (_08196_, _07146_, \uc8051golden_1.IRAM[15] [5]);
  and (_08197_, _08196_, _07148_);
  nand (_08198_, _08197_, _08195_);
  nand (_08199_, _07146_, \uc8051golden_1.IRAM[13] [5]);
  nand (_08200_, _07053_, \uc8051golden_1.IRAM[12] [5]);
  and (_08201_, _08200_, _07141_);
  nand (_08202_, _08201_, _08199_);
  nand (_08203_, _08202_, _08198_);
  nand (_08204_, _08203_, _07155_);
  nand (_08205_, _08204_, _08194_);
  nand (_08206_, _08205_, _07172_);
  nand (_08207_, _08206_, _08184_);
  or (_08208_, _08207_, _06194_);
  and (_08209_, _07999_, \uc8051golden_1.IP [5]);
  and (_08210_, _07988_, \uc8051golden_1.PSW [5]);
  nor (_08211_, _08210_, _08209_);
  and (_08212_, _07970_, \uc8051golden_1.P1 [5]);
  and (_08213_, _07992_, \uc8051golden_1.B [5]);
  nor (_08214_, _08213_, _08212_);
  and (_08215_, _08214_, _08211_);
  and (_08216_, _07980_, \uc8051golden_1.TH1 [5]);
  and (_08217_, _07995_, \uc8051golden_1.ACC [5]);
  nor (_08218_, _08217_, _08216_);
  and (_08219_, _07976_, \uc8051golden_1.TL1 [5]);
  and (_08220_, _07945_, \uc8051golden_1.P3 [5]);
  nor (_08221_, _08220_, _08219_);
  and (_08222_, _08221_, _08218_);
  and (_08223_, _07972_, \uc8051golden_1.SCON [5]);
  and (_08224_, _07948_, \uc8051golden_1.IE [5]);
  nor (_08225_, _08224_, _08223_);
  and (_08226_, _07940_, \uc8051golden_1.SBUF [5]);
  and (_08227_, _07931_, \uc8051golden_1.P2 [5]);
  nor (_08228_, _08227_, _08226_);
  and (_08229_, _08228_, _08225_);
  and (_08230_, _08229_, _08222_);
  and (_08231_, _08230_, _08215_);
  and (_08232_, _08019_, \uc8051golden_1.P0 [5]);
  not (_08233_, _08232_);
  and (_08234_, _07962_, \uc8051golden_1.DPL [5]);
  and (_08235_, _07938_, _06693_);
  and (_08236_, _07959_, _08235_);
  and (_08237_, _08236_, \uc8051golden_1.SP [5]);
  nor (_08238_, _08237_, _08234_);
  and (_08239_, _08238_, _08233_);
  and (_08240_, _08010_, \uc8051golden_1.TL0 [5]);
  and (_08241_, _08013_, \uc8051golden_1.TH0 [5]);
  nor (_08242_, _08241_, _08240_);
  and (_08243_, _08017_, \uc8051golden_1.TCON [5]);
  and (_08244_, _08006_, \uc8051golden_1.TMOD [5]);
  nor (_08245_, _08244_, _08243_);
  and (_08246_, _08245_, _08242_);
  and (_08247_, _08002_, \uc8051golden_1.PCON [5]);
  and (_08248_, _07964_, _06693_);
  and (_08249_, _08248_, _07959_);
  and (_08250_, _08249_, \uc8051golden_1.DPH [5]);
  nor (_08251_, _08250_, _08247_);
  and (_08252_, _08251_, _08246_);
  and (_08253_, _08252_, _08239_);
  and (_08254_, _08253_, _08231_);
  and (_08255_, _08254_, _08208_);
  not (_08256_, _08255_);
  nand (_08257_, _07146_, \uc8051golden_1.IRAM[1] [4]);
  nand (_08258_, _07053_, \uc8051golden_1.IRAM[0] [4]);
  and (_08259_, _08258_, _07141_);
  nand (_08260_, _08259_, _08257_);
  nand (_08261_, _07053_, \uc8051golden_1.IRAM[2] [4]);
  nand (_08262_, _07146_, \uc8051golden_1.IRAM[3] [4]);
  and (_08263_, _08262_, _07148_);
  nand (_08264_, _08263_, _08261_);
  nand (_08265_, _08264_, _08260_);
  nand (_08266_, _08265_, _06805_);
  nand (_08267_, _07053_, \uc8051golden_1.IRAM[6] [4]);
  nand (_08268_, _07146_, \uc8051golden_1.IRAM[7] [4]);
  and (_08269_, _08268_, _07148_);
  nand (_08270_, _08269_, _08267_);
  nand (_08271_, _07146_, \uc8051golden_1.IRAM[5] [4]);
  nand (_08272_, _07053_, \uc8051golden_1.IRAM[4] [4]);
  and (_08273_, _08272_, _07141_);
  nand (_08274_, _08273_, _08271_);
  nand (_08275_, _08274_, _08270_);
  nand (_08276_, _08275_, _07155_);
  nand (_08277_, _08276_, _08266_);
  nand (_08278_, _08277_, _06618_);
  nand (_08279_, _07053_, \uc8051golden_1.IRAM[10] [4]);
  nand (_08280_, _07146_, \uc8051golden_1.IRAM[11] [4]);
  and (_08281_, _08280_, _07148_);
  nand (_08282_, _08281_, _08279_);
  nand (_08283_, _07146_, \uc8051golden_1.IRAM[9] [4]);
  nand (_08284_, _07053_, \uc8051golden_1.IRAM[8] [4]);
  and (_08285_, _08284_, _07141_);
  nand (_08286_, _08285_, _08283_);
  nand (_08287_, _08286_, _08282_);
  nand (_08288_, _08287_, _06805_);
  nand (_08289_, _07053_, \uc8051golden_1.IRAM[14] [4]);
  nand (_08290_, _07146_, \uc8051golden_1.IRAM[15] [4]);
  and (_08291_, _08290_, _07148_);
  nand (_08292_, _08291_, _08289_);
  nand (_08293_, _07146_, \uc8051golden_1.IRAM[13] [4]);
  nand (_08294_, _07053_, \uc8051golden_1.IRAM[12] [4]);
  and (_08295_, _08294_, _07141_);
  nand (_08296_, _08295_, _08293_);
  nand (_08297_, _08296_, _08292_);
  nand (_08298_, _08297_, _07155_);
  nand (_08299_, _08298_, _08288_);
  nand (_08300_, _08299_, _07172_);
  nand (_08301_, _08300_, _08278_);
  or (_08302_, _08301_, _06194_);
  and (_08303_, _07945_, \uc8051golden_1.P3 [4]);
  and (_08304_, _07995_, \uc8051golden_1.ACC [4]);
  or (_08305_, _08304_, _08303_);
  and (_08306_, _07988_, \uc8051golden_1.PSW [4]);
  and (_08307_, _07992_, \uc8051golden_1.B [4]);
  or (_08308_, _08307_, _08306_);
  or (_08309_, _08308_, _08305_);
  and (_08310_, _07970_, \uc8051golden_1.P1 [4]);
  and (_08311_, _07972_, \uc8051golden_1.SCON [4]);
  nor (_08312_, _08311_, _08310_);
  and (_08313_, _08010_, \uc8051golden_1.TL0 [4]);
  and (_08314_, _07999_, \uc8051golden_1.IP [4]);
  nor (_08315_, _08314_, _08313_);
  nand (_08316_, _08315_, _08312_);
  and (_08317_, _08017_, \uc8051golden_1.TCON [4]);
  and (_08318_, _07980_, \uc8051golden_1.TH1 [4]);
  or (_08319_, _08318_, _08317_);
  and (_08320_, _08013_, \uc8051golden_1.TH0 [4]);
  and (_08321_, _07931_, \uc8051golden_1.P2 [4]);
  or (_08322_, _08321_, _08320_);
  or (_08323_, _08322_, _08319_);
  or (_08324_, _08323_, _08316_);
  or (_08325_, _08324_, _08309_);
  and (_08326_, _07962_, \uc8051golden_1.DPL [4]);
  and (_08327_, _08019_, \uc8051golden_1.P0 [4]);
  and (_08328_, _08249_, \uc8051golden_1.DPH [4]);
  or (_08329_, _08328_, _08327_);
  or (_08330_, _08329_, _08326_);
  and (_08331_, _08006_, \uc8051golden_1.TMOD [4]);
  and (_08332_, _07940_, \uc8051golden_1.SBUF [4]);
  or (_08333_, _08332_, _08331_);
  and (_08334_, _07976_, \uc8051golden_1.TL1 [4]);
  and (_08335_, _07948_, \uc8051golden_1.IE [4]);
  or (_08336_, _08335_, _08334_);
  or (_08337_, _08336_, _08333_);
  and (_08338_, _08002_, \uc8051golden_1.PCON [4]);
  and (_08339_, _08236_, \uc8051golden_1.SP [4]);
  or (_08340_, _08339_, _08338_);
  or (_08341_, _08340_, _08337_);
  or (_08342_, _08341_, _08330_);
  nor (_08343_, _08342_, _08325_);
  and (_08344_, _08343_, _08302_);
  not (_08345_, _08344_);
  or (_08346_, _07775_, _06194_);
  and (_08347_, _08019_, \uc8051golden_1.P0 [3]);
  and (_08348_, _07956_, \uc8051golden_1.SP [3]);
  and (_08349_, _07962_, \uc8051golden_1.DPL [3]);
  and (_08350_, _07966_, \uc8051golden_1.DPH [3]);
  and (_08351_, _08002_, \uc8051golden_1.PCON [3]);
  and (_08352_, _08017_, \uc8051golden_1.TCON [3]);
  and (_08353_, _08006_, \uc8051golden_1.TMOD [3]);
  and (_08354_, _08010_, \uc8051golden_1.TL0 [3]);
  and (_08355_, _08013_, \uc8051golden_1.TH0 [3]);
  and (_08356_, _07976_, \uc8051golden_1.TL1 [3]);
  and (_08357_, _07980_, \uc8051golden_1.TH1 [3]);
  and (_08358_, _07970_, \uc8051golden_1.P1 [3]);
  and (_08359_, _07972_, \uc8051golden_1.SCON [3]);
  and (_08360_, _07940_, \uc8051golden_1.SBUF [3]);
  and (_08361_, _07931_, \uc8051golden_1.P2 [3]);
  and (_08362_, _07948_, \uc8051golden_1.IE [3]);
  and (_08363_, _07945_, \uc8051golden_1.P3 [3]);
  and (_08364_, _07999_, \uc8051golden_1.IP [3]);
  and (_08365_, _07988_, \uc8051golden_1.PSW [3]);
  and (_08366_, _07995_, \uc8051golden_1.ACC [3]);
  and (_08367_, _07992_, \uc8051golden_1.B [3]);
  or (_08368_, _08367_, _08366_);
  or (_08369_, _08368_, _08365_);
  or (_08370_, _08369_, _08364_);
  or (_08371_, _08370_, _08363_);
  or (_08372_, _08371_, _08362_);
  or (_08373_, _08372_, _08361_);
  or (_08374_, _08373_, _08360_);
  or (_08375_, _08374_, _08359_);
  or (_08376_, _08375_, _08358_);
  or (_08377_, _08376_, _08357_);
  or (_08378_, _08377_, _08356_);
  or (_08379_, _08378_, _08355_);
  or (_08380_, _08379_, _08354_);
  or (_08381_, _08380_, _08353_);
  or (_08382_, _08381_, _08352_);
  or (_08383_, _08382_, _08351_);
  or (_08384_, _08383_, _08350_);
  or (_08385_, _08384_, _08349_);
  or (_08386_, _08385_, _08348_);
  nor (_08387_, _08386_, _08347_);
  and (_08388_, _08387_, _08346_);
  not (_08389_, _08388_);
  or (_08390_, _07623_, _06194_);
  and (_08391_, _08019_, \uc8051golden_1.P0 [2]);
  and (_08392_, _07956_, \uc8051golden_1.SP [2]);
  and (_08393_, _07962_, \uc8051golden_1.DPL [2]);
  and (_08394_, _07966_, \uc8051golden_1.DPH [2]);
  and (_08395_, _08002_, \uc8051golden_1.PCON [2]);
  and (_08396_, _08017_, \uc8051golden_1.TCON [2]);
  and (_08397_, _08006_, \uc8051golden_1.TMOD [2]);
  and (_08398_, _08010_, \uc8051golden_1.TL0 [2]);
  and (_08399_, _08013_, \uc8051golden_1.TH0 [2]);
  and (_08400_, _07976_, \uc8051golden_1.TL1 [2]);
  and (_08401_, _07980_, \uc8051golden_1.TH1 [2]);
  and (_08402_, _07970_, \uc8051golden_1.P1 [2]);
  and (_08403_, _07972_, \uc8051golden_1.SCON [2]);
  and (_08404_, _07940_, \uc8051golden_1.SBUF [2]);
  and (_08405_, _07931_, \uc8051golden_1.P2 [2]);
  and (_08406_, _07948_, \uc8051golden_1.IE [2]);
  and (_08407_, _07945_, \uc8051golden_1.P3 [2]);
  and (_08408_, _07999_, \uc8051golden_1.IP [2]);
  and (_08409_, _07988_, \uc8051golden_1.PSW [2]);
  and (_08410_, _07992_, \uc8051golden_1.B [2]);
  and (_08411_, _07995_, \uc8051golden_1.ACC [2]);
  or (_08412_, _08411_, _08410_);
  or (_08413_, _08412_, _08409_);
  or (_08414_, _08413_, _08408_);
  or (_08415_, _08414_, _08407_);
  or (_08416_, _08415_, _08406_);
  or (_08417_, _08416_, _08405_);
  or (_08418_, _08417_, _08404_);
  or (_08419_, _08418_, _08403_);
  or (_08420_, _08419_, _08402_);
  or (_08421_, _08420_, _08401_);
  or (_08422_, _08421_, _08400_);
  or (_08423_, _08422_, _08399_);
  or (_08424_, _08423_, _08398_);
  or (_08425_, _08424_, _08397_);
  or (_08426_, _08425_, _08396_);
  or (_08427_, _08426_, _08395_);
  or (_08428_, _08427_, _08394_);
  or (_08429_, _08428_, _08393_);
  or (_08430_, _08429_, _08392_);
  nor (_08431_, _08430_, _08391_);
  and (_08432_, _08431_, _08390_);
  not (_08433_, _08432_);
  or (_08434_, _07196_, _06194_);
  and (_08435_, _07940_, \uc8051golden_1.SBUF [1]);
  and (_08436_, _07931_, \uc8051golden_1.P2 [1]);
  and (_08437_, _07945_, \uc8051golden_1.P3 [1]);
  and (_08438_, _07948_, \uc8051golden_1.IE [1]);
  or (_08439_, _08438_, _08437_);
  or (_08440_, _08439_, _08436_);
  nor (_08441_, _08440_, _08435_);
  and (_08442_, _07970_, \uc8051golden_1.P1 [1]);
  and (_08443_, _07972_, \uc8051golden_1.SCON [1]);
  nor (_08444_, _08443_, _08442_);
  and (_08445_, _07980_, \uc8051golden_1.TH1 [1]);
  and (_08446_, _07976_, \uc8051golden_1.TL1 [1]);
  nor (_08447_, _08446_, _08445_);
  and (_08448_, _08447_, _08444_);
  and (_08449_, _08448_, _08441_);
  and (_08450_, _07999_, \uc8051golden_1.IP [1]);
  and (_08451_, _07995_, \uc8051golden_1.ACC [1]);
  and (_08452_, _07992_, \uc8051golden_1.B [1]);
  or (_08453_, _08452_, _08451_);
  nor (_08454_, _08453_, _08450_);
  and (_08455_, _07988_, \uc8051golden_1.PSW [1]);
  and (_08456_, _08002_, \uc8051golden_1.PCON [1]);
  nor (_08457_, _08456_, _08455_);
  and (_08458_, _08457_, _08454_);
  and (_08459_, _08006_, \uc8051golden_1.TMOD [1]);
  and (_08460_, _08010_, \uc8051golden_1.TL0 [1]);
  and (_08461_, _08013_, \uc8051golden_1.TH0 [1]);
  or (_08462_, _08461_, _08460_);
  nor (_08463_, _08462_, _08459_);
  and (_08464_, _08017_, \uc8051golden_1.TCON [1]);
  and (_08465_, _07962_, \uc8051golden_1.DPL [1]);
  and (_08466_, _07966_, \uc8051golden_1.DPH [1]);
  or (_08467_, _08466_, _08465_);
  and (_08468_, _08019_, \uc8051golden_1.P0 [1]);
  and (_08469_, _07956_, \uc8051golden_1.SP [1]);
  or (_08470_, _08469_, _08468_);
  or (_08471_, _08470_, _08467_);
  nor (_08472_, _08471_, _08464_);
  and (_08473_, _08472_, _08463_);
  and (_08474_, _08473_, _08458_);
  and (_08475_, _08474_, _08449_);
  and (_08476_, _08475_, _08434_);
  not (_08477_, _08476_);
  or (_08478_, _07485_, _06194_);
  and (_08479_, _07970_, \uc8051golden_1.P1 [0]);
  and (_08480_, _07992_, \uc8051golden_1.B [0]);
  nor (_08481_, _08480_, _08479_);
  and (_08482_, _07988_, \uc8051golden_1.PSW [0]);
  and (_08483_, _07995_, \uc8051golden_1.ACC [0]);
  nor (_08484_, _08483_, _08482_);
  and (_08485_, _08484_, _08481_);
  and (_08486_, _08013_, \uc8051golden_1.TH0 [0]);
  and (_08487_, _07976_, \uc8051golden_1.TL1 [0]);
  nor (_08488_, _08487_, _08486_);
  and (_08489_, _07940_, \uc8051golden_1.SBUF [0]);
  and (_08490_, _07945_, \uc8051golden_1.P3 [0]);
  nor (_08491_, _08490_, _08489_);
  and (_08492_, _08491_, _08488_);
  and (_08493_, _07972_, \uc8051golden_1.SCON [0]);
  and (_08494_, _07931_, \uc8051golden_1.P2 [0]);
  nor (_08495_, _08494_, _08493_);
  and (_08496_, _08006_, \uc8051golden_1.TMOD [0]);
  and (_08497_, _07948_, \uc8051golden_1.IE [0]);
  nor (_08498_, _08497_, _08496_);
  and (_08499_, _08498_, _08495_);
  and (_08500_, _08499_, _08492_);
  and (_08501_, _08500_, _08485_);
  and (_08502_, _08019_, \uc8051golden_1.P0 [0]);
  not (_08503_, _08502_);
  nand (_08504_, _08249_, \uc8051golden_1.DPH [0]);
  nand (_08505_, _08236_, \uc8051golden_1.SP [0]);
  and (_08506_, _08505_, _08504_);
  and (_08507_, _08506_, _08503_);
  and (_08508_, _08010_, \uc8051golden_1.TL0 [0]);
  and (_08509_, _07980_, \uc8051golden_1.TH1 [0]);
  nor (_08510_, _08509_, _08508_);
  and (_08511_, _08017_, \uc8051golden_1.TCON [0]);
  and (_08512_, _07999_, \uc8051golden_1.IP [0]);
  nor (_08513_, _08512_, _08511_);
  and (_08514_, _08513_, _08510_);
  and (_08515_, _07962_, \uc8051golden_1.DPL [0]);
  and (_08516_, _08002_, \uc8051golden_1.PCON [0]);
  nor (_08517_, _08516_, _08515_);
  and (_08518_, _08517_, _08514_);
  and (_08519_, _08518_, _08507_);
  and (_08520_, _08519_, _08501_);
  nand (_08521_, _08520_, _08478_);
  and (_08522_, _08521_, _08477_);
  and (_08523_, _08522_, _08433_);
  and (_08524_, _08523_, _08389_);
  and (_08525_, _08524_, _08345_);
  and (_08526_, _08525_, _08256_);
  and (_08527_, _08526_, _08162_);
  or (_08528_, _08527_, _08073_);
  nand (_08529_, _08527_, _08073_);
  and (_08530_, _08529_, _08528_);
  and (_08531_, _08530_, _06197_);
  and (_08532_, \uc8051golden_1.PC [5], \uc8051golden_1.PC [4]);
  and (_08533_, _08532_, \uc8051golden_1.PC [6]);
  and (_08534_, _05689_, \uc8051golden_1.PC [2]);
  and (_08535_, _08534_, \uc8051golden_1.PC [3]);
  and (_08536_, _08535_, _08533_);
  and (_08537_, _08536_, \uc8051golden_1.PC [7]);
  nor (_08538_, _08536_, \uc8051golden_1.PC [7]);
  nor (_08539_, _08538_, _08537_);
  not (_08540_, _08539_);
  nand (_08541_, _08540_, _06465_);
  and (_08542_, _07378_, _05968_);
  not (_08543_, _08542_);
  and (_08544_, _06462_, _05968_);
  nor (_08545_, _07694_, _08544_);
  and (_08546_, _08545_, _08543_);
  not (_08547_, _07300_);
  not (_08548_, _08070_);
  and (_08549_, _08301_, _08207_);
  and (_08550_, _07775_, _07623_);
  and (_08551_, _07485_, _07196_);
  and (_08552_, _08551_, _08550_);
  and (_08553_, _08552_, _08549_);
  and (_08554_, _08553_, _08118_);
  or (_08555_, _08554_, _08548_);
  nand (_08556_, _08554_, _08548_);
  and (_08557_, _08556_, _08555_);
  and (_08558_, _08557_, _08547_);
  or (_08559_, _08558_, _08546_);
  and (_08560_, _06508_, _04587_);
  and (_08561_, _06512_, _04585_);
  nor (_08562_, _08561_, _08560_);
  and (_08563_, _06516_, _04559_);
  and (_08564_, _06555_, _04575_);
  nor (_08565_, _08564_, _08563_);
  and (_08566_, _08565_, _08562_);
  and (_08567_, _06526_, _04561_);
  and (_08568_, _06528_, _04578_);
  nor (_08569_, _08568_, _08567_);
  and (_08570_, _06532_, _04595_);
  and (_08571_, _06552_, _04602_);
  nor (_08572_, _08571_, _08570_);
  and (_08573_, _08572_, _08569_);
  and (_08574_, _08573_, _08566_);
  and (_08575_, _06539_, _04507_);
  and (_08576_, _06541_, _04556_);
  nor (_08577_, _08576_, _08575_);
  and (_08578_, _06544_, _04554_);
  and (_08579_, _06546_, _04571_);
  nor (_08580_, _08579_, _08578_);
  and (_08581_, _08580_, _08577_);
  and (_08582_, _06550_, _04568_);
  and (_08583_, _06534_, _04583_);
  nor (_08584_, _08583_, _08582_);
  and (_08585_, _06520_, _04592_);
  and (_08586_, _06557_, _04599_);
  nor (_08587_, _08586_, _08585_);
  and (_08588_, _08587_, _08584_);
  and (_08589_, _08588_, _08581_);
  and (_08590_, _08589_, _08574_);
  nor (_08591_, _08590_, _08072_);
  and (_08592_, _08591_, _07280_);
  not (_08593_, _08001_);
  not (_08594_, _06808_);
  nor (_08595_, _08594_, _06266_);
  nor (_08596_, _06651_, _06374_);
  and (_08597_, _08596_, _08595_);
  and (_08598_, _08597_, _07944_);
  and (_08599_, _08598_, \uc8051golden_1.P3 [7]);
  not (_08600_, _06651_);
  and (_08601_, _08600_, _06374_);
  and (_08602_, _08601_, _08595_);
  and (_08603_, _08602_, _07930_);
  and (_08604_, _08603_, \uc8051golden_1.IE [7]);
  nor (_08605_, _08604_, _08599_);
  and (_08606_, _08602_, _07936_);
  and (_08607_, _08606_, \uc8051golden_1.SCON [7]);
  and (_08608_, _08597_, _07930_);
  and (_08609_, _08608_, \uc8051golden_1.P2 [7]);
  nor (_08610_, _08609_, _08607_);
  and (_08611_, _08610_, _08605_);
  and (_08612_, _08597_, _07987_);
  and (_08613_, _08612_, \uc8051golden_1.PSW [7]);
  and (_08614_, _08602_, _07944_);
  and (_08615_, _08614_, \uc8051golden_1.IP [7]);
  and (_08616_, _08597_, _07994_);
  and (_08617_, _08616_, \uc8051golden_1.ACC [7]);
  and (_08618_, _08597_, _07991_);
  and (_08619_, _08618_, \uc8051golden_1.B [7]);
  or (_08620_, _08619_, _08617_);
  or (_08621_, _08620_, _08615_);
  nor (_08622_, _08621_, _08613_);
  and (_08623_, _08602_, _07954_);
  and (_08624_, _08623_, \uc8051golden_1.TCON [7]);
  and (_08625_, _07959_, \uc8051golden_1.P0 [7]);
  and (_08626_, _08597_, _07936_);
  and (_08627_, _08626_, \uc8051golden_1.P1 [7]);
  or (_08628_, _08627_, _08625_);
  nor (_08629_, _08628_, _08624_);
  and (_08630_, _08629_, _08622_);
  and (_08631_, _08630_, _08611_);
  and (_08632_, _08631_, _08071_);
  nor (_08633_, _08632_, _08593_);
  not (_08634_, _08633_);
  nand (_08635_, _08632_, _08593_);
  and (_08636_, _08635_, _08634_);
  and (_08637_, _08636_, _07246_);
  not (_08638_, _07239_);
  nor (_08639_, _08632_, _08001_);
  or (_08640_, _08639_, _08638_);
  not (_08641_, _07218_);
  or (_08642_, _08635_, _08641_);
  nor (_08643_, _05996_, _06012_);
  not (_08644_, _08643_);
  or (_08645_, _08644_, _08557_);
  and (_08646_, _08533_, _06122_);
  and (_08647_, _08646_, \uc8051golden_1.PC [7]);
  nor (_08648_, _08646_, \uc8051golden_1.PC [7]);
  nor (_08649_, _08648_, _08647_);
  and (_08650_, _08649_, _06790_);
  not (_08651_, \uc8051golden_1.ACC [7]);
  nor (_08652_, _06790_, _08651_);
  or (_08653_, _08652_, _08650_);
  or (_08654_, _07355_, _07631_);
  or (_08655_, _08654_, _08653_);
  or (_08656_, _08655_, _07633_);
  and (_08657_, _08656_, _08645_);
  or (_08658_, _08657_, _07212_);
  not (_08659_, _07212_);
  nor (_08660_, \uc8051golden_1.SP [1], \uc8051golden_1.SP [0]);
  and (_08661_, _08660_, _06738_);
  nor (_08662_, _08661_, _06398_);
  nor (_08663_, \uc8051golden_1.SP [2], \uc8051golden_1.SP [1]);
  and (_08664_, _08663_, _06398_);
  and (_08665_, _08664_, _06270_);
  nor (_08666_, _08665_, _08662_);
  nor (_08667_, _06588_, _06305_);
  nor (_08668_, _08667_, _08666_);
  not (_08669_, _07257_);
  and (_08670_, _07775_, _08669_);
  and (_08671_, _07257_, _06372_);
  not (_08672_, _08671_);
  nand (_08673_, _08672_, _08667_);
  nor (_08674_, _08673_, _08670_);
  nor (_08675_, _08674_, _08668_);
  nor (_08676_, _08660_, _06738_);
  nor (_08677_, _08676_, _08661_);
  nor (_08678_, _08677_, _08667_);
  not (_08679_, _08678_);
  nand (_08680_, _07623_, _08669_);
  and (_08681_, _07257_, _06693_);
  not (_08682_, _08681_);
  and (_08683_, _08682_, _08667_);
  nand (_08684_, _08683_, _08680_);
  and (_08685_, _08684_, _08679_);
  nor (_08686_, _07257_, _07196_);
  nor (_08687_, _08669_, _06228_);
  or (_08688_, _08687_, _08686_);
  nand (_08689_, _08688_, _08667_);
  nor (_08690_, _08667_, _06273_);
  not (_08691_, _08690_);
  and (_08692_, _08691_, _08689_);
  or (_08693_, _07473_, _07257_);
  and (_08694_, _07257_, _06840_);
  not (_08695_, _08694_);
  and (_08696_, _08695_, _08667_);
  nand (_08697_, _08696_, _08693_);
  nor (_08698_, _08667_, \uc8051golden_1.SP [0]);
  not (_08699_, _08698_);
  and (_08700_, _08699_, _08697_);
  or (_08701_, _08700_, _08025_);
  nand (_08702_, _08700_, \uc8051golden_1.IRAM[0] [7]);
  nand (_08703_, _08702_, _08701_);
  and (_08704_, _08703_, _08692_);
  not (_08705_, _08700_);
  or (_08706_, _08705_, \uc8051golden_1.IRAM[2] [7]);
  nor (_08707_, _08700_, \uc8051golden_1.IRAM[3] [7]);
  nor (_08708_, _08707_, _08692_);
  and (_08709_, _08708_, _08706_);
  nor (_08710_, _08709_, _08704_);
  nand (_08711_, _08710_, _08685_);
  not (_08712_, _08685_);
  or (_08713_, _08700_, \uc8051golden_1.IRAM[5] [7]);
  or (_08714_, _08705_, \uc8051golden_1.IRAM[4] [7]);
  and (_08715_, _08714_, _08692_);
  and (_08716_, _08715_, _08713_);
  or (_08717_, _08705_, \uc8051golden_1.IRAM[6] [7]);
  nor (_08718_, _08700_, \uc8051golden_1.IRAM[7] [7]);
  nor (_08719_, _08718_, _08692_);
  and (_08720_, _08719_, _08717_);
  nor (_08721_, _08720_, _08716_);
  nand (_08722_, _08721_, _08712_);
  nand (_08723_, _08722_, _08711_);
  nand (_08724_, _08723_, _08675_);
  not (_08725_, _08675_);
  or (_08726_, _08705_, \uc8051golden_1.IRAM[8] [7]);
  or (_08727_, _08700_, \uc8051golden_1.IRAM[9] [7]);
  nand (_08728_, _08727_, _08726_);
  nand (_08729_, _08728_, _08692_);
  not (_08730_, _08692_);
  or (_08731_, _08705_, \uc8051golden_1.IRAM[10] [7]);
  or (_08732_, _08700_, \uc8051golden_1.IRAM[11] [7]);
  nand (_08733_, _08732_, _08731_);
  nand (_08734_, _08733_, _08730_);
  nand (_08735_, _08734_, _08729_);
  nand (_08736_, _08735_, _08685_);
  or (_08737_, _08705_, \uc8051golden_1.IRAM[12] [7]);
  or (_08738_, _08700_, \uc8051golden_1.IRAM[13] [7]);
  nand (_08739_, _08738_, _08737_);
  nand (_08740_, _08739_, _08692_);
  nand (_08741_, _08700_, \uc8051golden_1.IRAM[14] [7]);
  or (_08742_, _08700_, _05652_);
  and (_08743_, _08742_, _08741_);
  nand (_08744_, _08743_, _08730_);
  nand (_08745_, _08744_, _08740_);
  nand (_08746_, _08745_, _08712_);
  nand (_08747_, _08746_, _08736_);
  nand (_08748_, _08747_, _08725_);
  and (_08749_, _08748_, _08724_);
  or (_08750_, _08749_, _08659_);
  and (_08751_, _08750_, _08658_);
  or (_08752_, _08751_, _07211_);
  not (_08753_, _07211_);
  and (_08754_, _08344_, _08255_);
  or (_08755_, _08521_, _08477_);
  or (_08756_, _08755_, _08433_);
  nor (_08757_, _08756_, _08389_);
  and (_08758_, _08757_, _08754_);
  and (_08759_, _08758_, _08161_);
  or (_08760_, _08759_, _08073_);
  nand (_08761_, _08759_, _08073_);
  and (_08762_, _08761_, _08760_);
  or (_08763_, _08762_, _08753_);
  and (_08764_, _08763_, _08752_);
  or (_08765_, _08764_, _07218_);
  and (_08766_, _08765_, _08642_);
  or (_08767_, _08766_, _07351_);
  nor (_08768_, _08649_, _05997_);
  nor (_08769_, _08768_, _07222_);
  and (_08770_, _08769_, _08767_);
  and (_08771_, _08548_, _07222_);
  or (_08772_, _08771_, _07239_);
  or (_08773_, _08772_, _08770_);
  and (_08774_, _08773_, _08640_);
  or (_08775_, _08774_, _06419_);
  nand (_08776_, _08072_, _06419_);
  and (_08777_, _08776_, _07423_);
  and (_08778_, _08777_, _08775_);
  or (_08779_, _08778_, _08637_);
  and (_08780_, _08779_, _05994_);
  not (_08781_, _08649_);
  or (_08782_, _08781_, _05994_);
  nand (_08783_, _08782_, _06383_);
  or (_08784_, _08783_, _08780_);
  nand (_08785_, _08072_, _06384_);
  and (_08786_, _08785_, _08784_);
  or (_08787_, _08786_, _07257_);
  and (_08788_, _08749_, _06309_);
  nand (_08789_, _08024_, _07257_);
  or (_08790_, _08789_, _08788_);
  and (_08791_, _08790_, _07777_);
  and (_08792_, _08791_, _08787_);
  and (_08793_, _08001_, \uc8051golden_1.PSW [7]);
  or (_08794_, _08793_, _08639_);
  and (_08795_, _08794_, _07256_);
  or (_08796_, _08795_, _06017_);
  or (_08797_, _08796_, _08792_);
  nor (_08798_, _06293_, _06194_);
  and (_08799_, _08781_, _06017_);
  nor (_08800_, _08799_, _08798_);
  and (_08801_, _08800_, _08797_);
  nor (_08802_, _06282_, _06194_);
  not (_08803_, _08798_);
  nor (_08804_, _08803_, _08070_);
  or (_08805_, _08804_, _08802_);
  or (_08806_, _08805_, _08801_);
  nor (_08807_, _06194_, _06279_);
  not (_08808_, _08807_);
  not (_08809_, _08802_);
  or (_08810_, _08809_, _08749_);
  and (_08811_, _08810_, _08808_);
  and (_08812_, _08811_, _08806_);
  not (_08813_, _08590_);
  nor (_08814_, _08813_, _08070_);
  not (_08815_, _06562_);
  and (_08816_, _06736_, _08815_);
  not (_08817_, _06943_);
  and (_08818_, _07090_, _08817_);
  and (_08819_, _08818_, _08816_);
  and (_08820_, _06539_, _05012_);
  and (_08821_, _06508_, _05000_);
  nor (_08822_, _08821_, _08820_);
  and (_08823_, _06526_, _04991_);
  and (_08824_, _06534_, _05002_);
  nor (_08825_, _08824_, _08823_);
  and (_08826_, _08825_, _08822_);
  and (_08827_, _06528_, _04987_);
  and (_08828_, _06512_, _04998_);
  nor (_08829_, _08828_, _08827_);
  and (_08830_, _06555_, _05014_);
  and (_08831_, _06532_, _04976_);
  nor (_08832_, _08831_, _08830_);
  and (_08833_, _08832_, _08829_);
  and (_08834_, _08833_, _08826_);
  and (_08835_, _06552_, _04983_);
  and (_08836_, _06557_, _04981_);
  nor (_08837_, _08836_, _08835_);
  and (_08838_, _06544_, _05010_);
  and (_08839_, _06550_, _04989_);
  nor (_08840_, _08839_, _08838_);
  and (_08841_, _08840_, _08837_);
  and (_08842_, _06541_, _04996_);
  and (_08843_, _06546_, _05006_);
  nor (_08844_, _08843_, _08842_);
  and (_08845_, _06516_, _05008_);
  and (_08846_, _06520_, _04978_);
  nor (_08847_, _08846_, _08845_);
  and (_08848_, _08847_, _08844_);
  and (_08849_, _08848_, _08841_);
  and (_08850_, _08849_, _08834_);
  and (_08851_, _08850_, _08813_);
  and (_08852_, _06526_, _04897_);
  and (_08853_, _06534_, _04893_);
  nor (_08854_, _08853_, _08852_);
  and (_08855_, _06520_, _04910_);
  and (_08856_, _06557_, _04913_);
  nor (_08857_, _08856_, _08855_);
  and (_08858_, _08857_, _08854_);
  and (_08859_, _06550_, _04886_);
  and (_08860_, _06546_, _04922_);
  nor (_08861_, _08860_, _08859_);
  and (_08862_, _06541_, _04884_);
  and (_08863_, _06512_, _04888_);
  nor (_08864_, _08863_, _08862_);
  and (_08865_, _08864_, _08861_);
  and (_08866_, _08865_, _08858_);
  and (_08867_, _06539_, _04915_);
  and (_08868_, _06516_, _04904_);
  nor (_08869_, _08868_, _08867_);
  and (_08870_, _06555_, _04917_);
  and (_08871_, _06532_, _04908_);
  nor (_08872_, _08871_, _08870_);
  and (_08873_, _08872_, _08869_);
  and (_08874_, _06528_, _04924_);
  and (_08875_, _06552_, _04899_);
  nor (_08876_, _08875_, _08874_);
  and (_08877_, _06544_, _04902_);
  and (_08878_, _06508_, _04891_);
  nor (_08879_, _08878_, _08877_);
  and (_08880_, _08879_, _08876_);
  and (_08881_, _08880_, _08873_);
  and (_08882_, _08881_, _08866_);
  not (_08883_, _08882_);
  and (_08884_, _06539_, _04966_);
  and (_08885_, _06552_, _04937_);
  nor (_08886_, _08885_, _08884_);
  and (_08887_, _06544_, _04964_);
  and (_08888_, _06528_, _04952_);
  nor (_08889_, _08888_, _08887_);
  and (_08890_, _08889_, _08886_);
  and (_08892_, _06532_, _04940_);
  and (_08893_, _06520_, _04935_);
  nor (_08894_, _08893_, _08892_);
  and (_08895_, _06526_, _04954_);
  and (_08896_, _06555_, _04968_);
  nor (_08897_, _08896_, _08895_);
  and (_08898_, _08897_, _08894_);
  and (_08899_, _08898_, _08890_);
  and (_08900_, _06541_, _04950_);
  and (_08901_, _06516_, _04962_);
  nor (_08903_, _08901_, _08900_);
  and (_08904_, _06546_, _04960_);
  and (_08905_, _06512_, _04930_);
  nor (_08906_, _08905_, _08904_);
  and (_08907_, _08906_, _08903_);
  and (_08908_, _06550_, _04956_);
  and (_08909_, _06557_, _04942_);
  nor (_08910_, _08909_, _08908_);
  and (_08911_, _06508_, _04932_);
  and (_08912_, _06534_, _04946_);
  nor (_08914_, _08912_, _08911_);
  and (_08915_, _08914_, _08910_);
  and (_08916_, _08915_, _08907_);
  and (_08917_, _08916_, _08899_);
  and (_08918_, _08917_, _08883_);
  and (_08919_, _08918_, _08851_);
  and (_08920_, _08919_, _08819_);
  and (_08921_, _08920_, \uc8051golden_1.SBUF [7]);
  and (_08922_, _07090_, _06943_);
  and (_08923_, _06736_, _06562_);
  and (_08925_, _08923_, _08922_);
  nor (_08926_, _08850_, _08590_);
  and (_08927_, _08926_, _08925_);
  and (_08928_, _08927_, _08918_);
  and (_08929_, _08928_, \uc8051golden_1.PSW [7]);
  or (_08930_, _08929_, _08921_);
  and (_08931_, _08917_, _08882_);
  and (_08932_, _08931_, _08851_);
  and (_08933_, _08922_, _08816_);
  and (_08934_, _08933_, _08932_);
  and (_08936_, _08934_, \uc8051golden_1.TCON [7]);
  not (_08937_, _07090_);
  and (_08938_, _08937_, _06943_);
  and (_08939_, _08938_, _08816_);
  and (_08940_, _08939_, _08932_);
  and (_08941_, _08940_, \uc8051golden_1.TL0 [7]);
  or (_08942_, _08941_, _08936_);
  or (_08943_, _08942_, _08930_);
  and (_08944_, _08932_, _08819_);
  and (_08945_, _08944_, \uc8051golden_1.TMOD [7]);
  and (_08947_, _08933_, _08919_);
  and (_08948_, _08947_, \uc8051golden_1.SCON [7]);
  or (_08949_, _08948_, _08945_);
  and (_08950_, _08925_, _08919_);
  and (_08951_, _08950_, \uc8051golden_1.P1 [7]);
  nor (_08952_, _08917_, _08882_);
  and (_08953_, _08952_, _08927_);
  and (_08954_, _08953_, \uc8051golden_1.B [7]);
  or (_08955_, _08954_, _08951_);
  or (_08956_, _08955_, _08949_);
  not (_08958_, _08917_);
  and (_08959_, _08958_, _08882_);
  and (_08960_, _08959_, _08851_);
  and (_08961_, _08960_, _08925_);
  and (_08962_, _08961_, \uc8051golden_1.P2 [7]);
  and (_08963_, _08952_, _08851_);
  and (_08964_, _08963_, _08933_);
  and (_08965_, _08964_, \uc8051golden_1.IP [7]);
  or (_08966_, _08965_, _08962_);
  and (_08967_, _08960_, _08933_);
  and (_08968_, _08967_, \uc8051golden_1.IE [7]);
  and (_08969_, _08963_, _08925_);
  and (_08970_, _08969_, \uc8051golden_1.P3 [7]);
  or (_08971_, _08970_, _08968_);
  or (_08972_, _08971_, _08966_);
  and (_08973_, _08932_, _08925_);
  and (_08974_, _08973_, \uc8051golden_1.P0 [7]);
  and (_08975_, _08959_, _08927_);
  and (_08976_, _08975_, \uc8051golden_1.ACC [7]);
  or (_08977_, _08976_, _08974_);
  or (_08978_, _08977_, _08972_);
  or (_08979_, _08978_, _08956_);
  or (_08980_, _08979_, _08943_);
  nor (_08981_, _06736_, _06562_);
  and (_08982_, _08981_, _08932_);
  and (_08983_, _08982_, _08818_);
  and (_08984_, _08983_, \uc8051golden_1.TH1 [7]);
  nor (_08985_, _07090_, _06943_);
  and (_08986_, _08985_, _08932_);
  and (_08987_, _08986_, _08816_);
  and (_08988_, _08987_, \uc8051golden_1.TL1 [7]);
  and (_08989_, _08932_, _08923_);
  and (_08990_, _08989_, _08818_);
  and (_08991_, _08990_, \uc8051golden_1.SP [7]);
  or (_08992_, _08991_, _08988_);
  or (_08993_, _08992_, _08984_);
  not (_08994_, _06736_);
  and (_08995_, _08994_, _06562_);
  and (_08996_, _08995_, _08986_);
  and (_08997_, _08996_, \uc8051golden_1.PCON [7]);
  and (_08998_, _08986_, _08923_);
  and (_08999_, _08998_, \uc8051golden_1.DPH [7]);
  or (_09000_, _08999_, _08997_);
  and (_09001_, _08989_, _08938_);
  and (_09002_, _09001_, \uc8051golden_1.DPL [7]);
  and (_09003_, _08982_, _08922_);
  and (_09004_, _09003_, \uc8051golden_1.TH0 [7]);
  or (_09005_, _09004_, _09002_);
  or (_09006_, _09005_, _09000_);
  or (_09007_, _09006_, _08993_);
  or (_09008_, _09007_, _08980_);
  or (_09009_, _09008_, _08814_);
  and (_09010_, _09009_, _08807_);
  and (_09011_, _05942_, _05805_);
  nor (_09012_, _09011_, _07268_);
  not (_09013_, _09012_);
  or (_09014_, _09013_, _09010_);
  or (_09015_, _09014_, _08812_);
  nor (_09016_, _09012_, _06194_);
  nor (_09017_, _09016_, _06277_);
  and (_09018_, _09017_, _09015_);
  and (_09019_, _08813_, _06277_);
  or (_09020_, _09019_, _05943_);
  or (_09021_, _09020_, _09018_);
  and (_09022_, _08781_, _05943_);
  nor (_09023_, _09022_, _07283_);
  and (_09024_, _09023_, _09021_);
  not (_09025_, _08591_);
  nand (_09026_, _08590_, _08072_);
  and (_09027_, _09026_, _09025_);
  nor (_09028_, _09027_, _07285_);
  nor (_09029_, _09028_, _07286_);
  or (_09030_, _09029_, _09024_);
  not (_09031_, _07285_);
  nor (_09032_, _08072_, _08651_);
  and (_09033_, _08072_, _08651_);
  nor (_09034_, _09033_, _09032_);
  or (_09035_, _09034_, _09031_);
  and (_09036_, _09035_, _07281_);
  and (_09037_, _09036_, _09030_);
  or (_09038_, _09037_, _08592_);
  and (_09039_, _09038_, _07278_);
  and (_09040_, _09032_, _07277_);
  or (_09041_, _09040_, _05956_);
  or (_09042_, _09041_, _09039_);
  not (_09043_, _06479_);
  nor (_09044_, _09043_, _06194_);
  and (_09045_, _08781_, _05956_);
  nor (_09046_, _09045_, _09044_);
  and (_09047_, _09046_, _09042_);
  not (_09048_, _06572_);
  nor (_09049_, _09048_, _06194_);
  and (_09050_, _09026_, _09044_);
  or (_09051_, _09050_, _09049_);
  or (_09052_, _09051_, _09047_);
  nand (_09053_, _09033_, _09049_);
  and (_09054_, _09053_, _05967_);
  and (_09055_, _09054_, _09052_);
  and (_09056_, _06955_, _05968_);
  not (_09057_, _09056_);
  and (_09058_, _07103_, _05968_);
  nor (_09059_, _09058_, _08544_);
  and (_09060_, _09059_, _09057_);
  and (_09061_, _09060_, _08543_);
  nand (_09062_, _08649_, _05966_);
  nand (_09063_, _09062_, _09061_);
  or (_09064_, _09063_, _09055_);
  and (_09065_, _09064_, _08559_);
  and (_09066_, _06452_, _05968_);
  and (_09067_, _06466_, _05968_);
  nor (_09068_, _09067_, _09066_);
  not (_09069_, _09068_);
  and (_09070_, _08557_, _09069_);
  or (_09071_, _09070_, _07305_);
  or (_09072_, _09071_, _09065_);
  not (_09073_, _07304_);
  not (_09074_, _07305_);
  nand (_09075_, _08748_, _08724_);
  or (_09076_, _08700_, \uc8051golden_1.IRAM[1] [6]);
  or (_09077_, _08705_, \uc8051golden_1.IRAM[0] [6]);
  and (_09078_, _09077_, _08692_);
  and (_09079_, _09078_, _09076_);
  or (_09080_, _08705_, \uc8051golden_1.IRAM[2] [6]);
  nor (_09081_, _08700_, \uc8051golden_1.IRAM[3] [6]);
  nor (_09082_, _09081_, _08692_);
  and (_09083_, _09082_, _09080_);
  nor (_09084_, _09083_, _09079_);
  nand (_09085_, _09084_, _08685_);
  or (_09086_, _08700_, \uc8051golden_1.IRAM[5] [6]);
  or (_09087_, _08705_, \uc8051golden_1.IRAM[4] [6]);
  and (_09088_, _09087_, _08692_);
  and (_09089_, _09088_, _09086_);
  or (_09090_, _08705_, \uc8051golden_1.IRAM[6] [6]);
  nor (_09091_, _08700_, \uc8051golden_1.IRAM[7] [6]);
  nor (_09092_, _09091_, _08692_);
  and (_09093_, _09092_, _09090_);
  nor (_09094_, _09093_, _09089_);
  nand (_09095_, _09094_, _08712_);
  nand (_09096_, _09095_, _09085_);
  nand (_09097_, _09096_, _08675_);
  or (_09098_, _08705_, \uc8051golden_1.IRAM[8] [6]);
  or (_09099_, _08700_, \uc8051golden_1.IRAM[9] [6]);
  nand (_09100_, _09099_, _09098_);
  nand (_09101_, _09100_, _08692_);
  or (_09102_, _08705_, \uc8051golden_1.IRAM[10] [6]);
  or (_09103_, _08700_, \uc8051golden_1.IRAM[11] [6]);
  nand (_09104_, _09103_, _09102_);
  nand (_09105_, _09104_, _08730_);
  nand (_09106_, _09105_, _09101_);
  nand (_09107_, _09106_, _08685_);
  or (_09108_, _08705_, \uc8051golden_1.IRAM[12] [6]);
  or (_09109_, _08700_, \uc8051golden_1.IRAM[13] [6]);
  nand (_09110_, _09109_, _09108_);
  nand (_09111_, _09110_, _08692_);
  or (_09112_, _08705_, \uc8051golden_1.IRAM[14] [6]);
  or (_09113_, _08700_, \uc8051golden_1.IRAM[15] [6]);
  nand (_09114_, _09113_, _09112_);
  nand (_09115_, _09114_, _08730_);
  nand (_09116_, _09115_, _09111_);
  nand (_09117_, _09116_, _08712_);
  nand (_09118_, _09117_, _09107_);
  nand (_09119_, _09118_, _08725_);
  nand (_09120_, _09119_, _09097_);
  or (_09121_, _08700_, \uc8051golden_1.IRAM[1] [5]);
  or (_09122_, _08705_, \uc8051golden_1.IRAM[0] [5]);
  and (_09123_, _09122_, _08692_);
  and (_09124_, _09123_, _09121_);
  or (_09125_, _08705_, \uc8051golden_1.IRAM[2] [5]);
  nor (_09126_, _08700_, \uc8051golden_1.IRAM[3] [5]);
  nor (_09127_, _09126_, _08692_);
  and (_09128_, _09127_, _09125_);
  nor (_09129_, _09128_, _09124_);
  nand (_09130_, _09129_, _08685_);
  or (_09131_, _08700_, \uc8051golden_1.IRAM[5] [5]);
  or (_09132_, _08705_, \uc8051golden_1.IRAM[4] [5]);
  and (_09133_, _09132_, _08692_);
  and (_09134_, _09133_, _09131_);
  or (_09135_, _08705_, \uc8051golden_1.IRAM[6] [5]);
  nor (_09136_, _08700_, \uc8051golden_1.IRAM[7] [5]);
  nor (_09137_, _09136_, _08692_);
  and (_09138_, _09137_, _09135_);
  nor (_09139_, _09138_, _09134_);
  nand (_09140_, _09139_, _08712_);
  nand (_09141_, _09140_, _09130_);
  nand (_09142_, _09141_, _08675_);
  or (_09143_, _08705_, \uc8051golden_1.IRAM[8] [5]);
  or (_09144_, _08700_, \uc8051golden_1.IRAM[9] [5]);
  nand (_09145_, _09144_, _09143_);
  nand (_09146_, _09145_, _08692_);
  or (_09147_, _08705_, \uc8051golden_1.IRAM[10] [5]);
  or (_09148_, _08700_, \uc8051golden_1.IRAM[11] [5]);
  nand (_09149_, _09148_, _09147_);
  nand (_09150_, _09149_, _08730_);
  nand (_09151_, _09150_, _09146_);
  nand (_09152_, _09151_, _08685_);
  or (_09153_, _08705_, \uc8051golden_1.IRAM[12] [5]);
  or (_09154_, _08700_, \uc8051golden_1.IRAM[13] [5]);
  nand (_09155_, _09154_, _09153_);
  nand (_09156_, _09155_, _08692_);
  or (_09157_, _08705_, \uc8051golden_1.IRAM[14] [5]);
  or (_09158_, _08700_, \uc8051golden_1.IRAM[15] [5]);
  nand (_09159_, _09158_, _09157_);
  nand (_09160_, _09159_, _08730_);
  nand (_09161_, _09160_, _09156_);
  nand (_09162_, _09161_, _08712_);
  nand (_09163_, _09162_, _09152_);
  nand (_09164_, _09163_, _08725_);
  nand (_09165_, _09164_, _09142_);
  or (_09166_, _08700_, \uc8051golden_1.IRAM[1] [4]);
  or (_09167_, _08705_, \uc8051golden_1.IRAM[0] [4]);
  and (_09168_, _09167_, _08692_);
  and (_09169_, _09168_, _09166_);
  or (_09170_, _08705_, \uc8051golden_1.IRAM[2] [4]);
  nor (_09171_, _08700_, \uc8051golden_1.IRAM[3] [4]);
  nor (_09172_, _09171_, _08692_);
  and (_09173_, _09172_, _09170_);
  nor (_09174_, _09173_, _09169_);
  nand (_09175_, _09174_, _08685_);
  or (_09176_, _08700_, \uc8051golden_1.IRAM[5] [4]);
  or (_09177_, _08705_, \uc8051golden_1.IRAM[4] [4]);
  and (_09178_, _09177_, _08692_);
  and (_09179_, _09178_, _09176_);
  or (_09180_, _08705_, \uc8051golden_1.IRAM[6] [4]);
  nor (_09181_, _08700_, \uc8051golden_1.IRAM[7] [4]);
  nor (_09182_, _09181_, _08692_);
  and (_09183_, _09182_, _09180_);
  nor (_09184_, _09183_, _09179_);
  nand (_09185_, _09184_, _08712_);
  nand (_09186_, _09185_, _09175_);
  nand (_09187_, _09186_, _08675_);
  or (_09188_, _08705_, \uc8051golden_1.IRAM[8] [4]);
  or (_09189_, _08700_, \uc8051golden_1.IRAM[9] [4]);
  nand (_09190_, _09189_, _09188_);
  nand (_09191_, _09190_, _08692_);
  or (_09192_, _08705_, \uc8051golden_1.IRAM[10] [4]);
  or (_09193_, _08700_, \uc8051golden_1.IRAM[11] [4]);
  nand (_09194_, _09193_, _09192_);
  nand (_09195_, _09194_, _08730_);
  nand (_09196_, _09195_, _09191_);
  nand (_09197_, _09196_, _08685_);
  or (_09198_, _08705_, \uc8051golden_1.IRAM[12] [4]);
  or (_09199_, _08700_, \uc8051golden_1.IRAM[13] [4]);
  nand (_09200_, _09199_, _09198_);
  nand (_09201_, _09200_, _08692_);
  or (_09202_, _08705_, \uc8051golden_1.IRAM[14] [4]);
  or (_09203_, _08700_, \uc8051golden_1.IRAM[15] [4]);
  nand (_09204_, _09203_, _09202_);
  nand (_09205_, _09204_, _08730_);
  nand (_09206_, _09205_, _09201_);
  nand (_09207_, _09206_, _08712_);
  nand (_09208_, _09207_, _09197_);
  nand (_09209_, _09208_, _08725_);
  nand (_09210_, _09209_, _09187_);
  or (_09211_, _08700_, \uc8051golden_1.IRAM[1] [3]);
  or (_09212_, _08705_, \uc8051golden_1.IRAM[0] [3]);
  and (_09213_, _09212_, _08692_);
  and (_09214_, _09213_, _09211_);
  or (_09215_, _08705_, \uc8051golden_1.IRAM[2] [3]);
  nor (_09216_, _08700_, \uc8051golden_1.IRAM[3] [3]);
  nor (_09217_, _09216_, _08692_);
  and (_09218_, _09217_, _09215_);
  nor (_09219_, _09218_, _09214_);
  nand (_09220_, _09219_, _08685_);
  or (_09221_, _08700_, \uc8051golden_1.IRAM[5] [3]);
  or (_09222_, _08705_, \uc8051golden_1.IRAM[4] [3]);
  and (_09223_, _09222_, _08692_);
  and (_09224_, _09223_, _09221_);
  or (_09225_, _08705_, \uc8051golden_1.IRAM[6] [3]);
  nor (_09226_, _08700_, \uc8051golden_1.IRAM[7] [3]);
  nor (_09227_, _09226_, _08692_);
  and (_09228_, _09227_, _09225_);
  nor (_09229_, _09228_, _09224_);
  nand (_09230_, _09229_, _08712_);
  nand (_09231_, _09230_, _09220_);
  nand (_09232_, _09231_, _08675_);
  or (_09233_, _08705_, \uc8051golden_1.IRAM[8] [3]);
  or (_09234_, _08700_, \uc8051golden_1.IRAM[9] [3]);
  nand (_09235_, _09234_, _09233_);
  nand (_09236_, _09235_, _08692_);
  or (_09237_, _08705_, \uc8051golden_1.IRAM[10] [3]);
  or (_09238_, _08700_, \uc8051golden_1.IRAM[11] [3]);
  nand (_09239_, _09238_, _09237_);
  nand (_09240_, _09239_, _08730_);
  nand (_09241_, _09240_, _09236_);
  nand (_09242_, _09241_, _08685_);
  nand (_09243_, _08700_, _07767_);
  or (_09244_, _08700_, \uc8051golden_1.IRAM[13] [3]);
  nand (_09245_, _09244_, _09243_);
  nand (_09246_, _09245_, _08692_);
  nand (_09247_, _08700_, _07757_);
  or (_09248_, _08700_, \uc8051golden_1.IRAM[15] [3]);
  nand (_09249_, _09248_, _09247_);
  nand (_09250_, _09249_, _08730_);
  nand (_09251_, _09250_, _09246_);
  nand (_09252_, _09251_, _08712_);
  nand (_09253_, _09252_, _09242_);
  nand (_09254_, _09253_, _08725_);
  nand (_09255_, _09254_, _09232_);
  or (_09256_, _08700_, \uc8051golden_1.IRAM[1] [2]);
  or (_09257_, _08705_, \uc8051golden_1.IRAM[0] [2]);
  and (_09258_, _09257_, _08692_);
  and (_09259_, _09258_, _09256_);
  or (_09260_, _08705_, \uc8051golden_1.IRAM[2] [2]);
  nor (_09261_, _08700_, \uc8051golden_1.IRAM[3] [2]);
  nor (_09262_, _09261_, _08692_);
  and (_09263_, _09262_, _09260_);
  nor (_09264_, _09263_, _09259_);
  nand (_09265_, _09264_, _08685_);
  or (_09266_, _08700_, \uc8051golden_1.IRAM[5] [2]);
  nand (_09267_, _08700_, _07591_);
  and (_09268_, _09267_, _08692_);
  and (_09269_, _09268_, _09266_);
  or (_09270_, _08705_, \uc8051golden_1.IRAM[6] [2]);
  nor (_09271_, _08700_, \uc8051golden_1.IRAM[7] [2]);
  nor (_09272_, _09271_, _08692_);
  and (_09273_, _09272_, _09270_);
  nor (_09274_, _09273_, _09269_);
  nand (_09275_, _09274_, _08712_);
  nand (_09276_, _09275_, _09265_);
  nand (_09277_, _09276_, _08675_);
  or (_09278_, _08705_, \uc8051golden_1.IRAM[8] [2]);
  or (_09279_, _08700_, \uc8051golden_1.IRAM[9] [2]);
  nand (_09280_, _09279_, _09278_);
  nand (_09281_, _09280_, _08692_);
  or (_09282_, _08705_, \uc8051golden_1.IRAM[10] [2]);
  or (_09283_, _08700_, \uc8051golden_1.IRAM[11] [2]);
  nand (_09284_, _09283_, _09282_);
  nand (_09285_, _09284_, _08730_);
  nand (_09286_, _09285_, _09281_);
  nand (_09287_, _09286_, _08685_);
  or (_09288_, _08705_, \uc8051golden_1.IRAM[12] [2]);
  or (_09289_, _08700_, \uc8051golden_1.IRAM[13] [2]);
  nand (_09290_, _09289_, _09288_);
  nand (_09291_, _09290_, _08692_);
  nand (_09292_, _08700_, _07609_);
  or (_09293_, _08700_, \uc8051golden_1.IRAM[15] [2]);
  nand (_09294_, _09293_, _09292_);
  nand (_09295_, _09294_, _08730_);
  nand (_09296_, _09295_, _09291_);
  nand (_09297_, _09296_, _08712_);
  nand (_09298_, _09297_, _09287_);
  nand (_09299_, _09298_, _08725_);
  nand (_09300_, _09299_, _09277_);
  and (_09301_, _08700_, \uc8051golden_1.IRAM[0] [1]);
  nor (_09302_, _08700_, _06806_);
  or (_09303_, _09302_, _09301_);
  and (_09304_, _09303_, _08692_);
  nand (_09305_, _08700_, _07145_);
  nor (_09306_, _08700_, \uc8051golden_1.IRAM[3] [1]);
  nor (_09307_, _09306_, _08692_);
  and (_09308_, _09307_, _09305_);
  nor (_09309_, _09308_, _09304_);
  nand (_09310_, _09309_, _08685_);
  or (_09311_, _08700_, \uc8051golden_1.IRAM[5] [1]);
  nand (_09312_, _08700_, _07164_);
  and (_09313_, _09312_, _08692_);
  and (_09314_, _09313_, _09311_);
  nand (_09315_, _08700_, _07156_);
  nor (_09316_, _08700_, \uc8051golden_1.IRAM[7] [1]);
  nor (_09317_, _09316_, _08692_);
  and (_09318_, _09317_, _09315_);
  nor (_09319_, _09318_, _09314_);
  nand (_09320_, _09319_, _08712_);
  nand (_09321_, _09320_, _09310_);
  nand (_09322_, _09321_, _08675_);
  or (_09323_, _08705_, \uc8051golden_1.IRAM[8] [1]);
  or (_09324_, _08700_, \uc8051golden_1.IRAM[9] [1]);
  nand (_09325_, _09324_, _09323_);
  nand (_09326_, _09325_, _08692_);
  or (_09327_, _08705_, \uc8051golden_1.IRAM[10] [1]);
  or (_09328_, _08700_, \uc8051golden_1.IRAM[11] [1]);
  nand (_09329_, _09328_, _09327_);
  nand (_09330_, _09329_, _08730_);
  nand (_09331_, _09330_, _09326_);
  nand (_09332_, _09331_, _08685_);
  nand (_09333_, _08700_, \uc8051golden_1.IRAM[12] [1]);
  or (_09334_, _08700_, _07187_);
  and (_09335_, _09334_, _09333_);
  nand (_09336_, _09335_, _08692_);
  or (_09337_, _08705_, \uc8051golden_1.IRAM[14] [1]);
  or (_09338_, _08700_, \uc8051golden_1.IRAM[15] [1]);
  nand (_09339_, _09338_, _09337_);
  nand (_09340_, _09339_, _08730_);
  nand (_09341_, _09340_, _09336_);
  nand (_09342_, _09341_, _08712_);
  nand (_09343_, _09342_, _09332_);
  nand (_09344_, _09343_, _08725_);
  nand (_09345_, _09344_, _09322_);
  and (_09346_, _08700_, \uc8051golden_1.IRAM[0] [0]);
  nor (_09347_, _08700_, _07424_);
  or (_09348_, _09347_, _09346_);
  and (_09349_, _09348_, _08692_);
  nand (_09350_, _08700_, _07429_);
  nor (_09351_, _08700_, \uc8051golden_1.IRAM[3] [0]);
  nor (_09352_, _09351_, _08692_);
  and (_09353_, _09352_, _09350_);
  nor (_09354_, _09353_, _09349_);
  nand (_09355_, _09354_, _08685_);
  or (_09356_, _08700_, \uc8051golden_1.IRAM[5] [0]);
  nand (_09357_, _08700_, _07441_);
  and (_09358_, _09357_, _08692_);
  and (_09359_, _09358_, _09356_);
  or (_09360_, _08705_, \uc8051golden_1.IRAM[6] [0]);
  nor (_09361_, _08700_, \uc8051golden_1.IRAM[7] [0]);
  nor (_09362_, _09361_, _08692_);
  and (_09363_, _09362_, _09360_);
  nor (_09364_, _09363_, _09359_);
  nand (_09365_, _09364_, _08712_);
  nand (_09366_, _09365_, _09355_);
  nand (_09367_, _09366_, _08675_);
  or (_09368_, _08705_, \uc8051golden_1.IRAM[8] [0]);
  or (_09369_, _08700_, \uc8051golden_1.IRAM[9] [0]);
  nand (_09370_, _09369_, _09368_);
  nand (_09371_, _09370_, _08692_);
  or (_09372_, _08705_, \uc8051golden_1.IRAM[10] [0]);
  or (_09373_, _08700_, \uc8051golden_1.IRAM[11] [0]);
  nand (_09374_, _09373_, _09372_);
  nand (_09375_, _09374_, _08730_);
  nand (_09376_, _09375_, _09371_);
  nand (_09377_, _09376_, _08685_);
  nand (_09378_, _08700_, \uc8051golden_1.IRAM[12] [0]);
  or (_09379_, _08700_, _07464_);
  and (_09380_, _09379_, _09378_);
  nand (_09381_, _09380_, _08692_);
  nand (_09382_, _08700_, \uc8051golden_1.IRAM[14] [0]);
  or (_09383_, _08700_, _07460_);
  and (_09384_, _09383_, _09382_);
  nand (_09385_, _09384_, _08730_);
  nand (_09386_, _09385_, _09381_);
  nand (_09387_, _09386_, _08712_);
  nand (_09388_, _09387_, _09377_);
  nand (_09389_, _09388_, _08725_);
  nand (_09390_, _09389_, _09367_);
  and (_09391_, _09390_, _09345_);
  and (_09392_, _09391_, _09300_);
  and (_09393_, _09392_, _09255_);
  and (_09394_, _09393_, _09210_);
  and (_09395_, _09394_, _09165_);
  and (_09396_, _09395_, _09120_);
  nor (_09397_, _09396_, _09075_);
  and (_09398_, _09396_, _09075_);
  or (_09399_, _09398_, _09397_);
  or (_09400_, _09399_, _09074_);
  and (_09401_, _09400_, _09073_);
  and (_09402_, _09401_, _09072_);
  and (_09403_, _08762_, _07304_);
  or (_09404_, _09403_, _06465_);
  or (_09405_, _09404_, _09402_);
  and (_09406_, _09405_, _08541_);
  or (_09407_, _09406_, _05969_);
  and (_09408_, _08781_, _05969_);
  nor (_09409_, _09408_, _07311_);
  and (_09410_, _09409_, _09407_);
  and (_09411_, _08639_, _07311_);
  nor (_09412_, _06291_, _07363_);
  or (_09413_, _09412_, _09411_);
  or (_09414_, _09413_, _09410_);
  and (_09415_, _06285_, _05962_);
  not (_09416_, _09415_);
  not (_09417_, _09412_);
  not (_09418_, _08118_);
  not (_09419_, _08207_);
  not (_09420_, _08301_);
  not (_09421_, _07775_);
  not (_09422_, _07623_);
  nor (_09423_, _07485_, _07196_);
  and (_09424_, _09423_, _09422_);
  and (_09425_, _09424_, _09421_);
  and (_09426_, _09425_, _09420_);
  and (_09427_, _09426_, _09419_);
  and (_09428_, _09427_, _09418_);
  or (_09429_, _09428_, _08548_);
  nand (_09430_, _09428_, _08548_);
  and (_09431_, _09430_, _09429_);
  or (_09432_, _09431_, _09417_);
  and (_09433_, _09432_, _09416_);
  and (_09434_, _09433_, _09414_);
  and (_09435_, _09431_, _09415_);
  or (_09436_, _09435_, _07320_);
  or (_09437_, _09436_, _09434_);
  not (_09438_, _06197_);
  not (_09439_, _07320_);
  and (_09440_, _09119_, _09097_);
  and (_09441_, _09164_, _09142_);
  and (_09442_, _09209_, _09187_);
  and (_09443_, _09254_, _09232_);
  and (_09444_, _09299_, _09277_);
  and (_09445_, _09344_, _09322_);
  and (_09446_, _09389_, _09367_);
  and (_09447_, _09446_, _09445_);
  and (_09448_, _09447_, _09444_);
  and (_09449_, _09448_, _09443_);
  and (_09450_, _09449_, _09442_);
  and (_09451_, _09450_, _09441_);
  and (_09452_, _09451_, _09440_);
  nor (_09453_, _09452_, _09075_);
  and (_09454_, _09452_, _09075_);
  or (_09455_, _09454_, _09453_);
  or (_09456_, _09455_, _09439_);
  and (_09457_, _09456_, _09438_);
  and (_09458_, _09457_, _09437_);
  or (_09459_, _09458_, _08531_);
  and (_09460_, _09459_, _07415_);
  or (_09461_, _09460_, _07908_);
  and (_09462_, _09461_, _07923_);
  not (_09463_, _06465_);
  and (_09464_, \uc8051golden_1.PC [9], \uc8051golden_1.PC [8]);
  and (_09465_, _09464_, \uc8051golden_1.PC [10]);
  and (_09466_, _09465_, _08647_);
  and (_09467_, _09466_, \uc8051golden_1.PC [11]);
  and (_09468_, _09467_, \uc8051golden_1.PC [12]);
  and (_09469_, _09468_, \uc8051golden_1.PC [13]);
  and (_09470_, _09469_, \uc8051golden_1.PC [14]);
  nor (_09471_, _09470_, \uc8051golden_1.PC [15]);
  and (_09472_, _08647_, \uc8051golden_1.PC [8]);
  and (_09473_, _09472_, \uc8051golden_1.PC [9]);
  and (_09474_, _09473_, \uc8051golden_1.PC [10]);
  and (_09475_, _09474_, \uc8051golden_1.PC [11]);
  and (_09476_, _09475_, \uc8051golden_1.PC [12]);
  and (_09477_, _09476_, \uc8051golden_1.PC [13]);
  and (_09478_, _09477_, \uc8051golden_1.PC [14]);
  and (_09479_, _09478_, \uc8051golden_1.PC [15]);
  nor (_09480_, _09479_, _09471_);
  and (_09481_, _09480_, _09463_);
  and (_09482_, _09465_, _08537_);
  and (_09483_, _09482_, \uc8051golden_1.PC [11]);
  and (_09484_, _09483_, \uc8051golden_1.PC [12]);
  and (_09485_, _09484_, \uc8051golden_1.PC [13]);
  and (_09486_, _09485_, \uc8051golden_1.PC [14]);
  nor (_09487_, _09486_, \uc8051golden_1.PC [15]);
  and (_09488_, _08537_, \uc8051golden_1.PC [8]);
  and (_09489_, _09488_, \uc8051golden_1.PC [9]);
  and (_09490_, _09489_, \uc8051golden_1.PC [10]);
  and (_09491_, _09490_, \uc8051golden_1.PC [11]);
  and (_09492_, _09491_, \uc8051golden_1.PC [12]);
  and (_09493_, _09492_, \uc8051golden_1.PC [13]);
  and (_09494_, _09493_, \uc8051golden_1.PC [14]);
  and (_09495_, _09494_, \uc8051golden_1.PC [15]);
  nor (_09496_, _09495_, _09487_);
  and (_09497_, _09496_, _06465_);
  or (_09498_, _09497_, _09481_);
  and (_09499_, _09498_, _07918_);
  and (_09500_, _09499_, _07921_);
  or (_40322_, _09500_, _09462_);
  not (_09501_, \uc8051golden_1.B [7]);
  nor (_09502_, _01375_, _09501_);
  nor (_09503_, _07992_, _09501_);
  not (_09504_, _07992_);
  nor (_09505_, _09504_, _08070_);
  or (_09506_, _09505_, _09503_);
  or (_09508_, _09506_, _06293_);
  nor (_09509_, _08618_, _09501_);
  and (_09510_, _08639_, _08618_);
  or (_09511_, _09510_, _09509_);
  and (_09512_, _09511_, _06393_);
  and (_09513_, _08762_, _07992_);
  or (_09514_, _09513_, _09503_);
  or (_09515_, _09514_, _07210_);
  and (_09516_, _07992_, \uc8051golden_1.ACC [7]);
  or (_09517_, _09516_, _09503_);
  and (_09518_, _09517_, _07199_);
  nor (_09519_, _07199_, _09501_);
  or (_09520_, _09519_, _06401_);
  or (_09521_, _09520_, _09518_);
  and (_09522_, _09521_, _06396_);
  and (_09523_, _09522_, _09515_);
  and (_09524_, _08635_, _08618_);
  or (_09525_, _09524_, _09509_);
  and (_09526_, _09525_, _06395_);
  or (_09527_, _09526_, _06399_);
  or (_09529_, _09527_, _09523_);
  or (_09530_, _09506_, _07221_);
  and (_09531_, _09530_, _09529_);
  or (_09532_, _09531_, _06406_);
  or (_09533_, _09517_, _06414_);
  and (_09534_, _09533_, _06844_);
  and (_09535_, _09534_, _09532_);
  or (_09536_, _09535_, _09512_);
  and (_09537_, _09536_, _07245_);
  and (_09538_, _06481_, _06381_);
  or (_09539_, _09509_, _08634_);
  and (_09540_, _09539_, _06387_);
  and (_09541_, _09540_, _09525_);
  or (_09542_, _09541_, _09538_);
  or (_09543_, _09542_, _09537_);
  not (_09544_, _09538_);
  and (_09545_, \uc8051golden_1.B [1], \uc8051golden_1.ACC [7]);
  and (_09546_, \uc8051golden_1.B [0], \uc8051golden_1.ACC [6]);
  and (_09547_, _09546_, _09545_);
  and (_09548_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [2]);
  and (_09549_, \uc8051golden_1.B [0], \uc8051golden_1.ACC [7]);
  and (_09550_, \uc8051golden_1.B [1], \uc8051golden_1.ACC [6]);
  nor (_09551_, _09550_, _09549_);
  nor (_09552_, _09551_, _09547_);
  and (_09553_, _09552_, _09548_);
  nor (_09554_, _09553_, _09547_);
  and (_09555_, \uc8051golden_1.B [2], \uc8051golden_1.ACC [7]);
  and (_09556_, _09555_, _09550_);
  and (_09557_, \uc8051golden_1.B [2], \uc8051golden_1.ACC [6]);
  nor (_09558_, _09557_, _09545_);
  nor (_09559_, _09558_, _09556_);
  not (_09560_, _09559_);
  nor (_09561_, _09560_, _09554_);
  and (_09562_, \uc8051golden_1.B [5], \uc8051golden_1.ACC [3]);
  and (_09563_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [3]);
  and (_09564_, \uc8051golden_1.ACC [4], \uc8051golden_1.B [4]);
  and (_09565_, _09564_, _09563_);
  nor (_09566_, _09564_, _09563_);
  nor (_09567_, _09566_, _09565_);
  and (_09568_, _09567_, _09562_);
  nor (_09569_, _09567_, _09562_);
  nor (_09570_, _09569_, _09568_);
  and (_09571_, _09560_, _09554_);
  nor (_09572_, _09571_, _09561_);
  and (_09573_, _09572_, _09570_);
  nor (_09574_, _09573_, _09561_);
  not (_09575_, _09550_);
  and (_09576_, _09555_, _09575_);
  and (_09577_, \uc8051golden_1.ACC [4], \uc8051golden_1.B [5]);
  and (_09578_, \uc8051golden_1.B [4], \uc8051golden_1.ACC [6]);
  and (_09579_, _09578_, _09563_);
  and (_09580_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [4]);
  and (_09581_, \uc8051golden_1.B [3], \uc8051golden_1.ACC [6]);
  nor (_09582_, _09581_, _09580_);
  nor (_09583_, _09582_, _09579_);
  and (_09584_, _09583_, _09577_);
  nor (_09585_, _09583_, _09577_);
  nor (_09586_, _09585_, _09584_);
  and (_09587_, _09586_, _09576_);
  nor (_09588_, _09586_, _09576_);
  nor (_09589_, _09588_, _09587_);
  not (_09590_, _09589_);
  nor (_09591_, _09590_, _09574_);
  and (_09592_, \uc8051golden_1.B [6], \uc8051golden_1.ACC [2]);
  and (_09593_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [7]);
  and (_09594_, _09593_, _09592_);
  nor (_09595_, _09568_, _09565_);
  and (_09596_, \uc8051golden_1.ACC [2], \uc8051golden_1.B [7]);
  and (_09597_, \uc8051golden_1.B [6], \uc8051golden_1.ACC [3]);
  and (_09598_, _09597_, _09596_);
  nor (_09599_, _09597_, _09596_);
  nor (_09600_, _09599_, _09598_);
  not (_09601_, _09600_);
  nor (_09602_, _09601_, _09595_);
  and (_09603_, _09601_, _09595_);
  nor (_09604_, _09603_, _09602_);
  and (_09605_, _09604_, _09594_);
  nor (_09606_, _09604_, _09594_);
  nor (_09607_, _09606_, _09605_);
  and (_09608_, _09590_, _09574_);
  nor (_09609_, _09608_, _09591_);
  and (_09610_, _09609_, _09607_);
  nor (_09611_, _09610_, _09591_);
  nor (_09612_, _09584_, _09579_);
  and (_09613_, \uc8051golden_1.ACC [3], \uc8051golden_1.B [7]);
  and (_09614_, \uc8051golden_1.ACC [4], \uc8051golden_1.B [6]);
  and (_09615_, _09614_, _09613_);
  nor (_09616_, _09614_, _09613_);
  nor (_09617_, _09616_, _09615_);
  not (_09618_, _09617_);
  nor (_09619_, _09618_, _09612_);
  and (_09620_, _09618_, _09612_);
  nor (_09621_, _09620_, _09619_);
  and (_09622_, _09621_, _09598_);
  nor (_09623_, _09621_, _09598_);
  nor (_09624_, _09623_, _09622_);
  nor (_09625_, _09587_, _09556_);
  and (_09626_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [5]);
  and (_09627_, \uc8051golden_1.B [3], \uc8051golden_1.ACC [7]);
  and (_09628_, _09627_, _09578_);
  nor (_09629_, _09627_, _09578_);
  nor (_09630_, _09629_, _09628_);
  and (_09631_, _09630_, _09626_);
  nor (_09632_, _09630_, _09626_);
  nor (_09633_, _09632_, _09631_);
  not (_09634_, _09633_);
  nor (_09635_, _09634_, _09625_);
  and (_09636_, _09634_, _09625_);
  nor (_09637_, _09636_, _09635_);
  and (_09638_, _09637_, _09624_);
  nor (_09639_, _09637_, _09624_);
  nor (_09640_, _09639_, _09638_);
  not (_09641_, _09640_);
  nor (_09642_, _09641_, _09611_);
  nor (_09643_, _09605_, _09602_);
  not (_09644_, _09643_);
  and (_09645_, _09641_, _09611_);
  nor (_09646_, _09645_, _09642_);
  and (_09647_, _09646_, _09644_);
  nor (_09648_, _09647_, _09642_);
  nor (_09649_, _09622_, _09619_);
  not (_09650_, _09649_);
  nor (_09651_, _09638_, _09635_);
  not (_09652_, _09651_);
  and (_09653_, \uc8051golden_1.B [5], \uc8051golden_1.ACC [7]);
  and (_09654_, _09653_, _09578_);
  and (_09655_, \uc8051golden_1.B [4], \uc8051golden_1.ACC [7]);
  and (_09656_, \uc8051golden_1.B [5], \uc8051golden_1.ACC [6]);
  nor (_09657_, _09656_, _09655_);
  nor (_09658_, _09657_, _09654_);
  nor (_09659_, _09631_, _09628_);
  and (_09660_, \uc8051golden_1.ACC [4], \uc8051golden_1.B [7]);
  and (_09661_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [6]);
  and (_09662_, _09661_, _09660_);
  nor (_09663_, _09661_, _09660_);
  nor (_09664_, _09663_, _09662_);
  not (_09665_, _09664_);
  nor (_09666_, _09665_, _09659_);
  and (_09667_, _09665_, _09659_);
  nor (_09668_, _09667_, _09666_);
  and (_09669_, _09668_, _09615_);
  nor (_09670_, _09668_, _09615_);
  nor (_09671_, _09670_, _09669_);
  and (_09672_, _09671_, _09658_);
  nor (_09673_, _09671_, _09658_);
  nor (_09674_, _09673_, _09672_);
  and (_09675_, _09674_, _09652_);
  nor (_09676_, _09674_, _09652_);
  nor (_09677_, _09676_, _09675_);
  and (_09678_, _09677_, _09650_);
  nor (_09679_, _09677_, _09650_);
  nor (_09680_, _09679_, _09678_);
  not (_09681_, _09680_);
  nor (_09682_, _09681_, _09648_);
  nor (_09683_, _09678_, _09675_);
  nor (_09684_, _09669_, _09666_);
  not (_09685_, _09684_);
  and (_09686_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [7]);
  and (_09687_, \uc8051golden_1.B [6], \uc8051golden_1.ACC [6]);
  and (_09688_, _09687_, _09686_);
  nor (_09689_, _09687_, _09686_);
  nor (_09690_, _09689_, _09688_);
  and (_09691_, _09690_, _09654_);
  nor (_09692_, _09690_, _09654_);
  nor (_09693_, _09692_, _09691_);
  and (_09694_, _09693_, _09662_);
  nor (_09695_, _09693_, _09662_);
  nor (_09696_, _09695_, _09694_);
  and (_09697_, _09696_, _09653_);
  nor (_09698_, _09696_, _09653_);
  nor (_09699_, _09698_, _09697_);
  and (_09700_, _09699_, _09672_);
  nor (_09701_, _09699_, _09672_);
  nor (_09702_, _09701_, _09700_);
  and (_09703_, _09702_, _09685_);
  nor (_09704_, _09702_, _09685_);
  nor (_09705_, _09704_, _09703_);
  not (_09706_, _09705_);
  nor (_09707_, _09706_, _09683_);
  and (_09708_, _09706_, _09683_);
  nor (_09709_, _09708_, _09707_);
  and (_09710_, _09709_, _09682_);
  nor (_09711_, _09703_, _09700_);
  nor (_09712_, _09694_, _09691_);
  not (_09713_, _09712_);
  and (_09714_, \uc8051golden_1.ACC [6], \uc8051golden_1.B [7]);
  and (_09715_, \uc8051golden_1.B [6], \uc8051golden_1.ACC [7]);
  and (_09716_, _09715_, _09714_);
  nor (_09717_, _09715_, _09714_);
  nor (_09718_, _09717_, _09716_);
  and (_09719_, _09718_, _09688_);
  nor (_09720_, _09718_, _09688_);
  nor (_09721_, _09720_, _09719_);
  and (_09722_, _09721_, _09697_);
  nor (_09723_, _09721_, _09697_);
  nor (_09724_, _09723_, _09722_);
  and (_09725_, _09724_, _09713_);
  nor (_09726_, _09724_, _09713_);
  nor (_09727_, _09726_, _09725_);
  not (_09728_, _09727_);
  nor (_09729_, _09728_, _09711_);
  and (_09730_, _09728_, _09711_);
  nor (_09731_, _09730_, _09729_);
  and (_09732_, _09731_, _09707_);
  nor (_09733_, _09731_, _09707_);
  nor (_09734_, _09733_, _09732_);
  and (_09735_, _09734_, _09710_);
  nor (_09736_, _09734_, _09710_);
  and (_09737_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [0]);
  and (_09738_, _09737_, _09550_);
  and (_09739_, \uc8051golden_1.ACC [4], \uc8051golden_1.B [2]);
  and (_09740_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [1]);
  nor (_09741_, _09740_, _09546_);
  nor (_09742_, _09741_, _09738_);
  and (_09743_, _09742_, _09739_);
  nor (_09744_, _09743_, _09738_);
  not (_09745_, _09744_);
  nor (_09746_, _09552_, _09548_);
  nor (_09747_, _09746_, _09553_);
  and (_09748_, _09747_, _09745_);
  and (_09749_, \uc8051golden_1.B [5], \uc8051golden_1.ACC [2]);
  and (_09750_, \uc8051golden_1.ACC [4], \uc8051golden_1.B [3]);
  and (_09751_, \uc8051golden_1.B [4], \uc8051golden_1.ACC [3]);
  and (_09752_, _09751_, _09750_);
  nor (_09753_, _09751_, _09750_);
  nor (_09754_, _09753_, _09752_);
  and (_09755_, _09754_, _09749_);
  nor (_09756_, _09754_, _09749_);
  nor (_09757_, _09756_, _09755_);
  nor (_09758_, _09747_, _09745_);
  nor (_09759_, _09758_, _09748_);
  and (_09760_, _09759_, _09757_);
  nor (_09761_, _09760_, _09748_);
  nor (_09762_, _09572_, _09570_);
  nor (_09763_, _09762_, _09573_);
  not (_09764_, _09763_);
  nor (_09765_, _09764_, _09761_);
  and (_09766_, \uc8051golden_1.B [6], \uc8051golden_1.ACC [0]);
  and (_09767_, _09766_, _09593_);
  nor (_09768_, _09755_, _09752_);
  nor (_09769_, _09593_, _09592_);
  nor (_09770_, _09769_, _09594_);
  not (_09771_, _09770_);
  nor (_09772_, _09771_, _09768_);
  and (_09773_, _09771_, _09768_);
  nor (_09774_, _09773_, _09772_);
  and (_09775_, _09774_, _09767_);
  nor (_09776_, _09774_, _09767_);
  nor (_09777_, _09776_, _09775_);
  and (_09778_, _09764_, _09761_);
  nor (_09779_, _09778_, _09765_);
  and (_09780_, _09779_, _09777_);
  nor (_09781_, _09780_, _09765_);
  nor (_09782_, _09609_, _09607_);
  nor (_09783_, _09782_, _09610_);
  not (_09784_, _09783_);
  nor (_09785_, _09784_, _09781_);
  nor (_09786_, _09775_, _09772_);
  not (_09787_, _09786_);
  and (_09788_, _09784_, _09781_);
  nor (_09789_, _09788_, _09785_);
  and (_09790_, _09789_, _09787_);
  nor (_09791_, _09790_, _09785_);
  nor (_09792_, _09646_, _09644_);
  nor (_09793_, _09792_, _09647_);
  not (_09794_, _09793_);
  nor (_09795_, _09794_, _09791_);
  and (_09796_, _09681_, _09648_);
  nor (_09797_, _09796_, _09682_);
  and (_09798_, _09797_, _09795_);
  nor (_09799_, _09709_, _09682_);
  nor (_09800_, _09799_, _09710_);
  nand (_09801_, _09800_, _09798_);
  and (_09802_, \uc8051golden_1.ACC [4], \uc8051golden_1.B [1]);
  and (_09803_, _09802_, _09737_);
  and (_09804_, \uc8051golden_1.B [2], \uc8051golden_1.ACC [3]);
  nor (_09805_, _09802_, _09737_);
  nor (_09806_, _09805_, _09803_);
  and (_09807_, _09806_, _09804_);
  nor (_09808_, _09807_, _09803_);
  not (_09809_, _09808_);
  nor (_09810_, _09742_, _09739_);
  nor (_09811_, _09810_, _09743_);
  and (_09812_, _09811_, _09809_);
  and (_09813_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [5]);
  and (_09814_, \uc8051golden_1.B [3], \uc8051golden_1.ACC [3]);
  and (_09815_, \uc8051golden_1.B [4], \uc8051golden_1.ACC [2]);
  and (_09816_, _09815_, _09814_);
  nor (_09817_, _09815_, _09814_);
  nor (_09818_, _09817_, _09816_);
  and (_09819_, _09818_, _09813_);
  nor (_09820_, _09818_, _09813_);
  nor (_09821_, _09820_, _09819_);
  nor (_09822_, _09811_, _09809_);
  nor (_09823_, _09822_, _09812_);
  and (_09824_, _09823_, _09821_);
  nor (_09825_, _09824_, _09812_);
  not (_09826_, _09825_);
  nor (_09827_, _09759_, _09757_);
  nor (_09828_, _09827_, _09760_);
  and (_09829_, _09828_, _09826_);
  nor (_09830_, _09819_, _09816_);
  and (_09831_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [6]);
  and (_09832_, \uc8051golden_1.ACC [0], \uc8051golden_1.B [7]);
  nor (_09833_, _09832_, _09831_);
  nor (_09834_, _09833_, _09767_);
  not (_09835_, _09834_);
  nor (_09836_, _09835_, _09830_);
  and (_09837_, _09835_, _09830_);
  nor (_09838_, _09837_, _09836_);
  nor (_09839_, _09828_, _09826_);
  nor (_09840_, _09839_, _09829_);
  and (_09841_, _09840_, _09838_);
  nor (_09842_, _09841_, _09829_);
  nor (_09843_, _09779_, _09777_);
  nor (_09844_, _09843_, _09780_);
  not (_09845_, _09844_);
  nor (_09846_, _09845_, _09842_);
  and (_09847_, _09845_, _09842_);
  nor (_09848_, _09847_, _09846_);
  and (_09849_, _09848_, _09836_);
  nor (_09850_, _09849_, _09846_);
  nor (_09851_, _09789_, _09787_);
  nor (_09852_, _09851_, _09790_);
  not (_09853_, _09852_);
  nor (_09854_, _09853_, _09850_);
  and (_09855_, _09794_, _09791_);
  nor (_09856_, _09855_, _09795_);
  and (_09857_, _09856_, _09854_);
  nor (_09858_, _09797_, _09795_);
  nor (_09859_, _09858_, _09798_);
  and (_09860_, _09859_, _09857_);
  nor (_09861_, _09859_, _09857_);
  nor (_09862_, _09861_, _09860_);
  and (_09863_, \uc8051golden_1.ACC [4], \uc8051golden_1.B [0]);
  and (_09864_, \uc8051golden_1.B [1], \uc8051golden_1.ACC [3]);
  and (_09865_, _09864_, _09863_);
  and (_09866_, \uc8051golden_1.B [2], \uc8051golden_1.ACC [2]);
  nor (_09867_, _09864_, _09863_);
  nor (_09868_, _09867_, _09865_);
  and (_09869_, _09868_, _09866_);
  nor (_09870_, _09869_, _09865_);
  not (_09871_, _09870_);
  nor (_09872_, _09806_, _09804_);
  nor (_09873_, _09872_, _09807_);
  and (_09874_, _09873_, _09871_);
  and (_09875_, \uc8051golden_1.B [5], \uc8051golden_1.ACC [0]);
  and (_09876_, \uc8051golden_1.B [3], \uc8051golden_1.ACC [2]);
  and (_09877_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [4]);
  and (_09878_, _09877_, _09876_);
  nor (_09879_, _09877_, _09876_);
  nor (_09880_, _09879_, _09878_);
  and (_09881_, _09880_, _09875_);
  nor (_09882_, _09880_, _09875_);
  nor (_09883_, _09882_, _09881_);
  nor (_09884_, _09873_, _09871_);
  nor (_09885_, _09884_, _09874_);
  and (_09886_, _09885_, _09883_);
  nor (_09887_, _09886_, _09874_);
  not (_09888_, _09887_);
  nor (_09889_, _09823_, _09821_);
  nor (_09890_, _09889_, _09824_);
  and (_09891_, _09890_, _09888_);
  not (_09892_, _09766_);
  nor (_09893_, _09881_, _09878_);
  nor (_09894_, _09893_, _09892_);
  and (_09895_, _09893_, _09892_);
  nor (_09896_, _09895_, _09894_);
  nor (_09897_, _09890_, _09888_);
  nor (_09898_, _09897_, _09891_);
  and (_09899_, _09898_, _09896_);
  nor (_09900_, _09899_, _09891_);
  not (_09901_, _09900_);
  nor (_09902_, _09840_, _09838_);
  nor (_09903_, _09902_, _09841_);
  and (_09904_, _09903_, _09901_);
  nor (_09905_, _09903_, _09901_);
  nor (_09906_, _09905_, _09904_);
  and (_09907_, _09906_, _09894_);
  nor (_09908_, _09907_, _09904_);
  nor (_09909_, _09848_, _09836_);
  nor (_09910_, _09909_, _09849_);
  not (_09911_, _09910_);
  nor (_09912_, _09911_, _09908_);
  and (_09913_, _09853_, _09850_);
  nor (_09914_, _09913_, _09854_);
  and (_09915_, _09914_, _09912_);
  nor (_09916_, _09856_, _09854_);
  nor (_09917_, _09916_, _09857_);
  nand (_09918_, _09917_, _09915_);
  or (_09919_, _09917_, _09915_);
  and (_09920_, _09919_, _09918_);
  and (_09921_, \uc8051golden_1.B [0], \uc8051golden_1.ACC [3]);
  and (_09922_, \uc8051golden_1.B [1], \uc8051golden_1.ACC [2]);
  and (_09923_, _09922_, _09921_);
  and (_09924_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [2]);
  nor (_09925_, _09922_, _09921_);
  nor (_09926_, _09925_, _09923_);
  and (_09927_, _09926_, _09924_);
  nor (_09928_, _09927_, _09923_);
  not (_09929_, _09928_);
  nor (_09930_, _09868_, _09866_);
  nor (_09931_, _09930_, _09869_);
  and (_09932_, _09931_, _09929_);
  and (_09933_, \uc8051golden_1.B [3], \uc8051golden_1.ACC [0]);
  and (_09934_, _09933_, _09877_);
  and (_09935_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [3]);
  and (_09936_, \uc8051golden_1.B [4], \uc8051golden_1.ACC [0]);
  nor (_09937_, _09936_, _09935_);
  nor (_09938_, _09937_, _09934_);
  nor (_09939_, _09931_, _09929_);
  nor (_09940_, _09939_, _09932_);
  and (_09941_, _09940_, _09938_);
  nor (_09942_, _09941_, _09932_);
  not (_09943_, _09942_);
  nor (_09944_, _09885_, _09883_);
  nor (_09945_, _09944_, _09886_);
  and (_09946_, _09945_, _09943_);
  nor (_09947_, _09945_, _09943_);
  nor (_09948_, _09947_, _09946_);
  and (_09949_, _09948_, _09934_);
  nor (_09950_, _09949_, _09946_);
  not (_09951_, _09950_);
  nor (_09952_, _09898_, _09896_);
  nor (_09953_, _09952_, _09899_);
  and (_09954_, _09953_, _09951_);
  nor (_09955_, _09906_, _09894_);
  nor (_09956_, _09955_, _09907_);
  and (_09957_, _09956_, _09954_);
  and (_09958_, _09911_, _09908_);
  nor (_09959_, _09958_, _09912_);
  and (_09960_, _09959_, _09957_);
  nor (_09961_, _09914_, _09912_);
  nor (_09962_, _09961_, _09915_);
  and (_09963_, _09962_, _09960_);
  nor (_09964_, _09962_, _09960_);
  nor (_09965_, _09964_, _09963_);
  and (_09966_, \uc8051golden_1.B [0], \uc8051golden_1.ACC [2]);
  and (_09967_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [1]);
  and (_09968_, _09967_, _09966_);
  and (_09969_, \uc8051golden_1.B [2], \uc8051golden_1.ACC [0]);
  nor (_09970_, _09967_, _09966_);
  nor (_09971_, _09970_, _09968_);
  and (_09972_, _09971_, _09969_);
  nor (_09973_, _09972_, _09968_);
  not (_09974_, _09973_);
  nor (_09975_, _09926_, _09924_);
  nor (_09976_, _09975_, _09927_);
  and (_09977_, _09976_, _09974_);
  nor (_09978_, _09976_, _09974_);
  nor (_09979_, _09978_, _09977_);
  and (_09980_, _09979_, _09933_);
  nor (_09981_, _09980_, _09977_);
  not (_09982_, _09981_);
  nor (_09983_, _09940_, _09938_);
  nor (_09984_, _09983_, _09941_);
  and (_09985_, _09984_, _09982_);
  nor (_09986_, _09948_, _09934_);
  nor (_09987_, _09986_, _09949_);
  and (_09988_, _09987_, _09985_);
  nor (_09989_, _09953_, _09951_);
  nor (_09990_, _09989_, _09954_);
  and (_09991_, _09990_, _09988_);
  nor (_09992_, _09956_, _09954_);
  nor (_09993_, _09992_, _09957_);
  and (_09994_, _09993_, _09991_);
  nor (_09995_, _09959_, _09957_);
  nor (_09996_, _09995_, _09960_);
  and (_09997_, _09996_, _09994_);
  and (_09998_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [0]);
  and (_09999_, \uc8051golden_1.B [1], \uc8051golden_1.ACC [0]);
  and (_10000_, _09999_, _09998_);
  nor (_10001_, _09971_, _09969_);
  nor (_10002_, _10001_, _09972_);
  and (_10003_, _10002_, _10000_);
  nor (_10004_, _09979_, _09933_);
  nor (_10005_, _10004_, _09980_);
  and (_10006_, _10005_, _10003_);
  nor (_10007_, _09984_, _09982_);
  nor (_10008_, _10007_, _09985_);
  and (_10009_, _10008_, _10006_);
  nor (_10010_, _09987_, _09985_);
  nor (_10011_, _10010_, _09988_);
  and (_10012_, _10011_, _10009_);
  nor (_10013_, _09990_, _09988_);
  nor (_10014_, _10013_, _09991_);
  and (_10015_, _10014_, _10012_);
  nor (_10016_, _09993_, _09991_);
  nor (_10017_, _10016_, _09994_);
  and (_10018_, _10017_, _10015_);
  nor (_10019_, _09996_, _09994_);
  nor (_10020_, _10019_, _09997_);
  and (_10021_, _10020_, _10018_);
  nor (_10022_, _10021_, _09997_);
  not (_10023_, _10022_);
  and (_10024_, _10023_, _09965_);
  or (_10025_, _10024_, _09963_);
  nand (_10026_, _10025_, _09920_);
  and (_10027_, _10026_, _09918_);
  not (_10028_, _10027_);
  and (_10029_, _10028_, _09862_);
  or (_10030_, _10029_, _09860_);
  or (_10031_, _09800_, _09798_);
  and (_10032_, _10031_, _09801_);
  nand (_10033_, _10032_, _10030_);
  and (_10034_, _10033_, _09801_);
  nor (_10035_, _10034_, _09736_);
  or (_10036_, _10035_, _09735_);
  and (_10037_, \uc8051golden_1.ACC [7], \uc8051golden_1.B [7]);
  not (_10038_, _10037_);
  nor (_10039_, _10038_, _09687_);
  nor (_10040_, _10039_, _09719_);
  nor (_10041_, _09725_, _09722_);
  nor (_10042_, _10041_, _10040_);
  and (_10043_, _10041_, _10040_);
  nor (_10044_, _10043_, _10042_);
  nor (_10045_, _09732_, _09729_);
  and (_10046_, _10045_, _10044_);
  nor (_10047_, _10045_, _10044_);
  or (_10048_, _10047_, _10046_);
  and (_10049_, _10048_, _10036_);
  and (_10050_, _10044_, _09729_);
  or (_10051_, _10042_, _09716_);
  or (_10052_, _10051_, _10050_);
  and (_10053_, _10044_, _09732_);
  or (_10054_, _10053_, _10052_);
  or (_10055_, _10054_, _10049_);
  or (_10056_, _10055_, _09544_);
  and (_10057_, _10056_, _06446_);
  and (_10058_, _10057_, _09543_);
  not (_10059_, _06293_);
  and (_10060_, _08794_, _08618_);
  or (_10061_, _10060_, _09509_);
  and (_10062_, _10061_, _06300_);
  or (_10063_, _10062_, _10059_);
  or (_10064_, _10063_, _10058_);
  and (_10065_, _10064_, _09508_);
  or (_10066_, _10065_, _06281_);
  and (_10067_, _07992_, _08749_);
  or (_10068_, _09503_, _06282_);
  or (_10069_, _10068_, _10067_);
  and (_10070_, _10069_, _06279_);
  and (_10071_, _10070_, _10066_);
  and (_10072_, _06481_, _05935_);
  and (_10073_, _09009_, _07992_);
  or (_10074_, _10073_, _09503_);
  and (_10075_, _10074_, _06015_);
  or (_10076_, _10075_, _10072_);
  or (_10077_, _10076_, _10071_);
  not (_10078_, _10072_);
  not (_10079_, \uc8051golden_1.B [1]);
  nor (_10080_, \uc8051golden_1.B [6], \uc8051golden_1.B [5]);
  nor (_10081_, \uc8051golden_1.B [4], \uc8051golden_1.B [3]);
  and (_10082_, _10081_, _10080_);
  and (_10083_, _10082_, _10079_);
  not (_10084_, \uc8051golden_1.B [0]);
  and (_10085_, _10084_, \uc8051golden_1.ACC [7]);
  nor (_10086_, \uc8051golden_1.B [2], \uc8051golden_1.B [7]);
  and (_10087_, _10086_, _10085_);
  and (_10088_, _10087_, _10083_);
  not (_10089_, _10086_);
  and (_10090_, \uc8051golden_1.B [0], _08651_);
  nor (_10091_, _10090_, _10089_);
  and (_10092_, _10091_, _10083_);
  or (_10093_, _10092_, _08651_);
  not (_10094_, \uc8051golden_1.B [4]);
  not (_10095_, \uc8051golden_1.B [5]);
  nor (_10096_, \uc8051golden_1.B [6], \uc8051golden_1.B [7]);
  and (_10097_, _10096_, _10095_);
  and (_10098_, _10097_, _10094_);
  nor (_10099_, \uc8051golden_1.B [3], \uc8051golden_1.B [2]);
  and (_10100_, _10099_, _10098_);
  not (_10101_, \uc8051golden_1.ACC [6]);
  and (_10102_, \uc8051golden_1.B [0], _10101_);
  nor (_10103_, _10102_, _08651_);
  nor (_10104_, _10103_, _10079_);
  not (_10105_, _10104_);
  and (_10106_, _10105_, _10100_);
  nor (_10107_, _10106_, _10093_);
  nor (_10108_, _10107_, _10088_);
  and (_10109_, _10106_, \uc8051golden_1.B [0]);
  nor (_10110_, _10109_, _10101_);
  and (_10111_, _10110_, _10079_);
  nor (_10112_, _10110_, _10079_);
  nor (_10113_, _10112_, _10111_);
  nor (_10114_, \uc8051golden_1.ACC [5], \uc8051golden_1.B [0]);
  nor (_10115_, _10114_, _09737_);
  nor (_10116_, _10115_, \uc8051golden_1.ACC [4]);
  and (_10117_, \uc8051golden_1.ACC [4], _10084_);
  nor (_10118_, _10117_, \uc8051golden_1.ACC [5]);
  not (_10119_, \uc8051golden_1.ACC [4]);
  and (_10120_, _10119_, \uc8051golden_1.B [0]);
  nor (_10121_, _10120_, _10118_);
  nor (_10122_, _10121_, _10116_);
  not (_10123_, _10122_);
  and (_10124_, _10123_, _10113_);
  nor (_10125_, _10108_, \uc8051golden_1.B [2]);
  nor (_10126_, _10125_, _10111_);
  not (_10127_, _10126_);
  nor (_10128_, _10127_, _10124_);
  not (_10129_, _10128_);
  and (_10130_, \uc8051golden_1.B [2], _08651_);
  nor (_10131_, _10130_, \uc8051golden_1.B [7]);
  and (_10132_, _10131_, _10082_);
  and (_10133_, _10132_, _10129_);
  nor (_10134_, _10133_, _10108_);
  nor (_10135_, _10134_, _10088_);
  nor (_10136_, _10123_, _10113_);
  nor (_10137_, _10136_, _10124_);
  and (_10138_, _10137_, _10133_);
  not (_10139_, _10110_);
  nor (_10140_, _10133_, _10139_);
  nor (_10141_, _10140_, _10138_);
  nor (_10142_, _10141_, \uc8051golden_1.B [2]);
  and (_10143_, _10141_, \uc8051golden_1.B [2]);
  nor (_10144_, _10143_, _10142_);
  not (_10145_, \uc8051golden_1.ACC [5]);
  nor (_10146_, _10133_, _10145_);
  and (_10147_, _10133_, _10115_);
  or (_10148_, _10147_, _10146_);
  and (_10149_, _10148_, _10079_);
  nor (_10150_, _10148_, _10079_);
  nor (_10151_, _10150_, _10120_);
  nor (_10152_, _10151_, _10149_);
  not (_10153_, _10152_);
  and (_10154_, _10153_, _10144_);
  nor (_10155_, _10135_, \uc8051golden_1.B [3]);
  nor (_10156_, _10155_, _10142_);
  not (_10157_, _10156_);
  nor (_10158_, _10157_, _10154_);
  not (_10159_, _10158_);
  and (_10160_, \uc8051golden_1.B [3], _08651_);
  not (_10161_, _10160_);
  and (_10162_, _10161_, _10098_);
  and (_10163_, _10162_, _10159_);
  nor (_10164_, _10163_, _10135_);
  nor (_10165_, _10164_, _10088_);
  not (_10166_, \uc8051golden_1.B [3]);
  nor (_10167_, _10163_, _10141_);
  nor (_10168_, _10153_, _10144_);
  nor (_10169_, _10168_, _10154_);
  and (_10170_, _10169_, _10163_);
  or (_10171_, _10170_, _10167_);
  and (_10172_, _10171_, _10166_);
  nor (_10173_, _10171_, _10166_);
  nor (_10174_, _10173_, _10172_);
  not (_10175_, _10174_);
  nor (_10176_, _10163_, _10148_);
  nor (_10177_, _10150_, _10149_);
  and (_10178_, _10177_, _10120_);
  nor (_10179_, _10177_, _10120_);
  nor (_10180_, _10179_, _10178_);
  and (_10181_, _10180_, _10163_);
  or (_10182_, _10181_, _10176_);
  nor (_10183_, _10182_, \uc8051golden_1.B [2]);
  and (_10184_, _10182_, \uc8051golden_1.B [2]);
  nor (_10185_, _10120_, _10117_);
  and (_10186_, _10163_, _10185_);
  nor (_10187_, _10163_, \uc8051golden_1.ACC [4]);
  nor (_10188_, _10187_, _10186_);
  and (_10189_, _10188_, _10079_);
  nor (_10190_, \uc8051golden_1.B [0], \uc8051golden_1.ACC [3]);
  nor (_10191_, _10190_, _09921_);
  nor (_10192_, _10191_, \uc8051golden_1.ACC [2]);
  and (_10193_, _10084_, \uc8051golden_1.ACC [2]);
  nor (_10194_, _10193_, \uc8051golden_1.ACC [3]);
  not (_10195_, \uc8051golden_1.ACC [2]);
  and (_10196_, \uc8051golden_1.B [0], _10195_);
  nor (_10197_, _10196_, _10194_);
  nor (_10198_, _10197_, _10192_);
  not (_10199_, _10198_);
  nor (_10200_, _10188_, _10079_);
  nor (_10201_, _10200_, _10189_);
  and (_10202_, _10201_, _10199_);
  nor (_10203_, _10202_, _10189_);
  nor (_10204_, _10203_, _10184_);
  nor (_10205_, _10204_, _10183_);
  nor (_10206_, _10205_, _10175_);
  nor (_10207_, _10165_, \uc8051golden_1.B [4]);
  nor (_10208_, _10207_, _10172_);
  not (_10209_, _10208_);
  nor (_10210_, _10209_, _10206_);
  not (_10211_, _10210_);
  not (_10212_, _10097_);
  and (_10213_, \uc8051golden_1.B [4], _08651_);
  nor (_10214_, _10213_, _10212_);
  and (_10215_, _10214_, _10211_);
  nor (_10216_, _10215_, _10165_);
  nor (_10217_, _10216_, _10088_);
  and (_10218_, _10096_, \uc8051golden_1.ACC [7]);
  nor (_10219_, _10218_, _10097_);
  nor (_10220_, _10217_, \uc8051golden_1.B [5]);
  not (_10221_, _10215_);
  and (_10222_, _10205_, _10175_);
  nor (_10223_, _10222_, _10206_);
  nor (_10224_, _10223_, _10221_);
  nor (_10225_, _10215_, _10171_);
  nor (_10226_, _10225_, _10224_);
  and (_10227_, _10226_, _10094_);
  nor (_10228_, _10226_, _10094_);
  nor (_10229_, _10228_, _10227_);
  not (_10230_, _10229_);
  nor (_10231_, _10215_, _10182_);
  nor (_10232_, _10184_, _10183_);
  and (_10233_, _10232_, _10203_);
  nor (_10234_, _10232_, _10203_);
  nor (_10235_, _10234_, _10233_);
  nor (_10236_, _10235_, _10221_);
  nor (_10237_, _10236_, _10231_);
  nor (_10238_, _10237_, \uc8051golden_1.B [3]);
  and (_10239_, _10237_, \uc8051golden_1.B [3]);
  nor (_10240_, _10201_, _10199_);
  nor (_10241_, _10240_, _10202_);
  and (_10242_, _10241_, _10215_);
  and (_10243_, _10221_, _10188_);
  nor (_10244_, _10243_, _10242_);
  nor (_10245_, _10244_, \uc8051golden_1.B [2]);
  not (_10246_, \uc8051golden_1.ACC [3]);
  nor (_10247_, _10215_, _10246_);
  and (_10248_, _10215_, _10191_);
  or (_10249_, _10248_, _10247_);
  and (_10250_, _10249_, _10079_);
  nor (_10251_, _10249_, _10079_);
  nor (_10252_, _10251_, _10196_);
  nor (_10253_, _10252_, _10250_);
  not (_10254_, _10253_);
  and (_10255_, _10244_, \uc8051golden_1.B [2]);
  nor (_10256_, _10255_, _10245_);
  and (_10257_, _10256_, _10254_);
  nor (_10258_, _10257_, _10245_);
  nor (_10259_, _10258_, _10239_);
  nor (_10260_, _10259_, _10238_);
  nor (_10261_, _10260_, _10230_);
  or (_10262_, _10261_, _10227_);
  nor (_10263_, _10262_, _10220_);
  nor (_10264_, _10263_, _10219_);
  nor (_10265_, _10264_, _10217_);
  not (_10266_, _10264_);
  and (_10267_, _10260_, _10230_);
  nor (_10268_, _10267_, _10261_);
  nor (_10269_, _10268_, _10266_);
  nor (_10270_, _10264_, _10226_);
  nor (_10271_, _10270_, _10269_);
  and (_10272_, _10271_, _10095_);
  nor (_10273_, _10271_, _10095_);
  nor (_10274_, _10273_, _10272_);
  not (_10275_, _10274_);
  nor (_10276_, _10264_, _10237_);
  nor (_10277_, _10239_, _10238_);
  nor (_10278_, _10277_, _10258_);
  and (_10279_, _10277_, _10258_);
  or (_10280_, _10279_, _10278_);
  and (_10281_, _10280_, _10264_);
  or (_10282_, _10281_, _10276_);
  and (_10283_, _10282_, _10094_);
  nor (_10284_, _10282_, _10094_);
  nor (_10285_, _10264_, _10244_);
  nor (_10286_, _10256_, _10254_);
  nor (_10287_, _10286_, _10257_);
  and (_10288_, _10287_, _10264_);
  or (_10289_, _10288_, _10285_);
  and (_10290_, _10289_, _10166_);
  not (_10291_, \uc8051golden_1.B [2]);
  nor (_10292_, _10251_, _10250_);
  nor (_10293_, _10292_, _10196_);
  and (_10294_, _10292_, _10196_);
  or (_10295_, _10294_, _10293_);
  nor (_10296_, _10295_, _10266_);
  nor (_10297_, _10264_, _10249_);
  nor (_10298_, _10297_, _10296_);
  and (_10299_, _10298_, _10291_);
  nor (_10300_, _10298_, _10291_);
  nor (_10301_, _10196_, _10193_);
  and (_10302_, _10264_, _10301_);
  nor (_10303_, _10264_, \uc8051golden_1.ACC [2]);
  nor (_10304_, _10303_, _10302_);
  and (_10305_, _10304_, _10079_);
  and (_10306_, _05984_, \uc8051golden_1.B [0]);
  not (_10307_, _10306_);
  nor (_10308_, _10304_, _10079_);
  nor (_10309_, _10308_, _10305_);
  and (_10310_, _10309_, _10307_);
  nor (_10311_, _10310_, _10305_);
  nor (_10312_, _10311_, _10300_);
  nor (_10313_, _10312_, _10299_);
  nor (_10314_, _10289_, _10166_);
  nor (_10315_, _10314_, _10290_);
  not (_10316_, _10315_);
  nor (_10317_, _10316_, _10313_);
  nor (_10318_, _10317_, _10290_);
  nor (_10319_, _10318_, _10284_);
  nor (_10320_, _10319_, _10283_);
  nor (_10321_, _10320_, _10275_);
  nor (_10322_, _10321_, _10272_);
  and (_10323_, \uc8051golden_1.ACC [7], _09501_);
  nor (_10324_, _10323_, _10096_);
  nor (_10325_, _10324_, _10322_);
  not (_10326_, _10096_);
  nor (_10327_, _10265_, _10088_);
  nor (_10328_, _10327_, _10326_);
  nor (_10329_, _10328_, _10325_);
  and (_10330_, _10329_, _10265_);
  or (_10331_, _10330_, _10088_);
  nor (_10332_, _10331_, _09501_);
  nor (_10333_, _10331_, \uc8051golden_1.B [7]);
  nor (_10334_, _10333_, _10037_);
  not (_10335_, _10334_);
  not (_10336_, \uc8051golden_1.B [6]);
  and (_10337_, _10320_, _10275_);
  nor (_10338_, _10337_, _10321_);
  nor (_10339_, _10338_, _10329_);
  not (_10340_, _10329_);
  nor (_10341_, _10340_, _10271_);
  nor (_10342_, _10341_, _10339_);
  nor (_10343_, _10342_, _10336_);
  and (_10344_, _10342_, _10336_);
  nor (_10345_, _10284_, _10283_);
  nor (_10346_, _10345_, _10318_);
  and (_10347_, _10345_, _10318_);
  or (_10348_, _10347_, _10346_);
  nor (_10349_, _10348_, _10329_);
  nor (_10350_, _10340_, _10282_);
  nor (_10351_, _10350_, _10349_);
  nor (_10352_, _10351_, _10095_);
  and (_10353_, _10351_, _10095_);
  not (_10354_, _10353_);
  and (_10355_, _10316_, _10313_);
  nor (_10356_, _10355_, _10317_);
  nor (_10357_, _10356_, _10329_);
  nor (_10358_, _10340_, _10289_);
  nor (_10359_, _10358_, _10357_);
  nor (_10360_, _10359_, _10094_);
  and (_10361_, _10329_, _10298_);
  nor (_10362_, _10300_, _10299_);
  and (_10363_, _10362_, _10311_);
  nor (_10364_, _10362_, _10311_);
  nor (_10365_, _10364_, _10363_);
  nor (_10366_, _10365_, _10329_);
  or (_10367_, _10366_, _10361_);
  nor (_10368_, _10367_, _10166_);
  and (_10369_, _10367_, _10166_);
  nor (_10370_, _10369_, _10368_);
  nor (_10371_, _10309_, _10307_);
  nor (_10372_, _10371_, _10310_);
  nor (_10373_, _10372_, _10329_);
  nor (_10374_, _10340_, _10304_);
  nor (_10375_, _10374_, _10373_);
  nor (_10376_, _10375_, _10291_);
  and (_10377_, _10375_, _10291_);
  nor (_10378_, _10377_, _10376_);
  and (_10379_, _10378_, _10370_);
  and (_10380_, _10329_, _05984_);
  nor (_10381_, \uc8051golden_1.ACC [1], \uc8051golden_1.B [0]);
  nor (_10382_, _10381_, _09998_);
  nor (_10383_, _10329_, _10382_);
  nor (_10384_, _10383_, _10380_);
  and (_10385_, _10384_, _10079_);
  nor (_10386_, _10384_, _10079_);
  and (_10387_, _10084_, \uc8051golden_1.ACC [0]);
  not (_10388_, _10387_);
  nor (_10389_, _10388_, _10386_);
  nor (_10390_, _10389_, _10385_);
  and (_10391_, _10390_, _10379_);
  and (_10392_, _10376_, _10370_);
  nor (_10393_, _10392_, _10368_);
  not (_10394_, _10393_);
  nor (_10395_, _10394_, _10391_);
  and (_10396_, _10359_, _10094_);
  nor (_10397_, _10396_, _10395_);
  or (_10398_, _10397_, _10360_);
  and (_10399_, _10398_, _10354_);
  nor (_10400_, _10399_, _10352_);
  nor (_10401_, _10400_, _10344_);
  or (_10402_, _10401_, _10343_);
  and (_10403_, _10402_, _10335_);
  nor (_10404_, _10403_, _10332_);
  nor (_10405_, _10396_, _10360_);
  nor (_10406_, _10353_, _10352_);
  and (_10407_, _10406_, _10405_);
  nor (_10408_, _10344_, _10343_);
  and (_10409_, _10408_, _10335_);
  and (_10410_, _10409_, _10407_);
  nor (_10411_, _10386_, _10385_);
  and (_10412_, \uc8051golden_1.B [0], _06045_);
  not (_10413_, _10412_);
  and (_10414_, _10413_, _10411_);
  and (_10415_, _10414_, _10388_);
  and (_10416_, _10415_, _10379_);
  and (_10417_, _10416_, _10410_);
  nor (_10418_, _10417_, _10404_);
  or (_10419_, _10418_, _10088_);
  and (_10420_, _10419_, _10331_);
  or (_10421_, _10420_, _10078_);
  and (_10422_, _10421_, _10077_);
  or (_10423_, _10422_, _06275_);
  and (_10424_, _08813_, _07992_);
  or (_10425_, _10424_, _09503_);
  or (_10426_, _10425_, _06276_);
  and (_10427_, _10426_, _07282_);
  and (_10428_, _10427_, _10423_);
  and (_10429_, _09027_, _07992_);
  or (_10430_, _10429_, _09503_);
  and (_10431_, _10430_, _06474_);
  or (_10432_, _10431_, _06582_);
  or (_10433_, _10432_, _10428_);
  and (_10434_, _09034_, _07992_);
  or (_10435_, _10434_, _09503_);
  or (_10436_, _10435_, _07284_);
  and (_10437_, _10436_, _07279_);
  and (_10438_, _10437_, _10433_);
  or (_10439_, _09503_, _08073_);
  and (_10440_, _10425_, _06478_);
  and (_10441_, _10440_, _10439_);
  or (_10442_, _10441_, _10438_);
  and (_10443_, _10442_, _07276_);
  and (_10444_, _09517_, _06569_);
  and (_10445_, _10444_, _10439_);
  or (_10446_, _10445_, _06479_);
  or (_10447_, _10446_, _10443_);
  and (_10448_, _09026_, _07992_);
  or (_10449_, _09503_, _09043_);
  or (_10450_, _10449_, _10448_);
  and (_10451_, _10450_, _09048_);
  and (_10452_, _10451_, _10447_);
  nor (_10453_, _09033_, _09504_);
  or (_10454_, _10453_, _09503_);
  and (_10455_, _10454_, _06572_);
  or (_10456_, _10455_, _06606_);
  or (_10457_, _10456_, _10452_);
  or (_10458_, _09514_, _07037_);
  and (_10459_, _10458_, _06807_);
  and (_10460_, _10459_, _10457_);
  and (_10461_, _09511_, _06234_);
  or (_10462_, _10461_, _06195_);
  or (_10463_, _10462_, _10460_);
  and (_10464_, _08530_, _07992_);
  or (_10465_, _09503_, _06196_);
  or (_10466_, _10465_, _10464_);
  and (_10467_, _10466_, _01375_);
  and (_10468_, _10467_, _10463_);
  or (_10469_, _10468_, _09502_);
  and (_40323_, _10469_, _42545_);
  nor (_10470_, _01375_, _08651_);
  and (_10471_, _06280_, _05965_);
  not (_10472_, _10471_);
  and (_10473_, _09452_, \uc8051golden_1.PSW [7]);
  nor (_10474_, _10473_, _09075_);
  and (_10475_, _10473_, _09075_);
  nor (_10476_, _10475_, _10474_);
  and (_10477_, _10476_, \uc8051golden_1.ACC [7]);
  nor (_10478_, _10476_, \uc8051golden_1.ACC [7]);
  nor (_10479_, _10478_, _10477_);
  and (_10480_, _09451_, \uc8051golden_1.PSW [7]);
  nor (_10481_, _10480_, _09440_);
  nor (_10482_, _10481_, _10473_);
  nand (_10483_, _10482_, \uc8051golden_1.ACC [6]);
  nor (_10484_, _10482_, _10101_);
  and (_10485_, _10482_, _10101_);
  nor (_10486_, _10485_, _10484_);
  not (_10487_, _10486_);
  and (_10488_, _09450_, \uc8051golden_1.PSW [7]);
  nor (_10489_, _10488_, _09441_);
  nor (_10490_, _10489_, _10480_);
  and (_10491_, _10490_, \uc8051golden_1.ACC [5]);
  nor (_10492_, _10490_, _10145_);
  and (_10493_, _10490_, _10145_);
  nor (_10494_, _10493_, _10492_);
  and (_10495_, _09449_, \uc8051golden_1.PSW [7]);
  nor (_10496_, _10495_, _09442_);
  nor (_10497_, _10496_, _10488_);
  nand (_10498_, _10497_, \uc8051golden_1.ACC [4]);
  nor (_10499_, _10497_, _10119_);
  and (_10500_, _10497_, _10119_);
  or (_10501_, _10500_, _10499_);
  and (_10502_, _09448_, \uc8051golden_1.PSW [7]);
  nor (_10503_, _10502_, _09443_);
  nor (_10504_, _10503_, _10495_);
  and (_10505_, _10504_, \uc8051golden_1.ACC [3]);
  nor (_10506_, _10504_, _10246_);
  and (_10507_, _10504_, _10246_);
  nor (_10508_, _10507_, _10506_);
  and (_10509_, _09447_, \uc8051golden_1.PSW [7]);
  nor (_10510_, _10509_, _09444_);
  nor (_10511_, _10510_, _10502_);
  and (_10512_, _10511_, \uc8051golden_1.ACC [2]);
  nor (_10513_, _10511_, _10195_);
  and (_10514_, _10511_, _10195_);
  nor (_10515_, _10514_, _10513_);
  and (_10516_, _09446_, \uc8051golden_1.PSW [7]);
  nor (_10517_, _10516_, _09445_);
  nor (_10518_, _10517_, _10509_);
  and (_10519_, _10518_, \uc8051golden_1.ACC [1]);
  and (_10520_, _10518_, _05984_);
  nor (_10521_, _10518_, _05984_);
  nor (_10522_, _10521_, _10520_);
  not (_10523_, _10522_);
  not (_10524_, \uc8051golden_1.PSW [7]);
  and (_10525_, _09390_, _10524_);
  nor (_10526_, _10525_, _10516_);
  and (_10527_, _10526_, \uc8051golden_1.ACC [0]);
  and (_10528_, _10527_, _10523_);
  nor (_10529_, _10528_, _10519_);
  nor (_10530_, _10529_, _10515_);
  nor (_10531_, _10530_, _10512_);
  nor (_10532_, _10531_, _10508_);
  or (_10533_, _10532_, _10505_);
  nand (_10534_, _10533_, _10501_);
  and (_10535_, _10534_, _10498_);
  nor (_10536_, _10535_, _10494_);
  or (_10537_, _10536_, _10491_);
  nand (_10538_, _10537_, _10487_);
  and (_10539_, _10538_, _10483_);
  nor (_10540_, _10539_, _10479_);
  and (_10541_, _10539_, _10479_);
  nor (_10542_, _10541_, _10540_);
  or (_10543_, _10542_, _10472_);
  and (_10544_, _10543_, _06579_);
  nor (_10545_, _07995_, _08651_);
  and (_10546_, _09026_, _07995_);
  or (_10547_, _10546_, _10545_);
  and (_10548_, _10547_, _06479_);
  and (_10549_, _08070_, _08651_);
  and (_10550_, _06742_, _05946_);
  not (_10551_, _10550_);
  and (_10552_, _06751_, _05946_);
  and (_10553_, _07103_, _05946_);
  nor (_10554_, _10553_, _10552_);
  and (_10555_, _10554_, _10551_);
  not (_10556_, _10555_);
  nand (_10557_, _10556_, _10549_);
  and (_10558_, _08749_, \uc8051golden_1.ACC [7]);
  and (_10559_, _06280_, _05955_);
  not (_10560_, _10559_);
  or (_10561_, _10560_, _10558_);
  nor (_10562_, _08070_, _08651_);
  nor (_10563_, _10562_, _10549_);
  not (_10564_, _05951_);
  nor (_10565_, _06463_, _10564_);
  and (_10566_, _10565_, _10563_);
  or (_10567_, _06194_, _06021_);
  not (_10568_, _07995_);
  nor (_10569_, _10568_, _08070_);
  or (_10570_, _10569_, _10545_);
  or (_10571_, _10570_, _06293_);
  and (_10572_, _06481_, _06016_);
  not (_10573_, _10572_);
  and (_10574_, _08521_, \uc8051golden_1.PSW [7]);
  and (_10575_, _10574_, _08477_);
  and (_10576_, _10575_, _08433_);
  and (_10577_, _10576_, _08389_);
  and (_10578_, _10577_, _08345_);
  and (_10579_, _10578_, _08256_);
  and (_10580_, _10579_, _08162_);
  nor (_10581_, _10580_, _08072_);
  and (_10582_, _10580_, _08072_);
  nor (_10583_, _10582_, _10581_);
  and (_10584_, _10583_, \uc8051golden_1.ACC [7]);
  nor (_10585_, _10583_, \uc8051golden_1.ACC [7]);
  nor (_10586_, _10585_, _10584_);
  not (_10587_, _10586_);
  nor (_10588_, _10579_, _08162_);
  nor (_10589_, _10588_, _10580_);
  nor (_10590_, _10589_, _10101_);
  nor (_10591_, _10578_, _08256_);
  nor (_10592_, _10591_, _10579_);
  and (_10593_, _10592_, _10145_);
  nor (_10594_, _10592_, _10145_);
  nor (_10595_, _10577_, _08345_);
  nor (_10596_, _10595_, _10578_);
  nor (_10597_, _10596_, _10119_);
  nor (_10598_, _10597_, _10594_);
  nor (_10599_, _10598_, _10593_);
  nor (_10600_, _10594_, _10593_);
  not (_10601_, _10600_);
  and (_10602_, _10596_, _10119_);
  or (_10603_, _10602_, _10597_);
  or (_10604_, _10603_, _10601_);
  nor (_10605_, _10576_, _08389_);
  nor (_10606_, _10605_, _10577_);
  nor (_10607_, _10606_, _10246_);
  and (_10608_, _10606_, _10246_);
  nor (_10609_, _10608_, _10607_);
  nor (_10610_, _10575_, _08433_);
  nor (_10611_, _10610_, _10576_);
  nor (_10612_, _10611_, _10195_);
  and (_10613_, _10611_, _10195_);
  nor (_10614_, _10613_, _10612_);
  and (_10615_, _10614_, _10609_);
  nor (_10616_, _10574_, _08477_);
  nor (_10617_, _10616_, _10575_);
  nor (_10618_, _10617_, _05984_);
  and (_10619_, _10617_, _05984_);
  nor (_10620_, _08521_, \uc8051golden_1.PSW [7]);
  nor (_10621_, _10620_, _10574_);
  and (_10622_, _10621_, _06045_);
  nor (_10623_, _10622_, _10619_);
  or (_10624_, _10623_, _10618_);
  and (_10625_, _10624_, _10615_);
  and (_10626_, _10612_, _10609_);
  or (_10627_, _10626_, _10607_);
  nor (_10628_, _10627_, _10625_);
  nor (_10629_, _10628_, _10604_);
  nor (_10630_, _10629_, _10599_);
  and (_10631_, _10589_, _10101_);
  nor (_10632_, _10590_, _10631_);
  not (_10633_, _10632_);
  nor (_10634_, _10633_, _10630_);
  or (_10635_, _10634_, _10590_);
  and (_10636_, _10635_, _10587_);
  nor (_10637_, _10635_, _10587_);
  or (_10638_, _10637_, _10636_);
  or (_10639_, _10638_, _06442_);
  and (_10640_, _10639_, _10573_);
  and (_10641_, _06849_, _06016_);
  and (_10642_, _06481_, _06392_);
  nand (_10643_, _10642_, _10246_);
  nor (_10644_, _05999_, _06012_);
  nand (_10645_, _10644_, _08070_);
  nor (_10646_, _08616_, _08651_);
  and (_10647_, _08635_, _08616_);
  or (_10648_, _10647_, _10646_);
  or (_10649_, _10648_, _06396_);
  and (_10650_, _10649_, _07221_);
  and (_10651_, _08762_, _07995_);
  or (_10652_, _10651_, _10545_);
  and (_10653_, _10652_, _06401_);
  and (_10654_, _06481_, _06402_);
  not (_10655_, _10654_);
  or (_10656_, _10655_, _08749_);
  not (_10657_, _06285_);
  and (_10659_, _06463_, _10657_);
  not (_10660_, _07343_);
  and (_10661_, _06850_, _10660_);
  and (_10662_, _10661_, _10659_);
  nor (_10663_, _10662_, _06001_);
  not (_10664_, _10663_);
  nor (_10665_, _10664_, _08070_);
  or (_10666_, _06854_, \uc8051golden_1.ACC [7]);
  nand (_10667_, _06854_, \uc8051golden_1.ACC [7]);
  nand (_10668_, _10667_, _10666_);
  nor (_10670_, _10668_, _10663_);
  or (_10671_, _10670_, _10654_);
  or (_10672_, _10671_, _10665_);
  and (_10673_, _07210_, _06002_);
  and (_10674_, _10673_, _10672_);
  and (_10675_, _10674_, _10656_);
  or (_10676_, _10675_, _10653_);
  and (_10677_, _06481_, _06394_);
  not (_10678_, _10677_);
  and (_10679_, _10678_, _10676_);
  nor (_10681_, \uc8051golden_1.ACC [1], \uc8051golden_1.ACC [2]);
  nor (_10682_, _10681_, _10246_);
  and (_10683_, _10682_, \uc8051golden_1.ACC [4]);
  and (_10684_, _10683_, \uc8051golden_1.ACC [5]);
  and (_10685_, _10684_, \uc8051golden_1.ACC [6]);
  and (_10686_, _10685_, \uc8051golden_1.ACC [7]);
  nor (_10687_, _10685_, \uc8051golden_1.ACC [7]);
  nor (_10688_, _10687_, _10686_);
  nor (_10689_, _10683_, \uc8051golden_1.ACC [5]);
  nor (_10690_, _10689_, _10684_);
  nor (_10692_, _10684_, \uc8051golden_1.ACC [6]);
  nor (_10693_, _10692_, _10685_);
  nor (_10694_, _10693_, _10690_);
  not (_10695_, _10694_);
  and (_10696_, _10695_, _10688_);
  not (_10697_, _10696_);
  nor (_10698_, _10686_, \uc8051golden_1.PSW [7]);
  and (_10699_, _10698_, _10697_);
  nor (_10700_, _10699_, _10694_);
  or (_10701_, _10700_, _10688_);
  and (_10703_, _10697_, _10677_);
  and (_10704_, _10703_, _10701_);
  or (_10705_, _10704_, _06395_);
  or (_10706_, _10705_, _10679_);
  and (_10707_, _10706_, _10650_);
  and (_10708_, _10570_, _06399_);
  or (_10709_, _10708_, _10644_);
  or (_10710_, _10709_, _10707_);
  and (_10711_, _10710_, _10645_);
  or (_10712_, _10711_, _07233_);
  not (_10714_, _07233_);
  or (_10715_, _08749_, _10714_);
  and (_10716_, _10715_, _06414_);
  and (_10717_, _10716_, _10712_);
  nor (_10718_, _08072_, _06414_);
  or (_10719_, _10718_, _10642_);
  or (_10720_, _10719_, _10717_);
  and (_10721_, _10720_, _10643_);
  or (_10722_, _10721_, _06393_);
  and (_10723_, _08639_, _08616_);
  or (_10725_, _10723_, _10646_);
  or (_10726_, _10725_, _06844_);
  and (_10727_, _10726_, _07245_);
  and (_10728_, _10727_, _10722_);
  or (_10729_, _10646_, _08634_);
  and (_10730_, _10729_, _06387_);
  and (_10731_, _10730_, _10648_);
  or (_10732_, _10731_, _09538_);
  or (_10733_, _10732_, _10728_);
  nor (_10734_, _10017_, _10015_);
  nor (_10735_, _10734_, _10018_);
  or (_10736_, _10735_, _09544_);
  and (_10737_, _07632_, _06016_);
  nor (_10738_, _06290_, _07103_);
  nor (_10739_, _10738_, _06905_);
  nor (_10740_, _10739_, _10737_);
  and (_10741_, _10740_, _10736_);
  and (_10742_, _10741_, _10733_);
  and (_10743_, _09428_, \uc8051golden_1.PSW [7]);
  and (_10744_, _10743_, _08548_);
  nor (_10745_, _10743_, _08548_);
  or (_10746_, _10745_, _10744_);
  and (_10747_, _10746_, \uc8051golden_1.ACC [7]);
  nor (_10748_, _10746_, \uc8051golden_1.ACC [7]);
  nor (_10749_, _10748_, _10747_);
  not (_10750_, _10749_);
  and (_10751_, _09427_, \uc8051golden_1.PSW [7]);
  nor (_10752_, _10751_, _09418_);
  nor (_10753_, _10752_, _10743_);
  nor (_10754_, _10753_, _10101_);
  and (_10755_, _09426_, \uc8051golden_1.PSW [7]);
  nor (_10756_, _10755_, _09419_);
  nor (_10757_, _10756_, _10751_);
  and (_10758_, _10757_, _10145_);
  nor (_10759_, _10757_, _10145_);
  nor (_10760_, _10759_, _10758_);
  not (_10761_, _10760_);
  and (_10762_, _09425_, \uc8051golden_1.PSW [7]);
  nor (_10763_, _10762_, _09420_);
  nor (_10764_, _10763_, _10755_);
  nor (_10765_, _10764_, _10119_);
  and (_10766_, _10764_, _10119_);
  or (_10767_, _10766_, _10765_);
  or (_10768_, _10767_, _10761_);
  and (_10769_, _09424_, \uc8051golden_1.PSW [7]);
  nor (_10770_, _10769_, _09421_);
  nor (_10771_, _10770_, _10762_);
  nor (_10772_, _10771_, _10246_);
  and (_10773_, _10771_, _10246_);
  nor (_10774_, _10773_, _10772_);
  and (_10775_, _09423_, \uc8051golden_1.PSW [7]);
  nor (_10776_, _10775_, _09422_);
  nor (_10777_, _10776_, _10769_);
  nor (_10778_, _10777_, _10195_);
  and (_10779_, _10777_, _10195_);
  nor (_10780_, _10779_, _10778_);
  and (_10781_, _10780_, _10774_);
  not (_10782_, _07196_);
  and (_10783_, _07473_, \uc8051golden_1.PSW [7]);
  nor (_10784_, _10783_, _10782_);
  nor (_10785_, _10784_, _10775_);
  nor (_10786_, _10785_, _05984_);
  and (_10787_, _10785_, _05984_);
  and (_10788_, _07485_, _10524_);
  nor (_10789_, _10788_, _10783_);
  and (_10790_, _10789_, _06045_);
  nor (_10791_, _10790_, _10787_);
  or (_10792_, _10791_, _10786_);
  and (_10793_, _10792_, _10781_);
  and (_10794_, _10778_, _10774_);
  or (_10795_, _10794_, _10772_);
  nor (_10796_, _10795_, _10793_);
  nor (_10797_, _10796_, _10768_);
  and (_10798_, _10765_, _10760_);
  nor (_10799_, _10798_, _10759_);
  not (_10800_, _10799_);
  nor (_10801_, _10800_, _10797_);
  and (_10802_, _10753_, _10101_);
  nor (_10803_, _10754_, _10802_);
  not (_10804_, _10803_);
  nor (_10805_, _10804_, _10801_);
  or (_10806_, _10805_, _10754_);
  and (_10807_, _10806_, _10750_);
  nor (_10808_, _10806_, _10750_);
  nor (_10809_, _10808_, _10807_);
  nor (_10810_, _10809_, _10740_);
  nor (_10811_, _10810_, _10742_);
  and (_10812_, _07343_, _06016_);
  nor (_10813_, _10812_, _10811_);
  not (_10814_, _10479_);
  nor (_10815_, _10499_, _10492_);
  nor (_10816_, _10815_, _10493_);
  not (_10817_, _10494_);
  or (_10818_, _10501_, _10817_);
  and (_10819_, _10515_, _10508_);
  and (_10820_, _10526_, _06045_);
  nor (_10821_, _10820_, _10520_);
  or (_10822_, _10821_, _10521_);
  and (_10823_, _10822_, _10819_);
  and (_10824_, _10513_, _10508_);
  or (_10825_, _10824_, _10506_);
  nor (_10826_, _10825_, _10823_);
  nor (_10827_, _10826_, _10818_);
  nor (_10828_, _10827_, _10816_);
  nor (_10829_, _10828_, _10487_);
  or (_10830_, _10829_, _10484_);
  and (_10831_, _10830_, _10814_);
  nor (_10832_, _10830_, _10814_);
  or (_10833_, _10832_, _10831_);
  and (_10834_, _10833_, _10812_);
  nor (_10835_, _10834_, _10813_);
  nor (_10836_, _10835_, _10641_);
  and (_10837_, _10833_, _10641_);
  or (_10838_, _10837_, _10836_);
  or (_10839_, _10838_, _06437_);
  and (_10840_, _10839_, _10640_);
  and (_10841_, _07964_, \uc8051golden_1.PSW [7]);
  and (_10842_, _10841_, _07978_);
  and (_10843_, _10842_, _07943_);
  and (_10844_, _10843_, _07896_);
  and (_10845_, _10844_, _06309_);
  nor (_10846_, _10844_, _06309_);
  or (_10847_, _10846_, _10845_);
  nor (_10848_, _10847_, _08651_);
  and (_10849_, _10847_, _08651_);
  nor (_10850_, _10849_, _10848_);
  not (_10851_, _10850_);
  nor (_10852_, _10843_, _07896_);
  nor (_10853_, _10852_, _10844_);
  nor (_10854_, _10853_, _10101_);
  and (_10855_, _10842_, _07934_);
  nor (_10856_, _10855_, _07928_);
  nor (_10857_, _10856_, _10843_);
  and (_10858_, _10857_, _10145_);
  nor (_10859_, _10857_, _10145_);
  nor (_10860_, _10842_, _07934_);
  nor (_10861_, _10860_, _10855_);
  nor (_10862_, _10861_, _10119_);
  nor (_10863_, _10862_, _10859_);
  nor (_10864_, _10863_, _10858_);
  nor (_10865_, _10859_, _10858_);
  not (_10866_, _10865_);
  and (_10867_, _10861_, _10119_);
  or (_10868_, _10867_, _10862_);
  or (_10869_, _10868_, _10866_);
  nor (_10870_, _08793_, _06589_);
  nor (_10871_, _10870_, _10842_);
  and (_10872_, _10871_, _10246_);
  nor (_10873_, _10871_, _10246_);
  nor (_10874_, _10873_, _10872_);
  nor (_10875_, _10841_, _07573_);
  or (_10876_, _10875_, _08793_);
  nor (_10877_, _10876_, \uc8051golden_1.ACC [2]);
  and (_10878_, _10876_, \uc8051golden_1.ACC [2]);
  nor (_10879_, _10878_, _10877_);
  and (_10880_, _10879_, _10874_);
  nor (_10881_, _06840_, _10524_);
  nor (_10882_, _10881_, _06229_);
  nor (_10883_, _10882_, _10841_);
  nor (_10884_, _10883_, _05984_);
  and (_10885_, _10883_, _05984_);
  and (_10886_, _06840_, _10524_);
  nor (_10887_, _10886_, _10881_);
  and (_10888_, _10887_, _06045_);
  nor (_10889_, _10888_, _10885_);
  or (_10890_, _10889_, _10884_);
  and (_10891_, _10890_, _10880_);
  and (_10892_, _10878_, _10874_);
  or (_10893_, _10892_, _10873_);
  nor (_10894_, _10893_, _10891_);
  nor (_10895_, _10894_, _10869_);
  nor (_10896_, _10895_, _10864_);
  and (_10897_, _10853_, _10101_);
  nor (_10898_, _10854_, _10897_);
  not (_10899_, _10898_);
  nor (_10900_, _10899_, _10896_);
  or (_10901_, _10900_, _10854_);
  and (_10902_, _10901_, _10851_);
  nor (_10903_, _10901_, _10851_);
  or (_10904_, _10903_, _10902_);
  and (_10905_, _10904_, _10572_);
  or (_10906_, _10905_, _06022_);
  or (_10907_, _10906_, _10840_);
  or (_10908_, _06194_, _06023_);
  and (_10909_, _10908_, _06446_);
  and (_10910_, _10909_, _10907_);
  and (_10911_, _08794_, _08616_);
  or (_10912_, _10911_, _10646_);
  and (_10913_, _10912_, _06300_);
  or (_10914_, _10913_, _10059_);
  or (_10915_, _10914_, _10910_);
  and (_10916_, _10915_, _10571_);
  or (_10917_, _10916_, _06281_);
  and (_10918_, _07995_, _08749_);
  or (_10919_, _10545_, _06282_);
  or (_10920_, _10919_, _10918_);
  and (_10921_, _10920_, _06279_);
  and (_10922_, _10921_, _10917_);
  and (_10923_, _09009_, _07995_);
  or (_10924_, _10923_, _10545_);
  and (_10925_, _10924_, _06015_);
  or (_10926_, _10925_, _10072_);
  or (_10927_, _10926_, _10922_);
  or (_10928_, _10092_, _10078_);
  and (_10929_, _10928_, _10927_);
  or (_10930_, _10929_, _05982_);
  and (_10931_, _10930_, _10567_);
  or (_10932_, _10931_, _06275_);
  and (_10933_, _06481_, _05942_);
  not (_10934_, _10933_);
  and (_10935_, _08813_, _07995_);
  or (_10936_, _10935_, _10545_);
  or (_10937_, _10936_, _06276_);
  and (_10938_, _10937_, _10934_);
  and (_10939_, _10938_, _10932_);
  and (_10940_, _10933_, _06194_);
  and (_10941_, _07378_, _05951_);
  or (_10942_, _10941_, _10940_);
  or (_10943_, _10942_, _10939_);
  not (_10944_, _10565_);
  not (_10945_, _10941_);
  or (_10946_, _10945_, _10563_);
  and (_10947_, _10946_, _10944_);
  and (_10948_, _10947_, _10943_);
  or (_10949_, _10948_, _10566_);
  and (_10950_, _06285_, _05951_);
  not (_10951_, _10950_);
  and (_10952_, _10951_, _10949_);
  and (_10953_, _06280_, _05951_);
  and (_10954_, _10950_, _10563_);
  or (_10955_, _10954_, _10953_);
  or (_10956_, _10955_, _10952_);
  and (_10957_, _09075_, _08651_);
  nor (_10958_, _10957_, _10558_);
  not (_10959_, _10953_);
  or (_10960_, _10959_, _10958_);
  and (_10961_, _10960_, _10956_);
  or (_10962_, _10961_, _06580_);
  and (_10963_, _06481_, _05951_);
  not (_10964_, _10963_);
  or (_10965_, _09034_, _06581_);
  and (_10966_, _10965_, _10964_);
  and (_10967_, _10966_, _10962_);
  nor (_10968_, _06194_, \uc8051golden_1.ACC [7]);
  and (_10969_, _06194_, \uc8051golden_1.ACC [7]);
  nor (_10970_, _10969_, _10968_);
  and (_10971_, _10963_, _10970_);
  or (_10972_, _10971_, _06474_);
  or (_10973_, _10972_, _10967_);
  and (_10974_, _09027_, _07995_);
  or (_10975_, _10974_, _10545_);
  or (_10976_, _10975_, _07282_);
  and (_10977_, _10976_, _10973_);
  or (_10978_, _10977_, _06582_);
  or (_10979_, _10545_, _07284_);
  nand (_10980_, _05955_, _05805_);
  and (_10981_, _10980_, _10979_);
  and (_10982_, _10981_, _10978_);
  not (_10983_, _10980_);
  and (_10984_, _10983_, _10562_);
  or (_10985_, _10984_, _10559_);
  or (_10986_, _10985_, _10982_);
  and (_10987_, _10986_, _10561_);
  or (_10988_, _10987_, _06567_);
  and (_10989_, _06481_, _05955_);
  not (_10990_, _10989_);
  or (_10991_, _09032_, _06568_);
  and (_10992_, _10991_, _10990_);
  and (_10993_, _10992_, _10988_);
  and (_10994_, _10989_, _10969_);
  or (_10995_, _10994_, _10993_);
  and (_10996_, _10995_, _07279_);
  nand (_10997_, _10936_, _06478_);
  nor (_10998_, _10997_, _09033_);
  or (_10999_, _10998_, _10556_);
  or (_11000_, _10999_, _10996_);
  and (_11001_, _11000_, _10557_);
  or (_11002_, _06955_, _06466_);
  and (_11003_, _11002_, _05946_);
  or (_11004_, _11003_, _11001_);
  and (_11005_, _06452_, _05946_);
  not (_11006_, _11005_);
  nand (_11007_, _11003_, _10549_);
  and (_11008_, _11007_, _11006_);
  and (_11009_, _11008_, _11004_);
  nor (_11010_, _10549_, _11006_);
  and (_11011_, _06280_, _05946_);
  or (_11012_, _11011_, _11010_);
  or (_11013_, _11012_, _11009_);
  nand (_11014_, _11011_, _10957_);
  and (_11015_, _11014_, _06575_);
  and (_11016_, _11015_, _11013_);
  and (_11017_, _06481_, _05946_);
  nor (_11018_, _11017_, _06574_);
  not (_11019_, _11018_);
  not (_11020_, _11017_);
  nand (_11021_, _11020_, _09033_);
  and (_11022_, _11021_, _11019_);
  or (_11023_, _11022_, _11016_);
  nand (_11024_, _11017_, _10968_);
  and (_11025_, _11024_, _09043_);
  and (_11026_, _11025_, _11023_);
  or (_11027_, _11026_, _10548_);
  nand (_11028_, _05965_, _05805_);
  and (_11029_, _11028_, _11027_);
  not (_11030_, _11028_);
  and (_11031_, _10753_, \uc8051golden_1.ACC [6]);
  and (_11032_, _10757_, \uc8051golden_1.ACC [5]);
  nand (_11033_, _10764_, \uc8051golden_1.ACC [4]);
  and (_11034_, _10771_, \uc8051golden_1.ACC [3]);
  and (_11035_, _10777_, \uc8051golden_1.ACC [2]);
  and (_11036_, _10785_, \uc8051golden_1.ACC [1]);
  nor (_11037_, _10787_, _10786_);
  not (_11038_, _11037_);
  and (_11039_, _10789_, \uc8051golden_1.ACC [0]);
  and (_11040_, _11039_, _11038_);
  nor (_11041_, _11040_, _11036_);
  nor (_11042_, _11041_, _10780_);
  nor (_11043_, _11042_, _11035_);
  nor (_11044_, _11043_, _10774_);
  or (_11045_, _11044_, _11034_);
  nand (_11046_, _11045_, _10767_);
  and (_11047_, _11046_, _11033_);
  nor (_11048_, _11047_, _10760_);
  or (_11049_, _11048_, _11032_);
  and (_11050_, _11049_, _10804_);
  nor (_11051_, _11050_, _11031_);
  nor (_11052_, _11051_, _10749_);
  and (_11053_, _11051_, _10749_);
  nor (_11054_, _11053_, _11052_);
  and (_11055_, _11054_, _11030_);
  or (_11056_, _11055_, _10471_);
  or (_11057_, _11056_, _11029_);
  and (_11058_, _11057_, _10544_);
  and (_11059_, _06481_, _05965_);
  nor (_11060_, _11059_, _06578_);
  not (_11061_, _11060_);
  and (_11062_, _10589_, \uc8051golden_1.ACC [6]);
  and (_11063_, _10592_, \uc8051golden_1.ACC [5]);
  nand (_11064_, _10596_, \uc8051golden_1.ACC [4]);
  and (_11065_, _10606_, \uc8051golden_1.ACC [3]);
  and (_11066_, _10611_, \uc8051golden_1.ACC [2]);
  and (_11067_, _10617_, \uc8051golden_1.ACC [1]);
  nor (_11068_, _10619_, _10618_);
  not (_11069_, _11068_);
  and (_11070_, _10621_, \uc8051golden_1.ACC [0]);
  and (_11071_, _11070_, _11069_);
  nor (_11072_, _11071_, _11067_);
  nor (_11073_, _11072_, _10614_);
  nor (_11074_, _11073_, _11066_);
  nor (_11075_, _11074_, _10609_);
  or (_11076_, _11075_, _11065_);
  nand (_11077_, _11076_, _10603_);
  and (_11078_, _11077_, _11064_);
  nor (_11079_, _11078_, _10600_);
  or (_11080_, _11079_, _11063_);
  and (_11081_, _11080_, _10633_);
  nor (_11082_, _11081_, _11062_);
  nor (_11083_, _11082_, _10586_);
  and (_11084_, _11082_, _10586_);
  nor (_11085_, _11084_, _11083_);
  or (_11086_, _11085_, _11059_);
  and (_11087_, _11086_, _11061_);
  or (_11088_, _11087_, _11058_);
  and (_11089_, _05981_, _05965_);
  not (_11090_, _11089_);
  not (_11091_, _11059_);
  nand (_11092_, _10853_, \uc8051golden_1.ACC [6]);
  and (_11093_, _10857_, \uc8051golden_1.ACC [5]);
  nand (_11094_, _10861_, \uc8051golden_1.ACC [4]);
  and (_11095_, _10871_, \uc8051golden_1.ACC [3]);
  nor (_11096_, _10876_, _10195_);
  and (_11097_, _10883_, \uc8051golden_1.ACC [1]);
  nor (_11098_, _10885_, _10884_);
  not (_11099_, _11098_);
  and (_11100_, _10887_, \uc8051golden_1.ACC [0]);
  and (_11101_, _11100_, _11099_);
  nor (_11102_, _11101_, _11097_);
  nor (_11103_, _11102_, _10879_);
  nor (_11104_, _11103_, _11096_);
  nor (_11105_, _11104_, _10874_);
  or (_11106_, _11105_, _11095_);
  nand (_11107_, _11106_, _10868_);
  and (_11108_, _11107_, _11094_);
  nor (_11109_, _11108_, _10865_);
  or (_11110_, _11109_, _11093_);
  nand (_11111_, _11110_, _10899_);
  and (_11112_, _11111_, _11092_);
  nor (_11113_, _11112_, _10850_);
  and (_11114_, _11112_, _10850_);
  nor (_11115_, _11114_, _11113_);
  or (_11116_, _11115_, _11091_);
  and (_11117_, _11116_, _11090_);
  and (_11118_, _11117_, _11088_);
  and (_11119_, _11089_, \uc8051golden_1.ACC [6]);
  nand (_11120_, _05970_, _05805_);
  not (_11121_, _11120_);
  or (_11122_, _11121_, _11119_);
  or (_11123_, _11122_, _11118_);
  nor (_11124_, _08118_, _10101_);
  not (_11125_, _11124_);
  and (_11126_, _08118_, _10101_);
  nor (_11127_, _11126_, _11124_);
  nor (_11128_, _08207_, _10145_);
  and (_11129_, _08207_, _10145_);
  nor (_11130_, _11129_, _11128_);
  nor (_11131_, _08301_, _10119_);
  not (_11132_, _11131_);
  nand (_11133_, _08301_, _10119_);
  and (_11134_, _11133_, _11132_);
  nor (_11135_, _07775_, _10246_);
  and (_11136_, _07775_, _10246_);
  nor (_11137_, _07623_, _10195_);
  and (_11138_, _07623_, _10195_);
  nor (_11139_, _11138_, _11137_);
  nor (_11140_, _07196_, _05984_);
  and (_11141_, _07196_, _05984_);
  nor (_11142_, _11141_, _11140_);
  and (_11143_, _07473_, \uc8051golden_1.ACC [0]);
  and (_11144_, _11143_, _11142_);
  nor (_11145_, _11144_, _11140_);
  not (_11146_, _11145_);
  and (_11147_, _11146_, _11139_);
  nor (_11148_, _11147_, _11137_);
  nor (_11149_, _11148_, _11136_);
  or (_11150_, _11149_, _11135_);
  and (_11151_, _11150_, _11134_);
  nor (_11152_, _11151_, _11131_);
  not (_11153_, _11152_);
  and (_11154_, _11153_, _11130_);
  or (_11155_, _11154_, _11128_);
  nand (_11156_, _11155_, _11127_);
  and (_11157_, _11156_, _11125_);
  nor (_11158_, _11157_, _10563_);
  and (_11159_, _11157_, _10563_);
  or (_11160_, _11159_, _11158_);
  or (_11161_, _11160_, _11120_);
  and (_11162_, _11161_, _11123_);
  and (_11163_, _06280_, _05970_);
  or (_11164_, _11163_, _11162_);
  not (_11165_, _11163_);
  and (_11166_, _09440_, \uc8051golden_1.ACC [6]);
  not (_11167_, _11166_);
  or (_11168_, _09440_, \uc8051golden_1.ACC [6]);
  and (_11169_, _11167_, _11168_);
  and (_11170_, _09441_, \uc8051golden_1.ACC [5]);
  and (_11171_, _09165_, _10145_);
  and (_11172_, _09442_, \uc8051golden_1.ACC [4]);
  not (_11173_, _11172_);
  or (_11174_, _09442_, \uc8051golden_1.ACC [4]);
  and (_11175_, _11173_, _11174_);
  and (_11176_, _09443_, \uc8051golden_1.ACC [3]);
  and (_11177_, _09255_, _10246_);
  and (_11178_, _09444_, \uc8051golden_1.ACC [2]);
  and (_11179_, _09300_, _10195_);
  nor (_11180_, _11178_, _11179_);
  not (_11181_, _11180_);
  and (_11182_, _09445_, \uc8051golden_1.ACC [1]);
  or (_11183_, _09445_, \uc8051golden_1.ACC [1]);
  not (_11184_, _11182_);
  and (_11185_, _11184_, _11183_);
  and (_11186_, _09446_, \uc8051golden_1.ACC [0]);
  and (_11187_, _11186_, _11185_);
  nor (_11188_, _11187_, _11182_);
  nor (_11189_, _11188_, _11181_);
  nor (_11190_, _11189_, _11178_);
  nor (_11191_, _11190_, _11177_);
  or (_11192_, _11191_, _11176_);
  nand (_11193_, _11192_, _11175_);
  and (_11194_, _11193_, _11173_);
  nor (_11195_, _11194_, _11171_);
  or (_11196_, _11195_, _11170_);
  nand (_11197_, _11196_, _11169_);
  and (_11198_, _11197_, _11167_);
  and (_11199_, _11198_, _10958_);
  nor (_11200_, _11198_, _10958_);
  or (_11201_, _11200_, _11199_);
  or (_11202_, _11201_, _11165_);
  and (_11203_, _06481_, _05970_);
  nor (_11204_, _11203_, _06307_);
  and (_11205_, _11204_, _11202_);
  and (_11206_, _11205_, _11164_);
  nor (_11207_, _08161_, _10101_);
  not (_11208_, _11207_);
  and (_11209_, _08161_, _10101_);
  nor (_11210_, _11209_, _11207_);
  nor (_11211_, _08255_, _10145_);
  and (_11212_, _08255_, _10145_);
  nor (_11213_, _08344_, _10119_);
  not (_11214_, _11213_);
  and (_11215_, _08344_, _10119_);
  nor (_11216_, _11215_, _11213_);
  nor (_11217_, _08388_, _10246_);
  and (_11218_, _08388_, _10246_);
  nor (_11219_, _08432_, _10195_);
  and (_11220_, _08432_, _10195_);
  nor (_11221_, _11220_, _11219_);
  nor (_11222_, _08476_, _05984_);
  and (_11223_, _08476_, _05984_);
  nor (_11224_, _11223_, _11222_);
  and (_11225_, _08521_, \uc8051golden_1.ACC [0]);
  and (_11226_, _11225_, _11224_);
  nor (_11227_, _11226_, _11222_);
  not (_11228_, _11227_);
  and (_11229_, _11228_, _11221_);
  nor (_11230_, _11229_, _11219_);
  nor (_11231_, _11230_, _11218_);
  or (_11232_, _11231_, _11217_);
  nand (_11233_, _11232_, _11216_);
  and (_11234_, _11233_, _11214_);
  nor (_11235_, _11234_, _11212_);
  or (_11236_, _11235_, _11211_);
  nand (_11237_, _11236_, _11210_);
  and (_11238_, _11237_, _11208_);
  nor (_11239_, _11238_, _09034_);
  and (_11240_, _11238_, _09034_);
  or (_11241_, _11240_, _11239_);
  and (_11242_, _11241_, _06307_);
  and (_11243_, _05981_, _05970_);
  nor (_11244_, _06340_, _10101_);
  and (_11245_, _06340_, _10101_);
  nor (_11246_, _11244_, _11245_);
  nor (_11247_, _06650_, _10145_);
  and (_11248_, _06650_, _10145_);
  nor (_11249_, _06265_, _10119_);
  not (_11250_, _11249_);
  and (_11251_, _06265_, _10119_);
  nor (_11252_, _11249_, _11251_);
  nor (_11253_, _06372_, _10246_);
  and (_11254_, _06372_, _10246_);
  nor (_11255_, _06693_, _10195_);
  and (_11256_, _06693_, _10195_);
  nor (_11257_, _11255_, _11256_);
  nor (_11258_, _06228_, _05984_);
  and (_11259_, _06228_, _05984_);
  nor (_11260_, _11258_, _11259_);
  nor (_11261_, _06840_, _06045_);
  and (_11262_, _11261_, _11260_);
  nor (_11263_, _11262_, _11258_);
  not (_11264_, _11263_);
  and (_11265_, _11264_, _11257_);
  nor (_11266_, _11265_, _11255_);
  nor (_11267_, _11266_, _11254_);
  or (_11268_, _11267_, _11253_);
  nand (_11269_, _11268_, _11252_);
  and (_11270_, _11269_, _11250_);
  nor (_11271_, _11270_, _11248_);
  or (_11272_, _11271_, _11247_);
  and (_11273_, _11272_, _11246_);
  nor (_11274_, _11273_, _11244_);
  nor (_11275_, _11274_, _10970_);
  and (_11276_, _11274_, _10970_);
  or (_11277_, _11276_, _11275_);
  and (_11278_, _11277_, _11203_);
  or (_11279_, _11278_, _11243_);
  or (_11280_, _11279_, _11242_);
  or (_11281_, _11280_, _11206_);
  nand (_11282_, _11243_, _10101_);
  and (_11283_, _11282_, _11281_);
  or (_11284_, _11283_, _06606_);
  and (_11285_, _06481_, _05968_);
  not (_11286_, _11285_);
  or (_11287_, _10652_, _07037_);
  and (_11288_, _11287_, _11286_);
  and (_11289_, _11288_, _11284_);
  and (_11290_, _05981_, _05968_);
  and (_11291_, _10681_, _06045_);
  and (_11292_, _11291_, _10246_);
  and (_11293_, _11292_, _10119_);
  and (_11294_, _11293_, _10145_);
  and (_11295_, _11294_, _10101_);
  nor (_11296_, _11295_, _08651_);
  and (_11297_, _11295_, _08651_);
  or (_11298_, _11297_, _11296_);
  and (_11299_, _11298_, _11285_);
  or (_11300_, _11299_, _11290_);
  or (_11301_, _11300_, _11289_);
  nand (_11302_, _11290_, _10524_);
  and (_11303_, _11302_, _06807_);
  and (_11304_, _11303_, _11301_);
  and (_11305_, _10725_, _06234_);
  or (_11306_, _11305_, _06195_);
  or (_11307_, _11306_, _11304_);
  and (_11308_, _06481_, _05962_);
  not (_11309_, _11308_);
  and (_11310_, _08530_, _07995_);
  or (_11311_, _11310_, _10545_);
  or (_11312_, _11311_, _06196_);
  and (_11313_, _11312_, _11309_);
  and (_11314_, _11313_, _11307_);
  and (_11315_, _05981_, _05962_);
  and (_11316_, \uc8051golden_1.ACC [1], \uc8051golden_1.ACC [0]);
  and (_11317_, _11316_, \uc8051golden_1.ACC [2]);
  and (_11318_, _11317_, \uc8051golden_1.ACC [3]);
  and (_11319_, _11318_, \uc8051golden_1.ACC [4]);
  and (_11320_, _11319_, \uc8051golden_1.ACC [5]);
  and (_11321_, _11320_, \uc8051golden_1.ACC [6]);
  nor (_11322_, _11321_, _08651_);
  and (_11323_, _11321_, _08651_);
  or (_11324_, _11323_, _11322_);
  and (_11325_, _11324_, _11308_);
  or (_11326_, _11325_, _11315_);
  or (_11327_, _11326_, _11314_);
  nand (_11328_, _11315_, _06045_);
  and (_11329_, _11328_, _01375_);
  and (_11330_, _11329_, _11327_);
  or (_11331_, _11330_, _10470_);
  and (_40324_, _11331_, _42545_);
  not (_11332_, _08002_);
  and (_11333_, _11332_, \uc8051golden_1.PCON [7]);
  and (_11334_, _09034_, _08002_);
  or (_11335_, _11334_, _11333_);
  and (_11336_, _11335_, _06582_);
  nor (_11337_, _11332_, _08070_);
  or (_11338_, _11337_, _11333_);
  or (_11339_, _11338_, _06293_);
  and (_11340_, _08762_, _08002_);
  or (_11341_, _11340_, _11333_);
  or (_11342_, _11341_, _07210_);
  and (_11343_, _08002_, \uc8051golden_1.ACC [7]);
  or (_11344_, _11343_, _11333_);
  and (_11345_, _11344_, _07199_);
  and (_11346_, _07200_, \uc8051golden_1.PCON [7]);
  or (_11347_, _11346_, _06401_);
  or (_11348_, _11347_, _11345_);
  and (_11349_, _11348_, _07221_);
  and (_11350_, _11349_, _11342_);
  and (_11351_, _11338_, _06399_);
  or (_11352_, _11351_, _11350_);
  and (_11353_, _11352_, _06414_);
  and (_11354_, _11344_, _06406_);
  or (_11355_, _11354_, _10059_);
  or (_11356_, _11355_, _11353_);
  and (_11357_, _11356_, _11339_);
  or (_11358_, _11357_, _06281_);
  and (_11359_, _08002_, _08749_);
  or (_11360_, _11333_, _06282_);
  or (_11361_, _11360_, _11359_);
  and (_11362_, _11361_, _06279_);
  and (_11363_, _11362_, _11358_);
  and (_11364_, _09009_, _08002_);
  or (_11365_, _11364_, _11333_);
  and (_11366_, _11365_, _06015_);
  or (_11367_, _11366_, _06275_);
  or (_11368_, _11367_, _11363_);
  and (_11369_, _08813_, _08002_);
  or (_11370_, _11369_, _11333_);
  or (_11371_, _11370_, _06276_);
  and (_11372_, _11371_, _11368_);
  or (_11373_, _11372_, _06474_);
  and (_11374_, _09027_, _08002_);
  or (_11375_, _11374_, _11333_);
  or (_11376_, _11375_, _07282_);
  and (_11377_, _11376_, _07284_);
  and (_11378_, _11377_, _11373_);
  or (_11379_, _11378_, _11336_);
  and (_11380_, _11379_, _07279_);
  or (_11381_, _11333_, _08073_);
  and (_11382_, _11370_, _06478_);
  and (_11383_, _11382_, _11381_);
  or (_11384_, _11383_, _11380_);
  and (_11385_, _11384_, _07276_);
  and (_11386_, _11344_, _06569_);
  and (_11387_, _11386_, _11381_);
  or (_11388_, _11387_, _06479_);
  or (_11389_, _11388_, _11385_);
  and (_11390_, _09026_, _08002_);
  or (_11391_, _11333_, _09043_);
  or (_11392_, _11391_, _11390_);
  and (_11393_, _11392_, _09048_);
  and (_11394_, _11393_, _11389_);
  nor (_11395_, _09033_, _11332_);
  or (_11396_, _11395_, _11333_);
  and (_11397_, _11396_, _06572_);
  or (_11398_, _11397_, _06606_);
  or (_11399_, _11398_, _11394_);
  or (_11400_, _11341_, _07037_);
  and (_11401_, _11400_, _06196_);
  and (_11402_, _11401_, _11399_);
  and (_11403_, _08530_, _08002_);
  or (_11404_, _11403_, _11333_);
  and (_11405_, _11404_, _06195_);
  or (_11406_, _11405_, _01379_);
  or (_11407_, _11406_, _11402_);
  or (_11408_, _01375_, \uc8051golden_1.PCON [7]);
  and (_11409_, _11408_, _42545_);
  and (_40325_, _11409_, _11407_);
  not (_11410_, _08006_);
  and (_11411_, _11410_, \uc8051golden_1.TMOD [7]);
  and (_11412_, _09034_, _08006_);
  or (_11413_, _11412_, _11411_);
  and (_11414_, _11413_, _06582_);
  nor (_11415_, _11410_, _08070_);
  or (_11416_, _11415_, _11411_);
  or (_11417_, _11416_, _06293_);
  and (_11418_, _08762_, _08006_);
  or (_11419_, _11418_, _11411_);
  or (_11420_, _11419_, _07210_);
  and (_11421_, _08006_, \uc8051golden_1.ACC [7]);
  or (_11422_, _11421_, _11411_);
  and (_11423_, _11422_, _07199_);
  and (_11424_, _07200_, \uc8051golden_1.TMOD [7]);
  or (_11425_, _11424_, _06401_);
  or (_11426_, _11425_, _11423_);
  and (_11427_, _11426_, _07221_);
  and (_11428_, _11427_, _11420_);
  and (_11429_, _11416_, _06399_);
  or (_11430_, _11429_, _11428_);
  and (_11431_, _11430_, _06414_);
  and (_11432_, _11422_, _06406_);
  or (_11433_, _11432_, _10059_);
  or (_11434_, _11433_, _11431_);
  and (_11435_, _11434_, _11417_);
  or (_11436_, _11435_, _06281_);
  and (_11437_, _08006_, _08749_);
  or (_11438_, _11411_, _06282_);
  or (_11439_, _11438_, _11437_);
  and (_11440_, _11439_, _06279_);
  and (_11441_, _11440_, _11436_);
  and (_11442_, _09009_, _08006_);
  or (_11443_, _11442_, _11411_);
  and (_11444_, _11443_, _06015_);
  or (_11445_, _11444_, _06275_);
  or (_11446_, _11445_, _11441_);
  and (_11447_, _08813_, _08006_);
  or (_11448_, _11447_, _11411_);
  or (_11449_, _11448_, _06276_);
  and (_11450_, _11449_, _11446_);
  or (_11451_, _11450_, _06474_);
  and (_11452_, _09027_, _08006_);
  or (_11453_, _11452_, _11411_);
  or (_11454_, _11453_, _07282_);
  and (_11455_, _11454_, _07284_);
  and (_11456_, _11455_, _11451_);
  or (_11457_, _11456_, _11414_);
  and (_11458_, _11457_, _07279_);
  or (_11459_, _11411_, _08073_);
  and (_11460_, _11448_, _06478_);
  and (_11461_, _11460_, _11459_);
  or (_11462_, _11461_, _11458_);
  and (_11463_, _11462_, _07276_);
  and (_11464_, _11422_, _06569_);
  and (_11465_, _11464_, _11459_);
  or (_11466_, _11465_, _06479_);
  or (_11467_, _11466_, _11463_);
  and (_11468_, _09026_, _08006_);
  or (_11469_, _11411_, _09043_);
  or (_11470_, _11469_, _11468_);
  and (_11471_, _11470_, _09048_);
  and (_11472_, _11471_, _11467_);
  nor (_11473_, _09033_, _11410_);
  or (_11474_, _11473_, _11411_);
  and (_11475_, _11474_, _06572_);
  or (_11476_, _11475_, _06606_);
  or (_11477_, _11476_, _11472_);
  or (_11478_, _11419_, _07037_);
  and (_11479_, _11478_, _06196_);
  and (_11480_, _11479_, _11477_);
  and (_11481_, _08530_, _08006_);
  or (_11482_, _11481_, _11411_);
  and (_11483_, _11482_, _06195_);
  or (_11484_, _11483_, _01379_);
  or (_11485_, _11484_, _11480_);
  or (_11486_, _01375_, \uc8051golden_1.TMOD [7]);
  and (_11487_, _11486_, _42545_);
  and (_40326_, _11487_, _11485_);
  not (_11488_, \uc8051golden_1.DPL [7]);
  nor (_11489_, _07962_, _11488_);
  and (_11490_, _09034_, _07962_);
  or (_11491_, _11490_, _11489_);
  and (_11492_, _11491_, _06582_);
  not (_11493_, _07962_);
  nor (_11494_, _11493_, _08070_);
  or (_11495_, _11494_, _11489_);
  or (_11496_, _11495_, _06293_);
  and (_11497_, _08762_, _07962_);
  or (_11498_, _11497_, _11489_);
  or (_11499_, _11498_, _07210_);
  and (_11500_, _07962_, \uc8051golden_1.ACC [7]);
  or (_11501_, _11500_, _11489_);
  and (_11502_, _11501_, _07199_);
  nor (_11503_, _07199_, _11488_);
  or (_11504_, _11503_, _06401_);
  or (_11505_, _11504_, _11502_);
  and (_11506_, _11505_, _07221_);
  and (_11507_, _11506_, _11499_);
  and (_11508_, _11495_, _06399_);
  or (_11509_, _11508_, _06406_);
  or (_11510_, _11509_, _11507_);
  and (_11511_, _06381_, _05981_);
  not (_11512_, _11511_);
  or (_11513_, _11501_, _06414_);
  and (_11514_, _11513_, _11512_);
  and (_11515_, _11514_, _11510_);
  and (_11516_, \uc8051golden_1.DPL [1], \uc8051golden_1.DPL [0]);
  and (_11517_, _11516_, \uc8051golden_1.DPL [2]);
  and (_11518_, _11517_, \uc8051golden_1.DPL [3]);
  and (_11519_, _11518_, \uc8051golden_1.DPL [4]);
  and (_11520_, _11519_, \uc8051golden_1.DPL [5]);
  and (_11521_, _11520_, \uc8051golden_1.DPL [6]);
  nor (_11522_, _11521_, \uc8051golden_1.DPL [7]);
  and (_11523_, _11521_, \uc8051golden_1.DPL [7]);
  nor (_11524_, _11523_, _11522_);
  and (_11525_, _11524_, _11511_);
  or (_11526_, _11525_, _11515_);
  and (_11527_, _11526_, _06473_);
  nor (_11528_, _08590_, _06473_);
  or (_11529_, _11528_, _10059_);
  or (_11530_, _11529_, _11527_);
  and (_11531_, _11530_, _11496_);
  or (_11532_, _11531_, _06281_);
  and (_11533_, _07962_, _08749_);
  or (_11534_, _11489_, _06282_);
  or (_11535_, _11534_, _11533_);
  and (_11536_, _11535_, _06279_);
  and (_11537_, _11536_, _11532_);
  and (_11538_, _09009_, _07962_);
  or (_11539_, _11538_, _11489_);
  and (_11540_, _11539_, _06015_);
  or (_11541_, _11540_, _06275_);
  or (_11542_, _11541_, _11537_);
  and (_11543_, _08813_, _07962_);
  or (_11544_, _11543_, _11489_);
  or (_11545_, _11544_, _06276_);
  and (_11546_, _11545_, _11542_);
  or (_11547_, _11546_, _06474_);
  and (_11548_, _09027_, _07962_);
  or (_11549_, _11548_, _11489_);
  or (_11550_, _11549_, _07282_);
  and (_11551_, _11550_, _07284_);
  and (_11552_, _11551_, _11547_);
  or (_11553_, _11552_, _11492_);
  and (_11554_, _11553_, _07279_);
  or (_11555_, _11489_, _08073_);
  and (_11556_, _11544_, _06478_);
  and (_11557_, _11556_, _11555_);
  or (_11558_, _11557_, _11554_);
  and (_11559_, _11558_, _07276_);
  and (_11560_, _11501_, _06569_);
  and (_11561_, _11560_, _11555_);
  or (_11562_, _11561_, _06479_);
  or (_11563_, _11562_, _11559_);
  and (_11564_, _09026_, _07962_);
  or (_11565_, _11489_, _09043_);
  or (_11566_, _11565_, _11564_);
  and (_11567_, _11566_, _09048_);
  and (_11568_, _11567_, _11563_);
  nor (_11569_, _09033_, _11493_);
  or (_11570_, _11569_, _11489_);
  and (_11571_, _11570_, _06572_);
  or (_11572_, _11571_, _06606_);
  or (_11573_, _11572_, _11568_);
  or (_11574_, _11498_, _07037_);
  and (_11575_, _11574_, _06196_);
  and (_11576_, _11575_, _11573_);
  and (_11577_, _08530_, _07962_);
  or (_11578_, _11577_, _11489_);
  and (_11579_, _11578_, _06195_);
  or (_11580_, _11579_, _01379_);
  or (_11581_, _11580_, _11576_);
  or (_11582_, _01375_, \uc8051golden_1.DPL [7]);
  and (_11583_, _11582_, _42545_);
  and (_40328_, _11583_, _11581_);
  not (_11584_, \uc8051golden_1.DPH [7]);
  nor (_11585_, _07966_, _11584_);
  and (_11586_, _09034_, _08249_);
  or (_11587_, _11586_, _11585_);
  and (_11588_, _11587_, _06582_);
  not (_11589_, _08249_);
  nor (_11590_, _11589_, _08070_);
  or (_11591_, _11590_, _11585_);
  or (_11592_, _11591_, _06293_);
  and (_11593_, _08762_, _08249_);
  or (_11594_, _11593_, _11585_);
  or (_11595_, _11594_, _07210_);
  and (_11596_, _07966_, \uc8051golden_1.ACC [7]);
  or (_11597_, _11596_, _11585_);
  and (_11598_, _11597_, _07199_);
  nor (_11599_, _07199_, _11584_);
  or (_11600_, _11599_, _06401_);
  or (_11601_, _11600_, _11598_);
  and (_11602_, _11601_, _07221_);
  and (_11603_, _11602_, _11595_);
  and (_11604_, _11591_, _06399_);
  or (_11605_, _11604_, _06406_);
  or (_11606_, _11605_, _11603_);
  or (_11607_, _11597_, _06414_);
  and (_11608_, _11607_, _11512_);
  and (_11609_, _11608_, _11606_);
  and (_11610_, _11523_, \uc8051golden_1.DPH [0]);
  and (_11611_, _11610_, \uc8051golden_1.DPH [1]);
  and (_11612_, _11611_, \uc8051golden_1.DPH [2]);
  and (_11613_, _11612_, \uc8051golden_1.DPH [3]);
  and (_11614_, _11613_, \uc8051golden_1.DPH [4]);
  and (_11615_, _11614_, \uc8051golden_1.DPH [5]);
  and (_11616_, _11615_, \uc8051golden_1.DPH [6]);
  nor (_11617_, _11616_, _11584_);
  and (_11618_, _11616_, _11584_);
  or (_11619_, _11618_, _11617_);
  and (_11620_, _11619_, _11511_);
  or (_11621_, _11620_, _11609_);
  and (_11622_, _11621_, _06473_);
  and (_11623_, _06472_, _06194_);
  or (_11624_, _11623_, _10059_);
  or (_11625_, _11624_, _11622_);
  and (_11626_, _11625_, _11592_);
  or (_11627_, _11626_, _06281_);
  or (_11628_, _11585_, _06282_);
  and (_11629_, _07966_, _08749_);
  or (_11630_, _11629_, _11628_);
  and (_11631_, _11630_, _06279_);
  and (_11632_, _11631_, _11627_);
  and (_11633_, _09009_, _08249_);
  or (_11634_, _11633_, _11585_);
  and (_11635_, _11634_, _06015_);
  or (_11636_, _11635_, _06275_);
  or (_11637_, _11636_, _11632_);
  and (_11638_, _08813_, _07966_);
  or (_11639_, _11638_, _11585_);
  or (_11640_, _11639_, _06276_);
  and (_11641_, _11640_, _11637_);
  or (_11642_, _11641_, _06474_);
  and (_11643_, _09027_, _07966_);
  or (_11644_, _11643_, _11585_);
  or (_11645_, _11644_, _07282_);
  and (_11646_, _11645_, _07284_);
  and (_11647_, _11646_, _11642_);
  or (_11648_, _11647_, _11588_);
  and (_11649_, _11648_, _07279_);
  or (_11650_, _11585_, _08073_);
  and (_11651_, _11639_, _06478_);
  and (_11652_, _11651_, _11650_);
  or (_11653_, _11652_, _11649_);
  and (_11654_, _11653_, _07276_);
  and (_11655_, _11597_, _06569_);
  and (_11656_, _11655_, _11650_);
  or (_11657_, _11656_, _06479_);
  or (_11658_, _11657_, _11654_);
  and (_11659_, _09026_, _08249_);
  or (_11660_, _11585_, _09043_);
  or (_11661_, _11660_, _11659_);
  and (_11662_, _11661_, _09048_);
  and (_11663_, _11662_, _11658_);
  nor (_11664_, _09033_, _11589_);
  or (_11665_, _11664_, _11585_);
  and (_11666_, _11665_, _06572_);
  or (_11667_, _11666_, _06606_);
  or (_11668_, _11667_, _11663_);
  or (_11669_, _11594_, _07037_);
  and (_11670_, _11669_, _06196_);
  and (_11671_, _11670_, _11668_);
  and (_11672_, _08530_, _08249_);
  or (_11673_, _11672_, _11585_);
  and (_11674_, _11673_, _06195_);
  or (_11675_, _11674_, _01379_);
  or (_11676_, _11675_, _11671_);
  or (_11677_, _01375_, \uc8051golden_1.DPH [7]);
  and (_11678_, _11677_, _42545_);
  and (_40329_, _11678_, _11676_);
  not (_11679_, _07976_);
  and (_11680_, _11679_, \uc8051golden_1.TL1 [7]);
  and (_11681_, _09034_, _07976_);
  or (_11682_, _11681_, _11680_);
  and (_11683_, _11682_, _06582_);
  and (_11684_, _08762_, _07976_);
  or (_11685_, _11684_, _11680_);
  or (_11686_, _11685_, _07210_);
  and (_11687_, _07976_, \uc8051golden_1.ACC [7]);
  or (_11688_, _11687_, _11680_);
  and (_11689_, _11688_, _07199_);
  and (_11690_, _07200_, \uc8051golden_1.TL1 [7]);
  or (_11691_, _11690_, _06401_);
  or (_11692_, _11691_, _11689_);
  and (_11693_, _11692_, _07221_);
  and (_11694_, _11693_, _11686_);
  nor (_11695_, _11679_, _08070_);
  or (_11696_, _11695_, _11680_);
  and (_11697_, _11696_, _06399_);
  or (_11698_, _11697_, _11694_);
  and (_11699_, _11698_, _06414_);
  and (_11700_, _11688_, _06406_);
  or (_11701_, _11700_, _10059_);
  or (_11702_, _11701_, _11699_);
  or (_11703_, _11696_, _06293_);
  and (_11704_, _11703_, _11702_);
  or (_11705_, _11704_, _06281_);
  and (_11706_, _07976_, _08749_);
  or (_11707_, _11680_, _06282_);
  or (_11708_, _11707_, _11706_);
  and (_11709_, _11708_, _06279_);
  and (_11710_, _11709_, _11705_);
  and (_11711_, _09009_, _07976_);
  or (_11712_, _11711_, _11680_);
  and (_11713_, _11712_, _06015_);
  or (_11714_, _11713_, _06275_);
  or (_11715_, _11714_, _11710_);
  and (_11716_, _08813_, _07976_);
  or (_11717_, _11716_, _11680_);
  or (_11718_, _11717_, _06276_);
  and (_11719_, _11718_, _11715_);
  or (_11720_, _11719_, _06474_);
  and (_11721_, _09027_, _07976_);
  or (_11722_, _11721_, _11680_);
  or (_11723_, _11722_, _07282_);
  and (_11724_, _11723_, _07284_);
  and (_11725_, _11724_, _11720_);
  or (_11726_, _11725_, _11683_);
  and (_11727_, _11726_, _07279_);
  or (_11728_, _11680_, _08073_);
  and (_11729_, _11717_, _06478_);
  and (_11730_, _11729_, _11728_);
  or (_11731_, _11730_, _11727_);
  and (_11732_, _11731_, _07276_);
  and (_11733_, _11688_, _06569_);
  and (_11734_, _11733_, _11728_);
  or (_11735_, _11734_, _06479_);
  or (_11736_, _11735_, _11732_);
  and (_11737_, _09026_, _07976_);
  or (_11738_, _11680_, _09043_);
  or (_11739_, _11738_, _11737_);
  and (_11740_, _11739_, _09048_);
  and (_11741_, _11740_, _11736_);
  nor (_11742_, _09033_, _11679_);
  or (_11743_, _11742_, _11680_);
  and (_11744_, _11743_, _06572_);
  or (_11745_, _11744_, _06606_);
  or (_11746_, _11745_, _11741_);
  or (_11747_, _11685_, _07037_);
  and (_11748_, _11747_, _06196_);
  and (_11749_, _11748_, _11746_);
  and (_11750_, _08530_, _07976_);
  or (_11751_, _11750_, _11680_);
  and (_11752_, _11751_, _06195_);
  or (_11753_, _11752_, _01379_);
  or (_11754_, _11753_, _11749_);
  or (_11755_, _01375_, \uc8051golden_1.TL1 [7]);
  and (_11756_, _11755_, _42545_);
  and (_40330_, _11756_, _11754_);
  not (_11757_, _08010_);
  and (_11758_, _11757_, \uc8051golden_1.TL0 [7]);
  and (_11759_, _09034_, _08010_);
  or (_11760_, _11759_, _11758_);
  and (_11761_, _11760_, _06582_);
  nor (_11762_, _11757_, _08070_);
  or (_11763_, _11762_, _11758_);
  or (_11764_, _11763_, _06293_);
  and (_11765_, _08762_, _08010_);
  or (_11766_, _11765_, _11758_);
  or (_11767_, _11766_, _07210_);
  and (_11768_, _08010_, \uc8051golden_1.ACC [7]);
  or (_11769_, _11768_, _11758_);
  and (_11770_, _11769_, _07199_);
  and (_11771_, _07200_, \uc8051golden_1.TL0 [7]);
  or (_11772_, _11771_, _06401_);
  or (_11773_, _11772_, _11770_);
  and (_11774_, _11773_, _07221_);
  and (_11775_, _11774_, _11767_);
  and (_11776_, _11763_, _06399_);
  or (_11777_, _11776_, _11775_);
  and (_11778_, _11777_, _06414_);
  and (_11779_, _11769_, _06406_);
  or (_11780_, _11779_, _10059_);
  or (_11781_, _11780_, _11778_);
  and (_11782_, _11781_, _11764_);
  or (_11783_, _11782_, _06281_);
  and (_11784_, _08010_, _08749_);
  or (_11785_, _11758_, _06282_);
  or (_11786_, _11785_, _11784_);
  and (_11787_, _11786_, _06279_);
  and (_11788_, _11787_, _11783_);
  and (_11789_, _09009_, _08010_);
  or (_11790_, _11789_, _11758_);
  and (_11791_, _11790_, _06015_);
  or (_11792_, _11791_, _06275_);
  or (_11793_, _11792_, _11788_);
  and (_11794_, _08813_, _08010_);
  or (_11795_, _11794_, _11758_);
  or (_11796_, _11795_, _06276_);
  and (_11797_, _11796_, _11793_);
  or (_11798_, _11797_, _06474_);
  and (_11799_, _09027_, _08010_);
  or (_11800_, _11799_, _11758_);
  or (_11801_, _11800_, _07282_);
  and (_11802_, _11801_, _07284_);
  and (_11803_, _11802_, _11798_);
  or (_11804_, _11803_, _11761_);
  and (_11805_, _11804_, _07279_);
  or (_11806_, _11758_, _08073_);
  and (_11807_, _11795_, _06478_);
  and (_11808_, _11807_, _11806_);
  or (_11809_, _11808_, _11805_);
  and (_11810_, _11809_, _07276_);
  and (_11811_, _11769_, _06569_);
  and (_11812_, _11811_, _11806_);
  or (_11813_, _11812_, _06479_);
  or (_11814_, _11813_, _11810_);
  and (_11815_, _09026_, _08010_);
  or (_11816_, _11758_, _09043_);
  or (_11817_, _11816_, _11815_);
  and (_11818_, _11817_, _09048_);
  and (_11819_, _11818_, _11814_);
  nor (_11820_, _09033_, _11757_);
  or (_11821_, _11820_, _11758_);
  and (_11822_, _11821_, _06572_);
  or (_11823_, _11822_, _06606_);
  or (_11824_, _11823_, _11819_);
  or (_11825_, _11766_, _07037_);
  and (_11826_, _11825_, _06196_);
  and (_11827_, _11826_, _11824_);
  and (_11828_, _08530_, _08010_);
  or (_11829_, _11828_, _11758_);
  and (_11830_, _11829_, _06195_);
  or (_11831_, _11830_, _01379_);
  or (_11832_, _11831_, _11827_);
  or (_11833_, _01375_, \uc8051golden_1.TL0 [7]);
  and (_11834_, _11833_, _42545_);
  and (_40331_, _11834_, _11832_);
  and (_11835_, _01379_, \uc8051golden_1.TCON [7]);
  not (_11836_, _08017_);
  and (_11837_, _11836_, \uc8051golden_1.TCON [7]);
  and (_11838_, _09034_, _08017_);
  or (_11839_, _11838_, _11837_);
  and (_11840_, _11839_, _06582_);
  nor (_11841_, _11836_, _08070_);
  or (_11842_, _11841_, _11837_);
  or (_11843_, _11842_, _06293_);
  not (_11844_, _08623_);
  and (_11845_, _11844_, \uc8051golden_1.TCON [7]);
  and (_11846_, _08639_, _08623_);
  or (_11847_, _11846_, _11845_);
  and (_11848_, _11847_, _06393_);
  and (_11849_, _08762_, _08017_);
  or (_11850_, _11849_, _11837_);
  or (_11851_, _11850_, _07210_);
  and (_11852_, _08017_, \uc8051golden_1.ACC [7]);
  or (_11853_, _11852_, _11837_);
  and (_11854_, _11853_, _07199_);
  and (_11855_, _07200_, \uc8051golden_1.TCON [7]);
  or (_11856_, _11855_, _06401_);
  or (_11857_, _11856_, _11854_);
  and (_11858_, _11857_, _06396_);
  and (_11859_, _11858_, _11851_);
  and (_11860_, _08635_, _08623_);
  or (_11861_, _11860_, _11845_);
  and (_11862_, _11861_, _06395_);
  or (_11863_, _11862_, _06399_);
  or (_11864_, _11863_, _11859_);
  or (_11865_, _11842_, _07221_);
  and (_11866_, _11865_, _11864_);
  or (_11867_, _11866_, _06406_);
  or (_11868_, _11853_, _06414_);
  and (_11869_, _11868_, _06844_);
  and (_11870_, _11869_, _11867_);
  or (_11871_, _11870_, _11848_);
  and (_11872_, _11871_, _07245_);
  and (_11873_, _08636_, _08623_);
  or (_11874_, _11873_, _11845_);
  and (_11875_, _11874_, _06387_);
  or (_11876_, _11875_, _11872_);
  and (_11877_, _11876_, _06446_);
  and (_11878_, _08794_, _08623_);
  or (_11879_, _11878_, _11845_);
  and (_11880_, _11879_, _06300_);
  or (_11881_, _11880_, _10059_);
  or (_11882_, _11881_, _11877_);
  and (_11883_, _11882_, _11843_);
  or (_11884_, _11883_, _06281_);
  and (_11885_, _08017_, _08749_);
  or (_11886_, _11837_, _06282_);
  or (_11887_, _11886_, _11885_);
  and (_11888_, _11887_, _06279_);
  and (_11889_, _11888_, _11884_);
  and (_11890_, _09009_, _08017_);
  or (_11891_, _11890_, _11837_);
  and (_11892_, _11891_, _06015_);
  or (_11893_, _11892_, _06275_);
  or (_11894_, _11893_, _11889_);
  and (_11895_, _08813_, _08017_);
  or (_11896_, _11895_, _11837_);
  or (_11897_, _11896_, _06276_);
  and (_11898_, _11897_, _11894_);
  or (_11899_, _11898_, _06474_);
  and (_11900_, _09027_, _08017_);
  or (_11901_, _11900_, _11837_);
  or (_11902_, _11901_, _07282_);
  and (_11903_, _11902_, _07284_);
  and (_11904_, _11903_, _11899_);
  or (_11905_, _11904_, _11840_);
  and (_11906_, _11905_, _07279_);
  or (_11907_, _11837_, _08073_);
  and (_11908_, _11896_, _06478_);
  and (_11909_, _11908_, _11907_);
  or (_11910_, _11909_, _11906_);
  and (_11911_, _11910_, _07276_);
  and (_11912_, _11853_, _06569_);
  and (_11913_, _11912_, _11907_);
  or (_11914_, _11913_, _06479_);
  or (_11915_, _11914_, _11911_);
  and (_11916_, _09026_, _08017_);
  or (_11917_, _11837_, _09043_);
  or (_11918_, _11917_, _11916_);
  and (_11919_, _11918_, _09048_);
  and (_11920_, _11919_, _11915_);
  nor (_11921_, _09033_, _11836_);
  or (_11922_, _11921_, _11837_);
  and (_11923_, _11922_, _06572_);
  or (_11924_, _11923_, _06606_);
  or (_11925_, _11924_, _11920_);
  or (_11926_, _11850_, _07037_);
  and (_11927_, _11926_, _06807_);
  and (_11928_, _11927_, _11925_);
  and (_11929_, _11847_, _06234_);
  or (_11930_, _11929_, _06195_);
  or (_11931_, _11930_, _11928_);
  and (_11932_, _08530_, _08017_);
  or (_11933_, _11837_, _06196_);
  or (_11934_, _11933_, _11932_);
  and (_11935_, _11934_, _01375_);
  and (_11936_, _11935_, _11931_);
  or (_11937_, _11936_, _11835_);
  and (_40332_, _11937_, _42545_);
  not (_11938_, _07980_);
  and (_11939_, _11938_, \uc8051golden_1.TH1 [7]);
  and (_11940_, _09034_, _07980_);
  or (_11941_, _11940_, _11939_);
  and (_11942_, _11941_, _06582_);
  and (_11943_, _08762_, _07980_);
  or (_11944_, _11943_, _11939_);
  or (_11945_, _11944_, _07210_);
  and (_11946_, _07980_, \uc8051golden_1.ACC [7]);
  or (_11947_, _11946_, _11939_);
  and (_11948_, _11947_, _07199_);
  and (_11949_, _07200_, \uc8051golden_1.TH1 [7]);
  or (_11950_, _11949_, _06401_);
  or (_11951_, _11950_, _11948_);
  and (_11952_, _11951_, _07221_);
  and (_11953_, _11952_, _11945_);
  nor (_11954_, _11938_, _08070_);
  or (_11955_, _11954_, _11939_);
  and (_11956_, _11955_, _06399_);
  or (_11957_, _11956_, _11953_);
  and (_11958_, _11957_, _06414_);
  and (_11959_, _11947_, _06406_);
  or (_11960_, _11959_, _10059_);
  or (_11961_, _11960_, _11958_);
  or (_11962_, _11955_, _06293_);
  and (_11963_, _11962_, _11961_);
  or (_11964_, _11963_, _06281_);
  and (_11965_, _07980_, _08749_);
  or (_11966_, _11939_, _06282_);
  or (_11967_, _11966_, _11965_);
  and (_11968_, _11967_, _06279_);
  and (_11969_, _11968_, _11964_);
  and (_11970_, _09009_, _07980_);
  or (_11971_, _11970_, _11939_);
  and (_11972_, _11971_, _06015_);
  or (_11973_, _11972_, _06275_);
  or (_11974_, _11973_, _11969_);
  and (_11975_, _08813_, _07980_);
  or (_11976_, _11975_, _11939_);
  or (_11977_, _11976_, _06276_);
  and (_11978_, _11977_, _11974_);
  or (_11979_, _11978_, _06474_);
  and (_11980_, _09027_, _07980_);
  or (_11981_, _11980_, _11939_);
  or (_11982_, _11981_, _07282_);
  and (_11983_, _11982_, _07284_);
  and (_11984_, _11983_, _11979_);
  or (_11985_, _11984_, _11942_);
  and (_11986_, _11985_, _07279_);
  or (_11987_, _11939_, _08073_);
  and (_11988_, _11976_, _06478_);
  and (_11989_, _11988_, _11987_);
  or (_11990_, _11989_, _11986_);
  and (_11991_, _11990_, _07276_);
  and (_11992_, _11947_, _06569_);
  and (_11993_, _11992_, _11987_);
  or (_11994_, _11993_, _06479_);
  or (_11995_, _11994_, _11991_);
  and (_11996_, _09026_, _07980_);
  or (_11997_, _11939_, _09043_);
  or (_11998_, _11997_, _11996_);
  and (_11999_, _11998_, _09048_);
  and (_12000_, _11999_, _11995_);
  nor (_12001_, _09033_, _11938_);
  or (_12002_, _12001_, _11939_);
  and (_12003_, _12002_, _06572_);
  or (_12004_, _12003_, _06606_);
  or (_12005_, _12004_, _12000_);
  or (_12006_, _11944_, _07037_);
  and (_12007_, _12006_, _06196_);
  and (_12008_, _12007_, _12005_);
  and (_12009_, _08530_, _07980_);
  or (_12010_, _12009_, _11939_);
  and (_12011_, _12010_, _06195_);
  or (_12012_, _12011_, _01379_);
  or (_12013_, _12012_, _12008_);
  or (_12014_, _01375_, \uc8051golden_1.TH1 [7]);
  and (_12015_, _12014_, _42545_);
  and (_40334_, _12015_, _12013_);
  not (_12016_, _08013_);
  and (_12017_, _12016_, \uc8051golden_1.TH0 [7]);
  and (_12018_, _09034_, _08013_);
  or (_12019_, _12018_, _12017_);
  and (_12020_, _12019_, _06582_);
  and (_12021_, _08762_, _08013_);
  or (_12022_, _12021_, _12017_);
  or (_12023_, _12022_, _07210_);
  and (_12024_, _08013_, \uc8051golden_1.ACC [7]);
  or (_12025_, _12024_, _12017_);
  and (_12026_, _12025_, _07199_);
  and (_12027_, _07200_, \uc8051golden_1.TH0 [7]);
  or (_12028_, _12027_, _06401_);
  or (_12029_, _12028_, _12026_);
  and (_12030_, _12029_, _07221_);
  and (_12031_, _12030_, _12023_);
  nor (_12032_, _12016_, _08070_);
  or (_12033_, _12032_, _12017_);
  and (_12034_, _12033_, _06399_);
  or (_12035_, _12034_, _12031_);
  and (_12036_, _12035_, _06414_);
  and (_12037_, _12025_, _06406_);
  or (_12038_, _12037_, _10059_);
  or (_12039_, _12038_, _12036_);
  or (_12040_, _12033_, _06293_);
  and (_12041_, _12040_, _12039_);
  or (_12042_, _12041_, _06281_);
  and (_12043_, _08013_, _08749_);
  or (_12044_, _12017_, _06282_);
  or (_12045_, _12044_, _12043_);
  and (_12046_, _12045_, _06279_);
  and (_12047_, _12046_, _12042_);
  and (_12048_, _09009_, _08013_);
  or (_12049_, _12048_, _12017_);
  and (_12050_, _12049_, _06015_);
  or (_12051_, _12050_, _06275_);
  or (_12052_, _12051_, _12047_);
  and (_12053_, _08813_, _08013_);
  or (_12054_, _12053_, _12017_);
  or (_12055_, _12054_, _06276_);
  and (_12056_, _12055_, _12052_);
  or (_12057_, _12056_, _06474_);
  and (_12058_, _09027_, _08013_);
  or (_12059_, _12058_, _12017_);
  or (_12060_, _12059_, _07282_);
  and (_12061_, _12060_, _07284_);
  and (_12062_, _12061_, _12057_);
  or (_12063_, _12062_, _12020_);
  and (_12064_, _12063_, _07279_);
  or (_12065_, _12017_, _08073_);
  and (_12066_, _12054_, _06478_);
  and (_12067_, _12066_, _12065_);
  or (_12068_, _12067_, _12064_);
  and (_12069_, _12068_, _07276_);
  and (_12070_, _12025_, _06569_);
  and (_12071_, _12070_, _12065_);
  or (_12072_, _12071_, _06479_);
  or (_12073_, _12072_, _12069_);
  and (_12074_, _09026_, _08013_);
  or (_12075_, _12017_, _09043_);
  or (_12076_, _12075_, _12074_);
  and (_12077_, _12076_, _09048_);
  and (_12078_, _12077_, _12073_);
  nor (_12079_, _09033_, _12016_);
  or (_12080_, _12079_, _12017_);
  and (_12081_, _12080_, _06572_);
  or (_12082_, _12081_, _06606_);
  or (_12083_, _12082_, _12078_);
  or (_12084_, _12022_, _07037_);
  and (_12085_, _12084_, _06196_);
  and (_12086_, _12085_, _12083_);
  and (_12087_, _08530_, _08013_);
  or (_12088_, _12087_, _12017_);
  and (_12089_, _12088_, _06195_);
  or (_12090_, _12089_, _01379_);
  or (_12091_, _12090_, _12086_);
  or (_12092_, _01375_, \uc8051golden_1.TH0 [7]);
  and (_12093_, _12092_, _42545_);
  and (_40335_, _12093_, _12091_);
  not (_12094_, _11204_);
  not (_12095_, _05672_);
  and (_12096_, _08533_, _12095_);
  and (_12097_, _12096_, \uc8051golden_1.PC [7]);
  and (_12098_, _12097_, \uc8051golden_1.PC [8]);
  and (_12099_, _12098_, \uc8051golden_1.PC [9]);
  and (_12100_, _12099_, \uc8051golden_1.PC [10]);
  and (_12101_, _12100_, \uc8051golden_1.PC [11]);
  and (_12102_, _12101_, \uc8051golden_1.PC [12]);
  and (_12103_, _12102_, \uc8051golden_1.PC [13]);
  and (_12104_, _12103_, \uc8051golden_1.PC [14]);
  or (_12105_, _12104_, \uc8051golden_1.PC [15]);
  nand (_12106_, _12104_, \uc8051golden_1.PC [15]);
  and (_12107_, _12106_, _12105_);
  and (_12108_, _11165_, _11120_);
  or (_12109_, _12108_, _12107_);
  nor (_12110_, _09469_, \uc8051golden_1.PC [14]);
  nor (_12111_, _12110_, _09470_);
  and (_12112_, _12111_, _06194_);
  nor (_12113_, _12111_, _06194_);
  nor (_12114_, _12113_, _12112_);
  not (_12115_, _12114_);
  nor (_12116_, _09468_, \uc8051golden_1.PC [13]);
  nor (_12117_, _12116_, _09469_);
  and (_12118_, _12117_, _06194_);
  nor (_12119_, _12117_, _06194_);
  nor (_12120_, _09467_, \uc8051golden_1.PC [12]);
  nor (_12121_, _12120_, _09468_);
  and (_12122_, _12121_, _06194_);
  nor (_12123_, _09473_, \uc8051golden_1.PC [10]);
  nor (_12124_, _12123_, _09466_);
  and (_12125_, _12124_, _06194_);
  not (_12126_, _12125_);
  nor (_12127_, _09474_, \uc8051golden_1.PC [11]);
  nor (_12128_, _12127_, _09475_);
  and (_12129_, _12128_, _06194_);
  nor (_12130_, _12128_, _06194_);
  nor (_12131_, _12130_, _12129_);
  nor (_12132_, _12124_, _06194_);
  nor (_12133_, _12132_, _12125_);
  and (_12134_, _12133_, _12131_);
  nor (_12135_, _09472_, \uc8051golden_1.PC [9]);
  nor (_12136_, _12135_, _09473_);
  and (_12137_, _12136_, _06194_);
  nor (_12138_, _12136_, _06194_);
  nor (_12139_, _12138_, _12137_);
  and (_12140_, _08649_, _06194_);
  nor (_12141_, _08649_, _06194_);
  and (_12142_, _08532_, _06122_);
  nor (_12143_, _12142_, \uc8051golden_1.PC [6]);
  nor (_12144_, _12143_, _08646_);
  not (_12145_, _12144_);
  nor (_12146_, _12145_, _06340_);
  and (_12147_, _12145_, _06340_);
  nor (_12148_, _12147_, _12146_);
  and (_12149_, _06122_, \uc8051golden_1.PC [4]);
  nor (_12150_, _12149_, \uc8051golden_1.PC [5]);
  nor (_12151_, _12150_, _12142_);
  not (_12152_, _12151_);
  nor (_12153_, _12152_, _06650_);
  and (_12154_, _12152_, _06650_);
  nor (_12155_, _06122_, \uc8051golden_1.PC [4]);
  nor (_12156_, _12155_, _12149_);
  not (_12157_, _12156_);
  nor (_12158_, _12157_, _06265_);
  nor (_12159_, _06372_, _06134_);
  and (_12160_, _06372_, _06134_);
  nor (_12161_, _06693_, _06500_);
  nor (_12162_, _06228_, \uc8051golden_1.PC [1]);
  nor (_12163_, _06840_, _05685_);
  and (_12164_, _06228_, \uc8051golden_1.PC [1]);
  nor (_12165_, _12164_, _12162_);
  and (_12166_, _12165_, _12163_);
  nor (_12167_, _12166_, _12162_);
  and (_12168_, _06693_, _06500_);
  nor (_12169_, _12168_, _12161_);
  not (_12170_, _12169_);
  nor (_12171_, _12170_, _12167_);
  nor (_12172_, _12171_, _12161_);
  nor (_12173_, _12172_, _12160_);
  nor (_12174_, _12173_, _12159_);
  and (_12175_, _12157_, _06265_);
  nor (_12176_, _12175_, _12158_);
  not (_12177_, _12176_);
  nor (_12178_, _12177_, _12174_);
  nor (_12179_, _12178_, _12158_);
  nor (_12180_, _12179_, _12154_);
  nor (_12181_, _12180_, _12153_);
  not (_12182_, _12181_);
  and (_12183_, _12182_, _12148_);
  nor (_12184_, _12183_, _12146_);
  nor (_12185_, _12184_, _12141_);
  or (_12186_, _12185_, _12140_);
  nor (_12187_, _08647_, \uc8051golden_1.PC [8]);
  nor (_12188_, _12187_, _09472_);
  and (_12189_, _12188_, _06194_);
  nor (_12190_, _12188_, _06194_);
  nor (_12191_, _12190_, _12189_);
  and (_12192_, _12191_, _12186_);
  and (_12193_, _12192_, _12139_);
  and (_12194_, _12193_, _12134_);
  nor (_12195_, _12189_, _12137_);
  not (_12196_, _12195_);
  and (_12197_, _12196_, _12134_);
  or (_12198_, _12197_, _12129_);
  nor (_12199_, _12198_, _12194_);
  and (_12200_, _12199_, _12126_);
  nor (_12201_, _12121_, _06194_);
  nor (_12202_, _12201_, _12122_);
  not (_12203_, _12202_);
  nor (_12204_, _12203_, _12200_);
  nor (_12205_, _12204_, _12122_);
  nor (_12206_, _12205_, _12119_);
  nor (_12207_, _12206_, _12118_);
  nor (_12208_, _12207_, _12115_);
  nor (_12209_, _12208_, _12112_);
  nor (_12210_, _09480_, _06194_);
  and (_12211_, _09480_, _06194_);
  nor (_12212_, _12211_, _12210_);
  and (_12213_, _12212_, _12209_);
  nor (_12214_, _12212_, _12209_);
  or (_12215_, _12214_, _12213_);
  or (_12216_, _12215_, _10524_);
  and (_12217_, _06233_, _05946_);
  or (_12218_, _09480_, \uc8051golden_1.PSW [7]);
  and (_12219_, _12218_, _12217_);
  and (_12220_, _12219_, _12216_);
  not (_12221_, _05946_);
  nor (_12222_, _06288_, _06280_);
  and (_12223_, _12222_, _06379_);
  nor (_12224_, _12223_, _12221_);
  not (_12225_, _12224_);
  or (_12226_, _12225_, _12107_);
  nor (_12227_, _10963_, _06580_);
  not (_12228_, _12227_);
  and (_12229_, _06466_, _05951_);
  nor (_12230_, _12229_, _10565_);
  nor (_12231_, _10953_, _06959_);
  and (_12232_, _12231_, _10945_);
  and (_12233_, _12232_, _12230_);
  or (_12234_, _12233_, _12107_);
  or (_12235_, _09480_, _09012_);
  and (_12236_, _09496_, _06015_);
  and (_12237_, _06386_, _05981_);
  not (_12238_, _12237_);
  nor (_12239_, _11253_, _11254_);
  nor (_12240_, _12239_, _11257_);
  and (_12241_, _06840_, _06045_);
  nor (_12242_, _12241_, _11261_);
  nor (_12243_, _12242_, _11260_);
  and (_12244_, _12243_, _12240_);
  nor (_12245_, _11247_, _11248_);
  nor (_12246_, _12245_, _11252_);
  nor (_12247_, _11246_, _10970_);
  and (_12248_, _12247_, _12246_);
  and (_12249_, _12248_, _12244_);
  nor (_12250_, _09485_, \uc8051golden_1.PC [14]);
  nor (_12251_, _12250_, _09486_);
  not (_12252_, _12251_);
  nor (_12253_, _12252_, _08590_);
  and (_12254_, _12252_, _08590_);
  nor (_12255_, _12254_, _12253_);
  not (_12256_, _12255_);
  nor (_12257_, _09484_, \uc8051golden_1.PC [13]);
  nor (_12258_, _12257_, _09485_);
  and (_12259_, _12258_, _08813_);
  nor (_12260_, _12258_, _08813_);
  nor (_12261_, _09483_, \uc8051golden_1.PC [12]);
  nor (_12262_, _12261_, _09484_);
  not (_12263_, _12262_);
  nor (_12264_, _12263_, _08590_);
  not (_12265_, \uc8051golden_1.PC [11]);
  nor (_12266_, _09482_, _12265_);
  and (_12267_, _09482_, _12265_);
  or (_12268_, _12267_, _12266_);
  not (_12269_, _12268_);
  nor (_12270_, _12269_, _08590_);
  and (_12271_, _12269_, _08590_);
  nor (_12272_, _12271_, _12270_);
  nor (_12273_, _09489_, \uc8051golden_1.PC [10]);
  nor (_12274_, _12273_, _09482_);
  not (_12275_, _12274_);
  nor (_12276_, _12275_, _08590_);
  and (_12277_, _12275_, _08590_);
  nor (_12278_, _12277_, _12276_);
  and (_12279_, _12278_, _12272_);
  nor (_12280_, _09488_, \uc8051golden_1.PC [9]);
  nor (_12281_, _12280_, _09489_);
  not (_12282_, _12281_);
  nor (_12283_, _12282_, _08590_);
  and (_12284_, _12282_, _08590_);
  nor (_12285_, _12284_, _12283_);
  nor (_12286_, _08590_, _08540_);
  and (_12287_, _08590_, _08540_);
  nor (_12288_, _12287_, _12286_);
  not (_12289_, _12288_);
  and (_12290_, _08535_, _08532_);
  nor (_12291_, _12290_, \uc8051golden_1.PC [6]);
  nor (_12292_, _12291_, _08536_);
  not (_12293_, _12292_);
  nor (_12294_, _12293_, _08850_);
  and (_12295_, _12293_, _08850_);
  nor (_12296_, _12295_, _12294_);
  and (_12297_, _08535_, \uc8051golden_1.PC [4]);
  nor (_12298_, _12297_, \uc8051golden_1.PC [5]);
  nor (_12299_, _12298_, _12290_);
  not (_12300_, _12299_);
  nor (_12301_, _12300_, _08917_);
  and (_12302_, _12300_, _08917_);
  nor (_12303_, _08535_, \uc8051golden_1.PC [4]);
  nor (_12304_, _12303_, _12297_);
  not (_12305_, _12304_);
  nor (_12306_, _12305_, _08882_);
  nor (_12307_, _08534_, \uc8051golden_1.PC [3]);
  nor (_12308_, _12307_, _08535_);
  not (_12309_, _12308_);
  nor (_12310_, _12309_, _06562_);
  and (_12311_, _12309_, _06562_);
  nor (_12312_, _05689_, \uc8051golden_1.PC [2]);
  nor (_12313_, _12312_, _08534_);
  not (_12314_, _12313_);
  nor (_12315_, _12314_, _06736_);
  nor (_12316_, _07090_, _06024_);
  nor (_12317_, _06943_, \uc8051golden_1.PC [0]);
  and (_12318_, _07090_, _06024_);
  nor (_12319_, _12318_, _12316_);
  and (_12320_, _12319_, _12317_);
  nor (_12321_, _12320_, _12316_);
  and (_12322_, _12314_, _06736_);
  nor (_12323_, _12322_, _12315_);
  not (_12324_, _12323_);
  nor (_12325_, _12324_, _12321_);
  nor (_12326_, _12325_, _12315_);
  nor (_12327_, _12326_, _12311_);
  nor (_12328_, _12327_, _12310_);
  and (_12329_, _12305_, _08882_);
  nor (_12330_, _12329_, _12306_);
  not (_12331_, _12330_);
  nor (_12332_, _12331_, _12328_);
  nor (_12333_, _12332_, _12306_);
  nor (_12334_, _12333_, _12302_);
  or (_12335_, _12334_, _12301_);
  and (_12336_, _12335_, _12296_);
  nor (_12337_, _12336_, _12294_);
  nor (_12338_, _12337_, _12289_);
  nor (_12339_, _12338_, _12286_);
  nor (_12340_, _08537_, \uc8051golden_1.PC [8]);
  nor (_12341_, _12340_, _09488_);
  not (_12342_, _12341_);
  nor (_12343_, _12342_, _08590_);
  and (_12344_, _12342_, _08590_);
  nor (_12345_, _12344_, _12343_);
  not (_12346_, _12345_);
  nor (_12347_, _12346_, _12339_);
  and (_12348_, _12347_, _12285_);
  and (_12349_, _12348_, _12279_);
  nor (_12350_, _12343_, _12283_);
  not (_12351_, _12350_);
  and (_12352_, _12351_, _12279_);
  or (_12353_, _12352_, _12276_);
  or (_12354_, _12353_, _12349_);
  nor (_12355_, _12354_, _12270_);
  and (_12356_, _12263_, _08590_);
  nor (_12357_, _12356_, _12264_);
  not (_12358_, _12357_);
  nor (_12359_, _12358_, _12355_);
  nor (_12360_, _12359_, _12264_);
  nor (_12361_, _12360_, _12260_);
  nor (_12362_, _12361_, _12259_);
  nor (_12363_, _12362_, _12256_);
  nor (_12364_, _12363_, _12253_);
  not (_12365_, _09496_);
  and (_12366_, _12365_, _08590_);
  nor (_12367_, _12365_, _08590_);
  nor (_12368_, _12367_, _12366_);
  and (_12369_, _12368_, _12364_);
  nor (_12370_, _12368_, _12364_);
  or (_12371_, _12370_, _12369_);
  or (_12372_, _12371_, _12249_);
  nand (_12373_, _12249_, _12365_);
  and (_12374_, _12373_, _06482_);
  and (_12375_, _12374_, _12372_);
  and (_12376_, _09075_, _06194_);
  nor (_12377_, _12376_, _08788_);
  or (_12378_, _09440_, _06340_);
  or (_12379_, _09120_, _07896_);
  and (_12380_, _12379_, _12378_);
  and (_12381_, _12380_, _12377_);
  or (_12382_, _09165_, _07928_);
  or (_12383_, _09441_, _06650_);
  and (_12384_, _12383_, _12382_);
  or (_12385_, _09210_, _07934_);
  or (_12386_, _09442_, _06265_);
  and (_12387_, _12386_, _12385_);
  and (_12388_, _12387_, _12384_);
  and (_12389_, _12388_, _12381_);
  or (_12390_, _09443_, _06372_);
  or (_12391_, _09255_, _06589_);
  and (_12392_, _12391_, _12390_);
  or (_12393_, _09444_, _06693_);
  or (_12394_, _09300_, _07573_);
  and (_12395_, _12394_, _12393_);
  and (_12396_, _12395_, _12392_);
  or (_12397_, _09446_, _06840_);
  or (_12398_, _09390_, _06967_);
  or (_12399_, _09345_, _06229_);
  or (_12400_, _09445_, _06228_);
  and (_12401_, _12400_, _12399_);
  and (_12402_, _12401_, _12398_);
  and (_12403_, _12402_, _12397_);
  and (_12404_, _12403_, _12396_);
  and (_12405_, _12404_, _12389_);
  or (_12406_, _12405_, _12371_);
  nand (_12407_, _12404_, _12389_);
  or (_12408_, _12407_, _09496_);
  and (_12409_, _12408_, _06457_);
  and (_12410_, _12409_, _12406_);
  not (_12411_, _06457_);
  not (_12412_, _08071_);
  and (_12413_, _08070_, _06194_);
  nor (_12414_, _12413_, _12412_);
  nor (_12415_, _08118_, _07896_);
  and (_12416_, _08118_, _07896_);
  nor (_12417_, _12416_, _12415_);
  and (_12418_, _12417_, _12414_);
  and (_12419_, _08207_, _07928_);
  not (_12420_, _12419_);
  or (_12421_, _08207_, _07928_);
  and (_12422_, _12421_, _12420_);
  and (_12423_, _08301_, _07934_);
  nor (_12424_, _08301_, _07934_);
  nor (_12425_, _12424_, _12423_);
  and (_12426_, _12425_, _12422_);
  and (_12427_, _12426_, _12418_);
  and (_12428_, _07775_, _06589_);
  not (_12429_, _12428_);
  or (_12430_, _07775_, _06589_);
  and (_12431_, _12430_, _12429_);
  nor (_12432_, _07623_, _07573_);
  and (_12433_, _07623_, _07573_);
  nor (_12434_, _12433_, _12432_);
  and (_12435_, _12434_, _12431_);
  or (_12436_, _07485_, _06967_);
  nor (_12437_, _07196_, _06229_);
  and (_12438_, _07196_, _06229_);
  nor (_12439_, _12438_, _12437_);
  and (_12440_, _12439_, _12436_);
  or (_12441_, _07473_, _06840_);
  and (_12442_, _12441_, _12440_);
  and (_12443_, _12442_, _12435_);
  and (_12444_, _12443_, _12427_);
  nand (_12445_, _12444_, _12365_);
  and (_12446_, _06285_, _06386_);
  and (_12447_, _07378_, _06386_);
  nor (_12448_, _12447_, _12446_);
  and (_12449_, _12448_, _06464_);
  not (_12450_, _12449_);
  or (_12451_, _12444_, _12371_);
  and (_12452_, _12451_, _12450_);
  and (_12453_, _12452_, _12445_);
  and (_12454_, _09480_, _06406_);
  and (_12455_, _06407_, _05997_);
  or (_12456_, _12455_, _09480_);
  and (_12457_, _06394_, _05981_);
  nor (_12458_, _12457_, _10677_);
  and (_12459_, _08161_, _08072_);
  and (_12460_, _12459_, _08754_);
  and (_12461_, _08521_, _08476_);
  and (_12462_, _08432_, _08388_);
  and (_12463_, _12462_, _12461_);
  nand (_12464_, _12463_, _12460_);
  or (_12465_, _12464_, _09496_);
  and (_12466_, _12463_, _12460_);
  or (_12467_, _12466_, _12371_);
  and (_12468_, _12467_, _06401_);
  and (_12469_, _12468_, _12465_);
  and (_12470_, _08118_, _08070_);
  and (_12471_, _12470_, _08549_);
  and (_12472_, _07473_, _07196_);
  and (_12473_, _12472_, _08550_);
  nand (_12474_, _12473_, _12471_);
  and (_12475_, _12474_, _12215_);
  and (_12476_, _12473_, _12471_);
  and (_12477_, _12476_, _09480_);
  or (_12478_, _12477_, _08644_);
  or (_12479_, _12478_, _12475_);
  nor (_12480_, _07329_, _06001_);
  or (_12481_, _12480_, _10663_);
  nor (_12482_, _07199_, _06790_);
  or (_12483_, _12482_, _09480_);
  nand (_12484_, _06742_, _06402_);
  not (_12485_, _12484_);
  or (_12486_, _06790_, \uc8051golden_1.PC [15]);
  or (_12487_, _12486_, _12485_);
  or (_12488_, _12487_, _07332_);
  and (_12489_, _12488_, _12483_);
  or (_12490_, _12489_, _12481_);
  not (_12491_, _12481_);
  nor (_12492_, _07332_, _06854_);
  and (_12493_, _12492_, _12491_);
  or (_12494_, _12493_, _12107_);
  and (_12495_, _12494_, _12490_);
  or (_12496_, _12495_, _08643_);
  nor (_12497_, _07212_, _06401_);
  and (_12498_, _12497_, _12496_);
  and (_12499_, _12498_, _12479_);
  or (_12500_, _12499_, _12469_);
  and (_12501_, _12500_, _12458_);
  not (_12502_, _12455_);
  and (_12503_, _12458_, _08659_);
  not (_12504_, _12503_);
  and (_12505_, _12504_, _12107_);
  or (_12506_, _12505_, _12502_);
  or (_12507_, _12506_, _12501_);
  and (_12508_, _12507_, _12456_);
  nor (_12509_, _10644_, _07233_);
  not (_12510_, _12509_);
  or (_12511_, _12510_, _12508_);
  or (_12512_, _12509_, _12107_);
  and (_12513_, _12512_, _06414_);
  and (_12514_, _12513_, _12511_);
  or (_12515_, _12514_, _12454_);
  and (_12516_, _06392_, _05981_);
  nor (_12517_, _12516_, _10642_);
  and (_12518_, _12517_, _12515_);
  not (_12519_, _12517_);
  and (_12520_, _12519_, _12107_);
  not (_12521_, _06000_);
  nor (_12522_, _06419_, _12521_);
  and (_12523_, _12522_, _06844_);
  not (_12524_, _12523_);
  or (_12525_, _12524_, _12520_);
  or (_12526_, _12525_, _12518_);
  or (_12527_, _12523_, _09480_);
  and (_12528_, _12527_, _12449_);
  and (_12529_, _12528_, _12526_);
  or (_12530_, _12529_, _12453_);
  and (_12531_, _12530_, _12411_);
  or (_12532_, _12531_, _06420_);
  or (_12533_, _12532_, _12410_);
  not (_12534_, _06482_);
  nor (_12535_, _11218_, _11217_);
  nor (_12536_, _12535_, _11221_);
  not (_12537_, _11224_);
  nor (_12538_, _08521_, \uc8051golden_1.ACC [0]);
  or (_12539_, _12538_, _11225_);
  and (_12540_, _12539_, _12537_);
  and (_12541_, _12540_, _12536_);
  nor (_12542_, _11212_, _11211_);
  nor (_12543_, _12542_, _11216_);
  nor (_12544_, _11210_, _09034_);
  and (_12545_, _12544_, _12543_);
  and (_12546_, _12545_, _12541_);
  and (_12547_, _12546_, _09496_);
  not (_12548_, _12546_);
  and (_12549_, _12548_, _12371_);
  or (_12550_, _12549_, _06842_);
  or (_12551_, _12550_, _12547_);
  and (_12552_, _12551_, _12534_);
  and (_12553_, _12552_, _12533_);
  or (_12554_, _12553_, _12375_);
  and (_12555_, _12554_, _12238_);
  nand (_12556_, _12237_, _12107_);
  nor (_12557_, _06387_, _07349_);
  nor (_12558_, _07326_, _06006_);
  nor (_12559_, _12558_, _07252_);
  and (_12560_, _07103_, _06381_);
  and (_12561_, _06955_, _06381_);
  nor (_12562_, _12561_, _12560_);
  not (_12563_, _06388_);
  and (_12564_, _06483_, _06381_);
  and (_12565_, _06451_, _06381_);
  nor (_12566_, _12565_, _12564_);
  and (_12567_, _12566_, _12563_);
  and (_12568_, _12567_, _12562_);
  and (_12569_, _12568_, _12559_);
  and (_12570_, _12569_, _12557_);
  nand (_12571_, _12570_, _12556_);
  or (_12572_, _12571_, _12555_);
  and (_12573_, _06014_, _06381_);
  not (_12574_, _12573_);
  nor (_12575_, _11511_, _09538_);
  and (_12576_, _12575_, _12574_);
  or (_12577_, _12570_, _09480_);
  and (_12578_, _12577_, _12576_);
  and (_12579_, _12578_, _12572_);
  not (_12580_, _12576_);
  and (_12581_, _12580_, _12107_);
  and (_12582_, _06434_, _06007_);
  not (_12583_, _12582_);
  or (_12584_, _12583_, _12581_);
  or (_12585_, _12584_, _12579_);
  and (_12586_, _06280_, _06016_);
  not (_12587_, _12586_);
  and (_12588_, _10740_, _12587_);
  or (_12589_, _12582_, _09480_);
  and (_12590_, _12589_, _12588_);
  and (_12591_, _12590_, _12585_);
  nor (_12592_, _10572_, _06437_);
  not (_12593_, _12592_);
  not (_12594_, _12588_);
  and (_12595_, _12594_, _12107_);
  or (_12596_, _12595_, _12593_);
  or (_12597_, _12596_, _12591_);
  or (_12598_, _12592_, _09480_);
  and (_12599_, _12598_, _06023_);
  and (_12600_, _12599_, _12597_);
  and (_12601_, _12107_, _06022_);
  nor (_12602_, _06300_, _06017_);
  not (_12603_, _12602_);
  or (_12604_, _12603_, _12601_);
  or (_12605_, _12604_, _12600_);
  or (_12606_, _12602_, _09480_);
  and (_12607_, _12606_, _06473_);
  and (_12608_, _12607_, _12605_);
  nand (_12609_, _09496_, _06472_);
  nand (_12610_, _12609_, _06294_);
  or (_12611_, _12610_, _12608_);
  or (_12612_, _09480_, _06294_);
  and (_12613_, _12612_, _06279_);
  and (_12614_, _12613_, _12611_);
  or (_12615_, _12614_, _12236_);
  nor (_12616_, _10072_, _05982_);
  and (_12617_, _12616_, _12615_);
  nor (_12618_, _06376_, _05936_);
  not (_12619_, _12618_);
  not (_12620_, _12616_);
  and (_12621_, _12620_, _12107_);
  or (_12622_, _12621_, _12619_);
  or (_12623_, _12622_, _12617_);
  and (_12624_, _06233_, _05935_);
  not (_12625_, _12624_);
  or (_12626_, _12618_, _09480_);
  and (_12627_, _12626_, _12625_);
  and (_12628_, _12627_, _12623_);
  and (_12629_, _12624_, _12215_);
  or (_12630_, _12629_, _09013_);
  or (_12631_, _12630_, _12628_);
  and (_12632_, _12631_, _12235_);
  or (_12633_, _12632_, _06275_);
  or (_12634_, _09496_, _06276_);
  and (_12635_, _12634_, _10934_);
  and (_12636_, _12635_, _12633_);
  and (_12637_, _10933_, _09480_);
  or (_12638_, _12637_, _12636_);
  and (_12639_, _05981_, _05942_);
  not (_12640_, _12639_);
  and (_12641_, _12640_, _12638_);
  not (_12642_, \uc8051golden_1.DPH [0]);
  and (_12643_, \uc8051golden_1.DPL [7], \uc8051golden_1.ACC [7]);
  nor (_12644_, \uc8051golden_1.DPL [7], \uc8051golden_1.ACC [7]);
  and (_12645_, \uc8051golden_1.DPL [6], \uc8051golden_1.ACC [6]);
  nor (_12646_, \uc8051golden_1.DPL [6], \uc8051golden_1.ACC [6]);
  nor (_12647_, _12646_, _12645_);
  and (_12648_, \uc8051golden_1.DPL [5], \uc8051golden_1.ACC [5]);
  nor (_12649_, \uc8051golden_1.DPL [5], \uc8051golden_1.ACC [5]);
  and (_12650_, \uc8051golden_1.DPL [4], \uc8051golden_1.ACC [4]);
  nor (_12651_, _06115_, _06111_);
  nor (_12652_, \uc8051golden_1.DPL [4], \uc8051golden_1.ACC [4]);
  nor (_12653_, _12652_, _12650_);
  not (_12654_, _12653_);
  nor (_12655_, _12654_, _12651_);
  nor (_12656_, _12655_, _12650_);
  nor (_12657_, _12656_, _12649_);
  nor (_12658_, _12657_, _12648_);
  not (_12659_, _12658_);
  and (_12660_, _12659_, _12647_);
  nor (_12661_, _12660_, _12645_);
  nor (_12662_, _12661_, _12644_);
  nor (_12663_, _12662_, _12643_);
  nor (_12664_, _12663_, _12642_);
  and (_12665_, _12664_, \uc8051golden_1.DPH [1]);
  and (_12666_, _12665_, \uc8051golden_1.DPH [2]);
  and (_12667_, _12666_, \uc8051golden_1.DPH [3]);
  and (_12668_, _12667_, \uc8051golden_1.DPH [4]);
  and (_12669_, _12668_, \uc8051golden_1.DPH [5]);
  and (_12670_, _12669_, \uc8051golden_1.DPH [6]);
  nand (_12671_, _12670_, \uc8051golden_1.DPH [7]);
  or (_12672_, _12670_, \uc8051golden_1.DPH [7]);
  and (_12673_, _12672_, _12639_);
  and (_12674_, _12673_, _12671_);
  nor (_12676_, _06375_, _05943_);
  not (_12677_, _12676_);
  or (_12678_, _12677_, _12674_);
  or (_12679_, _12678_, _12641_);
  and (_12680_, _06233_, _05942_);
  not (_12681_, _12680_);
  or (_12682_, _12676_, _09480_);
  and (_12683_, _12682_, _12681_);
  and (_12684_, _12683_, _12679_);
  not (_12685_, _12233_);
  or (_12686_, _12215_, _11297_);
  not (_12687_, _11297_);
  or (_12688_, _12687_, _09480_);
  and (_12689_, _12688_, _12680_);
  and (_12690_, _12689_, _12686_);
  or (_12691_, _12690_, _12685_);
  or (_12692_, _12691_, _12684_);
  and (_12693_, _12692_, _12234_);
  or (_12694_, _12693_, _12228_);
  or (_12695_, _12227_, _09480_);
  and (_12697_, _12695_, _07282_);
  and (_12698_, _12697_, _12694_);
  and (_12699_, _09496_, _06474_);
  nor (_12700_, _06582_, _05952_);
  not (_12701_, _12700_);
  or (_12702_, _12701_, _12699_);
  or (_12703_, _12702_, _12698_);
  and (_12704_, _06233_, _05951_);
  not (_12705_, _12704_);
  or (_12706_, _12700_, _09480_);
  and (_12707_, _12706_, _12705_);
  and (_12708_, _12707_, _12703_);
  or (_12709_, _12215_, _12687_);
  or (_12710_, _11297_, _09480_);
  and (_12711_, _12710_, _12704_);
  and (_12712_, _12711_, _12709_);
  or (_12713_, _12712_, _12708_);
  not (_12714_, _05955_);
  or (_12715_, _10738_, _12714_);
  and (_12716_, _06285_, _05955_);
  nor (_12717_, _12716_, _06972_);
  and (_12718_, _12717_, _10560_);
  and (_12719_, _12718_, _12715_);
  and (_12720_, _12719_, _12713_);
  nor (_12721_, _10989_, _06567_);
  not (_12722_, _12721_);
  not (_12723_, _12719_);
  and (_12724_, _12723_, _12107_);
  or (_12725_, _12724_, _12722_);
  or (_12726_, _12725_, _12720_);
  or (_12727_, _12721_, _09480_);
  and (_12728_, _12727_, _07279_);
  and (_12729_, _12728_, _12726_);
  and (_12730_, _09496_, _06478_);
  nor (_12731_, _06569_, _05956_);
  not (_12732_, _12731_);
  or (_12733_, _12732_, _12730_);
  or (_12734_, _12733_, _12729_);
  and (_12735_, _06233_, _05955_);
  not (_12736_, _12735_);
  or (_12737_, _12731_, _09480_);
  and (_12738_, _12737_, _12736_);
  and (_12739_, _12738_, _12734_);
  or (_12740_, _12215_, \uc8051golden_1.PSW [7]);
  or (_12741_, _09480_, _10524_);
  and (_12742_, _12741_, _12735_);
  and (_12743_, _12742_, _12740_);
  or (_12744_, _12743_, _12224_);
  or (_12745_, _12744_, _12739_);
  and (_12746_, _12745_, _12226_);
  or (_12747_, _12746_, _11019_);
  or (_12748_, _11018_, _09480_);
  and (_12749_, _12748_, _09043_);
  and (_12750_, _12749_, _12747_);
  and (_12751_, _09496_, _06479_);
  nor (_12752_, _06572_, _05947_);
  not (_12753_, _12752_);
  or (_12754_, _12753_, _12751_);
  or (_12755_, _12754_, _12750_);
  not (_12756_, _12217_);
  or (_12757_, _12752_, _09480_);
  and (_12758_, _12757_, _12756_);
  and (_12759_, _12758_, _12755_);
  or (_12760_, _12759_, _12220_);
  and (_12761_, _11028_, _10472_);
  and (_12762_, _12761_, _12760_);
  not (_12763_, _12761_);
  and (_12764_, _12763_, _12107_);
  or (_12765_, _12764_, _11061_);
  or (_12766_, _12765_, _12762_);
  or (_12767_, _11060_, _09480_);
  and (_12768_, _12767_, _11090_);
  and (_12769_, _12768_, _12766_);
  and (_12770_, _12107_, _11089_);
  or (_12771_, _12770_, _06588_);
  or (_12772_, _12771_, _12769_);
  nand (_12773_, _08070_, _06588_);
  and (_12774_, _12773_, _12772_);
  or (_12775_, _12774_, _05966_);
  or (_12776_, _09480_, _05967_);
  and (_12777_, _12776_, _06596_);
  and (_12778_, _12777_, _12775_);
  not (_12779_, _12108_);
  not (_12780_, _07961_);
  and (_12781_, _08598_, \uc8051golden_1.P3 [2]);
  and (_12782_, _08603_, \uc8051golden_1.IE [2]);
  nor (_12783_, _12782_, _12781_);
  and (_12784_, _08606_, \uc8051golden_1.SCON [2]);
  and (_12785_, _08608_, \uc8051golden_1.P2 [2]);
  nor (_12786_, _12785_, _12784_);
  and (_12787_, _12786_, _12783_);
  and (_12788_, _08614_, \uc8051golden_1.IP [2]);
  and (_12789_, _08612_, \uc8051golden_1.PSW [2]);
  and (_12790_, _08618_, \uc8051golden_1.B [2]);
  and (_12791_, _08616_, \uc8051golden_1.ACC [2]);
  or (_12792_, _12791_, _12790_);
  or (_12793_, _12792_, _12789_);
  nor (_12794_, _12793_, _12788_);
  and (_12795_, _08623_, \uc8051golden_1.TCON [2]);
  and (_12796_, _07959_, \uc8051golden_1.P0 [2]);
  and (_12797_, _08626_, \uc8051golden_1.P1 [2]);
  or (_12798_, _12797_, _12796_);
  nor (_12799_, _12798_, _12795_);
  and (_12800_, _12799_, _12794_);
  and (_12801_, _12800_, _12787_);
  and (_12802_, _12801_, _08390_);
  nor (_12803_, _12802_, _12780_);
  not (_12804_, _08235_);
  and (_12805_, _08608_, \uc8051golden_1.P2 [1]);
  and (_12806_, _08598_, \uc8051golden_1.P3 [1]);
  and (_12807_, _08603_, \uc8051golden_1.IE [1]);
  or (_12808_, _12807_, _12806_);
  nor (_12809_, _12808_, _12805_);
  and (_12810_, _08623_, \uc8051golden_1.TCON [1]);
  and (_12811_, _08626_, \uc8051golden_1.P1 [1]);
  and (_12812_, _07959_, \uc8051golden_1.P0 [1]);
  or (_12813_, _12812_, _12811_);
  nor (_12814_, _12813_, _12810_);
  and (_12815_, _08612_, \uc8051golden_1.PSW [1]);
  and (_12816_, _08616_, \uc8051golden_1.ACC [1]);
  and (_12817_, _08618_, \uc8051golden_1.B [1]);
  or (_12818_, _12817_, _12816_);
  nor (_12819_, _12818_, _12815_);
  and (_12820_, _08606_, \uc8051golden_1.SCON [1]);
  and (_12821_, _08614_, \uc8051golden_1.IP [1]);
  nor (_12822_, _12821_, _12820_);
  and (_12823_, _12822_, _12819_);
  and (_12824_, _12823_, _12814_);
  and (_12825_, _12824_, _12809_);
  and (_12826_, _12825_, _08434_);
  nor (_12827_, _12826_, _12804_);
  nor (_12828_, _12827_, _12803_);
  and (_12829_, _08606_, \uc8051golden_1.SCON [4]);
  and (_12830_, _08598_, \uc8051golden_1.P3 [4]);
  and (_12831_, _08603_, \uc8051golden_1.IE [4]);
  or (_12832_, _12831_, _12830_);
  nor (_12833_, _12832_, _12829_);
  and (_12834_, _08623_, \uc8051golden_1.TCON [4]);
  and (_12835_, _08626_, \uc8051golden_1.P1 [4]);
  and (_12836_, _07959_, \uc8051golden_1.P0 [4]);
  or (_12837_, _12836_, _12835_);
  nor (_12838_, _12837_, _12834_);
  and (_12839_, _08612_, \uc8051golden_1.PSW [4]);
  and (_12840_, _08618_, \uc8051golden_1.B [4]);
  and (_12841_, _08616_, \uc8051golden_1.ACC [4]);
  or (_12842_, _12841_, _12840_);
  nor (_12843_, _12842_, _12839_);
  and (_12844_, _08608_, \uc8051golden_1.P2 [4]);
  and (_12845_, _08614_, \uc8051golden_1.IP [4]);
  nor (_12846_, _12845_, _12844_);
  and (_12847_, _12846_, _12843_);
  and (_12848_, _12847_, _12838_);
  and (_12849_, _12848_, _12833_);
  and (_12850_, _12849_, _08302_);
  and (_12851_, _07924_, _07573_);
  not (_12852_, _12851_);
  nor (_12853_, _12852_, _12850_);
  nor (_12854_, _12853_, _08633_);
  and (_12855_, _12854_, _12828_);
  and (_12856_, _07924_, _06693_);
  not (_12857_, _12856_);
  and (_12858_, _08598_, \uc8051golden_1.P3 [0]);
  and (_12859_, _08603_, \uc8051golden_1.IE [0]);
  nor (_12860_, _12859_, _12858_);
  and (_12861_, _08606_, \uc8051golden_1.SCON [0]);
  and (_12862_, _08608_, \uc8051golden_1.P2 [0]);
  nor (_12863_, _12862_, _12861_);
  and (_12864_, _12863_, _12860_);
  and (_12865_, _08614_, \uc8051golden_1.IP [0]);
  and (_12866_, _08612_, \uc8051golden_1.PSW [0]);
  and (_12867_, _08616_, \uc8051golden_1.ACC [0]);
  and (_12868_, _08618_, \uc8051golden_1.B [0]);
  or (_12869_, _12868_, _12867_);
  or (_12870_, _12869_, _12866_);
  nor (_12871_, _12870_, _12865_);
  and (_12872_, _08623_, \uc8051golden_1.TCON [0]);
  and (_12873_, _07959_, \uc8051golden_1.P0 [0]);
  and (_12874_, _08626_, \uc8051golden_1.P1 [0]);
  or (_12875_, _12874_, _12873_);
  nor (_12876_, _12875_, _12872_);
  and (_12877_, _12876_, _12871_);
  and (_12878_, _12877_, _12864_);
  and (_12879_, _12878_, _08478_);
  nor (_12880_, _12879_, _12857_);
  and (_12881_, _07959_, \uc8051golden_1.P0 [6]);
  and (_12882_, _08623_, \uc8051golden_1.TCON [6]);
  and (_12883_, _08626_, \uc8051golden_1.P1 [6]);
  and (_12884_, _08606_, \uc8051golden_1.SCON [6]);
  and (_12885_, _08608_, \uc8051golden_1.P2 [6]);
  and (_12886_, _08603_, \uc8051golden_1.IE [6]);
  and (_12887_, _08598_, \uc8051golden_1.P3 [6]);
  and (_12888_, _08614_, \uc8051golden_1.IP [6]);
  and (_12889_, _08612_, \uc8051golden_1.PSW [6]);
  and (_12890_, _08616_, \uc8051golden_1.ACC [6]);
  and (_12891_, _08618_, \uc8051golden_1.B [6]);
  or (_12892_, _12891_, _12890_);
  or (_12893_, _12892_, _12889_);
  or (_12894_, _12893_, _12888_);
  or (_12895_, _12894_, _12887_);
  or (_12896_, _12895_, _12886_);
  or (_12897_, _12896_, _12885_);
  or (_12898_, _12897_, _12884_);
  or (_12899_, _12898_, _12883_);
  or (_12900_, _12899_, _12882_);
  nor (_12901_, _12900_, _12881_);
  and (_12902_, _12901_, _08119_);
  and (_12903_, _07960_, _07573_);
  not (_12904_, _12903_);
  nor (_12905_, _12904_, _12902_);
  nor (_12906_, _12905_, _12880_);
  not (_12907_, _08248_);
  and (_12908_, _08598_, \uc8051golden_1.P3 [3]);
  and (_12909_, _08603_, \uc8051golden_1.IE [3]);
  nor (_12910_, _12909_, _12908_);
  and (_12911_, _08606_, \uc8051golden_1.SCON [3]);
  and (_12912_, _08608_, \uc8051golden_1.P2 [3]);
  nor (_12913_, _12912_, _12911_);
  and (_12914_, _12913_, _12910_);
  and (_12915_, _08614_, \uc8051golden_1.IP [3]);
  and (_12916_, _08612_, \uc8051golden_1.PSW [3]);
  and (_12917_, _08616_, \uc8051golden_1.ACC [3]);
  and (_12918_, _08618_, \uc8051golden_1.B [3]);
  or (_12919_, _12918_, _12917_);
  or (_12920_, _12919_, _12916_);
  nor (_12921_, _12920_, _12915_);
  and (_12922_, _08623_, \uc8051golden_1.TCON [3]);
  and (_12923_, _07959_, \uc8051golden_1.P0 [3]);
  and (_12924_, _08626_, \uc8051golden_1.P1 [3]);
  or (_12925_, _12924_, _12923_);
  nor (_12926_, _12925_, _12922_);
  and (_12927_, _12926_, _12921_);
  and (_12928_, _12927_, _12914_);
  and (_12929_, _12928_, _08346_);
  nor (_12930_, _12929_, _12907_);
  and (_12931_, _08612_, \uc8051golden_1.PSW [5]);
  and (_12932_, _08606_, \uc8051golden_1.SCON [5]);
  nor (_12933_, _12932_, _12931_);
  and (_12934_, _08614_, \uc8051golden_1.IP [5]);
  and (_12935_, _08616_, \uc8051golden_1.ACC [5]);
  and (_12936_, _08618_, \uc8051golden_1.B [5]);
  or (_12937_, _12936_, _12935_);
  nor (_12938_, _12937_, _12934_);
  and (_12939_, _08623_, \uc8051golden_1.TCON [5]);
  and (_12940_, _08626_, \uc8051golden_1.P1 [5]);
  and (_12941_, _07959_, \uc8051golden_1.P0 [5]);
  or (_12942_, _12941_, _12940_);
  nor (_12943_, _12942_, _12939_);
  and (_12944_, _08608_, \uc8051golden_1.P2 [5]);
  and (_12945_, _08603_, \uc8051golden_1.IE [5]);
  and (_12946_, _08598_, \uc8051golden_1.P3 [5]);
  or (_12947_, _12946_, _12945_);
  nor (_12948_, _12947_, _12944_);
  and (_12949_, _12948_, _12943_);
  and (_12950_, _12949_, _12938_);
  and (_12951_, _12950_, _12933_);
  and (_12952_, _12951_, _08208_);
  and (_12953_, _07938_, _07573_);
  not (_12954_, _12953_);
  nor (_12955_, _12954_, _12952_);
  nor (_12956_, _12955_, _12930_);
  and (_12957_, _12956_, _12906_);
  and (_12958_, _12957_, _12855_);
  not (_12959_, _12958_);
  or (_12960_, _12371_, _12959_);
  or (_12961_, _09496_, _12958_);
  and (_12962_, _12961_, _06460_);
  and (_12963_, _12962_, _12960_);
  or (_12964_, _12963_, _12779_);
  or (_12965_, _12964_, _12778_);
  and (_12966_, _12965_, _12109_);
  or (_12967_, _12966_, _12094_);
  not (_12968_, _11243_);
  or (_12969_, _11204_, _09480_);
  and (_12970_, _12969_, _12968_);
  and (_12971_, _12970_, _12967_);
  and (_12972_, _12107_, _11243_);
  or (_12973_, _12972_, _06305_);
  or (_12974_, _12973_, _12971_);
  nand (_12975_, _08070_, _06305_);
  and (_12976_, _12975_, _12974_);
  or (_12977_, _12976_, _05971_);
  not (_12978_, _06487_);
  not (_12979_, _05971_);
  or (_12980_, _09480_, _12979_);
  and (_12981_, _12980_, _12978_);
  and (_12982_, _12981_, _12977_);
  or (_12983_, _12371_, _12958_);
  nand (_12984_, _12365_, _12958_);
  and (_12985_, _12984_, _12983_);
  and (_12986_, _12985_, _06487_);
  and (_12987_, _08546_, _09074_);
  not (_12988_, _12987_);
  or (_12989_, _12988_, _12986_);
  or (_12990_, _12989_, _12982_);
  or (_12991_, _12987_, _12107_);
  and (_12992_, _12991_, _07037_);
  and (_12993_, _12992_, _12990_);
  nor (_12994_, _11290_, _11285_);
  not (_12995_, _12994_);
  and (_12996_, _09480_, _06606_);
  or (_12997_, _12996_, _12995_);
  or (_12998_, _12997_, _12993_);
  or (_12999_, _12107_, _12994_);
  and (_13000_, _12999_, _09463_);
  and (_13001_, _13000_, _12998_);
  and (_13002_, _06465_, _06194_);
  or (_13003_, _13002_, _05969_);
  or (_13004_, _13003_, _13001_);
  not (_13005_, _05969_);
  or (_13006_, _09480_, _13005_);
  and (_13007_, _13006_, _06807_);
  and (_13008_, _13007_, _13004_);
  and (_13009_, _12985_, _06234_);
  and (_13010_, _05962_, _05805_);
  nor (_13011_, _13010_, _07320_);
  not (_13012_, _13011_);
  or (_13013_, _13012_, _13009_);
  or (_13014_, _13013_, _13008_);
  or (_13015_, _13011_, _12107_);
  and (_13016_, _13015_, _06196_);
  and (_13017_, _13016_, _13014_);
  and (_13018_, _09480_, _06195_);
  nor (_13019_, _11315_, _11308_);
  not (_13020_, _13019_);
  or (_13021_, _13020_, _13018_);
  or (_13022_, _13021_, _13017_);
  not (_13023_, _06475_);
  or (_13024_, _13019_, _12107_);
  and (_13025_, _13024_, _13023_);
  and (_13026_, _13025_, _13022_);
  and (_13027_, _06475_, _06194_);
  or (_13028_, _13027_, _05963_);
  or (_13029_, _13028_, _13026_);
  and (_13030_, _06233_, _05962_);
  not (_13031_, _13030_);
  or (_13032_, _09480_, _05964_);
  and (_13033_, _13032_, _13031_);
  and (_13034_, _13033_, _13029_);
  and (_13035_, _13030_, _12107_);
  or (_13036_, _13035_, _13034_);
  or (_13037_, _13036_, _01379_);
  or (_13038_, _01375_, \uc8051golden_1.PC [15]);
  and (_13039_, _13038_, _42545_);
  and (_40336_, _13039_, _13037_);
  not (_13040_, _07931_);
  and (_13041_, _13040_, \uc8051golden_1.P2 [7]);
  and (_13042_, _09034_, _07931_);
  or (_13043_, _13042_, _13041_);
  and (_13044_, _13043_, _06582_);
  nor (_13045_, _13040_, _08070_);
  or (_13046_, _13045_, _13041_);
  or (_13047_, _13046_, _06293_);
  not (_13048_, _08608_);
  and (_13049_, _13048_, \uc8051golden_1.P2 [7]);
  and (_13050_, _08639_, _08608_);
  or (_13051_, _13050_, _13049_);
  and (_13052_, _13051_, _06393_);
  and (_13053_, _08762_, _07931_);
  or (_13054_, _13053_, _13041_);
  or (_13055_, _13054_, _07210_);
  and (_13056_, _07931_, \uc8051golden_1.ACC [7]);
  or (_13057_, _13056_, _13041_);
  and (_13058_, _13057_, _07199_);
  and (_13059_, _07200_, \uc8051golden_1.P2 [7]);
  or (_13060_, _13059_, _06401_);
  or (_13061_, _13060_, _13058_);
  and (_13062_, _13061_, _06396_);
  and (_13063_, _13062_, _13055_);
  and (_13064_, _08635_, _08608_);
  or (_13065_, _13064_, _13049_);
  and (_13066_, _13065_, _06395_);
  or (_13067_, _13066_, _06399_);
  or (_13068_, _13067_, _13063_);
  or (_13069_, _13046_, _07221_);
  and (_13070_, _13069_, _13068_);
  or (_13071_, _13070_, _06406_);
  or (_13072_, _13057_, _06414_);
  and (_13073_, _13072_, _06844_);
  and (_13074_, _13073_, _13071_);
  or (_13075_, _13074_, _13052_);
  and (_13076_, _13075_, _07245_);
  or (_13077_, _13049_, _08634_);
  and (_13078_, _13077_, _06387_);
  and (_13079_, _13078_, _13065_);
  or (_13080_, _13079_, _13076_);
  and (_13081_, _13080_, _06446_);
  and (_13082_, _08794_, _08608_);
  or (_13083_, _13082_, _13049_);
  and (_13084_, _13083_, _06300_);
  or (_13085_, _13084_, _10059_);
  or (_13086_, _13085_, _13081_);
  and (_13087_, _13086_, _13047_);
  or (_13088_, _13087_, _06281_);
  and (_13089_, _07931_, _08749_);
  or (_13090_, _13041_, _06282_);
  or (_13091_, _13090_, _13089_);
  and (_13092_, _13091_, _06279_);
  and (_13093_, _13092_, _13088_);
  and (_13094_, _09009_, _07931_);
  or (_13095_, _13094_, _13041_);
  and (_13096_, _13095_, _06015_);
  or (_13097_, _13096_, _06275_);
  or (_13098_, _13097_, _13093_);
  and (_13099_, _08813_, _07931_);
  or (_13100_, _13099_, _13041_);
  or (_13101_, _13100_, _06276_);
  and (_13102_, _13101_, _13098_);
  or (_13103_, _13102_, _06474_);
  and (_13104_, _09027_, _07931_);
  or (_13105_, _13104_, _13041_);
  or (_13106_, _13105_, _07282_);
  and (_13107_, _13106_, _07284_);
  and (_13108_, _13107_, _13103_);
  or (_13109_, _13108_, _13044_);
  and (_13110_, _13109_, _07279_);
  or (_13111_, _13041_, _08073_);
  and (_13112_, _13100_, _06478_);
  and (_13113_, _13112_, _13111_);
  or (_13114_, _13113_, _13110_);
  and (_13115_, _13114_, _07276_);
  and (_13116_, _13057_, _06569_);
  and (_13117_, _13116_, _13111_);
  or (_13118_, _13117_, _06479_);
  or (_13119_, _13118_, _13115_);
  and (_13120_, _09026_, _07931_);
  or (_13121_, _13041_, _09043_);
  or (_13122_, _13121_, _13120_);
  and (_13123_, _13122_, _09048_);
  and (_13124_, _13123_, _13119_);
  nor (_13125_, _09033_, _13040_);
  or (_13126_, _13125_, _13041_);
  and (_13127_, _13126_, _06572_);
  or (_13128_, _13127_, _06606_);
  or (_13129_, _13128_, _13124_);
  or (_13130_, _13054_, _07037_);
  and (_13131_, _13130_, _06807_);
  and (_13132_, _13131_, _13129_);
  and (_13133_, _13051_, _06234_);
  or (_13134_, _13133_, _06195_);
  or (_13135_, _13134_, _13132_);
  and (_13136_, _08530_, _07931_);
  or (_13137_, _13041_, _06196_);
  or (_13138_, _13137_, _13136_);
  and (_13139_, _13138_, _01375_);
  and (_13140_, _13139_, _13135_);
  nor (_13141_, \uc8051golden_1.P2 [7], rst);
  nor (_13142_, _13141_, _01382_);
  or (_40337_, _13142_, _13140_);
  not (_13143_, _07945_);
  and (_13144_, _13143_, \uc8051golden_1.P3 [7]);
  and (_13145_, _09034_, _07945_);
  or (_13146_, _13145_, _13144_);
  and (_13147_, _13146_, _06582_);
  nor (_13148_, _13143_, _08070_);
  or (_13149_, _13148_, _13144_);
  or (_13150_, _13149_, _06293_);
  not (_13151_, _08598_);
  and (_13152_, _13151_, \uc8051golden_1.P3 [7]);
  and (_13153_, _08639_, _08598_);
  or (_13154_, _13153_, _13152_);
  and (_13155_, _13154_, _06393_);
  and (_13156_, _08762_, _07945_);
  or (_13157_, _13156_, _13144_);
  or (_13158_, _13157_, _07210_);
  and (_13159_, _07945_, \uc8051golden_1.ACC [7]);
  or (_13160_, _13159_, _13144_);
  and (_13161_, _13160_, _07199_);
  and (_13162_, _07200_, \uc8051golden_1.P3 [7]);
  or (_13163_, _13162_, _06401_);
  or (_13164_, _13163_, _13161_);
  and (_13165_, _13164_, _06396_);
  and (_13166_, _13165_, _13158_);
  and (_13167_, _08635_, _08598_);
  or (_13168_, _13167_, _13152_);
  and (_13169_, _13168_, _06395_);
  or (_13170_, _13169_, _06399_);
  or (_13171_, _13170_, _13166_);
  or (_13172_, _13149_, _07221_);
  and (_13173_, _13172_, _13171_);
  or (_13174_, _13173_, _06406_);
  or (_13175_, _13160_, _06414_);
  and (_13176_, _13175_, _06844_);
  and (_13177_, _13176_, _13174_);
  or (_13178_, _13177_, _13155_);
  and (_13179_, _13178_, _07245_);
  and (_13180_, _08636_, _08598_);
  or (_13181_, _13180_, _13152_);
  and (_13182_, _13181_, _06387_);
  or (_13183_, _13182_, _13179_);
  and (_13184_, _13183_, _06446_);
  and (_13185_, _08794_, _08598_);
  or (_13186_, _13185_, _13152_);
  and (_13187_, _13186_, _06300_);
  or (_13188_, _13187_, _10059_);
  or (_13189_, _13188_, _13184_);
  and (_13190_, _13189_, _13150_);
  or (_13191_, _13190_, _06281_);
  and (_13192_, _07945_, _08749_);
  or (_13193_, _13144_, _06282_);
  or (_13194_, _13193_, _13192_);
  and (_13195_, _13194_, _06279_);
  and (_13196_, _13195_, _13191_);
  and (_13197_, _09009_, _07945_);
  or (_13198_, _13197_, _13144_);
  and (_13199_, _13198_, _06015_);
  or (_13200_, _13199_, _06275_);
  or (_13201_, _13200_, _13196_);
  and (_13202_, _08813_, _07945_);
  or (_13203_, _13202_, _13144_);
  or (_13204_, _13203_, _06276_);
  and (_13205_, _13204_, _13201_);
  or (_13206_, _13205_, _06474_);
  and (_13207_, _09027_, _07945_);
  or (_13208_, _13207_, _13144_);
  or (_13209_, _13208_, _07282_);
  and (_13210_, _13209_, _07284_);
  and (_13211_, _13210_, _13206_);
  or (_13212_, _13211_, _13147_);
  and (_13213_, _13212_, _07279_);
  or (_13214_, _13144_, _08073_);
  and (_13215_, _13203_, _06478_);
  and (_13216_, _13215_, _13214_);
  or (_13217_, _13216_, _13213_);
  and (_13218_, _13217_, _07276_);
  and (_13219_, _13160_, _06569_);
  and (_13220_, _13219_, _13214_);
  or (_13221_, _13220_, _06479_);
  or (_13222_, _13221_, _13218_);
  and (_13223_, _09026_, _07945_);
  or (_13224_, _13144_, _09043_);
  or (_13225_, _13224_, _13223_);
  and (_13226_, _13225_, _09048_);
  and (_13227_, _13226_, _13222_);
  nor (_13228_, _09033_, _13143_);
  or (_13229_, _13228_, _13144_);
  and (_13230_, _13229_, _06572_);
  or (_13231_, _13230_, _06606_);
  or (_13232_, _13231_, _13227_);
  or (_13233_, _13157_, _07037_);
  and (_13234_, _13233_, _06807_);
  and (_13235_, _13234_, _13232_);
  and (_13236_, _13154_, _06234_);
  or (_13237_, _13236_, _06195_);
  or (_13238_, _13237_, _13235_);
  and (_13239_, _08530_, _07945_);
  or (_13240_, _13144_, _06196_);
  or (_13241_, _13240_, _13239_);
  and (_13242_, _13241_, _01375_);
  and (_13243_, _13242_, _13238_);
  nor (_13244_, \uc8051golden_1.P3 [7], rst);
  nor (_13245_, _13244_, _01382_);
  or (_40338_, _13245_, _13243_);
  not (_13246_, _08019_);
  and (_13247_, _13246_, \uc8051golden_1.P0 [7]);
  and (_13248_, _09034_, _08019_);
  or (_13249_, _13248_, _13247_);
  and (_13250_, _13249_, _06582_);
  nor (_13251_, _13246_, _08070_);
  or (_13252_, _13251_, _13247_);
  or (_13253_, _13252_, _06293_);
  not (_13254_, _07959_);
  and (_13255_, _13254_, \uc8051golden_1.P0 [7]);
  and (_13256_, _08639_, _07959_);
  or (_13257_, _13256_, _13255_);
  and (_13258_, _13257_, _06393_);
  and (_13259_, _08762_, _08019_);
  or (_13260_, _13259_, _13247_);
  or (_13261_, _13260_, _07210_);
  and (_13262_, _08019_, \uc8051golden_1.ACC [7]);
  or (_13263_, _13262_, _13247_);
  and (_13264_, _13263_, _07199_);
  and (_13265_, _07200_, \uc8051golden_1.P0 [7]);
  or (_13266_, _13265_, _06401_);
  or (_13267_, _13266_, _13264_);
  and (_13268_, _13267_, _06396_);
  and (_13269_, _13268_, _13261_);
  and (_13270_, _08635_, _07959_);
  or (_13271_, _13270_, _13255_);
  and (_13272_, _13271_, _06395_);
  or (_13273_, _13272_, _06399_);
  or (_13274_, _13273_, _13269_);
  or (_13275_, _13252_, _07221_);
  and (_13276_, _13275_, _13274_);
  or (_13277_, _13276_, _06406_);
  or (_13278_, _13263_, _06414_);
  and (_13279_, _13278_, _06844_);
  and (_13280_, _13279_, _13277_);
  or (_13281_, _13280_, _13258_);
  and (_13282_, _13281_, _07245_);
  and (_13283_, _08636_, _07959_);
  or (_13284_, _13283_, _13255_);
  and (_13285_, _13284_, _06387_);
  or (_13286_, _13285_, _13282_);
  and (_13287_, _13286_, _06446_);
  and (_13288_, _08794_, _07959_);
  or (_13289_, _13288_, _13255_);
  and (_13290_, _13289_, _06300_);
  or (_13291_, _13290_, _10059_);
  or (_13292_, _13291_, _13287_);
  and (_13293_, _13292_, _13253_);
  or (_13294_, _13293_, _06281_);
  and (_13295_, _08019_, _08749_);
  or (_13296_, _13247_, _06282_);
  or (_13297_, _13296_, _13295_);
  and (_13298_, _13297_, _06279_);
  and (_13299_, _13298_, _13294_);
  and (_13300_, _09009_, _08019_);
  or (_13301_, _13300_, _13247_);
  and (_13302_, _13301_, _06015_);
  or (_13303_, _13302_, _06275_);
  or (_13304_, _13303_, _13299_);
  and (_13305_, _08813_, _08019_);
  or (_13306_, _13305_, _13247_);
  or (_13307_, _13306_, _06276_);
  and (_13308_, _13307_, _13304_);
  or (_13309_, _13308_, _06474_);
  and (_13310_, _09027_, _08019_);
  or (_13311_, _13310_, _13247_);
  or (_13312_, _13311_, _07282_);
  and (_13313_, _13312_, _07284_);
  and (_13314_, _13313_, _13309_);
  or (_13315_, _13314_, _13250_);
  and (_13316_, _13315_, _07279_);
  or (_13317_, _13247_, _08073_);
  and (_13318_, _13306_, _06478_);
  and (_13319_, _13318_, _13317_);
  or (_13320_, _13319_, _13316_);
  and (_13321_, _13320_, _07276_);
  and (_13322_, _13263_, _06569_);
  and (_13323_, _13322_, _13317_);
  or (_13324_, _13323_, _06479_);
  or (_13325_, _13324_, _13321_);
  and (_13326_, _09026_, _08019_);
  or (_13327_, _13247_, _09043_);
  or (_13328_, _13327_, _13326_);
  and (_13329_, _13328_, _09048_);
  and (_13330_, _13329_, _13325_);
  nor (_13331_, _09033_, _13246_);
  or (_13332_, _13331_, _13247_);
  and (_13333_, _13332_, _06572_);
  or (_13334_, _13333_, _06606_);
  or (_13335_, _13334_, _13330_);
  or (_13336_, _13260_, _07037_);
  and (_13337_, _13336_, _06807_);
  and (_13338_, _13337_, _13335_);
  and (_13339_, _13257_, _06234_);
  or (_13340_, _13339_, _06195_);
  or (_13341_, _13340_, _13338_);
  and (_13342_, _08530_, _08019_);
  or (_13343_, _13247_, _06196_);
  or (_13344_, _13343_, _13342_);
  and (_13345_, _13344_, _01375_);
  and (_13346_, _13345_, _13341_);
  nor (_13347_, \uc8051golden_1.P0 [7], rst);
  nor (_13348_, _13347_, _01382_);
  or (_40339_, _13348_, _13346_);
  nor (_13349_, \uc8051golden_1.P1 [7], rst);
  nor (_13350_, _13349_, _01382_);
  not (_13351_, _07970_);
  and (_13352_, _13351_, \uc8051golden_1.P1 [7]);
  and (_13353_, _09034_, _07970_);
  or (_13354_, _13353_, _13352_);
  and (_13355_, _13354_, _06582_);
  nor (_13356_, _13351_, _08070_);
  or (_13357_, _13356_, _13352_);
  or (_13358_, _13357_, _06293_);
  not (_13359_, _08626_);
  and (_13360_, _13359_, \uc8051golden_1.P1 [7]);
  and (_13361_, _08639_, _08626_);
  or (_13362_, _13361_, _13360_);
  and (_13363_, _13362_, _06393_);
  and (_13364_, _08762_, _07970_);
  or (_13365_, _13364_, _13352_);
  or (_13366_, _13365_, _07210_);
  and (_13367_, _07970_, \uc8051golden_1.ACC [7]);
  or (_13368_, _13367_, _13352_);
  and (_13369_, _13368_, _07199_);
  and (_13370_, _07200_, \uc8051golden_1.P1 [7]);
  or (_13371_, _13370_, _06401_);
  or (_13372_, _13371_, _13369_);
  and (_13373_, _13372_, _06396_);
  and (_13374_, _13373_, _13366_);
  and (_13375_, _08635_, _08626_);
  or (_13376_, _13375_, _13360_);
  and (_13377_, _13376_, _06395_);
  or (_13378_, _13377_, _06399_);
  or (_13379_, _13378_, _13374_);
  or (_13380_, _13357_, _07221_);
  and (_13381_, _13380_, _13379_);
  or (_13382_, _13381_, _06406_);
  or (_13383_, _13368_, _06414_);
  and (_13384_, _13383_, _06844_);
  and (_13385_, _13384_, _13382_);
  or (_13386_, _13385_, _13363_);
  and (_13387_, _13386_, _07245_);
  or (_13388_, _13360_, _08634_);
  and (_13389_, _13388_, _06387_);
  and (_13390_, _13389_, _13376_);
  or (_13391_, _13390_, _13387_);
  and (_13392_, _13391_, _06446_);
  and (_13393_, _08794_, _08626_);
  or (_13394_, _13393_, _13360_);
  and (_13395_, _13394_, _06300_);
  or (_13396_, _13395_, _10059_);
  or (_13397_, _13396_, _13392_);
  and (_13398_, _13397_, _13358_);
  or (_13399_, _13398_, _06281_);
  and (_13400_, _07970_, _08749_);
  or (_13401_, _13352_, _06282_);
  or (_13402_, _13401_, _13400_);
  and (_13403_, _13402_, _06279_);
  and (_13404_, _13403_, _13399_);
  and (_13405_, _09009_, _07970_);
  or (_13406_, _13405_, _13352_);
  and (_13407_, _13406_, _06015_);
  or (_13408_, _13407_, _06275_);
  or (_13409_, _13408_, _13404_);
  and (_13410_, _08813_, _07970_);
  or (_13411_, _13410_, _13352_);
  or (_13412_, _13411_, _06276_);
  and (_13413_, _13412_, _13409_);
  or (_13414_, _13413_, _06474_);
  and (_13415_, _09027_, _07970_);
  or (_13416_, _13415_, _13352_);
  or (_13417_, _13416_, _07282_);
  and (_13418_, _13417_, _07284_);
  and (_13419_, _13418_, _13414_);
  or (_13420_, _13419_, _13355_);
  and (_13421_, _13420_, _07279_);
  or (_13422_, _13352_, _08073_);
  and (_13423_, _13411_, _06478_);
  and (_13424_, _13423_, _13422_);
  or (_13425_, _13424_, _13421_);
  and (_13426_, _13425_, _07276_);
  and (_13427_, _13368_, _06569_);
  and (_13428_, _13427_, _13422_);
  or (_13429_, _13428_, _06479_);
  or (_13430_, _13429_, _13426_);
  and (_13431_, _09026_, _07970_);
  or (_13432_, _13352_, _09043_);
  or (_13433_, _13432_, _13431_);
  and (_13434_, _13433_, _09048_);
  and (_13435_, _13434_, _13430_);
  nor (_13436_, _09033_, _13351_);
  or (_13437_, _13436_, _13352_);
  and (_13438_, _13437_, _06572_);
  or (_13439_, _13438_, _06606_);
  or (_13440_, _13439_, _13435_);
  or (_13441_, _13365_, _07037_);
  and (_13442_, _13441_, _06807_);
  and (_13443_, _13442_, _13440_);
  and (_13444_, _13362_, _06234_);
  or (_13445_, _13444_, _06195_);
  or (_13446_, _13445_, _13443_);
  and (_13447_, _08530_, _07970_);
  or (_13448_, _13352_, _06196_);
  or (_13449_, _13448_, _13447_);
  and (_13450_, _13449_, _01375_);
  and (_13451_, _13450_, _13446_);
  or (_40340_, _13451_, _13350_);
  and (_13452_, _01379_, \uc8051golden_1.IP [7]);
  not (_13453_, _07999_);
  and (_13454_, _13453_, \uc8051golden_1.IP [7]);
  and (_13455_, _09034_, _07999_);
  or (_13456_, _13455_, _13454_);
  and (_13457_, _13456_, _06582_);
  nor (_13458_, _13453_, _08070_);
  or (_13459_, _13458_, _13454_);
  or (_13460_, _13459_, _06293_);
  not (_13461_, _08614_);
  and (_13462_, _13461_, \uc8051golden_1.IP [7]);
  and (_13463_, _08639_, _08614_);
  or (_13464_, _13463_, _13462_);
  and (_13465_, _13464_, _06393_);
  and (_13466_, _08762_, _07999_);
  or (_13467_, _13466_, _13454_);
  or (_13468_, _13467_, _07210_);
  and (_13469_, _07999_, \uc8051golden_1.ACC [7]);
  or (_13470_, _13469_, _13454_);
  and (_13471_, _13470_, _07199_);
  and (_13472_, _07200_, \uc8051golden_1.IP [7]);
  or (_13473_, _13472_, _06401_);
  or (_13474_, _13473_, _13471_);
  and (_13475_, _13474_, _06396_);
  and (_13476_, _13475_, _13468_);
  and (_13477_, _08635_, _08614_);
  or (_13478_, _13477_, _13462_);
  and (_13479_, _13478_, _06395_);
  or (_13480_, _13479_, _06399_);
  or (_13481_, _13480_, _13476_);
  or (_13482_, _13459_, _07221_);
  and (_13483_, _13482_, _13481_);
  or (_13484_, _13483_, _06406_);
  or (_13485_, _13470_, _06414_);
  and (_13486_, _13485_, _06844_);
  and (_13487_, _13486_, _13484_);
  or (_13488_, _13487_, _13465_);
  and (_13489_, _13488_, _07245_);
  and (_13490_, _08636_, _08614_);
  or (_13491_, _13490_, _13462_);
  and (_13492_, _13491_, _06387_);
  or (_13493_, _13492_, _13489_);
  and (_13494_, _13493_, _06446_);
  and (_13495_, _08794_, _08614_);
  or (_13496_, _13495_, _13462_);
  and (_13497_, _13496_, _06300_);
  or (_13498_, _13497_, _10059_);
  or (_13499_, _13498_, _13494_);
  and (_13500_, _13499_, _13460_);
  or (_13501_, _13500_, _06281_);
  and (_13502_, _07999_, _08749_);
  or (_13503_, _13454_, _06282_);
  or (_13504_, _13503_, _13502_);
  and (_13505_, _13504_, _06279_);
  and (_13506_, _13505_, _13501_);
  and (_13507_, _09009_, _07999_);
  or (_13508_, _13507_, _13454_);
  and (_13509_, _13508_, _06015_);
  or (_13510_, _13509_, _06275_);
  or (_13511_, _13510_, _13506_);
  and (_13512_, _08813_, _07999_);
  or (_13513_, _13512_, _13454_);
  or (_13514_, _13513_, _06276_);
  and (_13515_, _13514_, _13511_);
  or (_13516_, _13515_, _06474_);
  and (_13517_, _09027_, _07999_);
  or (_13518_, _13517_, _13454_);
  or (_13519_, _13518_, _07282_);
  and (_13520_, _13519_, _07284_);
  and (_13521_, _13520_, _13516_);
  or (_13522_, _13521_, _13457_);
  and (_13523_, _13522_, _07279_);
  or (_13524_, _13454_, _08073_);
  and (_13525_, _13513_, _06478_);
  and (_13526_, _13525_, _13524_);
  or (_13527_, _13526_, _13523_);
  and (_13528_, _13527_, _07276_);
  and (_13529_, _13470_, _06569_);
  and (_13530_, _13529_, _13524_);
  or (_13531_, _13530_, _06479_);
  or (_13532_, _13531_, _13528_);
  and (_13533_, _09026_, _07999_);
  or (_13534_, _13454_, _09043_);
  or (_13535_, _13534_, _13533_);
  and (_13536_, _13535_, _09048_);
  and (_13537_, _13536_, _13532_);
  nor (_13538_, _09033_, _13453_);
  or (_13539_, _13538_, _13454_);
  and (_13540_, _13539_, _06572_);
  or (_13541_, _13540_, _06606_);
  or (_13542_, _13541_, _13537_);
  or (_13543_, _13467_, _07037_);
  and (_13544_, _13543_, _06807_);
  and (_13545_, _13544_, _13542_);
  and (_13546_, _13464_, _06234_);
  or (_13547_, _13546_, _06195_);
  or (_13548_, _13547_, _13545_);
  and (_13549_, _08530_, _07999_);
  or (_13550_, _13454_, _06196_);
  or (_13551_, _13550_, _13549_);
  and (_13552_, _13551_, _01375_);
  and (_13553_, _13552_, _13548_);
  or (_13554_, _13553_, _13452_);
  and (_40341_, _13554_, _42545_);
  and (_13555_, _01379_, \uc8051golden_1.IE [7]);
  not (_13556_, _07948_);
  and (_13557_, _13556_, \uc8051golden_1.IE [7]);
  and (_13558_, _09034_, _07948_);
  or (_13559_, _13558_, _13557_);
  and (_13560_, _13559_, _06582_);
  nor (_13561_, _13556_, _08070_);
  or (_13562_, _13561_, _13557_);
  or (_13563_, _13562_, _06293_);
  not (_13564_, _08603_);
  and (_13565_, _13564_, \uc8051golden_1.IE [7]);
  and (_13566_, _08639_, _08603_);
  or (_13567_, _13566_, _13565_);
  and (_13568_, _13567_, _06393_);
  and (_13569_, _08762_, _07948_);
  or (_13570_, _13569_, _13557_);
  or (_13571_, _13570_, _07210_);
  and (_13572_, _07948_, \uc8051golden_1.ACC [7]);
  or (_13573_, _13572_, _13557_);
  and (_13574_, _13573_, _07199_);
  and (_13575_, _07200_, \uc8051golden_1.IE [7]);
  or (_13576_, _13575_, _06401_);
  or (_13577_, _13576_, _13574_);
  and (_13578_, _13577_, _06396_);
  and (_13579_, _13578_, _13571_);
  and (_13580_, _08635_, _08603_);
  or (_13581_, _13580_, _13565_);
  and (_13582_, _13581_, _06395_);
  or (_13583_, _13582_, _06399_);
  or (_13584_, _13583_, _13579_);
  or (_13585_, _13562_, _07221_);
  and (_13586_, _13585_, _13584_);
  or (_13587_, _13586_, _06406_);
  or (_13588_, _13573_, _06414_);
  and (_13589_, _13588_, _06844_);
  and (_13590_, _13589_, _13587_);
  or (_13591_, _13590_, _13568_);
  and (_13592_, _13591_, _07245_);
  and (_13593_, _08636_, _08603_);
  or (_13594_, _13593_, _13565_);
  and (_13595_, _13594_, _06387_);
  or (_13596_, _13595_, _13592_);
  and (_13597_, _13596_, _06446_);
  and (_13598_, _08794_, _08603_);
  or (_13599_, _13598_, _13565_);
  and (_13600_, _13599_, _06300_);
  or (_13601_, _13600_, _10059_);
  or (_13602_, _13601_, _13597_);
  and (_13603_, _13602_, _13563_);
  or (_13604_, _13603_, _06281_);
  and (_13605_, _07948_, _08749_);
  or (_13606_, _13557_, _06282_);
  or (_13607_, _13606_, _13605_);
  and (_13608_, _13607_, _06279_);
  and (_13609_, _13608_, _13604_);
  and (_13610_, _09009_, _07948_);
  or (_13612_, _13610_, _13557_);
  and (_13613_, _13612_, _06015_);
  or (_13614_, _13613_, _06275_);
  or (_13615_, _13614_, _13609_);
  and (_13616_, _08813_, _07948_);
  or (_13617_, _13616_, _13557_);
  or (_13618_, _13617_, _06276_);
  and (_13619_, _13618_, _13615_);
  or (_13620_, _13619_, _06474_);
  and (_13621_, _09027_, _07948_);
  or (_13623_, _13621_, _13557_);
  or (_13624_, _13623_, _07282_);
  and (_13625_, _13624_, _07284_);
  and (_13626_, _13625_, _13620_);
  or (_13627_, _13626_, _13560_);
  and (_13628_, _13627_, _07279_);
  or (_13629_, _13557_, _08073_);
  and (_13630_, _13617_, _06478_);
  and (_13631_, _13630_, _13629_);
  or (_13632_, _13631_, _13628_);
  and (_13634_, _13632_, _07276_);
  and (_13635_, _13573_, _06569_);
  and (_13636_, _13635_, _13629_);
  or (_13637_, _13636_, _06479_);
  or (_13638_, _13637_, _13634_);
  and (_13639_, _09026_, _07948_);
  or (_13640_, _13557_, _09043_);
  or (_13641_, _13640_, _13639_);
  and (_13642_, _13641_, _09048_);
  and (_13643_, _13642_, _13638_);
  nor (_13645_, _09033_, _13556_);
  or (_13646_, _13645_, _13557_);
  and (_13647_, _13646_, _06572_);
  or (_13648_, _13647_, _06606_);
  or (_13649_, _13648_, _13643_);
  or (_13650_, _13570_, _07037_);
  and (_13651_, _13650_, _06807_);
  and (_13652_, _13651_, _13649_);
  and (_13653_, _13567_, _06234_);
  or (_13654_, _13653_, _06195_);
  or (_13656_, _13654_, _13652_);
  and (_13657_, _08530_, _07948_);
  or (_13658_, _13557_, _06196_);
  or (_13659_, _13658_, _13657_);
  and (_13660_, _13659_, _01375_);
  and (_13661_, _13660_, _13656_);
  or (_13662_, _13661_, _13555_);
  and (_40342_, _13662_, _42545_);
  and (_13663_, _01379_, \uc8051golden_1.SCON [7]);
  not (_13664_, _07972_);
  and (_13666_, _13664_, \uc8051golden_1.SCON [7]);
  and (_13667_, _09034_, _07972_);
  or (_13668_, _13667_, _13666_);
  and (_13669_, _13668_, _06582_);
  nor (_13670_, _13664_, _08070_);
  or (_13671_, _13670_, _13666_);
  or (_13672_, _13671_, _06293_);
  not (_13673_, _08606_);
  and (_13674_, _13673_, \uc8051golden_1.SCON [7]);
  and (_13675_, _08639_, _08606_);
  or (_13677_, _13675_, _13674_);
  and (_13678_, _13677_, _06393_);
  and (_13679_, _08762_, _07972_);
  or (_13680_, _13679_, _13666_);
  or (_13681_, _13680_, _07210_);
  and (_13682_, _07972_, \uc8051golden_1.ACC [7]);
  or (_13683_, _13682_, _13666_);
  and (_13684_, _13683_, _07199_);
  and (_13685_, _07200_, \uc8051golden_1.SCON [7]);
  or (_13686_, _13685_, _06401_);
  or (_13688_, _13686_, _13684_);
  and (_13689_, _13688_, _06396_);
  and (_13690_, _13689_, _13681_);
  and (_13691_, _08635_, _08606_);
  or (_13692_, _13691_, _13674_);
  and (_13693_, _13692_, _06395_);
  or (_13694_, _13693_, _06399_);
  or (_13695_, _13694_, _13690_);
  or (_13696_, _13671_, _07221_);
  and (_13697_, _13696_, _13695_);
  or (_13699_, _13697_, _06406_);
  or (_13700_, _13683_, _06414_);
  and (_13701_, _13700_, _06844_);
  and (_13702_, _13701_, _13699_);
  or (_13703_, _13702_, _13678_);
  and (_13704_, _13703_, _07245_);
  and (_13705_, _08636_, _08606_);
  or (_13706_, _13705_, _13674_);
  and (_13707_, _13706_, _06387_);
  or (_13708_, _13707_, _13704_);
  and (_13710_, _13708_, _06446_);
  and (_13711_, _08794_, _08606_);
  or (_13712_, _13711_, _13674_);
  and (_13713_, _13712_, _06300_);
  or (_13714_, _13713_, _10059_);
  or (_13715_, _13714_, _13710_);
  and (_13716_, _13715_, _13672_);
  or (_13717_, _13716_, _06281_);
  and (_13718_, _07972_, _08749_);
  or (_13719_, _13666_, _06282_);
  or (_13721_, _13719_, _13718_);
  and (_13722_, _13721_, _06279_);
  and (_13723_, _13722_, _13717_);
  and (_13724_, _09009_, _07972_);
  or (_13725_, _13724_, _13666_);
  and (_13726_, _13725_, _06015_);
  or (_13727_, _13726_, _06275_);
  or (_13728_, _13727_, _13723_);
  and (_13729_, _08813_, _07972_);
  or (_13730_, _13729_, _13666_);
  or (_13732_, _13730_, _06276_);
  and (_13733_, _13732_, _13728_);
  or (_13734_, _13733_, _06474_);
  and (_13735_, _09027_, _07972_);
  or (_13736_, _13735_, _13666_);
  or (_13737_, _13736_, _07282_);
  and (_13738_, _13737_, _07284_);
  and (_13739_, _13738_, _13734_);
  or (_13740_, _13739_, _13669_);
  and (_13741_, _13740_, _07279_);
  or (_13743_, _13666_, _08073_);
  and (_13744_, _13730_, _06478_);
  and (_13745_, _13744_, _13743_);
  or (_13746_, _13745_, _13741_);
  and (_13747_, _13746_, _07276_);
  and (_13748_, _13683_, _06569_);
  and (_13749_, _13748_, _13743_);
  or (_13750_, _13749_, _06479_);
  or (_13751_, _13750_, _13747_);
  and (_13752_, _09026_, _07972_);
  or (_13754_, _13666_, _09043_);
  or (_13755_, _13754_, _13752_);
  and (_13756_, _13755_, _09048_);
  and (_13757_, _13756_, _13751_);
  nor (_13758_, _09033_, _13664_);
  or (_13759_, _13758_, _13666_);
  and (_13760_, _13759_, _06572_);
  or (_13761_, _13760_, _06606_);
  or (_13762_, _13761_, _13757_);
  or (_13763_, _13680_, _07037_);
  and (_13764_, _13763_, _06807_);
  and (_13765_, _13764_, _13762_);
  and (_13766_, _13677_, _06234_);
  or (_13767_, _13766_, _06195_);
  or (_13768_, _13767_, _13765_);
  and (_13769_, _08530_, _07972_);
  or (_13770_, _13666_, _06196_);
  or (_13771_, _13770_, _13769_);
  and (_13772_, _13771_, _01375_);
  and (_13773_, _13772_, _13768_);
  or (_13774_, _13773_, _13663_);
  and (_40343_, _13774_, _42545_);
  not (_13775_, \uc8051golden_1.SP [7]);
  nor (_13776_, _01375_, _13775_);
  and (_13777_, _07781_, \uc8051golden_1.SP [4]);
  and (_13778_, _13777_, \uc8051golden_1.SP [5]);
  and (_13779_, _13778_, \uc8051golden_1.SP [6]);
  or (_13780_, _13779_, \uc8051golden_1.SP [7]);
  nand (_13781_, _13779_, \uc8051golden_1.SP [7]);
  and (_13782_, _13781_, _13780_);
  or (_13783_, _13782_, _07312_);
  nor (_13784_, _07956_, _13775_);
  and (_13785_, _09034_, _08236_);
  or (_13786_, _13785_, _13784_);
  and (_13787_, _13786_, _06582_);
  not (_13788_, _06294_);
  not (_13789_, _08236_);
  nor (_13790_, _13789_, _08070_);
  or (_13791_, _13784_, _06281_);
  or (_13792_, _13791_, _13790_);
  and (_13793_, _13792_, _13788_);
  and (_13794_, _08762_, _08236_);
  or (_13795_, _13794_, _13784_);
  or (_13796_, _13795_, _07210_);
  and (_13797_, _07956_, \uc8051golden_1.ACC [7]);
  or (_13798_, _13797_, _13784_);
  or (_13799_, _13798_, _07200_);
  or (_13800_, _07199_, \uc8051golden_1.SP [7]);
  and (_13801_, _13800_, _07366_);
  and (_13802_, _13801_, _13799_);
  and (_13803_, _13782_, _06790_);
  or (_13804_, _13803_, _06401_);
  or (_13805_, _13804_, _13802_);
  and (_13806_, _13805_, _05997_);
  and (_13807_, _13806_, _13796_);
  and (_13808_, _13782_, _07351_);
  or (_13809_, _13808_, _06399_);
  or (_13810_, _13809_, _13807_);
  not (_13811_, \uc8051golden_1.SP [6]);
  not (_13812_, \uc8051golden_1.SP [5]);
  not (_13813_, \uc8051golden_1.SP [4]);
  and (_13814_, _08664_, _13813_);
  and (_13815_, _13814_, _13812_);
  and (_13816_, _13815_, _13811_);
  and (_13817_, _13816_, _06270_);
  nor (_13818_, _13817_, _13775_);
  and (_13819_, _13817_, _13775_);
  nor (_13820_, _13819_, _13818_);
  nand (_13821_, _13820_, _06399_);
  and (_13822_, _13821_, _13810_);
  or (_13823_, _13822_, _06406_);
  or (_13824_, _13798_, _06414_);
  and (_13825_, _13824_, _07785_);
  and (_13826_, _13825_, _13823_);
  and (_13827_, _13778_, \uc8051golden_1.SP [0]);
  and (_13828_, _13827_, \uc8051golden_1.SP [6]);
  nor (_13829_, _13828_, _13775_);
  and (_13830_, _13828_, _13775_);
  or (_13831_, _13830_, _13829_);
  nand (_13832_, _13831_, _06419_);
  nand (_13833_, _13832_, _07350_);
  or (_13834_, _13833_, _13826_);
  or (_13835_, _13782_, _07350_);
  and (_13836_, _13835_, _06293_);
  and (_13837_, _13836_, _13834_);
  or (_13838_, _13837_, _13793_);
  or (_13839_, _13784_, _06282_);
  and (_13840_, _07956_, _08749_);
  or (_13841_, _13840_, _13839_);
  and (_13842_, _13841_, _06279_);
  and (_13843_, _13842_, _13838_);
  and (_13844_, _09009_, _07956_);
  or (_13845_, _13844_, _13784_);
  and (_13846_, _13845_, _06015_);
  or (_13847_, _13846_, _06275_);
  or (_13848_, _13847_, _13843_);
  and (_13849_, _08813_, _07956_);
  or (_13850_, _13849_, _13784_);
  or (_13851_, _13850_, _06276_);
  and (_13852_, _13851_, _13848_);
  or (_13853_, _13852_, _05943_);
  not (_13854_, _05943_);
  or (_13855_, _13782_, _13854_);
  and (_13856_, _13855_, _13853_);
  or (_13857_, _13856_, _06474_);
  and (_13858_, _09027_, _07956_);
  or (_13859_, _13858_, _13784_);
  or (_13860_, _13859_, _07282_);
  and (_13861_, _13860_, _07284_);
  and (_13862_, _13861_, _13857_);
  or (_13863_, _13862_, _13787_);
  and (_13864_, _13863_, _07279_);
  or (_13865_, _13784_, _08073_);
  and (_13866_, _13850_, _06478_);
  and (_13867_, _13866_, _13865_);
  or (_13868_, _13867_, _13864_);
  and (_13869_, _13868_, _12731_);
  and (_13870_, _13798_, _06569_);
  and (_13871_, _13870_, _13865_);
  and (_13872_, _13782_, _05956_);
  or (_13873_, _13872_, _06479_);
  or (_13874_, _13873_, _13871_);
  or (_13875_, _13874_, _13869_);
  and (_13876_, _09026_, _07956_);
  or (_13877_, _13876_, _13784_);
  or (_13878_, _13877_, _09043_);
  and (_13879_, _13878_, _13875_);
  or (_13880_, _13879_, _06572_);
  not (_13881_, _06588_);
  nor (_13882_, _09033_, _13789_);
  or (_13883_, _13784_, _09048_);
  or (_13884_, _13883_, _13882_);
  and (_13885_, _13884_, _13881_);
  and (_13886_, _13885_, _13880_);
  or (_13887_, _13816_, \uc8051golden_1.SP [7]);
  nand (_13888_, _13816_, \uc8051golden_1.SP [7]);
  and (_13889_, _13888_, _13887_);
  and (_13890_, _13889_, _06588_);
  or (_13891_, _13890_, _05966_);
  or (_13892_, _13891_, _13886_);
  or (_13893_, _13782_, _05967_);
  and (_13894_, _13893_, _13892_);
  or (_13895_, _13894_, _06305_);
  or (_13896_, _13889_, _06306_);
  and (_13897_, _13896_, _07037_);
  and (_13898_, _13897_, _13895_);
  and (_13899_, _13795_, _06606_);
  or (_13900_, _13899_, _07887_);
  or (_13901_, _13900_, _13898_);
  and (_13902_, _13901_, _13783_);
  or (_13903_, _13902_, _06195_);
  and (_13904_, _08530_, _08236_);
  or (_13905_, _13784_, _06196_);
  or (_13906_, _13905_, _13904_);
  and (_13907_, _13906_, _01375_);
  and (_13908_, _13907_, _13903_);
  or (_13909_, _13908_, _13776_);
  and (_40345_, _13909_, _42545_);
  not (_13910_, _07940_);
  and (_13911_, _13910_, \uc8051golden_1.SBUF [7]);
  and (_13912_, _09034_, _07940_);
  or (_13913_, _13912_, _13911_);
  and (_13914_, _13913_, _06582_);
  and (_13915_, _08762_, _07940_);
  or (_13916_, _13915_, _13911_);
  or (_13917_, _13916_, _07210_);
  and (_13918_, _07940_, \uc8051golden_1.ACC [7]);
  or (_13919_, _13918_, _13911_);
  and (_13920_, _13919_, _07199_);
  and (_13921_, _07200_, \uc8051golden_1.SBUF [7]);
  or (_13922_, _13921_, _06401_);
  or (_13923_, _13922_, _13920_);
  and (_13924_, _13923_, _07221_);
  and (_13925_, _13924_, _13917_);
  nor (_13926_, _13910_, _08070_);
  or (_13927_, _13926_, _13911_);
  and (_13928_, _13927_, _06399_);
  or (_13929_, _13928_, _13925_);
  and (_13930_, _13929_, _06414_);
  and (_13931_, _13919_, _06406_);
  or (_13932_, _13931_, _10059_);
  or (_13933_, _13932_, _13930_);
  or (_13934_, _13927_, _06293_);
  and (_13935_, _13934_, _13933_);
  or (_13936_, _13935_, _06281_);
  and (_13937_, _07940_, _08749_);
  or (_13938_, _13911_, _06282_);
  or (_13939_, _13938_, _13937_);
  and (_13940_, _13939_, _06279_);
  and (_13941_, _13940_, _13936_);
  and (_13942_, _09009_, _07940_);
  or (_13943_, _13942_, _13911_);
  and (_13944_, _13943_, _06015_);
  or (_13945_, _13944_, _06275_);
  or (_13946_, _13945_, _13941_);
  and (_13947_, _08813_, _07940_);
  or (_13948_, _13947_, _13911_);
  or (_13949_, _13948_, _06276_);
  and (_13950_, _13949_, _13946_);
  or (_13951_, _13950_, _06474_);
  and (_13952_, _09027_, _07940_);
  or (_13953_, _13952_, _13911_);
  or (_13954_, _13953_, _07282_);
  and (_13955_, _13954_, _07284_);
  and (_13956_, _13955_, _13951_);
  or (_13957_, _13956_, _13914_);
  and (_13958_, _13957_, _07279_);
  or (_13959_, _13911_, _08073_);
  and (_13960_, _13948_, _06478_);
  and (_13961_, _13960_, _13959_);
  or (_13962_, _13961_, _13958_);
  and (_13963_, _13962_, _07276_);
  and (_13964_, _13919_, _06569_);
  and (_13965_, _13964_, _13959_);
  or (_13966_, _13965_, _06479_);
  or (_13967_, _13966_, _13963_);
  and (_13968_, _09026_, _07940_);
  or (_13969_, _13911_, _09043_);
  or (_13970_, _13969_, _13968_);
  and (_13971_, _13970_, _09048_);
  and (_13972_, _13971_, _13967_);
  nor (_13973_, _09033_, _13910_);
  or (_13974_, _13973_, _13911_);
  and (_13975_, _13974_, _06572_);
  or (_13976_, _13975_, _06606_);
  or (_13977_, _13976_, _13972_);
  or (_13978_, _13916_, _07037_);
  and (_13979_, _13978_, _06196_);
  and (_13980_, _13979_, _13977_);
  and (_13981_, _08530_, _07940_);
  or (_13982_, _13981_, _13911_);
  and (_13983_, _13982_, _06195_);
  or (_13984_, _13983_, _01379_);
  or (_13985_, _13984_, _13980_);
  or (_13986_, _01375_, \uc8051golden_1.SBUF [7]);
  and (_13987_, _13986_, _42545_);
  and (_40346_, _13987_, _13985_);
  nor (_13988_, _01375_, _10524_);
  nor (_13989_, _08612_, _10524_);
  and (_13990_, _08639_, _08612_);
  or (_13991_, _13990_, _13989_);
  or (_13992_, _13991_, _06807_);
  nor (_13993_, _07988_, _10524_);
  not (_13994_, _07988_);
  nor (_13995_, _09033_, _13994_);
  or (_13996_, _13995_, _13993_);
  and (_13997_, _13996_, _06572_);
  and (_13998_, _09034_, _07988_);
  or (_13999_, _13998_, _13993_);
  and (_14000_, _13999_, _06582_);
  and (_14001_, _09009_, _07988_);
  or (_14002_, _14001_, _13993_);
  and (_14003_, _14002_, _06015_);
  nor (_14004_, _13994_, _08070_);
  or (_14005_, _14004_, _13993_);
  or (_14006_, _14005_, _06293_);
  and (_14007_, _10580_, _08073_);
  and (_14008_, _10590_, _10586_);
  nor (_14009_, _14008_, _10584_);
  nand (_14010_, _10632_, _10586_);
  or (_14011_, _14010_, _10630_);
  and (_14012_, _14011_, _14009_);
  or (_14013_, _14012_, _14007_);
  and (_14014_, _14013_, _06437_);
  not (_14015_, _06432_);
  not (_14016_, _06433_);
  nor (_14017_, _12958_, _14016_);
  and (_14018_, _08635_, _08612_);
  or (_14019_, _14018_, _13989_);
  or (_14020_, _13989_, _08634_);
  and (_14021_, _14020_, _06387_);
  and (_14022_, _14021_, _14019_);
  nand (_14023_, _08388_, \uc8051golden_1.ACC [3]);
  nor (_14024_, _08388_, \uc8051golden_1.ACC [3]);
  nor (_14025_, _08432_, \uc8051golden_1.ACC [2]);
  or (_14026_, _14025_, _14024_);
  and (_14027_, _14026_, _14023_);
  nor (_14028_, _08476_, \uc8051golden_1.ACC [1]);
  nor (_14029_, _08521_, _06045_);
  nor (_14030_, _14029_, _11224_);
  or (_14031_, _14030_, _14028_);
  and (_14032_, _14031_, _12536_);
  or (_14033_, _14032_, _14027_);
  and (_14034_, _14033_, _12545_);
  nand (_14035_, _08255_, \uc8051golden_1.ACC [5]);
  nor (_14036_, _08255_, \uc8051golden_1.ACC [5]);
  nor (_14037_, _08344_, \uc8051golden_1.ACC [4]);
  or (_14038_, _14037_, _14036_);
  and (_14039_, _14038_, _14035_);
  and (_14040_, _14039_, _12544_);
  nor (_14041_, _08072_, \uc8051golden_1.ACC [7]);
  or (_14042_, _08161_, \uc8051golden_1.ACC [6]);
  nor (_14043_, _14042_, _09034_);
  or (_14044_, _14043_, _14041_);
  or (_14045_, _14044_, _14040_);
  or (_14046_, _14045_, _14034_);
  nor (_14047_, _12546_, _06842_);
  and (_14048_, _14047_, _14046_);
  and (_14049_, _08762_, _07988_);
  or (_14050_, _14049_, _13993_);
  or (_14051_, _14050_, _07210_);
  and (_14052_, _07988_, \uc8051golden_1.ACC [7]);
  or (_14053_, _14052_, _13993_);
  and (_14054_, _14053_, _07199_);
  nor (_14055_, _07199_, _10524_);
  or (_14056_, _14055_, _06401_);
  or (_14057_, _14056_, _14054_);
  and (_14058_, _14057_, _10678_);
  and (_14059_, _14058_, _14051_);
  nor (_14060_, _10699_, _10678_);
  not (_14061_, _12457_);
  nand (_14062_, _14061_, _06407_);
  or (_14063_, _14062_, _14060_);
  or (_14064_, _14063_, _14059_);
  or (_14065_, _14019_, _06396_);
  or (_14066_, _14005_, _07221_);
  and (_14067_, _14066_, _14065_);
  and (_14068_, _14067_, _14064_);
  or (_14069_, _14068_, _06406_);
  or (_14070_, _14053_, _06414_);
  nor (_14071_, _12516_, _06393_);
  and (_14072_, _14071_, _14070_);
  and (_14073_, _14072_, _14069_);
  and (_14074_, _13991_, _06393_);
  or (_14075_, _14074_, _12450_);
  or (_14076_, _14075_, _14073_);
  not (_14077_, _12444_);
  or (_14078_, _12416_, _12413_);
  and (_14079_, _14078_, _08071_);
  or (_14080_, _12423_, _12419_);
  and (_14081_, _12421_, _14080_);
  and (_14082_, _14081_, _12418_);
  or (_14083_, _14082_, _14079_);
  or (_14084_, _12440_, _12438_);
  and (_14085_, _14084_, _12435_);
  and (_14086_, _12433_, _12430_);
  or (_14087_, _14086_, _12428_);
  or (_14088_, _14087_, _14085_);
  and (_14089_, _14088_, _12427_);
  or (_14090_, _14089_, _14083_);
  and (_14091_, _14090_, _14077_);
  or (_14092_, _14091_, _12449_);
  and (_14093_, _14092_, _12411_);
  and (_14094_, _14093_, _14076_);
  not (_14095_, _12400_);
  or (_14096_, _12402_, _14095_);
  and (_14097_, _14096_, _12396_);
  not (_14098_, _12393_);
  nand (_14099_, _12391_, _14098_);
  nand (_14100_, _14099_, _12390_);
  or (_14101_, _14100_, _14097_);
  and (_14102_, _14101_, _12389_);
  nor (_14103_, _12378_, _08788_);
  or (_14104_, _14103_, _12376_);
  nand (_14105_, _12386_, _12383_);
  and (_14106_, _12381_, _14105_);
  and (_14107_, _14106_, _12382_);
  or (_14108_, _14107_, _14104_);
  or (_14109_, _14108_, _14102_);
  and (_14110_, _12407_, _06457_);
  and (_14111_, _14110_, _14109_);
  or (_14112_, _14111_, _14094_);
  and (_14113_, _14112_, _06842_);
  or (_14114_, _14113_, _14048_);
  and (_14115_, _14114_, _12534_);
  nor (_14116_, _06228_, \uc8051golden_1.ACC [1]);
  and (_14117_, _06228_, \uc8051golden_1.ACC [1]);
  and (_14118_, _06840_, \uc8051golden_1.ACC [0]);
  nor (_14119_, _14118_, _14117_);
  or (_14120_, _14119_, _14116_);
  and (_14121_, _14120_, _12240_);
  nand (_14122_, _06372_, \uc8051golden_1.ACC [3]);
  nor (_14123_, _06372_, \uc8051golden_1.ACC [3]);
  nor (_14124_, _06693_, \uc8051golden_1.ACC [2]);
  or (_14125_, _14124_, _14123_);
  and (_14126_, _14125_, _14122_);
  or (_14127_, _14126_, _14121_);
  and (_14128_, _14127_, _12248_);
  nand (_14129_, _06650_, \uc8051golden_1.ACC [5]);
  nor (_14130_, _06650_, \uc8051golden_1.ACC [5]);
  nor (_14131_, _06265_, \uc8051golden_1.ACC [4]);
  or (_14132_, _14131_, _14130_);
  and (_14133_, _14132_, _14129_);
  and (_14134_, _14133_, _12247_);
  and (_14135_, _06194_, _08651_);
  or (_14136_, _06340_, \uc8051golden_1.ACC [6]);
  nor (_14137_, _14136_, _10970_);
  or (_14138_, _14137_, _14135_);
  or (_14139_, _14138_, _14134_);
  or (_14140_, _14139_, _14128_);
  nor (_14141_, _12249_, _12534_);
  and (_14142_, _14141_, _14140_);
  or (_14143_, _14142_, _12237_);
  or (_14144_, _14143_, _14115_);
  nand (_14145_, _12237_, \uc8051golden_1.PSW [7]);
  and (_14146_, _14145_, _07245_);
  and (_14147_, _14146_, _14144_);
  or (_14148_, _14147_, _14022_);
  and (_14149_, _14148_, _12563_);
  and (_14150_, _06388_, \uc8051golden_1.PSW [7]);
  and (_14151_, _14150_, _12958_);
  or (_14152_, _14151_, _14149_);
  nor (_14153_, _09538_, _06433_);
  and (_14154_, _14153_, _14152_);
  or (_14155_, _14154_, _14017_);
  and (_14156_, _14155_, _14015_);
  not (_14157_, _10740_);
  or (_14158_, _12958_, \uc8051golden_1.PSW [7]);
  and (_14159_, _14158_, _06432_);
  or (_14160_, _14159_, _14157_);
  or (_14161_, _14160_, _14156_);
  and (_14162_, _10754_, _10749_);
  nor (_14163_, _14162_, _10747_);
  nand (_14164_, _10803_, _10749_);
  or (_14165_, _14164_, _10801_);
  and (_14166_, _14165_, _14163_);
  or (_14167_, _10744_, _10740_);
  or (_14168_, _14167_, _14166_);
  and (_14169_, _14168_, _14161_);
  or (_14170_, _14169_, _12586_);
  and (_14171_, _10484_, _10479_);
  nor (_14172_, _14171_, _10477_);
  nand (_14173_, _10486_, _10479_);
  or (_14174_, _14173_, _10828_);
  and (_14175_, _14174_, _14172_);
  and (_14176_, _10480_, _09440_);
  and (_14177_, _14176_, _08749_);
  or (_14178_, _12587_, _14177_);
  or (_14179_, _14178_, _14175_);
  and (_14180_, _14179_, _06442_);
  and (_14181_, _14180_, _14170_);
  or (_14182_, _14181_, _14014_);
  and (_14183_, _14182_, _10573_);
  and (_14184_, _10842_, _07991_);
  and (_14185_, _10854_, _10850_);
  nor (_14186_, _14185_, _10848_);
  nand (_14187_, _10898_, _10850_);
  or (_14188_, _14187_, _10896_);
  and (_14189_, _14188_, _14186_);
  or (_14190_, _14189_, _14184_);
  and (_14191_, _14190_, _10572_);
  or (_14192_, _14191_, _10059_);
  or (_14193_, _14192_, _14183_);
  and (_14194_, _14193_, _14006_);
  or (_14195_, _14194_, _06281_);
  and (_14196_, _07988_, _08749_);
  or (_14197_, _13993_, _06282_);
  or (_14198_, _14197_, _14196_);
  and (_14199_, _14198_, _06279_);
  and (_14200_, _14199_, _14195_);
  or (_14201_, _14200_, _14003_);
  nor (_14202_, _10072_, _06376_);
  and (_14203_, _14202_, _14201_);
  nor (_14204_, _12958_, _10524_);
  and (_14205_, _14204_, _06376_);
  or (_14206_, _14205_, _06275_);
  or (_14207_, _14206_, _14203_);
  and (_14208_, _08813_, _07988_);
  or (_14209_, _14208_, _13993_);
  or (_14210_, _14209_, _06276_);
  and (_14211_, _14210_, _14207_);
  or (_14212_, _14211_, _06375_);
  nand (_14213_, _12958_, _10524_);
  or (_14214_, _14213_, _06952_);
  and (_14215_, _14214_, _14212_);
  or (_14216_, _14215_, _06474_);
  and (_14217_, _09027_, _07988_);
  or (_14218_, _14217_, _13993_);
  or (_14219_, _14218_, _07282_);
  and (_14220_, _14219_, _07284_);
  and (_14221_, _14220_, _14216_);
  or (_14222_, _14221_, _14000_);
  and (_14223_, _14222_, _07279_);
  or (_14224_, _13993_, _08073_);
  and (_14225_, _14209_, _06478_);
  and (_14226_, _14225_, _14224_);
  or (_14227_, _14226_, _14223_);
  and (_14228_, _14227_, _07276_);
  and (_14229_, _14053_, _06569_);
  and (_14230_, _14229_, _14224_);
  or (_14231_, _14230_, _06479_);
  or (_14232_, _14231_, _14228_);
  and (_14233_, _09026_, _07988_);
  or (_14234_, _13993_, _09043_);
  or (_14235_, _14234_, _14233_);
  and (_14236_, _14235_, _09048_);
  and (_14237_, _14236_, _14232_);
  or (_14238_, _14237_, _13997_);
  and (_14239_, _14238_, _11028_);
  nor (_14240_, _10746_, _08651_);
  or (_14241_, _14240_, _11052_);
  or (_14242_, _14241_, _10744_);
  and (_14243_, _14242_, _11030_);
  or (_14244_, _14243_, _10471_);
  or (_14245_, _14244_, _14239_);
  nor (_14246_, _10476_, _08651_);
  or (_14247_, _14246_, _10540_);
  or (_14248_, _14177_, _10472_);
  or (_14249_, _14248_, _14247_);
  and (_14250_, _14249_, _06579_);
  and (_14251_, _14250_, _14245_);
  nor (_14252_, _10583_, _08651_);
  or (_14253_, _14252_, _11083_);
  or (_14254_, _14253_, _14007_);
  and (_14255_, _14254_, _06578_);
  or (_14256_, _14255_, _14251_);
  or (_14257_, _14256_, _11059_);
  and (_14258_, _10847_, \uc8051golden_1.ACC [7]);
  or (_14259_, _14258_, _11113_);
  or (_14260_, _11091_, _14184_);
  or (_14261_, _14260_, _14259_);
  and (_14262_, _14261_, _11090_);
  and (_14263_, _14262_, _14257_);
  and (_14264_, _11089_, \uc8051golden_1.ACC [7]);
  or (_14265_, _14264_, _11121_);
  or (_14266_, _14265_, _14263_);
  not (_14267_, _10563_);
  nor (_14268_, _11156_, _14267_);
  nor (_14269_, _11124_, _10562_);
  nor (_14270_, _14269_, _10549_);
  or (_14271_, _14270_, _11120_);
  or (_14272_, _14271_, _14268_);
  and (_14273_, _14272_, _14266_);
  or (_14274_, _14273_, _11163_);
  not (_14275_, _10558_);
  nor (_14276_, _11198_, _10957_);
  nor (_14277_, _14276_, _11165_);
  nand (_14278_, _14277_, _14275_);
  and (_14279_, _14278_, _06308_);
  and (_14280_, _14279_, _14274_);
  not (_14281_, _09033_);
  not (_14282_, _09032_);
  nand (_14283_, _11238_, _14282_);
  and (_14284_, _14283_, _06307_);
  and (_14285_, _14284_, _14281_);
  or (_14286_, _14285_, _11203_);
  or (_14287_, _14286_, _14280_);
  not (_14288_, _10969_);
  not (_14289_, _11203_);
  nor (_14290_, _11274_, _10968_);
  nor (_14291_, _14290_, _14289_);
  nand (_14292_, _14291_, _14288_);
  and (_14293_, _14292_, _14287_);
  or (_14294_, _14293_, _06606_);
  nor (_14295_, _14050_, _07037_);
  nor (_14296_, _14295_, _11290_);
  and (_14297_, _14296_, _14294_);
  and (_14298_, _11290_, \uc8051golden_1.ACC [0]);
  or (_14299_, _14298_, _06234_);
  or (_14300_, _14299_, _14297_);
  and (_14301_, _14300_, _13992_);
  or (_14302_, _14301_, _06195_);
  and (_14303_, _08530_, _07988_);
  or (_14304_, _13993_, _06196_);
  or (_14305_, _14304_, _14303_);
  and (_14306_, _14305_, _01375_);
  and (_14307_, _14306_, _14302_);
  or (_14308_, _14307_, _13988_);
  and (_40347_, _14308_, _42545_);
  nor (_14309_, _07565_, _07417_);
  nor (_14310_, _07906_, _07416_);
  nor (_14311_, _14310_, _07713_);
  and (_14312_, _14311_, _07415_);
  and (_14313_, _14312_, _14309_);
  or (_14314_, _14313_, \uc8051golden_1.IRAM[0] [0]);
  not (_14315_, _14313_);
  or (_14316_, _07485_, _07320_);
  and (_14317_, _14316_, _13012_);
  and (_14318_, _05969_, \uc8051golden_1.PC [0]);
  not (_14319_, _09049_);
  or (_14320_, _08521_, _08817_);
  and (_14321_, _14320_, _09044_);
  and (_14322_, _08521_, _08817_);
  not (_14323_, _14322_);
  and (_14324_, _14323_, _14320_);
  and (_14325_, _14324_, _07283_);
  or (_14326_, _08521_, _07785_);
  nor (_14327_, _12879_, _12856_);
  or (_14328_, _14327_, _08638_);
  or (_14329_, _08644_, _07485_);
  nand (_14330_, _06790_, _05685_);
  or (_14331_, _06790_, \uc8051golden_1.ACC [0]);
  and (_14332_, _14331_, _14330_);
  nor (_14333_, _14332_, _08643_);
  nor (_14334_, _14333_, _07211_);
  and (_14335_, _14334_, _14329_);
  nor (_14336_, _08521_, _08753_);
  or (_14337_, _14336_, _14335_);
  and (_14338_, _14337_, _08641_);
  nand (_14339_, _12879_, _12857_);
  and (_14340_, _14339_, _07218_);
  or (_14341_, _14340_, _07351_);
  or (_14342_, _14341_, _14338_);
  nor (_14343_, _05997_, \uc8051golden_1.PC [0]);
  nor (_14344_, _14343_, _07222_);
  and (_14345_, _14344_, _14342_);
  and (_14346_, _07473_, _07222_);
  or (_14347_, _14346_, _07239_);
  or (_14348_, _14347_, _14345_);
  and (_14349_, _14348_, _14328_);
  or (_14350_, _14349_, _06419_);
  and (_14351_, _14350_, _14326_);
  or (_14352_, _14351_, _07246_);
  not (_14353_, _12880_);
  and (_14354_, _14339_, _14353_);
  or (_14355_, _14354_, _07423_);
  and (_14356_, _14355_, _05994_);
  and (_14357_, _14356_, _14352_);
  or (_14358_, _05994_, _05685_);
  nand (_14359_, _06383_, _14358_);
  or (_14360_, _14359_, _14357_);
  or (_14361_, _08521_, _06383_);
  and (_14362_, _14361_, _14360_);
  or (_14363_, _14362_, _07257_);
  or (_14364_, _09390_, _06194_);
  and (_14365_, _08520_, _07257_);
  nand (_14366_, _14365_, _14364_);
  and (_14367_, _14366_, _07777_);
  and (_14368_, _14367_, _14363_);
  and (_14369_, _07924_, \uc8051golden_1.PSW [7]);
  and (_14370_, _14369_, _06693_);
  or (_14371_, _14370_, _14327_);
  and (_14372_, _14371_, _07256_);
  or (_14373_, _14372_, _06017_);
  or (_14374_, _14373_, _14368_);
  and (_14375_, _06017_, _05685_);
  nor (_14376_, _14375_, _08798_);
  and (_14377_, _14376_, _14374_);
  and (_14378_, _08798_, _07473_);
  or (_14379_, _14378_, _08802_);
  or (_14380_, _14379_, _14377_);
  or (_14381_, _08809_, _09446_);
  and (_14382_, _14381_, _08808_);
  and (_14383_, _14382_, _14380_);
  and (_14384_, _08590_, _07473_);
  and (_14385_, _08973_, \uc8051golden_1.P0 [0]);
  and (_14386_, _08975_, \uc8051golden_1.ACC [0]);
  or (_14387_, _14386_, _14385_);
  and (_14388_, _08950_, \uc8051golden_1.P1 [0]);
  and (_14389_, _08920_, \uc8051golden_1.SBUF [0]);
  or (_14390_, _14389_, _14388_);
  or (_14391_, _14390_, _14387_);
  and (_14392_, _08934_, \uc8051golden_1.TCON [0]);
  and (_14393_, _08947_, \uc8051golden_1.SCON [0]);
  or (_14394_, _14393_, _14392_);
  and (_14395_, _08944_, \uc8051golden_1.TMOD [0]);
  and (_14396_, _08928_, \uc8051golden_1.PSW [0]);
  or (_14397_, _14396_, _14395_);
  or (_14398_, _14397_, _14394_);
  and (_14399_, _08961_, \uc8051golden_1.P2 [0]);
  and (_14400_, _08967_, \uc8051golden_1.IE [0]);
  or (_14401_, _14400_, _14399_);
  and (_14402_, _08969_, \uc8051golden_1.P3 [0]);
  and (_14403_, _08964_, \uc8051golden_1.IP [0]);
  or (_14404_, _14403_, _14402_);
  or (_14405_, _14404_, _14401_);
  and (_14406_, _08940_, \uc8051golden_1.TL0 [0]);
  and (_14407_, _08953_, \uc8051golden_1.B [0]);
  or (_14408_, _14407_, _14406_);
  or (_14409_, _14408_, _14405_);
  or (_14410_, _14409_, _14398_);
  or (_14411_, _14410_, _14391_);
  and (_14412_, _09001_, \uc8051golden_1.DPL [0]);
  and (_14413_, _09003_, \uc8051golden_1.TH0 [0]);
  and (_14414_, _08998_, \uc8051golden_1.DPH [0]);
  or (_14415_, _14414_, _14413_);
  or (_14416_, _14415_, _14412_);
  and (_14417_, _08996_, \uc8051golden_1.PCON [0]);
  and (_14418_, _08987_, \uc8051golden_1.TL1 [0]);
  or (_14419_, _14418_, _14417_);
  and (_14420_, _08983_, \uc8051golden_1.TH1 [0]);
  and (_14421_, _08990_, \uc8051golden_1.SP [0]);
  or (_14422_, _14421_, _14420_);
  or (_14423_, _14422_, _14419_);
  or (_14424_, _14423_, _14416_);
  or (_14425_, _14424_, _14411_);
  or (_14426_, _14425_, _14384_);
  and (_14427_, _14426_, _08807_);
  or (_14428_, _14427_, _09013_);
  or (_14429_, _14428_, _14383_);
  and (_14430_, _09013_, _06840_);
  nor (_14431_, _14430_, _06277_);
  and (_14432_, _14431_, _14429_);
  and (_14433_, _08817_, _06277_);
  or (_14434_, _14433_, _05943_);
  or (_14435_, _14434_, _14432_);
  and (_14436_, _05943_, _05685_);
  nor (_14437_, _14436_, _07283_);
  and (_14438_, _14437_, _14435_);
  or (_14439_, _14438_, _14325_);
  and (_14440_, _14439_, _09031_);
  nor (_14441_, _12539_, _09031_);
  or (_14442_, _14441_, _14440_);
  and (_14443_, _14442_, _07281_);
  and (_14444_, _14322_, _07280_);
  or (_14445_, _14444_, _14443_);
  and (_14446_, _14445_, _07278_);
  and (_14447_, _11225_, _07277_);
  or (_14448_, _14447_, _05956_);
  or (_14449_, _14448_, _14446_);
  and (_14450_, _05956_, _05685_);
  nor (_14451_, _14450_, _09044_);
  and (_14452_, _14451_, _14449_);
  or (_14453_, _14452_, _14321_);
  and (_14454_, _14453_, _14319_);
  nor (_14455_, _12538_, _14319_);
  or (_14456_, _14455_, _05966_);
  or (_14457_, _14456_, _14454_);
  nand (_14458_, _05966_, _05685_);
  and (_14459_, _14458_, _08546_);
  and (_14460_, _14459_, _14457_);
  not (_14461_, _08546_);
  and (_14462_, _14461_, _07485_);
  or (_14463_, _14462_, _14460_);
  and (_14464_, _14463_, _09074_);
  and (_14465_, _09390_, _07305_);
  or (_14466_, _14465_, _07304_);
  or (_14467_, _14466_, _14464_);
  nand (_14468_, _08521_, _07304_);
  and (_14469_, _14468_, _07312_);
  and (_14470_, _14469_, _14467_);
  and (_14471_, _06465_, _05685_);
  or (_14472_, _14471_, _14470_);
  or (_14473_, _14472_, _14318_);
  or (_14474_, _14473_, _07311_);
  not (_14475_, _13010_);
  or (_14476_, _14327_, _07418_);
  and (_14477_, _14476_, _14475_);
  and (_14478_, _14477_, _14474_);
  or (_14479_, _14478_, _14317_);
  or (_14480_, _09390_, _09439_);
  and (_14481_, _14480_, _14479_);
  or (_14482_, _14481_, _06197_);
  nand (_14483_, _08521_, _06197_);
  and (_14484_, _14483_, _07415_);
  and (_14485_, _14484_, _14482_);
  or (_14486_, _14485_, _14315_);
  and (_14487_, _14486_, _14314_);
  and (_14488_, _07918_, _07912_);
  nor (_14489_, _07919_, _14488_);
  and (_14490_, _14489_, _07918_);
  nand (_14491_, _14490_, _06271_);
  and (_14492_, _14491_, _14487_);
  nor (_14493_, _08664_, _07781_);
  not (_14494_, _14493_);
  and (_14495_, _14494_, _07918_);
  and (_14496_, _14495_, _06271_);
  not (_14497_, _12188_);
  nor (_14498_, _14497_, _06465_);
  and (_14499_, _12341_, _06465_);
  or (_14500_, _14499_, _14498_);
  and (_14501_, _14500_, _14496_);
  or (_40361_, _14501_, _14492_);
  nor (_14502_, _09423_, _08551_);
  nand (_14503_, _14502_, _06783_);
  nand (_14504_, _08476_, _07090_);
  nor (_14505_, _08476_, _07090_);
  not (_14506_, _14505_);
  and (_14507_, _14506_, _14504_);
  and (_14508_, _14507_, _07283_);
  nand (_14509_, _08798_, _07196_);
  or (_14510_, _09345_, _06194_);
  nand (_14511_, _14510_, _08475_);
  and (_14512_, _14511_, _07257_);
  not (_14513_, _12827_);
  nand (_14514_, _12826_, _12804_);
  and (_14515_, _14514_, _07246_);
  and (_14516_, _14515_, _14513_);
  nor (_14517_, _12826_, _08235_);
  or (_14518_, _14517_, _08638_);
  nand (_14519_, _14502_, _08643_);
  or (_14520_, _06462_, _07103_);
  and (_14521_, _14520_, _06394_);
  and (_14522_, _06790_, _05653_);
  and (_14523_, _07378_, _06394_);
  or (_14524_, _07633_, _14523_);
  nor (_14525_, _06790_, _05984_);
  or (_14526_, _14525_, _14524_);
  or (_14527_, _14526_, _14522_);
  or (_14528_, _14527_, _14521_);
  and (_14529_, _14528_, _14519_);
  and (_14530_, _14529_, _08753_);
  not (_14531_, _08522_);
  and (_14532_, _14531_, _08755_);
  nor (_14533_, _14532_, _08753_);
  or (_14534_, _14533_, _14530_);
  or (_14535_, _14534_, _07218_);
  or (_14536_, _14514_, _08641_);
  and (_14537_, _14536_, _14535_);
  or (_14538_, _14537_, _07351_);
  nor (_14539_, _05997_, _05653_);
  nor (_14540_, _14539_, _07222_);
  and (_14541_, _14540_, _14538_);
  and (_14542_, _07222_, _10782_);
  or (_14543_, _14542_, _07239_);
  or (_14544_, _14543_, _14541_);
  and (_14545_, _14544_, _14518_);
  or (_14546_, _14545_, _06419_);
  nand (_14547_, _08476_, _06419_);
  and (_14548_, _14547_, _07423_);
  and (_14549_, _14548_, _14546_);
  or (_14550_, _14549_, _14516_);
  and (_14551_, _14550_, _05994_);
  or (_14552_, _05994_, \uc8051golden_1.PC [1]);
  nand (_14553_, _06383_, _14552_);
  or (_14554_, _14553_, _14551_);
  nand (_14555_, _08476_, _06384_);
  and (_14556_, _14555_, _08669_);
  and (_14557_, _14556_, _14554_);
  or (_14558_, _14557_, _14512_);
  and (_14559_, _14558_, _07777_);
  nand (_14560_, _08235_, _10524_);
  and (_14561_, _14560_, _07256_);
  and (_14562_, _14561_, _14514_);
  or (_14563_, _14562_, _14559_);
  and (_14564_, _14563_, _07846_);
  and (_14565_, _06017_, _05653_);
  or (_14566_, _08798_, _14565_);
  or (_14567_, _14566_, _14564_);
  and (_14568_, _14567_, _14509_);
  or (_14569_, _14568_, _08802_);
  or (_14570_, _08809_, _09445_);
  and (_14571_, _14570_, _08808_);
  and (_14572_, _14571_, _14569_);
  nor (_14573_, _08813_, _07196_);
  and (_14574_, _08934_, \uc8051golden_1.TCON [1]);
  and (_14575_, _08920_, \uc8051golden_1.SBUF [1]);
  or (_14576_, _14575_, _14574_);
  and (_14577_, _08973_, \uc8051golden_1.P0 [1]);
  and (_14578_, _08947_, \uc8051golden_1.SCON [1]);
  or (_14579_, _14578_, _14577_);
  or (_14580_, _14579_, _14576_);
  and (_14581_, _08940_, \uc8051golden_1.TL0 [1]);
  and (_14582_, _08953_, \uc8051golden_1.B [1]);
  or (_14583_, _14582_, _14581_);
  and (_14584_, _08950_, \uc8051golden_1.P1 [1]);
  and (_14585_, _08928_, \uc8051golden_1.PSW [1]);
  or (_14586_, _14585_, _14584_);
  or (_14587_, _14586_, _14583_);
  and (_14588_, _08961_, \uc8051golden_1.P2 [1]);
  and (_14589_, _08969_, \uc8051golden_1.P3 [1]);
  or (_14590_, _14589_, _14588_);
  and (_14591_, _08967_, \uc8051golden_1.IE [1]);
  and (_14592_, _08964_, \uc8051golden_1.IP [1]);
  or (_14593_, _14592_, _14591_);
  or (_14594_, _14593_, _14590_);
  and (_14595_, _08944_, \uc8051golden_1.TMOD [1]);
  and (_14596_, _08975_, \uc8051golden_1.ACC [1]);
  or (_14597_, _14596_, _14595_);
  or (_14598_, _14597_, _14594_);
  or (_14599_, _14598_, _14587_);
  or (_14600_, _14599_, _14580_);
  and (_14601_, _08983_, \uc8051golden_1.TH1 [1]);
  and (_14602_, _09001_, \uc8051golden_1.DPL [1]);
  and (_14603_, _08998_, \uc8051golden_1.DPH [1]);
  or (_14604_, _14603_, _14602_);
  or (_14605_, _14604_, _14601_);
  and (_14606_, _08996_, \uc8051golden_1.PCON [1]);
  and (_14607_, _08990_, \uc8051golden_1.SP [1]);
  or (_14608_, _14607_, _14606_);
  and (_14609_, _09003_, \uc8051golden_1.TH0 [1]);
  and (_14610_, _08987_, \uc8051golden_1.TL1 [1]);
  or (_14611_, _14610_, _14609_);
  or (_14612_, _14611_, _14608_);
  or (_14613_, _14612_, _14605_);
  or (_14614_, _14613_, _14600_);
  or (_14615_, _14614_, _14573_);
  and (_14616_, _14615_, _08807_);
  or (_14617_, _14616_, _09013_);
  or (_14618_, _14617_, _14572_);
  and (_14619_, _09013_, _06228_);
  nor (_14620_, _14619_, _06277_);
  and (_14621_, _14620_, _14618_);
  and (_14622_, _08937_, _06277_);
  or (_14623_, _14622_, _05943_);
  or (_14624_, _14623_, _14621_);
  and (_14625_, _05943_, \uc8051golden_1.PC [1]);
  nor (_14626_, _14625_, _07283_);
  and (_14627_, _14626_, _14624_);
  or (_14628_, _14627_, _14508_);
  and (_14629_, _14628_, _09031_);
  and (_14630_, _11224_, _07285_);
  or (_14631_, _14630_, _14629_);
  and (_14632_, _14631_, _07281_);
  and (_14633_, _14505_, _07280_);
  or (_14634_, _14633_, _14632_);
  and (_14635_, _14634_, _07278_);
  and (_14636_, _11222_, _07277_);
  or (_14637_, _14636_, _05956_);
  or (_14638_, _14637_, _14635_);
  and (_14639_, _05956_, \uc8051golden_1.PC [1]);
  nor (_14640_, _14639_, _09044_);
  and (_14641_, _14640_, _14638_);
  and (_14642_, _14504_, _09044_);
  or (_14643_, _14642_, _09049_);
  or (_14644_, _14643_, _14641_);
  nand (_14645_, _11223_, _09049_);
  and (_14646_, _14645_, _05967_);
  and (_14647_, _14646_, _14644_);
  and (_14648_, _05966_, _05653_);
  or (_14649_, _06783_, _14648_);
  or (_14650_, _14649_, _14647_);
  and (_14651_, _14650_, _14503_);
  or (_14652_, _14651_, _06772_);
  and (_14653_, _06289_, _05968_);
  not (_14654_, _14653_);
  nand (_14655_, _14502_, _06772_);
  and (_14656_, _14655_, _14654_);
  and (_14657_, _14656_, _14652_);
  nor (_14658_, _14502_, _14654_);
  or (_14659_, _14658_, _09069_);
  or (_14660_, _14659_, _14657_);
  nand (_14661_, _07305_, _05979_);
  nand (_14662_, _14502_, _07300_);
  and (_14663_, _14662_, _14661_);
  and (_14664_, _14663_, _14660_);
  not (_14665_, _07031_);
  nor (_14666_, _09391_, _09447_);
  nand (_14667_, _14666_, _14665_);
  and (_14668_, _14667_, _07305_);
  or (_14669_, _14668_, _14664_);
  nand (_14670_, _14666_, _07031_);
  and (_14671_, _14670_, _09073_);
  and (_14672_, _14671_, _14669_);
  nor (_14673_, _14532_, _09073_);
  or (_14674_, _14673_, _06465_);
  or (_14675_, _14674_, _14672_);
  nand (_14676_, _06465_, _06024_);
  and (_14677_, _14676_, _13005_);
  and (_14678_, _14677_, _14675_);
  and (_14679_, _05969_, _05653_);
  or (_14680_, _07311_, _14679_);
  or (_14681_, _14680_, _14678_);
  not (_14682_, _07379_);
  and (_14683_, _14682_, _07365_);
  or (_14684_, _14517_, _07418_);
  and (_14685_, _14684_, _14683_);
  and (_14686_, _14685_, _14681_);
  not (_14687_, _14683_);
  and (_14688_, _14502_, _14687_);
  or (_14689_, _14688_, _07048_);
  or (_14690_, _14689_, _14686_);
  not (_14691_, _07048_);
  or (_14692_, _14502_, _14691_);
  and (_14693_, _14692_, _09439_);
  and (_14694_, _14693_, _14690_);
  and (_14695_, _14666_, _07320_);
  or (_14696_, _14695_, _06197_);
  or (_14697_, _14696_, _14694_);
  or (_14698_, _14532_, _09438_);
  and (_14699_, _14698_, _07415_);
  and (_14700_, _14699_, _14697_);
  or (_14701_, _14700_, _14315_);
  or (_14702_, _14313_, \uc8051golden_1.IRAM[0] [1]);
  and (_14703_, _14702_, _14491_);
  and (_14704_, _14703_, _14701_);
  nor (_14705_, _07917_, _01379_);
  and (_14706_, _14705_, _42545_);
  nor (_14707_, _07917_, _06270_);
  and (_14708_, _14707_, _01375_);
  and (_14709_, _14708_, _42545_);
  nor (_14710_, _07917_, \uc8051golden_1.SP [1]);
  and (_14711_, _14710_, _01375_);
  and (_14712_, _14711_, _42545_);
  nor (_14713_, _14712_, _14709_);
  not (_14714_, _07912_);
  nor (_14715_, _07917_, _14714_);
  and (_14716_, _14715_, _01375_);
  and (_14717_, _14716_, _42545_);
  not (_14718_, _07915_);
  nor (_14719_, _07917_, _14718_);
  and (_14720_, _14719_, _01375_);
  and (_14721_, _14720_, _42545_);
  nor (_14722_, _14721_, _14717_);
  and (_14723_, _14722_, _14713_);
  and (_14724_, _14723_, _14706_);
  not (_14725_, _07917_);
  not (_14726_, _12136_);
  nor (_14727_, _14726_, _06465_);
  and (_14728_, _12281_, _06465_);
  or (_14729_, _14728_, _14727_);
  and (_14730_, _14729_, _14725_);
  and (_14731_, _14730_, _01375_);
  and (_14732_, _14731_, _42545_);
  and (_14733_, _14732_, _14724_);
  or (_40362_, _14733_, _14704_);
  nor (_14734_, _09423_, _09422_);
  nor (_14735_, _14734_, _09424_);
  and (_14736_, _14735_, _13010_);
  and (_14737_, _08551_, _07623_);
  nor (_14738_, _08551_, _07623_);
  or (_14739_, _14738_, _14737_);
  or (_14740_, _14739_, _08543_);
  nand (_14741_, _08432_, _06736_);
  nor (_14742_, _08432_, _06736_);
  not (_14743_, _14742_);
  and (_14744_, _14743_, _14741_);
  and (_14745_, _14744_, _07283_);
  or (_14746_, _09300_, _06194_);
  nand (_14747_, _14746_, _08431_);
  and (_14748_, _14747_, _07257_);
  nor (_14749_, _12802_, _07961_);
  or (_14750_, _14749_, _08638_);
  nand (_14751_, _12802_, _12780_);
  or (_14752_, _14751_, _08641_);
  nand (_14753_, _08755_, _08433_);
  nand (_14754_, _14753_, _08756_);
  and (_14755_, _14754_, _07211_);
  and (_14756_, _06790_, _06065_);
  nor (_14757_, _06790_, _10195_);
  or (_14758_, _14757_, _14756_);
  and (_14759_, _14758_, _08644_);
  and (_14760_, _14739_, _08643_);
  or (_14761_, _14760_, _14759_);
  and (_14762_, _14761_, _08753_);
  or (_14763_, _14762_, _07218_);
  or (_14764_, _14763_, _14755_);
  and (_14765_, _14764_, _14752_);
  or (_14766_, _14765_, _07351_);
  nor (_14767_, _06065_, _05997_);
  nor (_14768_, _14767_, _07222_);
  and (_14769_, _14768_, _14766_);
  and (_14770_, _09422_, _07222_);
  or (_14771_, _14770_, _07239_);
  or (_14772_, _14771_, _14769_);
  and (_14773_, _14772_, _14750_);
  or (_14774_, _14773_, _06419_);
  nand (_14775_, _08432_, _06419_);
  and (_14776_, _14775_, _07423_);
  and (_14777_, _14776_, _14774_);
  not (_14778_, _12803_);
  and (_14779_, _14751_, _14778_);
  and (_14780_, _14779_, _07246_);
  or (_14781_, _14780_, _14777_);
  and (_14782_, _14781_, _05994_);
  or (_14783_, _06500_, _05994_);
  nand (_14784_, _06383_, _14783_);
  or (_14785_, _14784_, _14782_);
  nand (_14786_, _08432_, _06384_);
  and (_14787_, _14786_, _08669_);
  and (_14788_, _14787_, _14785_);
  or (_14789_, _14788_, _14748_);
  and (_14790_, _14789_, _07777_);
  and (_14791_, _07960_, \uc8051golden_1.PSW [7]);
  and (_14792_, _14791_, _06693_);
  or (_14793_, _14792_, _14749_);
  and (_14794_, _14793_, _07256_);
  or (_14795_, _14794_, _06017_);
  or (_14796_, _14795_, _14790_);
  and (_14797_, _06500_, _06017_);
  nor (_14798_, _14797_, _08798_);
  and (_14799_, _14798_, _14796_);
  nor (_14800_, _08803_, _07623_);
  or (_14801_, _14800_, _08802_);
  or (_14802_, _14801_, _14799_);
  or (_14803_, _08809_, _09444_);
  and (_14804_, _14803_, _08808_);
  and (_14805_, _14804_, _14802_);
  nor (_14806_, _08813_, _07623_);
  and (_14807_, _08973_, \uc8051golden_1.P0 [2]);
  and (_14808_, _08975_, \uc8051golden_1.ACC [2]);
  or (_14809_, _14808_, _14807_);
  and (_14810_, _08920_, \uc8051golden_1.SBUF [2]);
  and (_14811_, _08953_, \uc8051golden_1.B [2]);
  or (_14812_, _14811_, _14810_);
  or (_14813_, _14812_, _14809_);
  and (_14814_, _08944_, \uc8051golden_1.TMOD [2]);
  and (_14815_, _08940_, \uc8051golden_1.TL0 [2]);
  or (_14816_, _14815_, _14814_);
  and (_14817_, _08950_, \uc8051golden_1.P1 [2]);
  and (_14818_, _08928_, \uc8051golden_1.PSW [2]);
  or (_14819_, _14818_, _14817_);
  or (_14820_, _14819_, _14816_);
  and (_14821_, _08967_, \uc8051golden_1.IE [2]);
  and (_14822_, _08969_, \uc8051golden_1.P3 [2]);
  or (_14823_, _14822_, _14821_);
  and (_14824_, _08961_, \uc8051golden_1.P2 [2]);
  and (_14825_, _08964_, \uc8051golden_1.IP [2]);
  or (_14826_, _14825_, _14824_);
  or (_14827_, _14826_, _14823_);
  and (_14828_, _08934_, \uc8051golden_1.TCON [2]);
  and (_14829_, _08947_, \uc8051golden_1.SCON [2]);
  or (_14830_, _14829_, _14828_);
  or (_14831_, _14830_, _14827_);
  or (_14832_, _14831_, _14820_);
  or (_14833_, _14832_, _14813_);
  and (_14834_, _08998_, \uc8051golden_1.DPH [2]);
  and (_14835_, _08996_, \uc8051golden_1.PCON [2]);
  and (_14836_, _09003_, \uc8051golden_1.TH0 [2]);
  or (_14837_, _14836_, _14835_);
  or (_14838_, _14837_, _14834_);
  and (_14839_, _09001_, \uc8051golden_1.DPL [2]);
  and (_14840_, _08987_, \uc8051golden_1.TL1 [2]);
  or (_14841_, _14840_, _14839_);
  and (_14842_, _08983_, \uc8051golden_1.TH1 [2]);
  and (_14843_, _08990_, \uc8051golden_1.SP [2]);
  or (_14844_, _14843_, _14842_);
  or (_14845_, _14844_, _14841_);
  or (_14846_, _14845_, _14838_);
  or (_14847_, _14846_, _14833_);
  or (_14848_, _14847_, _14806_);
  and (_14849_, _14848_, _08807_);
  or (_14850_, _14849_, _09013_);
  or (_14851_, _14850_, _14805_);
  and (_14852_, _09013_, _06693_);
  nor (_14853_, _14852_, _06277_);
  and (_14854_, _14853_, _14851_);
  and (_14855_, _08994_, _06277_);
  or (_14856_, _14855_, _05943_);
  or (_14857_, _14856_, _14854_);
  and (_14858_, _06500_, _05943_);
  nor (_14859_, _14858_, _07283_);
  and (_14860_, _14859_, _14857_);
  or (_14861_, _14860_, _14745_);
  and (_14862_, _14861_, _09031_);
  and (_14863_, _11221_, _07285_);
  or (_14864_, _14863_, _14862_);
  and (_14865_, _14864_, _07281_);
  and (_14866_, _14742_, _07280_);
  or (_14867_, _14866_, _14865_);
  and (_14868_, _14867_, _07278_);
  and (_14869_, _11219_, _07277_);
  or (_14870_, _14869_, _05956_);
  or (_14871_, _14870_, _14868_);
  and (_14872_, _06500_, _05956_);
  nor (_14873_, _14872_, _09044_);
  and (_14874_, _14873_, _14871_);
  and (_14875_, _14741_, _09044_);
  or (_14876_, _14875_, _09049_);
  or (_14877_, _14876_, _14874_);
  nand (_14878_, _11220_, _09049_);
  and (_14879_, _14878_, _05967_);
  and (_14880_, _14879_, _14877_);
  and (_14881_, _06065_, _05966_);
  or (_14882_, _08542_, _14881_);
  or (_14883_, _14882_, _14880_);
  nand (_14884_, _14883_, _14740_);
  nand (_14885_, _14884_, _08545_);
  or (_14886_, _14739_, _08545_);
  and (_14887_, _14886_, _14661_);
  and (_14888_, _14887_, _14885_);
  nor (_14889_, _09391_, _09300_);
  or (_14890_, _14889_, _09392_);
  or (_14891_, _14890_, _07031_);
  and (_14892_, _14891_, _07305_);
  or (_14893_, _14892_, _14888_);
  or (_14894_, _14890_, _14665_);
  and (_14895_, _14894_, _09073_);
  and (_14896_, _14895_, _14893_);
  and (_14897_, _14754_, _07304_);
  or (_14898_, _14897_, _06465_);
  or (_14899_, _14898_, _14896_);
  nand (_14900_, _12314_, _06465_);
  and (_14901_, _14900_, _13005_);
  and (_14902_, _14901_, _14899_);
  and (_14903_, _06065_, _05969_);
  or (_14904_, _07311_, _14903_);
  or (_14905_, _14904_, _14902_);
  or (_14906_, _14749_, _07418_);
  and (_14907_, _14906_, _14475_);
  and (_14908_, _14907_, _14905_);
  or (_14909_, _14908_, _14736_);
  and (_14910_, _14909_, _09439_);
  or (_14911_, _09447_, _09444_);
  nor (_14912_, _09448_, _09439_);
  and (_14913_, _14912_, _14911_);
  or (_14914_, _14913_, _06197_);
  or (_14915_, _14914_, _14910_);
  nor (_14916_, _08522_, _08433_);
  nor (_14917_, _14916_, _08523_);
  or (_14918_, _14917_, _09438_);
  and (_14919_, _14918_, _07415_);
  and (_14920_, _14919_, _14915_);
  or (_14921_, _14920_, _14315_);
  not (_14922_, _14496_);
  or (_14923_, _14313_, \uc8051golden_1.IRAM[0] [2]);
  and (_14924_, _14923_, _14922_);
  and (_14925_, _14924_, _14921_);
  and (_14926_, _12274_, _06465_);
  not (_14927_, _12124_);
  nor (_14928_, _14927_, _06465_);
  or (_14929_, _14928_, _14926_);
  and (_14930_, _14929_, _14496_);
  or (_40363_, _14930_, _14925_);
  nand (_14931_, _08388_, _06562_);
  nor (_14932_, _08388_, _06562_);
  not (_14933_, _14932_);
  and (_14934_, _14933_, _14931_);
  and (_14935_, _14934_, _07283_);
  nand (_14936_, _08798_, _07775_);
  nor (_14937_, _14737_, _07775_);
  or (_14938_, _14937_, _08552_);
  or (_14939_, _14938_, _08644_);
  and (_14940_, _06790_, _06124_);
  nor (_14941_, _06790_, _10246_);
  or (_14942_, _14941_, _08643_);
  or (_14943_, _14942_, _14940_);
  and (_14944_, _14943_, _14939_);
  and (_14945_, _14944_, _08753_);
  and (_14946_, _08756_, _08389_);
  or (_14947_, _14946_, _08757_);
  and (_14948_, _14947_, _07211_);
  or (_14949_, _14948_, _14945_);
  or (_14950_, _14949_, _07218_);
  nand (_14951_, _12929_, _12907_);
  or (_14952_, _14951_, _08641_);
  and (_14953_, _14952_, _14950_);
  or (_14954_, _14953_, _07351_);
  nor (_14955_, _06124_, _05997_);
  nor (_14956_, _14955_, _07222_);
  and (_14957_, _14956_, _14954_);
  and (_14958_, _09421_, _07222_);
  or (_14959_, _14958_, _07239_);
  or (_14960_, _14959_, _14957_);
  nor (_14961_, _12929_, _08248_);
  or (_14962_, _14961_, _08638_);
  and (_14963_, _14962_, _14960_);
  or (_14964_, _14963_, _06419_);
  nand (_14965_, _08388_, _06419_);
  and (_14966_, _14965_, _07423_);
  and (_14967_, _14966_, _14964_);
  not (_14968_, _12930_);
  and (_14969_, _14951_, _14968_);
  and (_14970_, _14969_, _07246_);
  or (_14971_, _14970_, _14967_);
  and (_14972_, _14971_, _05994_);
  or (_14973_, _06134_, _05994_);
  nand (_14974_, _06383_, _14973_);
  or (_14975_, _14974_, _14972_);
  nand (_14976_, _08388_, _06384_);
  and (_14977_, _14976_, _14975_);
  or (_14978_, _14977_, _07257_);
  and (_14979_, _09443_, _06309_);
  nand (_14980_, _08387_, _07257_);
  or (_14981_, _14980_, _14979_);
  and (_14982_, _14981_, _14978_);
  or (_14983_, _14982_, _07256_);
  and (_14984_, _08248_, \uc8051golden_1.PSW [7]);
  or (_14985_, _14961_, _14984_);
  or (_14986_, _14985_, _07777_);
  and (_14987_, _14986_, _07846_);
  and (_14988_, _14987_, _14983_);
  and (_14989_, _06124_, _06017_);
  or (_14990_, _08798_, _14989_);
  or (_14991_, _14990_, _14988_);
  and (_14992_, _14991_, _14936_);
  or (_14993_, _14992_, _08802_);
  or (_14994_, _08809_, _09443_);
  and (_14995_, _14994_, _08808_);
  and (_14996_, _14995_, _14993_);
  nor (_14997_, _08813_, _07775_);
  and (_14998_, _08944_, \uc8051golden_1.TMOD [3]);
  and (_14999_, _08950_, \uc8051golden_1.P1 [3]);
  or (_15000_, _14999_, _14998_);
  and (_15001_, _08973_, \uc8051golden_1.P0 [3]);
  and (_15002_, _08934_, \uc8051golden_1.TCON [3]);
  or (_15003_, _15002_, _15001_);
  or (_15004_, _15003_, _15000_);
  and (_15005_, _08975_, \uc8051golden_1.ACC [3]);
  and (_15006_, _08928_, \uc8051golden_1.PSW [3]);
  or (_15007_, _15006_, _15005_);
  and (_15008_, _08947_, \uc8051golden_1.SCON [3]);
  and (_15009_, _08920_, \uc8051golden_1.SBUF [3]);
  or (_15010_, _15009_, _15008_);
  or (_15011_, _15010_, _15007_);
  and (_15012_, _08969_, \uc8051golden_1.P3 [3]);
  and (_15013_, _08964_, \uc8051golden_1.IP [3]);
  or (_15014_, _15013_, _15012_);
  and (_15015_, _08961_, \uc8051golden_1.P2 [3]);
  and (_15016_, _08967_, \uc8051golden_1.IE [3]);
  or (_15017_, _15016_, _15015_);
  or (_15018_, _15017_, _15014_);
  and (_15019_, _08940_, \uc8051golden_1.TL0 [3]);
  and (_15020_, _08953_, \uc8051golden_1.B [3]);
  or (_15021_, _15020_, _15019_);
  or (_15022_, _15021_, _15018_);
  or (_15023_, _15022_, _15011_);
  or (_15024_, _15023_, _15004_);
  and (_15025_, _08983_, \uc8051golden_1.TH1 [3]);
  and (_15026_, _09001_, \uc8051golden_1.DPL [3]);
  and (_15027_, _08996_, \uc8051golden_1.PCON [3]);
  or (_15028_, _15027_, _15026_);
  or (_15029_, _15028_, _15025_);
  and (_15030_, _08987_, \uc8051golden_1.TL1 [3]);
  and (_15031_, _08998_, \uc8051golden_1.DPH [3]);
  or (_15032_, _15031_, _15030_);
  and (_15033_, _09003_, \uc8051golden_1.TH0 [3]);
  and (_15034_, _08990_, \uc8051golden_1.SP [3]);
  or (_15035_, _15034_, _15033_);
  or (_15036_, _15035_, _15032_);
  or (_15037_, _15036_, _15029_);
  or (_15038_, _15037_, _15024_);
  or (_15039_, _15038_, _14997_);
  and (_15040_, _15039_, _08807_);
  or (_15041_, _15040_, _09013_);
  or (_15042_, _15041_, _14996_);
  and (_15043_, _09013_, _06372_);
  nor (_15044_, _15043_, _06277_);
  and (_15045_, _15044_, _15042_);
  and (_15046_, _08815_, _06277_);
  or (_15047_, _15046_, _05943_);
  or (_15048_, _15047_, _15045_);
  and (_15049_, _06134_, _05943_);
  nor (_15050_, _15049_, _07283_);
  and (_15051_, _15050_, _15048_);
  or (_15052_, _15051_, _14935_);
  and (_15053_, _15052_, _09031_);
  and (_15054_, _12535_, _07285_);
  or (_15055_, _15054_, _15053_);
  and (_15056_, _15055_, _07281_);
  and (_15057_, _14932_, _07280_);
  or (_15058_, _15057_, _15056_);
  and (_15059_, _15058_, _07278_);
  and (_15060_, _11217_, _07277_);
  or (_15061_, _15060_, _05956_);
  or (_15062_, _15061_, _15059_);
  and (_15063_, _06134_, _05956_);
  nor (_15064_, _15063_, _09044_);
  and (_15065_, _15064_, _15062_);
  and (_15066_, _14931_, _09044_);
  or (_15067_, _15066_, _09049_);
  or (_15068_, _15067_, _15065_);
  nand (_15069_, _11218_, _09049_);
  and (_15070_, _15069_, _05967_);
  and (_15071_, _15070_, _15068_);
  and (_15072_, _06124_, _05966_);
  nor (_15073_, _07300_, _15072_);
  nand (_15074_, _15073_, _09061_);
  or (_15075_, _15074_, _15071_);
  or (_15076_, _14938_, _08546_);
  and (_15077_, _15076_, _14661_);
  and (_15078_, _15077_, _15075_);
  nor (_15079_, _09392_, _09255_);
  or (_15080_, _15079_, _09393_);
  or (_15081_, _15080_, _07031_);
  and (_15082_, _15081_, _07305_);
  or (_15083_, _15082_, _15078_);
  or (_15084_, _15080_, _14665_);
  and (_15085_, _15084_, _09073_);
  and (_15086_, _15085_, _15083_);
  and (_15087_, _14947_, _07304_);
  or (_15088_, _15087_, _06465_);
  or (_15089_, _15088_, _15086_);
  nand (_15090_, _12309_, _06465_);
  and (_15091_, _15090_, _13005_);
  and (_15092_, _15091_, _15089_);
  and (_15093_, _06124_, _05969_);
  or (_15094_, _07311_, _15093_);
  or (_15095_, _15094_, _15092_);
  or (_15096_, _14961_, _07418_);
  and (_15097_, _15096_, _14683_);
  and (_15098_, _15097_, _15095_);
  nor (_15099_, _09424_, _09421_);
  nor (_15100_, _15099_, _09425_);
  and (_15101_, _15100_, _14687_);
  or (_15102_, _15101_, _07048_);
  or (_15103_, _15102_, _15098_);
  or (_15104_, _15100_, _14691_);
  and (_15105_, _15104_, _09439_);
  and (_15106_, _15105_, _15103_);
  or (_15107_, _09448_, _09443_);
  nor (_15108_, _09449_, _09439_);
  and (_15109_, _15108_, _15107_);
  or (_15110_, _15109_, _06197_);
  or (_15111_, _15110_, _15106_);
  nor (_15112_, _08523_, _08389_);
  nor (_15113_, _15112_, _08524_);
  or (_15114_, _15113_, _09438_);
  and (_15115_, _15114_, _07415_);
  and (_15116_, _15115_, _15111_);
  or (_15117_, _15116_, _14315_);
  or (_15118_, _14313_, \uc8051golden_1.IRAM[0] [3]);
  and (_15119_, _15118_, _14922_);
  and (_15120_, _15119_, _15117_);
  and (_15121_, _12268_, _06465_);
  and (_15122_, _12128_, _09463_);
  or (_15123_, _15122_, _15121_);
  and (_15124_, _15123_, _14725_);
  and (_15125_, _15124_, _01375_);
  and (_15126_, _15125_, _42545_);
  and (_15127_, _15126_, _14724_);
  or (_40364_, _15127_, _15120_);
  and (_15128_, _08757_, _08344_);
  nor (_15129_, _08757_, _08344_);
  or (_15130_, _15129_, _15128_);
  or (_15131_, _15130_, _09073_);
  nor (_15132_, _08882_, _08344_);
  not (_15133_, _15132_);
  nand (_15134_, _08882_, _08344_);
  and (_15135_, _15134_, _15133_);
  and (_15136_, _15135_, _07283_);
  and (_15137_, _12156_, _06017_);
  not (_15138_, _12853_);
  nand (_15139_, _12852_, _12850_);
  and (_15140_, _15139_, _07246_);
  and (_15141_, _15140_, _15138_);
  or (_15142_, _15139_, _08641_);
  and (_15143_, _08552_, _08301_);
  nor (_15144_, _08552_, _08301_);
  or (_15145_, _15144_, _15143_);
  and (_15146_, _15145_, _08643_);
  nor (_15147_, _06790_, _10119_);
  and (_15148_, _12156_, _06790_);
  or (_15149_, _15148_, _15147_);
  and (_15150_, _15149_, _08644_);
  or (_15151_, _15150_, _07212_);
  or (_15152_, _15151_, _15146_);
  or (_15153_, _09442_, _08659_);
  and (_15154_, _15153_, _15152_);
  or (_15155_, _15154_, _07211_);
  or (_15157_, _15130_, _08753_);
  and (_15158_, _15157_, _15155_);
  or (_15159_, _15158_, _07218_);
  and (_15160_, _15159_, _15142_);
  or (_15161_, _15160_, _07351_);
  nor (_15162_, _12156_, _05997_);
  nor (_15163_, _15162_, _07222_);
  and (_15164_, _15163_, _15161_);
  and (_15165_, _09420_, _07222_);
  or (_15166_, _15165_, _07239_);
  or (_15167_, _15166_, _15164_);
  nor (_15168_, _12851_, _12850_);
  or (_15169_, _15168_, _08638_);
  and (_15170_, _15169_, _15167_);
  or (_15171_, _15170_, _06419_);
  nand (_15172_, _08344_, _06419_);
  and (_15173_, _15172_, _07423_);
  and (_15174_, _15173_, _15171_);
  or (_15175_, _15174_, _15141_);
  and (_15176_, _15175_, _05994_);
  or (_15177_, _12157_, _05994_);
  nand (_15178_, _15177_, _06383_);
  or (_15179_, _15178_, _15176_);
  nand (_15180_, _08344_, _06384_);
  and (_15181_, _15180_, _15179_);
  or (_15182_, _15181_, _07257_);
  and (_15183_, _09442_, _06309_);
  nand (_15184_, _08343_, _07257_);
  or (_15185_, _15184_, _15183_);
  and (_15186_, _15185_, _15182_);
  or (_15187_, _15186_, _07256_);
  and (_15188_, _14369_, _07573_);
  or (_15189_, _15188_, _15168_);
  or (_15190_, _15189_, _07777_);
  and (_15191_, _15190_, _07846_);
  and (_15192_, _15191_, _15187_);
  or (_15193_, _15192_, _15137_);
  and (_15194_, _15193_, _08803_);
  nor (_15195_, _08803_, _08301_);
  or (_15196_, _15195_, _08802_);
  or (_15197_, _15196_, _15194_);
  or (_15198_, _08809_, _09442_);
  and (_15199_, _15198_, _08808_);
  and (_15200_, _15199_, _15197_);
  nor (_15201_, _08813_, _08301_);
  and (_15202_, _08934_, \uc8051golden_1.TCON [4]);
  and (_15203_, _08947_, \uc8051golden_1.SCON [4]);
  or (_15204_, _15203_, _15202_);
  and (_15205_, _08944_, \uc8051golden_1.TMOD [4]);
  and (_15206_, _08950_, \uc8051golden_1.P1 [4]);
  or (_15207_, _15206_, _15205_);
  or (_15208_, _15207_, _15204_);
  and (_15209_, _08973_, \uc8051golden_1.P0 [4]);
  and (_15210_, _08928_, \uc8051golden_1.PSW [4]);
  or (_15211_, _15210_, _15209_);
  and (_15212_, _08920_, \uc8051golden_1.SBUF [4]);
  and (_15213_, _08953_, \uc8051golden_1.B [4]);
  or (_15214_, _15213_, _15212_);
  or (_15215_, _15214_, _15211_);
  and (_15216_, _08969_, \uc8051golden_1.P3 [4]);
  and (_15217_, _08964_, \uc8051golden_1.IP [4]);
  or (_15218_, _15217_, _15216_);
  and (_15219_, _08961_, \uc8051golden_1.P2 [4]);
  and (_15220_, _08967_, \uc8051golden_1.IE [4]);
  or (_15221_, _15220_, _15219_);
  or (_15222_, _15221_, _15218_);
  and (_15223_, _08940_, \uc8051golden_1.TL0 [4]);
  and (_15224_, _08975_, \uc8051golden_1.ACC [4]);
  or (_15225_, _15224_, _15223_);
  or (_15226_, _15225_, _15222_);
  or (_15227_, _15226_, _15215_);
  or (_15228_, _15227_, _15208_);
  and (_15229_, _08987_, \uc8051golden_1.TL1 [4]);
  and (_15230_, _09003_, \uc8051golden_1.TH0 [4]);
  and (_15231_, _08998_, \uc8051golden_1.DPH [4]);
  or (_15232_, _15231_, _15230_);
  or (_15233_, _15232_, _15229_);
  and (_15234_, _09001_, \uc8051golden_1.DPL [4]);
  and (_15235_, _08996_, \uc8051golden_1.PCON [4]);
  or (_15236_, _15235_, _15234_);
  and (_15237_, _08983_, \uc8051golden_1.TH1 [4]);
  and (_15238_, _08990_, \uc8051golden_1.SP [4]);
  or (_15239_, _15238_, _15237_);
  or (_15240_, _15239_, _15236_);
  or (_15241_, _15240_, _15233_);
  or (_15242_, _15241_, _15228_);
  or (_15243_, _15242_, _15201_);
  and (_15244_, _15243_, _08807_);
  or (_15245_, _15244_, _09013_);
  or (_15246_, _15245_, _15200_);
  and (_15247_, _09013_, _06265_);
  nor (_15248_, _15247_, _06277_);
  and (_15249_, _15248_, _15246_);
  and (_15250_, _08883_, _06277_);
  or (_15251_, _15250_, _05943_);
  or (_15252_, _15251_, _15249_);
  and (_15253_, _12157_, _05943_);
  nor (_15254_, _15253_, _07283_);
  and (_15255_, _15254_, _15252_);
  or (_15256_, _15255_, _15136_);
  and (_15257_, _15256_, _09031_);
  and (_15258_, _11216_, _07285_);
  or (_15259_, _15258_, _15257_);
  and (_15260_, _15259_, _07281_);
  and (_15261_, _15132_, _07280_);
  or (_15262_, _15261_, _15260_);
  and (_15263_, _15262_, _07278_);
  and (_15264_, _11213_, _07277_);
  or (_15265_, _15264_, _05956_);
  or (_15266_, _15265_, _15263_);
  and (_15267_, _12157_, _05956_);
  nor (_15268_, _15267_, _09044_);
  and (_15269_, _15268_, _15266_);
  and (_15270_, _15134_, _09044_);
  or (_15271_, _15270_, _09049_);
  or (_15272_, _15271_, _15269_);
  nand (_15273_, _11215_, _09049_);
  and (_15274_, _15273_, _05967_);
  and (_15275_, _15274_, _15272_);
  nand (_15276_, _12156_, _05966_);
  nand (_15277_, _15276_, _08546_);
  or (_15278_, _15277_, _15275_);
  or (_15279_, _15145_, _09061_);
  or (_15280_, _15145_, _08547_);
  and (_15281_, _15280_, _09074_);
  and (_15282_, _15281_, _15279_);
  and (_15283_, _15282_, _15278_);
  nor (_15284_, _09393_, _09210_);
  or (_15285_, _15284_, _09394_);
  and (_15286_, _15285_, _07305_);
  or (_15287_, _15286_, _07304_);
  or (_15288_, _15287_, _15283_);
  and (_15289_, _15288_, _15131_);
  or (_15290_, _15289_, _06465_);
  nand (_15291_, _12305_, _06465_);
  and (_15292_, _15291_, _13005_);
  and (_15293_, _15292_, _15290_);
  and (_15294_, _12156_, _05969_);
  or (_15295_, _15294_, _07311_);
  or (_15296_, _15295_, _15293_);
  or (_15297_, _15168_, _07418_);
  and (_15298_, _15297_, _14475_);
  and (_15299_, _15298_, _15296_);
  or (_15300_, _09425_, _09420_);
  nor (_15301_, _14475_, _09426_);
  and (_15302_, _15301_, _15300_);
  or (_15303_, _15302_, _07344_);
  or (_15304_, _15303_, _15299_);
  not (_15305_, _07344_);
  nor (_15306_, _09449_, _09442_);
  nor (_15307_, _15306_, _09450_);
  nor (_15308_, _15307_, _15305_);
  nor (_15309_, _15308_, _07045_);
  and (_15310_, _15309_, _15304_);
  and (_15311_, _15307_, _07045_);
  or (_15312_, _15311_, _06197_);
  or (_15313_, _15312_, _15310_);
  nor (_15314_, _08524_, _08345_);
  nor (_15315_, _15314_, _08525_);
  or (_15316_, _15315_, _09438_);
  and (_15317_, _15316_, _07415_);
  and (_15318_, _15317_, _15313_);
  or (_15319_, _15318_, _14315_);
  or (_15320_, _14313_, \uc8051golden_1.IRAM[0] [4]);
  and (_15321_, _15320_, _14922_);
  and (_15322_, _15321_, _15319_);
  not (_15323_, _12121_);
  nor (_15324_, _15323_, _06465_);
  and (_15325_, _12262_, _06465_);
  or (_15326_, _15325_, _15324_);
  and (_15327_, _15326_, _14725_);
  and (_15328_, _15327_, _01375_);
  and (_15329_, _15328_, _42545_);
  and (_15330_, _15329_, _14724_);
  or (_40366_, _15330_, _15322_);
  nor (_15331_, _09450_, _09441_);
  nor (_15332_, _15331_, _09451_);
  or (_15333_, _15332_, _09439_);
  and (_15334_, _12151_, _05966_);
  nand (_15335_, _08917_, _08255_);
  nor (_15336_, _08917_, _08255_);
  not (_15337_, _15336_);
  and (_15338_, _15337_, _15335_);
  and (_15339_, _15338_, _07283_);
  nand (_15340_, _08798_, _08207_);
  nand (_15341_, _12954_, _12952_);
  nand (_15342_, _12953_, _10524_);
  and (_15343_, _15342_, _07256_);
  and (_15344_, _15343_, _15341_);
  nor (_15345_, _12953_, _12952_);
  or (_15346_, _15345_, _08638_);
  nor (_15347_, _15128_, _08255_);
  or (_15348_, _15347_, _08758_);
  and (_15349_, _15348_, _07211_);
  or (_15350_, _09441_, _08659_);
  nor (_15351_, _15143_, _08207_);
  or (_15352_, _15351_, _08553_);
  and (_15353_, _15352_, _08643_);
  nand (_15354_, _12152_, _06790_);
  or (_15355_, _06790_, \uc8051golden_1.ACC [5]);
  and (_15356_, _15355_, _15354_);
  and (_15357_, _15356_, _08644_);
  or (_15358_, _15357_, _07212_);
  or (_15359_, _15358_, _15353_);
  and (_15360_, _15359_, _08753_);
  and (_15361_, _15360_, _15350_);
  or (_15362_, _15361_, _15349_);
  and (_15363_, _15362_, _08641_);
  and (_15364_, _15341_, _07218_);
  or (_15365_, _15364_, _07351_);
  or (_15366_, _15365_, _15363_);
  nor (_15367_, _12151_, _05997_);
  nor (_15368_, _15367_, _07222_);
  and (_15369_, _15368_, _15366_);
  and (_15370_, _09419_, _07222_);
  or (_15371_, _15370_, _07239_);
  or (_15372_, _15371_, _15369_);
  and (_15373_, _15372_, _15346_);
  or (_15374_, _15373_, _06419_);
  nand (_15375_, _08255_, _06419_);
  and (_15376_, _15375_, _07423_);
  and (_15377_, _15376_, _15374_);
  not (_15378_, _12955_);
  and (_15379_, _15341_, _07246_);
  and (_15380_, _15379_, _15378_);
  or (_15381_, _15380_, _15377_);
  and (_15382_, _15381_, _05994_);
  or (_15383_, _12152_, _05994_);
  nand (_15384_, _15383_, _06383_);
  or (_15385_, _15384_, _15382_);
  nand (_15386_, _08255_, _06384_);
  and (_15387_, _15386_, _15385_);
  or (_15388_, _15387_, _07257_);
  and (_15389_, _09441_, _06309_);
  nand (_15390_, _08254_, _07257_);
  or (_15391_, _15390_, _15389_);
  and (_15392_, _15391_, _07777_);
  and (_15393_, _15392_, _15388_);
  or (_15394_, _15393_, _15344_);
  and (_15395_, _15394_, _07846_);
  and (_15396_, _12151_, _06017_);
  or (_15397_, _15396_, _08798_);
  or (_15398_, _15397_, _15395_);
  and (_15399_, _15398_, _15340_);
  or (_15400_, _15399_, _08802_);
  or (_15401_, _08809_, _09441_);
  and (_15402_, _15401_, _08808_);
  and (_15403_, _15402_, _15400_);
  nor (_15404_, _08813_, _08207_);
  and (_15405_, _08973_, \uc8051golden_1.P0 [5]);
  and (_15406_, _08928_, \uc8051golden_1.PSW [5]);
  or (_15407_, _15406_, _15405_);
  and (_15408_, _08944_, \uc8051golden_1.TMOD [5]);
  and (_15409_, _08975_, \uc8051golden_1.ACC [5]);
  or (_15410_, _15409_, _15408_);
  or (_15411_, _15410_, _15407_);
  and (_15412_, _08934_, \uc8051golden_1.TCON [5]);
  and (_15413_, _08947_, \uc8051golden_1.SCON [5]);
  or (_15414_, _15413_, _15412_);
  and (_15415_, _08950_, \uc8051golden_1.P1 [5]);
  and (_15416_, _08953_, \uc8051golden_1.B [5]);
  or (_15417_, _15416_, _15415_);
  or (_15418_, _15417_, _15414_);
  and (_15419_, _08961_, \uc8051golden_1.P2 [5]);
  and (_15420_, _08967_, \uc8051golden_1.IE [5]);
  or (_15421_, _15420_, _15419_);
  and (_15422_, _08969_, \uc8051golden_1.P3 [5]);
  and (_15423_, _08964_, \uc8051golden_1.IP [5]);
  or (_15424_, _15423_, _15422_);
  or (_15425_, _15424_, _15421_);
  and (_15426_, _08940_, \uc8051golden_1.TL0 [5]);
  and (_15427_, _08920_, \uc8051golden_1.SBUF [5]);
  or (_15428_, _15427_, _15426_);
  or (_15429_, _15428_, _15425_);
  or (_15430_, _15429_, _15418_);
  or (_15431_, _15430_, _15411_);
  and (_15432_, _08987_, \uc8051golden_1.TL1 [5]);
  and (_15433_, _09001_, \uc8051golden_1.DPL [5]);
  and (_15434_, _08996_, \uc8051golden_1.PCON [5]);
  or (_15435_, _15434_, _15433_);
  or (_15436_, _15435_, _15432_);
  and (_15437_, _09003_, \uc8051golden_1.TH0 [5]);
  and (_15438_, _08983_, \uc8051golden_1.TH1 [5]);
  or (_15439_, _15438_, _15437_);
  and (_15440_, _08998_, \uc8051golden_1.DPH [5]);
  and (_15441_, _08990_, \uc8051golden_1.SP [5]);
  or (_15442_, _15441_, _15440_);
  or (_15443_, _15442_, _15439_);
  or (_15444_, _15443_, _15436_);
  or (_15445_, _15444_, _15431_);
  or (_15446_, _15445_, _15404_);
  and (_15447_, _15446_, _08807_);
  or (_15448_, _15447_, _09013_);
  or (_15449_, _15448_, _15403_);
  and (_15450_, _09013_, _06650_);
  nor (_15451_, _15450_, _06277_);
  and (_15452_, _15451_, _15449_);
  and (_15453_, _08958_, _06277_);
  or (_15454_, _15453_, _05943_);
  or (_15455_, _15454_, _15452_);
  and (_15456_, _12152_, _05943_);
  nor (_15457_, _15456_, _07283_);
  and (_15458_, _15457_, _15455_);
  or (_15459_, _15458_, _15339_);
  and (_15460_, _15459_, _09031_);
  and (_15461_, _12542_, _07285_);
  or (_15462_, _15461_, _15460_);
  and (_15463_, _15462_, _07281_);
  and (_15464_, _15336_, _07280_);
  or (_15465_, _15464_, _15463_);
  and (_15466_, _15465_, _07278_);
  and (_15467_, _11211_, _07277_);
  or (_15468_, _15467_, _05956_);
  or (_15469_, _15468_, _15466_);
  and (_15470_, _12152_, _05956_);
  nor (_15471_, _15470_, _09044_);
  and (_15472_, _15471_, _15469_);
  and (_15473_, _15335_, _09044_);
  or (_15474_, _15473_, _09049_);
  or (_15475_, _15474_, _15472_);
  nand (_15476_, _11212_, _09049_);
  and (_15477_, _15476_, _05967_);
  and (_15478_, _15477_, _15475_);
  or (_15479_, _15478_, _15334_);
  and (_15480_, _15479_, _08546_);
  and (_15481_, _15352_, _14461_);
  or (_15482_, _15481_, _15480_);
  and (_15483_, _15482_, _09074_);
  nor (_15484_, _09394_, _09165_);
  or (_15485_, _15484_, _09395_);
  and (_15486_, _15485_, _07305_);
  or (_15487_, _15486_, _15483_);
  and (_15488_, _15487_, _09073_);
  and (_15489_, _15348_, _07304_);
  or (_15490_, _15489_, _06465_);
  or (_15491_, _15490_, _15488_);
  nand (_15492_, _12300_, _06465_);
  and (_15493_, _15492_, _13005_);
  and (_15494_, _15493_, _15491_);
  and (_15495_, _12151_, _05969_);
  or (_15496_, _15495_, _07311_);
  or (_15497_, _15496_, _15494_);
  or (_15498_, _15345_, _07418_);
  and (_15499_, _15498_, _14475_);
  and (_15500_, _15499_, _15497_);
  nor (_15501_, _09426_, _09419_);
  or (_15502_, _15501_, _09427_);
  nor (_15503_, _15502_, _14475_);
  or (_15504_, _15503_, _07320_);
  or (_15505_, _15504_, _15500_);
  and (_15506_, _15505_, _15333_);
  or (_15507_, _15506_, _06197_);
  nor (_15508_, _08525_, _08256_);
  nor (_15509_, _15508_, _08526_);
  or (_15510_, _15509_, _09438_);
  and (_15511_, _15510_, _07415_);
  and (_15512_, _15511_, _15507_);
  or (_15513_, _15512_, _14315_);
  or (_15514_, _14313_, \uc8051golden_1.IRAM[0] [5]);
  and (_15515_, _15514_, _14922_);
  and (_15516_, _15515_, _15513_);
  and (_15517_, _12258_, _06465_);
  not (_15518_, _12117_);
  nor (_15519_, _15518_, _06465_);
  or (_15520_, _15519_, _15517_);
  and (_15521_, _15520_, _14725_);
  and (_15522_, _15521_, _01375_);
  and (_15523_, _15522_, _42545_);
  and (_15524_, _15523_, _14724_);
  or (_40367_, _15524_, _15516_);
  nor (_15525_, _09427_, _09418_);
  nor (_15526_, _15525_, _09428_);
  and (_15527_, _15526_, _09415_);
  nand (_15528_, _08850_, _08161_);
  nor (_15529_, _08850_, _08161_);
  not (_15530_, _15529_);
  and (_15531_, _15530_, _15528_);
  and (_15532_, _15531_, _07283_);
  and (_15533_, _12144_, _06017_);
  and (_15534_, _09418_, _07222_);
  nand (_15535_, _12904_, _12902_);
  or (_15536_, _15535_, _08641_);
  or (_15537_, _09440_, _08659_);
  nor (_15538_, _08553_, _08118_);
  or (_15539_, _15538_, _08554_);
  and (_15540_, _15539_, _08643_);
  nand (_15541_, _12145_, _06790_);
  or (_15542_, _06790_, \uc8051golden_1.ACC [6]);
  and (_15543_, _15542_, _15541_);
  and (_15544_, _15543_, _08644_);
  or (_15545_, _15544_, _07212_);
  or (_15546_, _15545_, _15540_);
  and (_15547_, _15546_, _15537_);
  or (_15548_, _15547_, _07211_);
  nor (_15549_, _08758_, _08161_);
  or (_15550_, _15549_, _08759_);
  or (_15551_, _15550_, _08753_);
  and (_15552_, _15551_, _15548_);
  or (_15553_, _15552_, _07218_);
  and (_15554_, _15553_, _15536_);
  or (_15555_, _15554_, _07351_);
  nor (_15556_, _12144_, _05997_);
  nor (_15557_, _15556_, _07222_);
  and (_15558_, _15557_, _15555_);
  or (_15559_, _15558_, _15534_);
  and (_15560_, _15559_, _08638_);
  nor (_15561_, _12903_, _12902_);
  and (_15562_, _15561_, _07239_);
  or (_15563_, _15562_, _06419_);
  or (_15564_, _15563_, _15560_);
  nand (_15565_, _08161_, _06419_);
  and (_15566_, _15565_, _07423_);
  and (_15567_, _15566_, _15564_);
  not (_15568_, _12905_);
  and (_15569_, _15535_, _15568_);
  and (_15570_, _15569_, _07246_);
  or (_15571_, _15570_, _15567_);
  and (_15572_, _15571_, _05994_);
  or (_15573_, _12145_, _05994_);
  nand (_15574_, _15573_, _06383_);
  or (_15575_, _15574_, _15572_);
  nand (_15576_, _08161_, _06384_);
  and (_15577_, _15576_, _08669_);
  and (_15578_, _15577_, _15575_);
  or (_15579_, _09120_, _06194_);
  nand (_15580_, _15579_, _08160_);
  and (_15581_, _15580_, _07257_);
  or (_15582_, _15581_, _07256_);
  or (_15583_, _15582_, _15578_);
  and (_15584_, _14791_, _07573_);
  or (_15585_, _15584_, _15561_);
  or (_15586_, _15585_, _07777_);
  and (_15587_, _15586_, _07846_);
  and (_15588_, _15587_, _15583_);
  or (_15589_, _15588_, _15533_);
  and (_15590_, _15589_, _08803_);
  nor (_15591_, _08803_, _08118_);
  or (_15592_, _15591_, _08802_);
  or (_15593_, _15592_, _15590_);
  or (_15594_, _08809_, _09440_);
  and (_15595_, _15594_, _08808_);
  and (_15596_, _15595_, _15593_);
  nor (_15597_, _08813_, _08118_);
  and (_15598_, _08940_, \uc8051golden_1.TL0 [6]);
  and (_15599_, _08953_, \uc8051golden_1.B [6]);
  or (_15600_, _15599_, _15598_);
  and (_15601_, _08950_, \uc8051golden_1.P1 [6]);
  and (_15602_, _08928_, \uc8051golden_1.PSW [6]);
  or (_15603_, _15602_, _15601_);
  or (_15604_, _15603_, _15600_);
  and (_15605_, _08944_, \uc8051golden_1.TMOD [6]);
  and (_15606_, _08975_, \uc8051golden_1.ACC [6]);
  or (_15607_, _15606_, _15605_);
  and (_15608_, _08973_, \uc8051golden_1.P0 [6]);
  and (_15609_, _08920_, \uc8051golden_1.SBUF [6]);
  or (_15610_, _15609_, _15608_);
  or (_15611_, _15610_, _15607_);
  and (_15612_, _08961_, \uc8051golden_1.P2 [6]);
  and (_15613_, _08964_, \uc8051golden_1.IP [6]);
  or (_15614_, _15613_, _15612_);
  and (_15615_, _08967_, \uc8051golden_1.IE [6]);
  and (_15616_, _08969_, \uc8051golden_1.P3 [6]);
  or (_15617_, _15616_, _15615_);
  or (_15618_, _15617_, _15614_);
  and (_15619_, _08934_, \uc8051golden_1.TCON [6]);
  and (_15620_, _08947_, \uc8051golden_1.SCON [6]);
  or (_15621_, _15620_, _15619_);
  or (_15622_, _15621_, _15618_);
  or (_15623_, _15622_, _15611_);
  or (_15624_, _15623_, _15604_);
  and (_15625_, _08983_, \uc8051golden_1.TH1 [6]);
  and (_15626_, _09003_, \uc8051golden_1.TH0 [6]);
  and (_15627_, _08998_, \uc8051golden_1.DPH [6]);
  or (_15628_, _15627_, _15626_);
  or (_15629_, _15628_, _15625_);
  and (_15630_, _08996_, \uc8051golden_1.PCON [6]);
  and (_15631_, _08990_, \uc8051golden_1.SP [6]);
  or (_15632_, _15631_, _15630_);
  and (_15633_, _09001_, \uc8051golden_1.DPL [6]);
  and (_15634_, _08987_, \uc8051golden_1.TL1 [6]);
  or (_15635_, _15634_, _15633_);
  or (_15636_, _15635_, _15632_);
  or (_15637_, _15636_, _15629_);
  or (_15638_, _15637_, _15624_);
  or (_15639_, _15638_, _15597_);
  and (_15640_, _15639_, _08807_);
  or (_15641_, _15640_, _09013_);
  or (_15642_, _15641_, _15596_);
  and (_15643_, _09013_, _06340_);
  nor (_15644_, _15643_, _06277_);
  and (_15645_, _15644_, _15642_);
  not (_15646_, _08850_);
  and (_15647_, _15646_, _06277_);
  or (_15648_, _15647_, _05943_);
  or (_15649_, _15648_, _15645_);
  and (_15650_, _12145_, _05943_);
  nor (_15651_, _15650_, _07283_);
  and (_15652_, _15651_, _15649_);
  or (_15653_, _15652_, _15532_);
  and (_15654_, _15653_, _09031_);
  and (_15655_, _11210_, _07285_);
  or (_15656_, _15655_, _15654_);
  and (_15657_, _15656_, _07281_);
  and (_15658_, _15529_, _07280_);
  or (_15659_, _15658_, _15657_);
  and (_15660_, _15659_, _07278_);
  and (_15661_, _11207_, _07277_);
  or (_15662_, _15661_, _05956_);
  or (_15663_, _15662_, _15660_);
  and (_15664_, _12145_, _05956_);
  nor (_15665_, _15664_, _09044_);
  and (_15666_, _15665_, _15663_);
  and (_15667_, _15528_, _09044_);
  or (_15668_, _15667_, _09049_);
  or (_15669_, _15668_, _15666_);
  nand (_15670_, _11209_, _09049_);
  and (_15671_, _15670_, _05967_);
  and (_15672_, _15671_, _15669_);
  and (_15673_, _12144_, _05966_);
  nor (_15674_, _15673_, _07300_);
  nand (_15675_, _15674_, _09061_);
  or (_15676_, _15675_, _15672_);
  or (_15677_, _15539_, _09068_);
  or (_15678_, _15539_, _09061_);
  and (_15679_, _15678_, _14661_);
  and (_15680_, _15679_, _15677_);
  and (_15681_, _15680_, _15676_);
  nor (_15682_, _09395_, _09120_);
  or (_15683_, _15682_, _09396_);
  or (_15684_, _15683_, _07031_);
  and (_15685_, _15684_, _07305_);
  or (_15686_, _15685_, _15681_);
  or (_15687_, _15683_, _14665_);
  and (_15688_, _15687_, _09073_);
  and (_15689_, _15688_, _15686_);
  and (_15690_, _15550_, _07304_);
  or (_15691_, _15690_, _06465_);
  or (_15692_, _15691_, _15689_);
  nand (_15693_, _12293_, _06465_);
  and (_15694_, _15693_, _13005_);
  and (_15695_, _15694_, _15692_);
  and (_15696_, _12144_, _05969_);
  or (_15697_, _15696_, _07311_);
  or (_15698_, _15697_, _15695_);
  or (_15699_, _15561_, _07418_);
  and (_15700_, _15699_, _15698_);
  or (_15701_, _15700_, _09412_);
  or (_15702_, _15526_, _09417_);
  and (_15703_, _15702_, _09416_);
  and (_15704_, _15703_, _15701_);
  or (_15705_, _15704_, _15527_);
  and (_15706_, _15705_, _09439_);
  or (_15707_, _09451_, _09440_);
  nor (_15708_, _09452_, _09439_);
  and (_15709_, _15708_, _15707_);
  or (_15710_, _15709_, _06197_);
  or (_15711_, _15710_, _15706_);
  nor (_15712_, _08526_, _08162_);
  nor (_15713_, _15712_, _08527_);
  or (_15714_, _15713_, _09438_);
  and (_15715_, _15714_, _07415_);
  and (_15716_, _15715_, _15711_);
  or (_15717_, _15716_, _14315_);
  or (_15718_, _14313_, \uc8051golden_1.IRAM[0] [6]);
  and (_15719_, _15718_, _14922_);
  and (_15720_, _15719_, _15717_);
  and (_15721_, _12251_, _06465_);
  not (_15722_, _12111_);
  nor (_15723_, _15722_, _06465_);
  or (_15724_, _15723_, _15721_);
  and (_15725_, _15724_, _14725_);
  and (_15726_, _15725_, _01375_);
  and (_15727_, _15726_, _42545_);
  and (_15728_, _15727_, _14724_);
  or (_40368_, _15728_, _15720_);
  or (_15729_, _14315_, _09460_);
  or (_15730_, _14313_, \uc8051golden_1.IRAM[0] [7]);
  and (_15731_, _15730_, _14922_);
  and (_15732_, _15731_, _15729_);
  and (_15733_, _09498_, _14725_);
  and (_15734_, _15733_, _01375_);
  and (_15735_, _15734_, _42545_);
  and (_15736_, _14724_, _15735_);
  or (_40370_, _15736_, _15732_);
  nand (_15737_, _14495_, _07568_);
  or (_15738_, _15737_, _14500_);
  and (_15739_, _07565_, _07324_);
  and (_15740_, _15739_, _14311_);
  and (_15741_, _15740_, _14485_);
  or (_15742_, _15740_, _07424_);
  nand (_15743_, _15742_, _15737_);
  or (_15744_, _15743_, _15741_);
  and (_40374_, _15744_, _15738_);
  nor (_15745_, _15740_, _06806_);
  and (_15746_, _15740_, _14700_);
  or (_15747_, _15746_, _15745_);
  and (_15748_, _15747_, _15737_);
  not (_15749_, _14712_);
  and (_15750_, _15749_, _14709_);
  and (_15751_, _15750_, _14722_);
  and (_15752_, _15751_, _14732_);
  or (_40375_, _15752_, _15748_);
  not (_15753_, _15740_);
  or (_15754_, _15753_, _14920_);
  or (_15755_, _15740_, \uc8051golden_1.IRAM[1] [2]);
  and (_15756_, _15755_, _15737_);
  and (_15757_, _15756_, _15754_);
  and (_15758_, _14495_, _07568_);
  and (_15759_, _15758_, _14929_);
  or (_40376_, _15759_, _15757_);
  or (_15760_, _15753_, _15116_);
  or (_15761_, _15740_, \uc8051golden_1.IRAM[1] [3]);
  and (_15762_, _15761_, _15737_);
  and (_15763_, _15762_, _15760_);
  and (_15764_, _15751_, _15126_);
  or (_40378_, _15764_, _15763_);
  or (_15765_, _15753_, _15318_);
  or (_15766_, _15740_, \uc8051golden_1.IRAM[1] [4]);
  and (_15767_, _15766_, _15737_);
  and (_15768_, _15767_, _15765_);
  and (_15769_, _15751_, _15329_);
  or (_40379_, _15769_, _15768_);
  or (_15770_, _15753_, _15512_);
  or (_15771_, _15740_, \uc8051golden_1.IRAM[1] [5]);
  and (_15772_, _15771_, _15737_);
  and (_15773_, _15772_, _15770_);
  and (_15774_, _15751_, _15523_);
  or (_40380_, _15774_, _15773_);
  or (_15775_, _15753_, _15716_);
  or (_15776_, _15740_, \uc8051golden_1.IRAM[1] [6]);
  and (_15777_, _15776_, _15737_);
  and (_15778_, _15777_, _15775_);
  and (_15779_, _15751_, _15727_);
  or (_40381_, _15779_, _15778_);
  or (_15780_, _15753_, _09460_);
  or (_15781_, _15740_, \uc8051golden_1.IRAM[1] [7]);
  and (_15782_, _15781_, _15737_);
  and (_15783_, _15782_, _15780_);
  and (_15784_, _15751_, _15735_);
  or (_40382_, _15784_, _15783_);
  and (_15785_, _14495_, _08660_);
  not (_15786_, _15785_);
  or (_15787_, _15786_, _14500_);
  and (_15788_, _07564_, _07417_);
  and (_15789_, _15788_, _14311_);
  and (_15790_, _15789_, _14485_);
  nor (_15791_, _15789_, _07429_);
  or (_15792_, _15791_, _15785_);
  or (_15793_, _15792_, _15790_);
  and (_40387_, _15793_, _15787_);
  nor (_15794_, _15789_, _07145_);
  and (_15795_, _15789_, _14700_);
  or (_15796_, _15795_, _15794_);
  and (_15797_, _15796_, _15786_);
  and (_15798_, _14729_, _07918_);
  and (_15799_, _15798_, _15785_);
  or (_40388_, _15799_, _15797_);
  not (_15800_, _15789_);
  or (_15801_, _15800_, _14920_);
  or (_15802_, _15789_, \uc8051golden_1.IRAM[2] [2]);
  and (_15803_, _15802_, _15786_);
  and (_15804_, _15803_, _15801_);
  and (_15805_, _15785_, _14929_);
  or (_40389_, _15805_, _15804_);
  or (_15806_, _15800_, _15116_);
  or (_15807_, _15789_, \uc8051golden_1.IRAM[2] [3]);
  and (_15808_, _15807_, _15786_);
  and (_15809_, _15808_, _15806_);
  and (_15810_, _15123_, _07918_);
  and (_15811_, _15810_, _15785_);
  or (_40390_, _15811_, _15809_);
  or (_15812_, _15800_, _15318_);
  or (_15813_, _15789_, \uc8051golden_1.IRAM[2] [4]);
  and (_15814_, _15813_, _15786_);
  and (_15815_, _15814_, _15812_);
  and (_15816_, _15326_, _07918_);
  and (_15817_, _15816_, _15785_);
  or (_40391_, _15817_, _15815_);
  or (_15818_, _15800_, _15512_);
  or (_15819_, _15789_, \uc8051golden_1.IRAM[2] [5]);
  and (_15820_, _15819_, _15786_);
  and (_15821_, _15820_, _15818_);
  and (_15822_, _15520_, _07918_);
  and (_15823_, _15822_, _15785_);
  or (_40392_, _15823_, _15821_);
  or (_15824_, _15800_, _15716_);
  or (_15825_, _15789_, \uc8051golden_1.IRAM[2] [6]);
  and (_15826_, _15825_, _15786_);
  and (_15827_, _15826_, _15824_);
  and (_15828_, _15724_, _07918_);
  and (_15829_, _15828_, _15785_);
  or (_40393_, _15829_, _15827_);
  or (_15830_, _15800_, _09460_);
  or (_15831_, _15789_, \uc8051golden_1.IRAM[2] [7]);
  and (_15832_, _15831_, _15786_);
  and (_15833_, _15832_, _15830_);
  and (_15834_, _15785_, _09499_);
  or (_40394_, _15834_, _15833_);
  and (_15835_, _14311_, _07566_);
  or (_15836_, _15835_, \uc8051golden_1.IRAM[3] [0]);
  not (_15837_, _15835_);
  or (_15838_, _15837_, _14485_);
  and (_15839_, _14495_, _06269_);
  not (_15840_, _15839_);
  and (_15841_, _15840_, _15838_);
  and (_15842_, _15841_, _15836_);
  and (_15843_, _14500_, _07918_);
  and (_15844_, _15843_, _15839_);
  or (_40398_, _15844_, _15842_);
  nor (_15845_, _15835_, _07149_);
  and (_15846_, _15835_, _14700_);
  or (_15847_, _15846_, _15845_);
  and (_15848_, _15847_, _15840_);
  and (_15849_, _15839_, _15798_);
  or (_40399_, _15849_, _15848_);
  and (_15850_, _14929_, _07918_);
  or (_15851_, _15850_, _15840_);
  and (_15852_, _15835_, _14920_);
  nor (_15853_, _15835_, _07580_);
  or (_15854_, _15853_, _15839_);
  or (_15855_, _15854_, _15852_);
  and (_40400_, _15855_, _15851_);
  or (_15856_, _15837_, _15116_);
  or (_15857_, _15835_, \uc8051golden_1.IRAM[3] [3]);
  and (_15858_, _15857_, _15840_);
  and (_15859_, _15858_, _15856_);
  and (_15860_, _15839_, _15810_);
  or (_40401_, _15860_, _15859_);
  or (_15861_, _15837_, _15318_);
  or (_15862_, _15835_, \uc8051golden_1.IRAM[3] [4]);
  and (_15863_, _15862_, _15840_);
  and (_15864_, _15863_, _15861_);
  and (_15865_, _15839_, _15816_);
  or (_40403_, _15865_, _15864_);
  or (_15866_, _15837_, _15512_);
  or (_15867_, _15835_, \uc8051golden_1.IRAM[3] [5]);
  and (_15868_, _15867_, _15840_);
  and (_15869_, _15868_, _15866_);
  and (_15870_, _15839_, _15822_);
  or (_40404_, _15870_, _15869_);
  or (_15871_, _15837_, _15716_);
  or (_15872_, _15835_, \uc8051golden_1.IRAM[3] [6]);
  and (_15873_, _15872_, _15840_);
  and (_15874_, _15873_, _15871_);
  and (_15875_, _15839_, _15828_);
  or (_40405_, _15875_, _15874_);
  or (_15876_, _15837_, _09460_);
  or (_15877_, _15835_, \uc8051golden_1.IRAM[3] [7]);
  and (_15878_, _15877_, _15840_);
  and (_15879_, _15878_, _15876_);
  and (_15880_, _15839_, _09499_);
  or (_40406_, _15880_, _15879_);
  and (_15881_, _07906_, _07713_);
  and (_15882_, _15881_, _14309_);
  not (_15883_, _15882_);
  or (_15884_, _15883_, _14485_);
  and (_15885_, _14488_, _14718_);
  and (_15886_, _15885_, _06271_);
  not (_15887_, _15886_);
  or (_15888_, _15882_, \uc8051golden_1.IRAM[4] [0]);
  and (_15889_, _15888_, _15887_);
  and (_15890_, _15889_, _15884_);
  and (_15891_, _15886_, _15843_);
  or (_40410_, _15891_, _15890_);
  or (_15892_, _15883_, _14700_);
  or (_15893_, _15882_, \uc8051golden_1.IRAM[4] [1]);
  and (_15894_, _15893_, _15887_);
  and (_15895_, _15894_, _15892_);
  and (_15896_, _15886_, _15798_);
  or (_40412_, _15896_, _15895_);
  or (_15897_, _15883_, _14920_);
  or (_15898_, _15882_, \uc8051golden_1.IRAM[4] [2]);
  and (_15899_, _15898_, _15887_);
  and (_15900_, _15899_, _15897_);
  and (_15901_, _15886_, _15850_);
  or (_40413_, _15901_, _15900_);
  or (_15902_, _15883_, _15116_);
  or (_15903_, _15882_, \uc8051golden_1.IRAM[4] [3]);
  and (_15904_, _15903_, _15887_);
  and (_15905_, _15904_, _15902_);
  and (_15906_, _15886_, _15810_);
  or (_40414_, _15906_, _15905_);
  or (_15907_, _15883_, _15318_);
  or (_15908_, _15882_, \uc8051golden_1.IRAM[4] [4]);
  and (_15909_, _15908_, _15887_);
  and (_15910_, _15909_, _15907_);
  and (_15911_, _15886_, _15816_);
  or (_40415_, _15911_, _15910_);
  or (_15912_, _15883_, _15512_);
  or (_15913_, _15882_, \uc8051golden_1.IRAM[4] [5]);
  and (_15914_, _15913_, _15887_);
  and (_15915_, _15914_, _15912_);
  and (_15916_, _15886_, _15822_);
  or (_40416_, _15916_, _15915_);
  or (_15917_, _15883_, _15716_);
  or (_15918_, _15882_, \uc8051golden_1.IRAM[4] [6]);
  and (_15919_, _15918_, _15887_);
  and (_15920_, _15919_, _15917_);
  and (_15921_, _15886_, _15828_);
  or (_40418_, _15921_, _15920_);
  or (_15922_, _15883_, _09460_);
  or (_15923_, _15882_, \uc8051golden_1.IRAM[4] [7]);
  and (_15924_, _15923_, _15887_);
  and (_15925_, _15924_, _15922_);
  and (_15926_, _15886_, _09499_);
  or (_40419_, _15926_, _15925_);
  and (_15927_, _15881_, _15739_);
  not (_15928_, _15927_);
  or (_15929_, _15928_, _14485_);
  and (_15930_, _15885_, _07568_);
  not (_15931_, _15930_);
  or (_15932_, _15927_, \uc8051golden_1.IRAM[5] [0]);
  and (_15933_, _15932_, _15931_);
  and (_15934_, _15933_, _15929_);
  and (_15935_, _15930_, _15843_);
  or (_40423_, _15935_, _15934_);
  or (_15936_, _15928_, _14700_);
  or (_15937_, _15927_, \uc8051golden_1.IRAM[5] [1]);
  and (_15938_, _15937_, _15931_);
  and (_15939_, _15938_, _15936_);
  and (_15940_, _15930_, _15798_);
  or (_40424_, _15940_, _15939_);
  or (_15941_, _15928_, _14920_);
  or (_15942_, _15927_, \uc8051golden_1.IRAM[5] [2]);
  and (_15943_, _15942_, _15931_);
  and (_15944_, _15943_, _15941_);
  and (_15945_, _15930_, _15850_);
  or (_40425_, _15945_, _15944_);
  or (_15946_, _15928_, _15116_);
  or (_15947_, _15927_, \uc8051golden_1.IRAM[5] [3]);
  and (_15948_, _15947_, _15931_);
  and (_15949_, _15948_, _15946_);
  and (_15950_, _15930_, _15810_);
  or (_40426_, _15950_, _15949_);
  or (_15951_, _15928_, _15318_);
  or (_15952_, _15927_, \uc8051golden_1.IRAM[5] [4]);
  and (_15953_, _15952_, _15931_);
  and (_15954_, _15953_, _15951_);
  and (_15955_, _15930_, _15816_);
  or (_40427_, _15955_, _15954_);
  or (_15956_, _15928_, _15512_);
  or (_15957_, _15927_, \uc8051golden_1.IRAM[5] [5]);
  and (_15958_, _15957_, _15931_);
  and (_15959_, _15958_, _15956_);
  and (_15960_, _15930_, _15822_);
  or (_40429_, _15960_, _15959_);
  or (_15961_, _15928_, _15716_);
  or (_15962_, _15927_, \uc8051golden_1.IRAM[5] [6]);
  and (_15963_, _15962_, _15931_);
  and (_15964_, _15963_, _15961_);
  and (_15965_, _15930_, _15828_);
  or (_40430_, _15965_, _15964_);
  or (_15966_, _15928_, _09460_);
  or (_15967_, _15927_, \uc8051golden_1.IRAM[5] [7]);
  and (_15968_, _15967_, _15931_);
  and (_15969_, _15968_, _15966_);
  and (_15970_, _15930_, _09499_);
  or (_40431_, _15970_, _15969_);
  not (_15971_, _07417_);
  nor (_15972_, _07565_, _15971_);
  and (_15973_, _15881_, _15972_);
  not (_15974_, _15973_);
  or (_15975_, _15974_, _14485_);
  and (_15976_, _15885_, _08660_);
  not (_15977_, _15976_);
  or (_15978_, _15973_, \uc8051golden_1.IRAM[6] [0]);
  and (_15979_, _15978_, _15977_);
  and (_15980_, _15979_, _15975_);
  and (_15981_, _15976_, _15843_);
  or (_40435_, _15981_, _15980_);
  or (_15982_, _15974_, _14700_);
  or (_15983_, _15973_, \uc8051golden_1.IRAM[6] [1]);
  and (_15984_, _15983_, _15977_);
  and (_15985_, _15984_, _15982_);
  and (_15986_, _15976_, _15798_);
  or (_40436_, _15986_, _15985_);
  or (_15987_, _15974_, _14920_);
  or (_15988_, _15973_, \uc8051golden_1.IRAM[6] [2]);
  and (_15989_, _15988_, _15977_);
  and (_15990_, _15989_, _15987_);
  and (_15991_, _15976_, _15850_);
  or (_40437_, _15991_, _15990_);
  or (_15992_, _15974_, _15116_);
  or (_15993_, _15973_, \uc8051golden_1.IRAM[6] [3]);
  and (_15994_, _15993_, _15977_);
  and (_15995_, _15994_, _15992_);
  and (_15996_, _15976_, _15810_);
  or (_40438_, _15996_, _15995_);
  or (_15997_, _15974_, _15318_);
  or (_15998_, _15973_, \uc8051golden_1.IRAM[6] [4]);
  and (_15999_, _15998_, _15977_);
  and (_16000_, _15999_, _15997_);
  and (_16001_, _15976_, _15816_);
  or (_40439_, _16001_, _16000_);
  or (_16002_, _15974_, _15512_);
  or (_16003_, _15973_, \uc8051golden_1.IRAM[6] [5]);
  and (_16004_, _16003_, _15977_);
  and (_16005_, _16004_, _16002_);
  and (_16006_, _15976_, _15822_);
  or (_40441_, _16006_, _16005_);
  or (_16007_, _15974_, _15716_);
  or (_16008_, _15973_, \uc8051golden_1.IRAM[6] [6]);
  and (_16009_, _16008_, _15977_);
  and (_16010_, _16009_, _16007_);
  and (_16011_, _15976_, _15828_);
  or (_40442_, _16011_, _16010_);
  or (_16012_, _15974_, _09460_);
  or (_16013_, _15973_, \uc8051golden_1.IRAM[6] [7]);
  and (_16014_, _16013_, _15977_);
  and (_16015_, _16014_, _16012_);
  and (_16016_, _15976_, _09499_);
  or (_40443_, _16016_, _16015_);
  and (_16017_, _15881_, _07566_);
  not (_16018_, _16017_);
  or (_16019_, _16018_, _14485_);
  and (_16020_, _15885_, _06269_);
  not (_16021_, _16020_);
  or (_16022_, _16017_, \uc8051golden_1.IRAM[7] [0]);
  and (_16023_, _16022_, _16021_);
  and (_16024_, _16023_, _16019_);
  and (_16025_, _16020_, _15843_);
  or (_40446_, _16025_, _16024_);
  or (_16026_, _16018_, _14700_);
  or (_16027_, _16017_, \uc8051golden_1.IRAM[7] [1]);
  and (_16028_, _16027_, _16021_);
  and (_16029_, _16028_, _16026_);
  and (_16030_, _16020_, _15798_);
  or (_40447_, _16030_, _16029_);
  or (_16031_, _16018_, _14920_);
  or (_16032_, _16017_, \uc8051golden_1.IRAM[7] [2]);
  and (_16033_, _16032_, _16021_);
  and (_16034_, _16033_, _16031_);
  and (_16035_, _16020_, _15850_);
  or (_40448_, _16035_, _16034_);
  or (_16036_, _16018_, _15116_);
  or (_16037_, _16017_, \uc8051golden_1.IRAM[7] [3]);
  and (_16038_, _16037_, _16021_);
  and (_16039_, _16038_, _16036_);
  and (_16040_, _16020_, _15810_);
  or (_40449_, _16040_, _16039_);
  or (_16041_, _16018_, _15318_);
  or (_16042_, _16017_, \uc8051golden_1.IRAM[7] [4]);
  and (_16043_, _16042_, _16021_);
  and (_16044_, _16043_, _16041_);
  and (_16045_, _16020_, _15816_);
  or (_40452_, _16045_, _16044_);
  or (_16046_, _16018_, _15512_);
  or (_16047_, _16017_, \uc8051golden_1.IRAM[7] [5]);
  and (_16048_, _16047_, _16021_);
  and (_16049_, _16048_, _16046_);
  and (_16050_, _16020_, _15822_);
  or (_40453_, _16050_, _16049_);
  or (_16051_, _16018_, _15716_);
  or (_16052_, _16017_, \uc8051golden_1.IRAM[7] [6]);
  and (_16053_, _16052_, _16021_);
  and (_16054_, _16053_, _16051_);
  and (_16055_, _16020_, _15828_);
  or (_40454_, _16055_, _16054_);
  or (_16056_, _16018_, _09460_);
  or (_16057_, _16017_, \uc8051golden_1.IRAM[7] [7]);
  and (_16058_, _16057_, _16021_);
  and (_16059_, _16058_, _16056_);
  and (_16060_, _16020_, _09499_);
  or (_40455_, _16060_, _16059_);
  and (_16061_, _14310_, _07712_);
  and (_16062_, _16061_, _14309_);
  not (_16063_, _16062_);
  nor (_16064_, _16063_, _14485_);
  nor (_16065_, _16062_, \uc8051golden_1.IRAM[8] [0]);
  or (_16066_, _16065_, _16064_);
  and (_16067_, _07919_, _14714_);
  and (_16068_, _16067_, _06271_);
  not (_16069_, _16068_);
  nand (_16070_, _16069_, _16066_);
  or (_16071_, _16069_, _15843_);
  and (_40458_, _16071_, _16070_);
  or (_16072_, _16063_, _14700_);
  or (_16073_, _16062_, \uc8051golden_1.IRAM[8] [1]);
  and (_16074_, _16073_, _16069_);
  and (_16075_, _16074_, _16072_);
  and (_16076_, _16068_, _15798_);
  or (_40461_, _16076_, _16075_);
  or (_16077_, _16063_, _14920_);
  or (_16078_, _16062_, \uc8051golden_1.IRAM[8] [2]);
  and (_16079_, _16078_, _16069_);
  and (_16080_, _16079_, _16077_);
  and (_16081_, _16068_, _15850_);
  or (_40462_, _16081_, _16080_);
  or (_16082_, _16063_, _15116_);
  or (_16083_, _16062_, \uc8051golden_1.IRAM[8] [3]);
  and (_16084_, _16083_, _16069_);
  and (_16085_, _16084_, _16082_);
  and (_16086_, _16068_, _15810_);
  or (_40463_, _16086_, _16085_);
  or (_16087_, _16063_, _15318_);
  or (_16088_, _16062_, \uc8051golden_1.IRAM[8] [4]);
  and (_16089_, _16088_, _16069_);
  and (_16090_, _16089_, _16087_);
  and (_16091_, _16068_, _15816_);
  or (_40464_, _16091_, _16090_);
  or (_16092_, _16063_, _15512_);
  or (_16093_, _16062_, \uc8051golden_1.IRAM[8] [5]);
  and (_16094_, _16093_, _16069_);
  and (_16095_, _16094_, _16092_);
  and (_16096_, _16068_, _15822_);
  or (_40465_, _16096_, _16095_);
  or (_16097_, _16063_, _15716_);
  or (_16098_, _16062_, \uc8051golden_1.IRAM[8] [6]);
  and (_16099_, _16098_, _16069_);
  and (_16100_, _16099_, _16097_);
  and (_16101_, _16068_, _15828_);
  or (_40467_, _16101_, _16100_);
  or (_16102_, _16063_, _09460_);
  or (_16103_, _16062_, \uc8051golden_1.IRAM[8] [7]);
  and (_16104_, _16103_, _16069_);
  and (_16105_, _16104_, _16102_);
  and (_16106_, _16068_, _09499_);
  or (_40468_, _16106_, _16105_);
  and (_16107_, _16061_, _15739_);
  not (_16108_, _16107_);
  or (_16109_, _16108_, _14485_);
  and (_16110_, _16067_, _07568_);
  not (_16111_, _16110_);
  or (_16112_, _16107_, \uc8051golden_1.IRAM[9] [0]);
  and (_16113_, _16112_, _16111_);
  and (_16114_, _16113_, _16109_);
  and (_16115_, _16110_, _15843_);
  or (_40472_, _16115_, _16114_);
  or (_16116_, _16108_, _14700_);
  or (_16117_, _16107_, \uc8051golden_1.IRAM[9] [1]);
  and (_16118_, _16117_, _16111_);
  and (_16119_, _16118_, _16116_);
  and (_16120_, _16110_, _15798_);
  or (_40473_, _16120_, _16119_);
  or (_16121_, _16108_, _14920_);
  or (_16122_, _16107_, \uc8051golden_1.IRAM[9] [2]);
  and (_16123_, _16122_, _16111_);
  and (_16124_, _16123_, _16121_);
  and (_16125_, _16110_, _15850_);
  or (_40474_, _16125_, _16124_);
  or (_16126_, _16108_, _15116_);
  or (_16127_, _16107_, \uc8051golden_1.IRAM[9] [3]);
  and (_16128_, _16127_, _16111_);
  and (_16129_, _16128_, _16126_);
  and (_16130_, _16110_, _15810_);
  or (_40475_, _16130_, _16129_);
  or (_16131_, _16108_, _15318_);
  or (_16132_, _16107_, \uc8051golden_1.IRAM[9] [4]);
  and (_16133_, _16132_, _16111_);
  and (_16134_, _16133_, _16131_);
  and (_16135_, _16110_, _15816_);
  or (_40476_, _16135_, _16134_);
  or (_16136_, _16108_, _15512_);
  or (_16137_, _16107_, \uc8051golden_1.IRAM[9] [5]);
  and (_16138_, _16137_, _16111_);
  and (_16139_, _16138_, _16136_);
  and (_16140_, _16110_, _15822_);
  or (_40478_, _16140_, _16139_);
  or (_16141_, _16108_, _15716_);
  or (_16142_, _16107_, \uc8051golden_1.IRAM[9] [6]);
  and (_16143_, _16142_, _16111_);
  and (_16144_, _16143_, _16141_);
  and (_16145_, _16110_, _15828_);
  or (_40479_, _16145_, _16144_);
  or (_16146_, _16108_, _09460_);
  or (_16147_, _16107_, \uc8051golden_1.IRAM[9] [7]);
  and (_16148_, _16147_, _16111_);
  and (_16149_, _16148_, _16146_);
  and (_16150_, _16110_, _09499_);
  or (_40480_, _16150_, _16149_);
  and (_16151_, _16061_, _15788_);
  not (_16152_, _16151_);
  or (_16153_, _16152_, _14485_);
  and (_16154_, _16067_, _08660_);
  not (_16155_, _16154_);
  or (_16156_, _16151_, \uc8051golden_1.IRAM[10] [0]);
  and (_16157_, _16156_, _16155_);
  and (_16158_, _16157_, _16153_);
  and (_16159_, _16154_, _15843_);
  or (_40484_, _16159_, _16158_);
  or (_16160_, _16152_, _14700_);
  or (_16161_, _16151_, \uc8051golden_1.IRAM[10] [1]);
  and (_16162_, _16161_, _16155_);
  and (_16163_, _16162_, _16160_);
  and (_16164_, _16154_, _15798_);
  or (_40485_, _16164_, _16163_);
  or (_16165_, _16152_, _14920_);
  or (_16166_, _16151_, \uc8051golden_1.IRAM[10] [2]);
  and (_16167_, _16166_, _16155_);
  and (_16168_, _16167_, _16165_);
  and (_16169_, _16154_, _15850_);
  or (_40486_, _16169_, _16168_);
  or (_16170_, _16152_, _15116_);
  or (_16171_, _16151_, \uc8051golden_1.IRAM[10] [3]);
  and (_16172_, _16171_, _16155_);
  and (_16173_, _16172_, _16170_);
  and (_16174_, _16154_, _15810_);
  or (_40487_, _16174_, _16173_);
  or (_16175_, _16152_, _15318_);
  or (_16176_, _16151_, \uc8051golden_1.IRAM[10] [4]);
  and (_16177_, _16176_, _16155_);
  and (_16178_, _16177_, _16175_);
  and (_16179_, _16154_, _15816_);
  or (_40488_, _16179_, _16178_);
  or (_16180_, _16152_, _15512_);
  or (_16181_, _16151_, \uc8051golden_1.IRAM[10] [5]);
  and (_16182_, _16181_, _16155_);
  and (_16183_, _16182_, _16180_);
  and (_16184_, _16154_, _15822_);
  or (_40490_, _16184_, _16183_);
  or (_16185_, _16152_, _15716_);
  or (_16186_, _16151_, \uc8051golden_1.IRAM[10] [6]);
  and (_16187_, _16186_, _16155_);
  and (_16188_, _16187_, _16185_);
  and (_16189_, _16154_, _15828_);
  or (_40491_, _16189_, _16188_);
  or (_16190_, _16152_, _09460_);
  or (_16191_, _16151_, \uc8051golden_1.IRAM[10] [7]);
  and (_16192_, _16191_, _16155_);
  and (_16193_, _16192_, _16190_);
  and (_16194_, _16154_, _09499_);
  or (_40492_, _16194_, _16193_);
  and (_16195_, _16061_, _07566_);
  not (_16196_, _16195_);
  or (_16197_, _16196_, _14485_);
  and (_16198_, _16067_, _06269_);
  not (_16199_, _16198_);
  or (_16200_, _16195_, \uc8051golden_1.IRAM[11] [0]);
  and (_16201_, _16200_, _16199_);
  and (_16202_, _16201_, _16197_);
  and (_16203_, _16198_, _15843_);
  or (_40495_, _16203_, _16202_);
  or (_16204_, _16196_, _14700_);
  or (_16205_, _16195_, \uc8051golden_1.IRAM[11] [1]);
  and (_16206_, _16205_, _16199_);
  and (_16207_, _16206_, _16204_);
  and (_16208_, _16198_, _15798_);
  or (_40496_, _16208_, _16207_);
  or (_16209_, _16196_, _14920_);
  or (_16210_, _16195_, \uc8051golden_1.IRAM[11] [2]);
  and (_16211_, _16210_, _16199_);
  and (_16212_, _16211_, _16209_);
  and (_16213_, _16198_, _15850_);
  or (_40497_, _16213_, _16212_);
  or (_16214_, _16196_, _15116_);
  or (_16215_, _16195_, \uc8051golden_1.IRAM[11] [3]);
  and (_16216_, _16215_, _16199_);
  and (_16217_, _16216_, _16214_);
  and (_16218_, _16198_, _15810_);
  or (_40498_, _16218_, _16217_);
  or (_16219_, _16196_, _15318_);
  or (_16220_, _16195_, \uc8051golden_1.IRAM[11] [4]);
  and (_16221_, _16220_, _16199_);
  and (_16222_, _16221_, _16219_);
  and (_16223_, _16198_, _15816_);
  or (_40501_, _16223_, _16222_);
  or (_16224_, _16196_, _15512_);
  or (_16225_, _16195_, \uc8051golden_1.IRAM[11] [5]);
  and (_16226_, _16225_, _16199_);
  and (_16227_, _16226_, _16224_);
  and (_16228_, _16198_, _15822_);
  or (_40502_, _16228_, _16227_);
  or (_16229_, _16196_, _15716_);
  or (_16230_, _16195_, \uc8051golden_1.IRAM[11] [6]);
  and (_16231_, _16230_, _16199_);
  and (_16232_, _16231_, _16229_);
  and (_16233_, _16198_, _15828_);
  or (_40503_, _16233_, _16232_);
  or (_16234_, _16196_, _09460_);
  or (_16235_, _16195_, \uc8051golden_1.IRAM[11] [7]);
  and (_16236_, _16235_, _16199_);
  and (_16237_, _16236_, _16234_);
  and (_16238_, _16198_, _09499_);
  or (_40504_, _16238_, _16237_);
  not (_16239_, _07712_);
  and (_16240_, _14310_, _16239_);
  and (_16241_, _14309_, _16240_);
  not (_16242_, _16241_);
  or (_16243_, _16242_, _14485_);
  and (_16244_, _07920_, _06271_);
  not (_16245_, _16244_);
  or (_16246_, _16241_, \uc8051golden_1.IRAM[12] [0]);
  and (_16247_, _16246_, _16245_);
  and (_16248_, _16247_, _16243_);
  and (_16249_, _16244_, _15843_);
  or (_40508_, _16249_, _16248_);
  or (_16250_, _16242_, _14700_);
  or (_16251_, _16241_, \uc8051golden_1.IRAM[12] [1]);
  and (_16252_, _16251_, _16245_);
  and (_16253_, _16252_, _16250_);
  and (_16254_, _16244_, _15798_);
  or (_40509_, _16254_, _16253_);
  or (_16255_, _16242_, _14920_);
  or (_16256_, _16241_, \uc8051golden_1.IRAM[12] [2]);
  and (_16257_, _16256_, _16245_);
  and (_16258_, _16257_, _16255_);
  and (_16259_, _16244_, _15850_);
  or (_40510_, _16259_, _16258_);
  nand (_16260_, _14309_, _07907_);
  nand (_16261_, _16260_, _07767_);
  and (_16262_, _16261_, _16245_);
  or (_16263_, _16260_, _15116_);
  and (_16264_, _16263_, _16262_);
  and (_16265_, _16244_, _15810_);
  or (_40512_, _16265_, _16264_);
  or (_16266_, _16241_, \uc8051golden_1.IRAM[12] [4]);
  and (_16267_, _16266_, _16245_);
  or (_16268_, _16242_, _15318_);
  and (_16269_, _16268_, _16267_);
  and (_16270_, _16244_, _15816_);
  or (_40513_, _16270_, _16269_);
  or (_16271_, _16241_, \uc8051golden_1.IRAM[12] [5]);
  and (_16272_, _16271_, _16245_);
  or (_16273_, _16242_, _15512_);
  and (_16274_, _16273_, _16272_);
  and (_16275_, _16244_, _15822_);
  or (_40514_, _16275_, _16274_);
  or (_16276_, _16241_, \uc8051golden_1.IRAM[12] [6]);
  and (_16277_, _16276_, _16245_);
  or (_16278_, _16242_, _15716_);
  and (_16279_, _16278_, _16277_);
  and (_16280_, _16244_, _15828_);
  or (_40515_, _16280_, _16279_);
  or (_16281_, _16241_, \uc8051golden_1.IRAM[12] [7]);
  and (_16282_, _16281_, _16245_);
  or (_16283_, _16242_, _09460_);
  and (_16284_, _16283_, _16282_);
  and (_16285_, _16244_, _09499_);
  or (_40516_, _16285_, _16284_);
  and (_16286_, _15739_, _07907_);
  and (_16287_, _16286_, _14485_);
  or (_16288_, _16286_, _07464_);
  not (_16289_, _07568_);
  nand (_16290_, _14488_, _07915_);
  or (_16291_, _16290_, _16289_);
  nand (_16292_, _16291_, _16288_);
  or (_16293_, _16292_, _16287_);
  and (_16294_, _07920_, _07568_);
  not (_16295_, _16294_);
  or (_16296_, _16295_, _15843_);
  and (_40520_, _16296_, _16293_);
  and (_16297_, _15739_, _16240_);
  not (_16298_, _16297_);
  or (_16299_, _16298_, _14700_);
  or (_16300_, _16297_, \uc8051golden_1.IRAM[13] [1]);
  and (_16301_, _16300_, _16295_);
  and (_16302_, _16301_, _16299_);
  and (_16303_, _16294_, _15798_);
  or (_40521_, _16303_, _16302_);
  or (_16304_, _16286_, \uc8051golden_1.IRAM[13] [2]);
  and (_16305_, _16304_, _16295_);
  or (_16306_, _16298_, _14920_);
  and (_16307_, _16306_, _16305_);
  and (_16308_, _16294_, _15850_);
  or (_40523_, _16308_, _16307_);
  or (_16309_, _16286_, \uc8051golden_1.IRAM[13] [3]);
  and (_16310_, _16309_, _16295_);
  or (_16311_, _16298_, _15116_);
  and (_16312_, _16311_, _16310_);
  and (_16313_, _16294_, _15810_);
  or (_40524_, _16313_, _16312_);
  or (_16314_, _16298_, _15318_);
  or (_16315_, _16286_, \uc8051golden_1.IRAM[13] [4]);
  and (_16316_, _16315_, _16295_);
  and (_16317_, _16316_, _16314_);
  and (_16318_, _16294_, _15816_);
  or (_40525_, _16318_, _16317_);
  or (_16319_, _16286_, \uc8051golden_1.IRAM[13] [5]);
  and (_16320_, _16319_, _16295_);
  or (_16321_, _16298_, _15512_);
  and (_16322_, _16321_, _16320_);
  and (_16323_, _16294_, _15822_);
  or (_40526_, _16323_, _16322_);
  or (_16324_, _16286_, \uc8051golden_1.IRAM[13] [6]);
  and (_16325_, _16324_, _16295_);
  or (_16326_, _16298_, _15716_);
  and (_16327_, _16326_, _16325_);
  and (_16328_, _16294_, _15828_);
  or (_40527_, _16328_, _16327_);
  or (_16329_, _16286_, \uc8051golden_1.IRAM[13] [7]);
  and (_16330_, _16329_, _16295_);
  or (_16331_, _16298_, _09460_);
  and (_16332_, _16331_, _16330_);
  and (_16333_, _16294_, _09499_);
  or (_40528_, _16333_, _16332_);
  and (_16334_, _15788_, _16240_);
  not (_16335_, _16334_);
  or (_16336_, _16335_, _14485_);
  and (_16337_, _08660_, _07920_);
  not (_16338_, _16337_);
  or (_16339_, _16334_, \uc8051golden_1.IRAM[14] [0]);
  and (_16340_, _16339_, _16338_);
  and (_16341_, _16340_, _16336_);
  and (_16342_, _16337_, _15843_);
  or (_40532_, _16342_, _16341_);
  or (_16343_, _16335_, _14700_);
  or (_16344_, _16334_, \uc8051golden_1.IRAM[14] [1]);
  and (_16345_, _16344_, _16338_);
  and (_16346_, _16345_, _16343_);
  and (_16347_, _16337_, _15798_);
  or (_40533_, _16347_, _16346_);
  nand (_16348_, _15788_, _07907_);
  nand (_16349_, _16348_, _07609_);
  and (_16350_, _16349_, _16338_);
  or (_16351_, _16348_, _14920_);
  and (_16352_, _16351_, _16350_);
  and (_16353_, _16337_, _15850_);
  or (_40535_, _16353_, _16352_);
  nand (_16354_, _16348_, _07757_);
  and (_16355_, _16354_, _16338_);
  or (_16356_, _16348_, _15116_);
  and (_16357_, _16356_, _16355_);
  and (_16358_, _16337_, _15810_);
  or (_40536_, _16358_, _16357_);
  or (_16359_, _16348_, _15318_);
  or (_16360_, _16334_, \uc8051golden_1.IRAM[14] [4]);
  and (_16361_, _16360_, _16338_);
  and (_16362_, _16361_, _16359_);
  and (_16363_, _16337_, _15816_);
  or (_40537_, _16363_, _16362_);
  or (_16364_, _16334_, \uc8051golden_1.IRAM[14] [5]);
  and (_16365_, _16364_, _16338_);
  or (_16366_, _16335_, _15512_);
  and (_16367_, _16366_, _16365_);
  and (_16368_, _16337_, _15822_);
  or (_40538_, _16368_, _16367_);
  or (_16369_, _16348_, _15716_);
  or (_16370_, _16334_, \uc8051golden_1.IRAM[14] [6]);
  and (_16371_, _16370_, _16338_);
  and (_16372_, _16371_, _16369_);
  and (_16373_, _16337_, _15828_);
  or (_40539_, _16373_, _16372_);
  or (_16374_, _16334_, \uc8051golden_1.IRAM[14] [7]);
  and (_16375_, _16374_, _16338_);
  or (_16376_, _16335_, _09460_);
  and (_16377_, _16376_, _16375_);
  and (_16378_, _16337_, _09499_);
  or (_40541_, _16378_, _16377_);
  and (_16379_, _16240_, _07566_);
  not (_16380_, _16379_);
  or (_16381_, _14485_, _16380_);
  nand (_16382_, _07908_, _07460_);
  and (_16383_, _16382_, _07922_);
  and (_16384_, _16383_, _16381_);
  and (_16385_, _15843_, _07921_);
  or (_40544_, _16385_, _16384_);
  or (_16386_, _14700_, _16380_);
  or (_16387_, _16379_, \uc8051golden_1.IRAM[15] [1]);
  and (_16388_, _16387_, _07922_);
  and (_16389_, _16388_, _16386_);
  and (_16390_, _15798_, _07921_);
  or (_40545_, _16390_, _16389_);
  nand (_16391_, _07908_, _07611_);
  and (_16392_, _16391_, _07922_);
  or (_16393_, _14920_, _07908_);
  and (_16394_, _16393_, _16392_);
  and (_16395_, _15850_, _07921_);
  or (_40547_, _16395_, _16394_);
  nand (_16396_, _07908_, _07760_);
  and (_16397_, _16396_, _07922_);
  or (_16398_, _15116_, _07908_);
  and (_16399_, _16398_, _16397_);
  and (_16400_, _15810_, _07921_);
  or (_40548_, _16400_, _16399_);
  or (_16401_, _16379_, \uc8051golden_1.IRAM[15] [4]);
  and (_16402_, _16401_, _07922_);
  or (_16403_, _15318_, _16380_);
  and (_16404_, _16403_, _16402_);
  and (_16405_, _15816_, _07921_);
  or (_40549_, _16405_, _16404_);
  or (_16406_, _16379_, \uc8051golden_1.IRAM[15] [5]);
  and (_16407_, _16406_, _07922_);
  or (_16408_, _15512_, _16380_);
  and (_16409_, _16408_, _16407_);
  and (_16410_, _15822_, _07921_);
  or (_40550_, _16410_, _16409_);
  or (_16411_, _15716_, _07908_);
  or (_16412_, _16379_, \uc8051golden_1.IRAM[15] [6]);
  and (_16413_, _16412_, _07922_);
  and (_16414_, _16413_, _16411_);
  and (_16415_, _15828_, _07921_);
  or (_40551_, _16415_, _16414_);
  nor (_16416_, _01375_, _10084_);
  and (_16417_, _07992_, \uc8051golden_1.ACC [0]);
  and (_16418_, _16417_, _08521_);
  nor (_16419_, _07992_, _10084_);
  or (_16420_, _16419_, _07276_);
  or (_16421_, _16420_, _16418_);
  and (_16422_, _07992_, _08817_);
  or (_16423_, _16422_, _16419_);
  or (_16424_, _16423_, _06276_);
  and (_16425_, _07992_, _07473_);
  or (_16426_, _16425_, _16419_);
  or (_16427_, _16426_, _06293_);
  nor (_16428_, _08521_, _09504_);
  or (_16429_, _16428_, _16419_);
  or (_16430_, _16429_, _07210_);
  or (_16431_, _16417_, _16419_);
  and (_16432_, _16431_, _07199_);
  nor (_16433_, _07199_, _10084_);
  or (_16434_, _16433_, _06401_);
  or (_16435_, _16434_, _16432_);
  and (_16436_, _16435_, _06396_);
  and (_16437_, _16436_, _16430_);
  and (_16438_, _14339_, _08618_);
  nor (_16439_, _08618_, _10084_);
  or (_16440_, _16439_, _16438_);
  and (_16441_, _16440_, _06395_);
  or (_16442_, _16441_, _16437_);
  and (_16443_, _16442_, _07221_);
  and (_16444_, _16426_, _06399_);
  or (_16445_, _16444_, _06406_);
  or (_16446_, _16445_, _16443_);
  or (_16447_, _16431_, _06414_);
  and (_16448_, _16447_, _06844_);
  and (_16449_, _16448_, _16446_);
  and (_16450_, _16419_, _06393_);
  or (_16451_, _16450_, _06387_);
  or (_16452_, _16451_, _16449_);
  or (_16453_, _16429_, _07245_);
  and (_16454_, _16453_, _16452_);
  or (_16455_, _16454_, _09538_);
  nor (_16456_, _10020_, _10018_);
  nor (_16457_, _16456_, _10021_);
  or (_16458_, _16457_, _09544_);
  and (_16459_, _16458_, _06446_);
  and (_16460_, _16459_, _16455_);
  and (_16461_, _14371_, _08618_);
  or (_16462_, _16461_, _16439_);
  and (_16463_, _16462_, _06300_);
  or (_16464_, _16463_, _10059_);
  or (_16465_, _16464_, _16460_);
  and (_16466_, _16465_, _16427_);
  or (_16467_, _16466_, _06281_);
  and (_16468_, _07992_, _09446_);
  or (_16469_, _16419_, _06282_);
  or (_16470_, _16469_, _16468_);
  and (_16471_, _16470_, _16467_);
  or (_16472_, _16471_, _06015_);
  and (_16473_, _14426_, _07992_);
  or (_16474_, _16419_, _06279_);
  or (_16475_, _16474_, _16473_);
  and (_16476_, _16475_, _10078_);
  and (_16477_, _16476_, _16472_);
  nand (_16478_, _10418_, _06045_);
  or (_16479_, _10412_, _10387_);
  or (_16480_, _10418_, _16479_);
  and (_16481_, _16480_, _10072_);
  and (_16482_, _16481_, _16478_);
  or (_16483_, _16482_, _06275_);
  or (_16484_, _16483_, _16477_);
  and (_16485_, _16484_, _16424_);
  or (_16486_, _16485_, _06474_);
  and (_16487_, _14324_, _07992_);
  or (_16488_, _16487_, _16419_);
  or (_16489_, _16488_, _07282_);
  and (_16490_, _16489_, _07284_);
  and (_16491_, _16490_, _16486_);
  nor (_16492_, _12538_, _09504_);
  or (_16493_, _16492_, _16419_);
  nor (_16494_, _16418_, _07284_);
  and (_16495_, _16494_, _16493_);
  or (_16496_, _16495_, _16491_);
  and (_16497_, _16496_, _07279_);
  nand (_16498_, _16423_, _06478_);
  nor (_16499_, _16498_, _16428_);
  or (_16500_, _16499_, _06569_);
  or (_16501_, _16500_, _16497_);
  and (_16502_, _16501_, _16421_);
  or (_16503_, _16502_, _06479_);
  and (_16504_, _14320_, _07992_);
  or (_16505_, _16419_, _09043_);
  or (_16506_, _16505_, _16504_);
  and (_16507_, _16506_, _09048_);
  and (_16508_, _16507_, _16503_);
  and (_16509_, _16493_, _06572_);
  or (_16510_, _16509_, _06606_);
  or (_16511_, _16510_, _16508_);
  or (_16512_, _16429_, _07037_);
  and (_16513_, _16512_, _16511_);
  or (_16514_, _16513_, _06234_);
  or (_16515_, _16419_, _06807_);
  and (_16516_, _16515_, _16514_);
  or (_16517_, _16516_, _06195_);
  or (_16518_, _16429_, _06196_);
  and (_16519_, _16518_, _01375_);
  and (_16520_, _16519_, _16517_);
  or (_16521_, _16520_, _16416_);
  and (_42889_, _16521_, _42545_);
  nor (_16522_, _01375_, _10079_);
  nor (_16523_, _07992_, _10079_);
  nor (_16524_, _11223_, _09504_);
  or (_16525_, _16524_, _16523_);
  or (_16526_, _16525_, _09048_);
  nand (_16527_, _07992_, _07090_);
  or (_16528_, _07992_, \uc8051golden_1.B [1]);
  and (_16529_, _16528_, _06275_);
  and (_16530_, _16529_, _16527_);
  nor (_16531_, _08618_, _10079_);
  and (_16532_, _14517_, _08618_);
  or (_16533_, _16532_, _16531_);
  and (_16534_, _16533_, _06393_);
  nor (_16535_, _09504_, _07196_);
  or (_16536_, _16535_, _16523_);
  or (_16537_, _16536_, _07221_);
  and (_16538_, _14532_, _07992_);
  not (_16539_, _16538_);
  and (_16540_, _16539_, _16528_);
  or (_16541_, _16540_, _07210_);
  and (_16542_, _07992_, \uc8051golden_1.ACC [1]);
  or (_16543_, _16542_, _16523_);
  and (_16544_, _16543_, _07199_);
  nor (_16545_, _07199_, _10079_);
  or (_16546_, _16545_, _06401_);
  or (_16547_, _16546_, _16544_);
  and (_16548_, _16547_, _06396_);
  and (_16549_, _16548_, _16541_);
  and (_16550_, _14514_, _08618_);
  or (_16551_, _16550_, _16531_);
  and (_16552_, _16551_, _06395_);
  or (_16553_, _16552_, _06399_);
  or (_16554_, _16553_, _16549_);
  and (_16555_, _16554_, _16537_);
  or (_16556_, _16555_, _06406_);
  or (_16557_, _16543_, _06414_);
  and (_16558_, _16557_, _06844_);
  and (_16559_, _16558_, _16556_);
  or (_16560_, _16559_, _16534_);
  and (_16561_, _16560_, _07245_);
  and (_16562_, _16550_, _14513_);
  or (_16563_, _16562_, _16531_);
  and (_16564_, _16563_, _06387_);
  or (_16565_, _16564_, _09538_);
  or (_16566_, _16565_, _16561_);
  nor (_16567_, _10023_, _09965_);
  nor (_16568_, _16567_, _10024_);
  or (_16569_, _16568_, _09544_);
  and (_16570_, _16569_, _06446_);
  and (_16571_, _16570_, _16566_);
  or (_16572_, _16531_, _14560_);
  and (_16573_, _16572_, _06300_);
  and (_16574_, _16573_, _16551_);
  or (_16575_, _16574_, _10059_);
  or (_16576_, _16575_, _16571_);
  or (_16577_, _16536_, _06293_);
  and (_16578_, _16577_, _16576_);
  or (_16579_, _16578_, _06281_);
  and (_16580_, _07992_, _09445_);
  or (_16581_, _16523_, _06282_);
  or (_16582_, _16581_, _16580_);
  and (_16583_, _16582_, _06279_);
  and (_16584_, _16583_, _16579_);
  or (_16585_, _14615_, _09504_);
  and (_16586_, _16528_, _06015_);
  and (_16587_, _16586_, _16585_);
  or (_16588_, _16587_, _10072_);
  or (_16589_, _16588_, _16584_);
  nor (_16590_, _10413_, _10411_);
  or (_16591_, _16590_, _10414_);
  nor (_16592_, _16591_, _10418_);
  and (_16593_, _10418_, _10384_);
  or (_16594_, _16593_, _16592_);
  or (_16595_, _16594_, _10078_);
  and (_16596_, _16595_, _06276_);
  and (_16597_, _16596_, _16589_);
  or (_16598_, _16597_, _16530_);
  and (_16599_, _16598_, _07282_);
  or (_16600_, _14507_, _09504_);
  and (_16601_, _16528_, _06474_);
  and (_16602_, _16601_, _16600_);
  or (_16603_, _16602_, _06582_);
  or (_16604_, _16603_, _16599_);
  and (_16605_, _11224_, _07992_);
  or (_16606_, _16605_, _16523_);
  or (_16607_, _16606_, _07284_);
  and (_16608_, _16607_, _07279_);
  and (_16609_, _16608_, _16604_);
  or (_16610_, _14505_, _09504_);
  and (_16611_, _16528_, _06478_);
  and (_16612_, _16611_, _16610_);
  or (_16613_, _16612_, _06569_);
  or (_16614_, _16613_, _16609_);
  and (_16615_, _16542_, _08477_);
  or (_16616_, _16523_, _07276_);
  or (_16617_, _16616_, _16615_);
  and (_16618_, _16617_, _09043_);
  and (_16619_, _16618_, _16614_);
  or (_16620_, _16527_, _08477_);
  and (_16621_, _16528_, _06479_);
  and (_16622_, _16621_, _16620_);
  or (_16623_, _16622_, _06572_);
  or (_16624_, _16623_, _16619_);
  and (_16625_, _16624_, _16526_);
  or (_16626_, _16625_, _06606_);
  or (_16627_, _16540_, _07037_);
  and (_16628_, _16627_, _06807_);
  and (_16629_, _16628_, _16626_);
  and (_16630_, _16533_, _06234_);
  or (_16631_, _16630_, _06195_);
  or (_16632_, _16631_, _16629_);
  or (_16633_, _16523_, _06196_);
  or (_16634_, _16633_, _16538_);
  and (_16635_, _16634_, _01375_);
  and (_16636_, _16635_, _16632_);
  or (_16637_, _16636_, _16522_);
  and (_42890_, _16637_, _42545_);
  nor (_16638_, _01375_, _10291_);
  nor (_16639_, _07992_, _10291_);
  and (_16640_, _07992_, _08994_);
  or (_16641_, _16640_, _16639_);
  or (_16642_, _16641_, _06276_);
  nor (_16643_, _09504_, _07623_);
  or (_16644_, _16643_, _16639_);
  or (_16645_, _16644_, _06293_);
  and (_16646_, _14751_, _08618_);
  and (_16647_, _16646_, _14778_);
  nor (_16648_, _08618_, _10291_);
  or (_16649_, _16648_, _07245_);
  or (_16650_, _16649_, _16647_);
  or (_16651_, _16644_, _07221_);
  and (_16652_, _14754_, _07992_);
  or (_16653_, _16652_, _16639_);
  or (_16654_, _16653_, _07210_);
  and (_16655_, _07992_, \uc8051golden_1.ACC [2]);
  or (_16656_, _16655_, _16639_);
  and (_16657_, _16656_, _07199_);
  nor (_16658_, _07199_, _10291_);
  or (_16659_, _16658_, _06401_);
  or (_16660_, _16659_, _16657_);
  and (_16661_, _16660_, _06396_);
  and (_16662_, _16661_, _16654_);
  or (_16663_, _16648_, _16646_);
  and (_16664_, _16663_, _06395_);
  or (_16665_, _16664_, _06399_);
  or (_16666_, _16665_, _16662_);
  and (_16667_, _16666_, _16651_);
  or (_16668_, _16667_, _06406_);
  or (_16669_, _16656_, _06414_);
  and (_16670_, _16669_, _06844_);
  and (_16671_, _16670_, _16668_);
  and (_16672_, _14749_, _08618_);
  or (_16673_, _16672_, _16648_);
  and (_16674_, _16673_, _06393_);
  or (_16675_, _16674_, _06387_);
  or (_16676_, _16675_, _16671_);
  and (_16677_, _16676_, _16650_);
  or (_16678_, _16677_, _09538_);
  or (_16679_, _10025_, _09920_);
  and (_16680_, _16679_, _10026_);
  or (_16681_, _16680_, _09544_);
  and (_16682_, _16681_, _06446_);
  and (_16683_, _16682_, _16678_);
  and (_16684_, _14793_, _08618_);
  or (_16685_, _16684_, _16648_);
  and (_16686_, _16685_, _06300_);
  or (_16687_, _16686_, _10059_);
  or (_16688_, _16687_, _16683_);
  and (_16689_, _16688_, _16645_);
  or (_16690_, _16689_, _06281_);
  and (_16691_, _07992_, _09444_);
  or (_16692_, _16639_, _06282_);
  or (_16693_, _16692_, _16691_);
  and (_16694_, _16693_, _16690_);
  or (_16695_, _16694_, _06015_);
  and (_16696_, _14848_, _07992_);
  or (_16697_, _16639_, _06279_);
  or (_16698_, _16697_, _16696_);
  and (_16699_, _16698_, _10078_);
  and (_16700_, _16699_, _16695_);
  not (_16701_, _10418_);
  or (_16702_, _16701_, _10375_);
  nor (_16703_, _10414_, _10385_);
  not (_16704_, _16703_);
  and (_16705_, _16704_, _10378_);
  nor (_16706_, _16704_, _10378_);
  nor (_16707_, _16706_, _16705_);
  or (_16708_, _16707_, _10418_);
  and (_16709_, _16708_, _10072_);
  and (_16710_, _16709_, _16702_);
  or (_16711_, _16710_, _06275_);
  or (_16712_, _16711_, _16700_);
  and (_16713_, _16712_, _16642_);
  or (_16714_, _16713_, _06474_);
  and (_16715_, _14744_, _07992_);
  or (_16716_, _16715_, _16639_);
  or (_16717_, _16716_, _07282_);
  and (_16718_, _16717_, _07284_);
  and (_16719_, _16718_, _16714_);
  and (_16720_, _11221_, _07992_);
  or (_16721_, _16720_, _16639_);
  and (_16722_, _16721_, _06582_);
  or (_16723_, _16722_, _16719_);
  and (_16724_, _16723_, _07279_);
  or (_16725_, _16639_, _08433_);
  and (_16726_, _16641_, _06478_);
  and (_16727_, _16726_, _16725_);
  or (_16728_, _16727_, _16724_);
  and (_16729_, _16728_, _07276_);
  and (_16730_, _16656_, _06569_);
  and (_16731_, _16730_, _16725_);
  or (_16732_, _16731_, _06479_);
  or (_16733_, _16732_, _16729_);
  and (_16734_, _14741_, _07992_);
  or (_16735_, _16639_, _09043_);
  or (_16736_, _16735_, _16734_);
  and (_16737_, _16736_, _09048_);
  and (_16738_, _16737_, _16733_);
  nor (_16739_, _11220_, _09504_);
  or (_16740_, _16739_, _16639_);
  and (_16741_, _16740_, _06572_);
  or (_16742_, _16741_, _06606_);
  or (_16743_, _16742_, _16738_);
  or (_16744_, _16653_, _07037_);
  and (_16745_, _16744_, _06807_);
  and (_16746_, _16745_, _16743_);
  and (_16747_, _16673_, _06234_);
  or (_16748_, _16747_, _06195_);
  or (_16749_, _16748_, _16746_);
  and (_16750_, _14917_, _07992_);
  or (_16751_, _16639_, _06196_);
  or (_16752_, _16751_, _16750_);
  and (_16753_, _16752_, _01375_);
  and (_16754_, _16753_, _16749_);
  or (_16755_, _16754_, _16638_);
  and (_42891_, _16755_, _42545_);
  nor (_16756_, _01375_, _10166_);
  nor (_16757_, _07992_, _10166_);
  and (_16758_, _07992_, _08815_);
  or (_16759_, _16758_, _16757_);
  or (_16760_, _16759_, _06276_);
  nor (_16761_, _09504_, _07775_);
  or (_16762_, _16761_, _16757_);
  or (_16763_, _16762_, _06293_);
  nor (_16764_, _08618_, _10166_);
  and (_16765_, _14951_, _08618_);
  or (_16766_, _16765_, _16764_);
  or (_16767_, _16764_, _14968_);
  and (_16768_, _16767_, _16766_);
  or (_16769_, _16768_, _07245_);
  and (_16770_, _14947_, _07992_);
  or (_16771_, _16770_, _16757_);
  or (_16772_, _16771_, _07210_);
  and (_16773_, _07992_, \uc8051golden_1.ACC [3]);
  or (_16774_, _16773_, _16757_);
  and (_16775_, _16774_, _07199_);
  nor (_16776_, _07199_, _10166_);
  or (_16777_, _16776_, _06401_);
  or (_16778_, _16777_, _16775_);
  and (_16779_, _16778_, _06396_);
  and (_16780_, _16779_, _16772_);
  and (_16781_, _16766_, _06395_);
  or (_16782_, _16781_, _06399_);
  or (_16783_, _16782_, _16780_);
  or (_16784_, _16762_, _07221_);
  and (_16785_, _16784_, _16783_);
  or (_16786_, _16785_, _06406_);
  or (_16787_, _16774_, _06414_);
  and (_16788_, _16787_, _06844_);
  and (_16789_, _16788_, _16786_);
  and (_16790_, _14961_, _08618_);
  or (_16791_, _16790_, _16764_);
  and (_16792_, _16791_, _06393_);
  or (_16793_, _16792_, _06387_);
  or (_16794_, _16793_, _16789_);
  and (_16795_, _16794_, _16769_);
  or (_16796_, _16795_, _09538_);
  nor (_16797_, _10028_, _09862_);
  nor (_16798_, _16797_, _10029_);
  or (_16799_, _16798_, _09544_);
  and (_16800_, _16799_, _06446_);
  and (_16801_, _16800_, _16796_);
  and (_16802_, _14985_, _08618_);
  or (_16803_, _16802_, _16764_);
  and (_16804_, _16803_, _06300_);
  or (_16805_, _16804_, _10059_);
  or (_16806_, _16805_, _16801_);
  and (_16807_, _16806_, _16763_);
  or (_16808_, _16807_, _06281_);
  and (_16809_, _07992_, _09443_);
  or (_16810_, _16757_, _06282_);
  or (_16811_, _16810_, _16809_);
  and (_16812_, _16811_, _16808_);
  or (_16813_, _16812_, _06015_);
  and (_16814_, _15039_, _07992_);
  or (_16815_, _16757_, _06279_);
  or (_16816_, _16815_, _16814_);
  and (_16817_, _16816_, _10078_);
  and (_16818_, _16817_, _16813_);
  nor (_16819_, _16705_, _10377_);
  nor (_16820_, _16819_, _10370_);
  and (_16821_, _16819_, _10370_);
  or (_16822_, _16821_, _16820_);
  or (_16823_, _16822_, _10418_);
  or (_16824_, _16701_, _10367_);
  and (_16825_, _16824_, _10072_);
  and (_16826_, _16825_, _16823_);
  or (_16827_, _16826_, _06275_);
  or (_16828_, _16827_, _16818_);
  and (_16829_, _16828_, _16760_);
  or (_16830_, _16829_, _06474_);
  and (_16831_, _14934_, _07992_);
  or (_16832_, _16831_, _16757_);
  or (_16833_, _16832_, _07282_);
  and (_16834_, _16833_, _07284_);
  and (_16835_, _16834_, _16830_);
  and (_16836_, _12535_, _07992_);
  or (_16837_, _16836_, _16757_);
  and (_16838_, _16837_, _06582_);
  or (_16839_, _16838_, _16835_);
  and (_16840_, _16839_, _07279_);
  or (_16841_, _16757_, _08389_);
  and (_16842_, _16759_, _06478_);
  and (_16843_, _16842_, _16841_);
  or (_16844_, _16843_, _16840_);
  and (_16845_, _16844_, _07276_);
  and (_16846_, _16774_, _06569_);
  and (_16847_, _16846_, _16841_);
  or (_16848_, _16847_, _06479_);
  or (_16849_, _16848_, _16845_);
  and (_16850_, _14931_, _07992_);
  or (_16851_, _16757_, _09043_);
  or (_16852_, _16851_, _16850_);
  and (_16853_, _16852_, _09048_);
  and (_16854_, _16853_, _16849_);
  nor (_16855_, _11218_, _09504_);
  or (_16856_, _16855_, _16757_);
  and (_16857_, _16856_, _06572_);
  or (_16858_, _16857_, _06606_);
  or (_16859_, _16858_, _16854_);
  or (_16860_, _16771_, _07037_);
  and (_16861_, _16860_, _06807_);
  and (_16862_, _16861_, _16859_);
  and (_16863_, _16791_, _06234_);
  or (_16864_, _16863_, _06195_);
  or (_16865_, _16864_, _16862_);
  and (_16866_, _15113_, _07992_);
  or (_16867_, _16757_, _06196_);
  or (_16868_, _16867_, _16866_);
  and (_16869_, _16868_, _01375_);
  and (_16870_, _16869_, _16865_);
  or (_16871_, _16870_, _16756_);
  and (_42892_, _16871_, _42545_);
  nor (_16872_, _01375_, _10094_);
  nor (_16873_, _07992_, _10094_);
  and (_16874_, _08883_, _07992_);
  or (_16875_, _16874_, _16873_);
  or (_16876_, _16875_, _06276_);
  and (_16877_, _15243_, _07992_);
  or (_16878_, _16877_, _16873_);
  and (_16879_, _16878_, _06015_);
  nor (_16880_, _08618_, _10094_);
  and (_16881_, _15168_, _08618_);
  or (_16882_, _16881_, _16880_);
  and (_16883_, _16882_, _06393_);
  and (_16884_, _15130_, _07992_);
  or (_16885_, _16884_, _16873_);
  or (_16886_, _16885_, _07210_);
  and (_16887_, _07992_, \uc8051golden_1.ACC [4]);
  or (_16888_, _16887_, _16873_);
  and (_16889_, _16888_, _07199_);
  nor (_16890_, _07199_, _10094_);
  or (_16891_, _16890_, _06401_);
  or (_16892_, _16891_, _16889_);
  and (_16893_, _16892_, _06396_);
  and (_16894_, _16893_, _16886_);
  and (_16895_, _15139_, _08618_);
  or (_16896_, _16895_, _16880_);
  and (_16897_, _16896_, _06395_);
  or (_16898_, _16897_, _06399_);
  or (_16899_, _16898_, _16894_);
  nor (_16900_, _09504_, _08301_);
  or (_16901_, _16900_, _16873_);
  or (_16902_, _16901_, _07221_);
  and (_16903_, _16902_, _16899_);
  or (_16904_, _16903_, _06406_);
  or (_16905_, _16888_, _06414_);
  and (_16906_, _16905_, _06844_);
  and (_16907_, _16906_, _16904_);
  or (_16908_, _16907_, _16883_);
  and (_16909_, _16908_, _07245_);
  or (_16910_, _16880_, _15138_);
  and (_16911_, _16910_, _06387_);
  and (_16912_, _16911_, _16896_);
  or (_16913_, _16912_, _09538_);
  or (_16914_, _16913_, _16909_);
  or (_16915_, _10032_, _10030_);
  and (_16916_, _16915_, _10033_);
  or (_16917_, _16916_, _09544_);
  and (_16918_, _16917_, _06446_);
  and (_16919_, _16918_, _16914_);
  and (_16920_, _15189_, _08618_);
  or (_16921_, _16920_, _16880_);
  and (_16922_, _16921_, _06300_);
  or (_16923_, _16922_, _10059_);
  or (_16924_, _16923_, _16919_);
  or (_16925_, _16901_, _06293_);
  and (_16926_, _16925_, _16924_);
  or (_16927_, _16926_, _06281_);
  and (_16928_, _07992_, _09442_);
  or (_16929_, _16873_, _06282_);
  or (_16930_, _16929_, _16928_);
  and (_16931_, _16930_, _06279_);
  and (_16932_, _16931_, _16927_);
  or (_16933_, _16932_, _16879_);
  and (_16934_, _16933_, _10078_);
  or (_16935_, _16701_, _10359_);
  nor (_16936_, _16819_, _10368_);
  or (_16937_, _16936_, _10369_);
  nand (_16938_, _16937_, _10405_);
  or (_16939_, _16937_, _10405_);
  and (_16940_, _16939_, _16938_);
  or (_16941_, _16940_, _10418_);
  and (_16942_, _16941_, _10072_);
  and (_16943_, _16942_, _16935_);
  or (_16944_, _16943_, _06275_);
  or (_16945_, _16944_, _16934_);
  and (_16946_, _16945_, _16876_);
  or (_16947_, _16946_, _06474_);
  and (_16948_, _15135_, _07992_);
  or (_16949_, _16948_, _16873_);
  or (_16950_, _16949_, _07282_);
  and (_16951_, _16950_, _07284_);
  and (_16952_, _16951_, _16947_);
  and (_16953_, _11216_, _07992_);
  or (_16954_, _16953_, _16873_);
  and (_16955_, _16954_, _06582_);
  or (_16956_, _16955_, _16952_);
  and (_16957_, _16956_, _07279_);
  or (_16958_, _16873_, _08345_);
  and (_16959_, _16875_, _06478_);
  and (_16960_, _16959_, _16958_);
  or (_16961_, _16960_, _16957_);
  and (_16962_, _16961_, _07276_);
  and (_16963_, _16888_, _06569_);
  and (_16964_, _16963_, _16958_);
  or (_16965_, _16964_, _06479_);
  or (_16966_, _16965_, _16962_);
  and (_16967_, _15134_, _07992_);
  or (_16968_, _16873_, _09043_);
  or (_16969_, _16968_, _16967_);
  and (_16970_, _16969_, _09048_);
  and (_16971_, _16970_, _16966_);
  nor (_16972_, _11215_, _09504_);
  or (_16973_, _16972_, _16873_);
  and (_16974_, _16973_, _06572_);
  or (_16975_, _16974_, _06606_);
  or (_16976_, _16975_, _16971_);
  or (_16977_, _16885_, _07037_);
  and (_16978_, _16977_, _06807_);
  and (_16979_, _16978_, _16976_);
  and (_16980_, _16882_, _06234_);
  or (_16981_, _16980_, _06195_);
  or (_16982_, _16981_, _16979_);
  and (_16983_, _15315_, _07992_);
  or (_16984_, _16873_, _06196_);
  or (_16985_, _16984_, _16983_);
  and (_16986_, _16985_, _01375_);
  and (_16987_, _16986_, _16982_);
  or (_16988_, _16987_, _16872_);
  and (_42893_, _16988_, _42545_);
  nor (_16989_, _01375_, _10095_);
  nor (_16990_, _07992_, _10095_);
  and (_16991_, _15446_, _07992_);
  or (_16992_, _16991_, _16990_);
  and (_16993_, _16992_, _06015_);
  nor (_16994_, _09504_, _08207_);
  or (_16995_, _16994_, _16990_);
  or (_16996_, _16995_, _06293_);
  nor (_16997_, _08618_, _10095_);
  and (_16998_, _15345_, _08618_);
  or (_16999_, _16998_, _16997_);
  and (_17000_, _16999_, _06393_);
  and (_17001_, _15348_, _07992_);
  or (_17002_, _17001_, _16990_);
  or (_17003_, _17002_, _07210_);
  and (_17004_, _07992_, \uc8051golden_1.ACC [5]);
  or (_17005_, _17004_, _16990_);
  and (_17006_, _17005_, _07199_);
  nor (_17007_, _07199_, _10095_);
  or (_17008_, _17007_, _06401_);
  or (_17009_, _17008_, _17006_);
  and (_17010_, _17009_, _06396_);
  and (_17011_, _17010_, _17003_);
  and (_17012_, _15341_, _08618_);
  or (_17013_, _17012_, _16997_);
  and (_17014_, _17013_, _06395_);
  or (_17015_, _17014_, _06399_);
  or (_17016_, _17015_, _17011_);
  or (_17017_, _16995_, _07221_);
  and (_17018_, _17017_, _17016_);
  or (_17019_, _17018_, _06406_);
  or (_17020_, _17005_, _06414_);
  and (_17021_, _17020_, _06844_);
  and (_17022_, _17021_, _17019_);
  or (_17023_, _17022_, _17000_);
  and (_17024_, _17023_, _07245_);
  or (_17025_, _16997_, _15378_);
  and (_17026_, _17025_, _06387_);
  and (_17027_, _17026_, _17013_);
  or (_17028_, _17027_, _09538_);
  or (_17029_, _17028_, _17024_);
  or (_17030_, _09735_, _09736_);
  and (_17031_, _17030_, _10034_);
  nor (_17032_, _17031_, _10035_);
  or (_17033_, _17032_, _09544_);
  and (_17034_, _17033_, _06446_);
  and (_17035_, _17034_, _17029_);
  or (_17036_, _16997_, _15342_);
  and (_17037_, _17036_, _06300_);
  and (_17038_, _17037_, _17013_);
  or (_17039_, _17038_, _10059_);
  or (_17040_, _17039_, _17035_);
  and (_17041_, _17040_, _16996_);
  or (_17042_, _17041_, _06281_);
  and (_17043_, _07992_, _09441_);
  or (_17044_, _16990_, _06282_);
  or (_17045_, _17044_, _17043_);
  and (_17046_, _17045_, _06279_);
  and (_17047_, _17046_, _17042_);
  or (_17048_, _17047_, _16993_);
  and (_17049_, _17048_, _10078_);
  or (_17050_, _16701_, _10351_);
  not (_17051_, _10396_);
  and (_17052_, _16938_, _17051_);
  nor (_17053_, _17052_, _10406_);
  and (_17054_, _17052_, _10406_);
  or (_17055_, _17054_, _17053_);
  or (_17056_, _17055_, _10418_);
  and (_17057_, _17056_, _10072_);
  and (_17058_, _17057_, _17050_);
  or (_17059_, _17058_, _06275_);
  or (_17060_, _17059_, _17049_);
  and (_17061_, _08958_, _07992_);
  or (_17062_, _17061_, _16990_);
  or (_17063_, _17062_, _06276_);
  and (_17064_, _17063_, _17060_);
  or (_17065_, _17064_, _06474_);
  and (_17066_, _15338_, _07992_);
  or (_17067_, _17066_, _16990_);
  or (_17068_, _17067_, _07282_);
  and (_17069_, _17068_, _07284_);
  and (_17070_, _17069_, _17065_);
  and (_17071_, _12542_, _07992_);
  or (_17072_, _17071_, _16990_);
  and (_17073_, _17072_, _06582_);
  or (_17074_, _17073_, _17070_);
  and (_17075_, _17074_, _07279_);
  or (_17076_, _16990_, _08256_);
  and (_17077_, _17062_, _06478_);
  and (_17078_, _17077_, _17076_);
  or (_17079_, _17078_, _17075_);
  and (_17080_, _17079_, _07276_);
  and (_17081_, _17005_, _06569_);
  and (_17082_, _17081_, _17076_);
  or (_17083_, _17082_, _06479_);
  or (_17084_, _17083_, _17080_);
  and (_17085_, _15335_, _07992_);
  or (_17086_, _16990_, _09043_);
  or (_17087_, _17086_, _17085_);
  and (_17088_, _17087_, _09048_);
  and (_17089_, _17088_, _17084_);
  nor (_17090_, _11212_, _09504_);
  or (_17091_, _17090_, _16990_);
  and (_17092_, _17091_, _06572_);
  or (_17093_, _17092_, _06606_);
  or (_17094_, _17093_, _17089_);
  or (_17095_, _17002_, _07037_);
  and (_17096_, _17095_, _06807_);
  and (_17097_, _17096_, _17094_);
  and (_17098_, _16999_, _06234_);
  or (_17099_, _17098_, _06195_);
  or (_17100_, _17099_, _17097_);
  and (_17101_, _15509_, _07992_);
  or (_17102_, _16990_, _06196_);
  or (_17103_, _17102_, _17101_);
  and (_17104_, _17103_, _01375_);
  and (_17105_, _17104_, _17100_);
  or (_17106_, _17105_, _16989_);
  and (_42894_, _17106_, _42545_);
  nor (_17107_, _01375_, _10336_);
  nor (_17108_, _07992_, _10336_);
  and (_17109_, _15646_, _07992_);
  or (_17110_, _17109_, _17108_);
  or (_17111_, _17110_, _06276_);
  and (_17112_, _15639_, _07992_);
  or (_17113_, _17112_, _17108_);
  and (_17114_, _17113_, _06015_);
  nor (_17115_, _09504_, _08118_);
  or (_17116_, _17115_, _17108_);
  or (_17117_, _17116_, _06293_);
  nor (_17118_, _08618_, _10336_);
  and (_17119_, _15561_, _08618_);
  or (_17120_, _17119_, _17118_);
  and (_17121_, _17120_, _06393_);
  and (_17122_, _15550_, _07992_);
  or (_17123_, _17122_, _17108_);
  or (_17124_, _17123_, _07210_);
  and (_17125_, _07992_, \uc8051golden_1.ACC [6]);
  or (_17126_, _17125_, _17108_);
  and (_17127_, _17126_, _07199_);
  nor (_17128_, _07199_, _10336_);
  or (_17129_, _17128_, _06401_);
  or (_17130_, _17129_, _17127_);
  and (_17131_, _17130_, _06396_);
  and (_17132_, _17131_, _17124_);
  and (_17133_, _15535_, _08618_);
  or (_17134_, _17133_, _17118_);
  and (_17135_, _17134_, _06395_);
  or (_17136_, _17135_, _06399_);
  or (_17137_, _17136_, _17132_);
  or (_17138_, _17116_, _07221_);
  and (_17139_, _17138_, _17137_);
  or (_17140_, _17139_, _06406_);
  or (_17141_, _17126_, _06414_);
  and (_17142_, _17141_, _06844_);
  and (_17143_, _17142_, _17140_);
  or (_17144_, _17143_, _17121_);
  and (_17145_, _17144_, _07245_);
  or (_17146_, _17118_, _15568_);
  and (_17147_, _17146_, _06387_);
  and (_17148_, _17147_, _17134_);
  or (_17149_, _17148_, _09538_);
  or (_17150_, _17149_, _17145_);
  nor (_17151_, _10048_, _10036_);
  nor (_17152_, _17151_, _10049_);
  or (_17153_, _17152_, _09544_);
  and (_17154_, _17153_, _06446_);
  and (_17155_, _17154_, _17150_);
  and (_17156_, _15585_, _08618_);
  or (_17157_, _17156_, _17118_);
  and (_17158_, _17157_, _06300_);
  or (_17159_, _17158_, _10059_);
  or (_17160_, _17159_, _17155_);
  and (_17161_, _17160_, _17117_);
  or (_17162_, _17161_, _06281_);
  and (_17163_, _07992_, _09440_);
  or (_17164_, _17108_, _06282_);
  or (_17165_, _17164_, _17163_);
  and (_17166_, _17165_, _06279_);
  and (_17167_, _17166_, _17162_);
  or (_17168_, _17167_, _17114_);
  and (_17169_, _17168_, _10078_);
  nor (_17170_, _17052_, _10352_);
  or (_17171_, _17170_, _10353_);
  or (_17172_, _17171_, _10408_);
  nand (_17173_, _17171_, _10408_);
  and (_17174_, _17173_, _17172_);
  or (_17175_, _17174_, _10418_);
  nor (_17176_, _10418_, _10078_);
  and (_17177_, _10342_, _10072_);
  or (_17178_, _17177_, _17176_);
  and (_17179_, _17178_, _17175_);
  or (_17180_, _17179_, _06275_);
  or (_17181_, _17180_, _17169_);
  and (_17182_, _17181_, _17111_);
  or (_17183_, _17182_, _06474_);
  and (_17184_, _15531_, _07992_);
  or (_17185_, _17184_, _17108_);
  or (_17186_, _17185_, _07282_);
  and (_17187_, _17186_, _07284_);
  and (_17188_, _17187_, _17183_);
  and (_17189_, _11210_, _07992_);
  or (_17190_, _17189_, _17108_);
  and (_17191_, _17190_, _06582_);
  or (_17192_, _17191_, _17188_);
  and (_17193_, _17192_, _07279_);
  or (_17194_, _17108_, _08162_);
  and (_17195_, _17110_, _06478_);
  and (_17196_, _17195_, _17194_);
  or (_17197_, _17196_, _17193_);
  and (_17198_, _17197_, _07276_);
  and (_17199_, _17126_, _06569_);
  and (_17200_, _17199_, _17194_);
  or (_17201_, _17200_, _06479_);
  or (_17202_, _17201_, _17198_);
  and (_17203_, _15528_, _07992_);
  or (_17204_, _17108_, _09043_);
  or (_17205_, _17204_, _17203_);
  and (_17206_, _17205_, _09048_);
  and (_17207_, _17206_, _17202_);
  nor (_17208_, _11209_, _09504_);
  or (_17209_, _17208_, _17108_);
  and (_17210_, _17209_, _06572_);
  or (_17211_, _17210_, _06606_);
  or (_17212_, _17211_, _17207_);
  or (_17213_, _17123_, _07037_);
  and (_17214_, _17213_, _06807_);
  and (_17215_, _17214_, _17212_);
  and (_17216_, _17120_, _06234_);
  or (_17217_, _17216_, _06195_);
  or (_17218_, _17217_, _17215_);
  and (_17219_, _15713_, _07992_);
  or (_17220_, _17108_, _06196_);
  or (_17221_, _17220_, _17219_);
  and (_17222_, _17221_, _01375_);
  and (_17223_, _17222_, _17218_);
  or (_17224_, _17223_, _17107_);
  and (_42895_, _17224_, _42545_);
  nor (_17225_, _01375_, _06045_);
  nand (_17226_, _11243_, _08651_);
  and (_17227_, _07485_, _06045_);
  nor (_17228_, _17227_, _11143_);
  and (_17229_, _11121_, _17228_);
  nor (_17230_, _10887_, _06045_);
  or (_17231_, _17230_, _10888_);
  or (_17232_, _11091_, _17231_);
  nand (_17233_, _11017_, _12241_);
  nand (_17234_, _12539_, _06580_);
  and (_17235_, _17234_, _10964_);
  nor (_17236_, _10950_, _10565_);
  not (_17237_, _17236_);
  and (_17238_, _17237_, _17228_);
  nand (_17239_, _06840_, _05982_);
  nor (_17240_, _07995_, _06045_);
  and (_17241_, _14426_, _07995_);
  or (_17242_, _17241_, _17240_);
  and (_17243_, _17242_, _06015_);
  and (_17244_, _07995_, _07473_);
  or (_17245_, _17244_, _17240_);
  or (_17246_, _17245_, _06293_);
  not (_17247_, _10644_);
  or (_17248_, _17247_, _07473_);
  nor (_17249_, _10654_, _07212_);
  or (_17250_, _17249_, _09446_);
  and (_17251_, _10663_, _07473_);
  or (_17252_, _06854_, \uc8051golden_1.ACC [0]);
  nand (_17253_, _06854_, \uc8051golden_1.ACC [0]);
  nand (_17254_, _17253_, _17252_);
  nor (_17255_, _17254_, _10663_);
  or (_17256_, _17255_, _10654_);
  or (_17257_, _17256_, _17251_);
  and (_17258_, _17257_, _06002_);
  or (_17259_, _17258_, _07212_);
  and (_17260_, _17259_, _07210_);
  and (_17261_, _17260_, _17250_);
  nor (_17262_, _08521_, _10568_);
  or (_17263_, _17262_, _17240_);
  and (_17264_, _17263_, _06401_);
  or (_17265_, _17264_, _06395_);
  or (_17266_, _17265_, _17261_);
  and (_17267_, _14339_, _08616_);
  nor (_17268_, _08616_, _06045_);
  or (_17269_, _17268_, _06396_);
  or (_17270_, _17269_, _17267_);
  and (_17271_, _17270_, _07221_);
  and (_17272_, _17271_, _17266_);
  and (_17273_, _17245_, _06399_);
  or (_17274_, _17273_, _10644_);
  or (_17275_, _17274_, _17272_);
  and (_17276_, _17275_, _17248_);
  or (_17277_, _17276_, _07233_);
  or (_17278_, _09446_, _10714_);
  and (_17279_, _17278_, _06414_);
  and (_17280_, _17279_, _17277_);
  and (_17281_, _08521_, _06406_);
  or (_17282_, _17281_, _10642_);
  or (_17283_, _17282_, _17280_);
  nand (_17284_, _10642_, _10119_);
  and (_17285_, _17284_, _17283_);
  or (_17286_, _17285_, _06393_);
  or (_17287_, _17240_, _06844_);
  and (_17288_, _17287_, _07245_);
  and (_17289_, _17288_, _17286_);
  and (_17290_, _17263_, _06387_);
  or (_17291_, _17290_, _09538_);
  or (_17292_, _17291_, _17289_);
  nand (_17293_, \uc8051golden_1.B [0], \uc8051golden_1.ACC [0]);
  nand (_17294_, _17293_, _09538_);
  and (_17295_, _17294_, _10740_);
  and (_17296_, _17295_, _17292_);
  nor (_17297_, _10789_, _06045_);
  or (_17298_, _17297_, _10790_);
  and (_17299_, _17298_, _14157_);
  or (_17300_, _17299_, _12586_);
  or (_17301_, _17300_, _17296_);
  nor (_17302_, _10526_, _06045_);
  or (_17303_, _17302_, _10820_);
  or (_17304_, _17303_, _12587_);
  and (_17305_, _17304_, _17301_);
  or (_17306_, _17305_, _06437_);
  nor (_17307_, _10621_, _06045_);
  or (_17308_, _17307_, _10622_);
  or (_17309_, _17308_, _06442_);
  and (_17310_, _17309_, _10573_);
  and (_17311_, _17310_, _17306_);
  and (_17312_, _17231_, _10572_);
  or (_17313_, _17312_, _06022_);
  or (_17314_, _17313_, _17311_);
  nand (_17315_, _06840_, _06022_);
  and (_17316_, _17315_, _06446_);
  and (_17317_, _17316_, _17314_);
  and (_17318_, _14371_, _08616_);
  or (_17319_, _17318_, _17268_);
  and (_17320_, _17319_, _06300_);
  or (_17321_, _17320_, _10059_);
  or (_17322_, _17321_, _17317_);
  and (_17323_, _17322_, _17246_);
  or (_17324_, _17323_, _06281_);
  and (_17325_, _07995_, _09446_);
  or (_17326_, _17240_, _06282_);
  or (_17327_, _17326_, _17325_);
  and (_17328_, _17327_, _06279_);
  and (_17329_, _17328_, _17324_);
  or (_17330_, _17329_, _17243_);
  and (_17331_, _17330_, _10078_);
  or (_17332_, _17176_, _05982_);
  or (_17333_, _17332_, _17331_);
  and (_17334_, _17333_, _17239_);
  or (_17335_, _17334_, _06275_);
  and (_17336_, _07995_, _08817_);
  or (_17338_, _17336_, _17240_);
  or (_17339_, _17338_, _06276_);
  and (_17340_, _17339_, _10934_);
  and (_17341_, _17340_, _17335_);
  nor (_17342_, _10934_, _06840_);
  or (_17343_, _17342_, _10941_);
  or (_17344_, _17343_, _17341_);
  or (_17345_, _10945_, _17228_);
  and (_17346_, _17345_, _17236_);
  and (_17347_, _17346_, _17344_);
  or (_17349_, _17347_, _17238_);
  and (_17350_, _17349_, _10959_);
  and (_17351_, _09390_, _06045_);
  nor (_17352_, _11186_, _17351_);
  and (_17353_, _10953_, _17352_);
  or (_17354_, _17353_, _06580_);
  or (_17355_, _17354_, _17350_);
  and (_17356_, _17355_, _17235_);
  and (_17357_, _10963_, _12242_);
  or (_17358_, _17357_, _06474_);
  or (_17360_, _17358_, _17356_);
  and (_17361_, _14324_, _07995_);
  or (_17362_, _17361_, _17240_);
  or (_17363_, _17362_, _07282_);
  and (_17364_, _17363_, _17360_);
  or (_17365_, _17364_, _06582_);
  or (_17366_, _17240_, _07284_);
  and (_17367_, _17366_, _10980_);
  and (_17368_, _17367_, _17365_);
  and (_17369_, _10983_, _11143_);
  or (_17371_, _17369_, _10559_);
  or (_17372_, _17371_, _17368_);
  or (_17373_, _11186_, _10560_);
  and (_17374_, _17373_, _06568_);
  and (_17375_, _17374_, _17372_);
  or (_17376_, _10989_, _11225_);
  and (_17377_, _17376_, _12722_);
  or (_17378_, _17377_, _17375_);
  or (_17379_, _10990_, _11261_);
  and (_17380_, _17379_, _07279_);
  and (_17382_, _17380_, _17378_);
  nand (_17383_, _17338_, _06478_);
  nor (_17384_, _17383_, _17262_);
  or (_17385_, _17384_, _17382_);
  and (_17386_, _17385_, _10555_);
  nor (_17387_, _17227_, _10555_);
  or (_17388_, _17387_, _11003_);
  or (_17389_, _17388_, _17386_);
  nand (_17390_, _11003_, _17227_);
  and (_17391_, _17390_, _11006_);
  and (_17393_, _17391_, _17389_);
  nor (_17394_, _17227_, _11006_);
  or (_17395_, _17394_, _11011_);
  or (_17396_, _17395_, _17393_);
  nand (_17397_, _11011_, _17351_);
  and (_17398_, _17397_, _06575_);
  and (_17399_, _17398_, _17396_);
  nand (_17400_, _11020_, _12538_);
  and (_17401_, _17400_, _11019_);
  or (_17402_, _17401_, _17399_);
  and (_17403_, _17402_, _17233_);
  or (_17404_, _17403_, _06479_);
  and (_17405_, _14320_, _07995_);
  or (_17406_, _17240_, _09043_);
  or (_17407_, _17406_, _17405_);
  and (_17408_, _17407_, _11028_);
  and (_17409_, _17408_, _17404_);
  and (_17410_, _11030_, _17298_);
  or (_17411_, _17410_, _10471_);
  or (_17412_, _17411_, _17409_);
  or (_17413_, _17303_, _10472_);
  and (_17414_, _17413_, _06579_);
  and (_17415_, _17414_, _17412_);
  or (_17416_, _11059_, _17308_);
  and (_17417_, _17416_, _11061_);
  or (_17418_, _17417_, _17415_);
  and (_17419_, _17418_, _17232_);
  or (_17420_, _17419_, _11089_);
  nand (_17421_, _11089_, _10524_);
  and (_17422_, _17421_, _11120_);
  and (_17423_, _17422_, _17420_);
  or (_17424_, _17423_, _17229_);
  and (_17425_, _17424_, _11165_);
  and (_17426_, _11163_, _17352_);
  or (_17427_, _17426_, _06307_);
  or (_17428_, _17427_, _17425_);
  nand (_17429_, _12539_, _06307_);
  and (_17430_, _17429_, _14289_);
  and (_17431_, _17430_, _17428_);
  and (_17432_, _11203_, _12242_);
  or (_17433_, _17432_, _11243_);
  or (_17434_, _17433_, _17431_);
  and (_17435_, _17434_, _17226_);
  or (_17436_, _17435_, _06606_);
  or (_17437_, _17263_, _07037_);
  and (_17438_, _17437_, _11286_);
  and (_17439_, _17438_, _17436_);
  nor (_17440_, _11290_, _06045_);
  nor (_17441_, _17440_, _12994_);
  or (_17442_, _17441_, _17439_);
  nand (_17443_, _11290_, _05984_);
  and (_17444_, _17443_, _06807_);
  and (_17445_, _17444_, _17442_);
  and (_17446_, _17240_, _06234_);
  or (_17447_, _17446_, _06195_);
  or (_17448_, _17447_, _17445_);
  or (_17449_, _17263_, _06196_);
  and (_17450_, _17449_, _11309_);
  and (_17451_, _17450_, _17448_);
  nor (_17452_, _11315_, _06045_);
  nor (_17453_, _17452_, _13019_);
  or (_17454_, _17453_, _17451_);
  nand (_17455_, _11315_, _05984_);
  and (_17456_, _17455_, _01375_);
  and (_17457_, _17456_, _17454_);
  or (_17458_, _17457_, _17225_);
  and (_42896_, _17458_, _42545_);
  nor (_17459_, _01375_, _05984_);
  or (_17460_, _11070_, _11069_);
  nor (_17461_, _11071_, _06579_);
  and (_17462_, _17461_, _17460_);
  and (_17463_, _07343_, _05965_);
  not (_17464_, _17463_);
  nor (_17465_, _10527_, _10523_);
  nor (_17466_, _17465_, _10528_);
  or (_17467_, _17466_, _17464_);
  not (_17468_, _07095_);
  nor (_17469_, _11141_, _17468_);
  or (_17470_, _11182_, _10560_);
  not (_17471_, _12715_);
  nor (_17472_, _07995_, _05984_);
  or (_17473_, _17472_, _07284_);
  or (_17474_, _11224_, _06581_);
  and (_17475_, _17474_, _10964_);
  nor (_17476_, _10568_, _07196_);
  or (_17477_, _17476_, _17472_);
  or (_17478_, _17477_, _06293_);
  nor (_17479_, _08616_, _05984_);
  and (_17480_, _14514_, _08616_);
  or (_17481_, _17480_, _17479_);
  or (_17482_, _17479_, _14513_);
  and (_17483_, _17482_, _06387_);
  and (_17484_, _17483_, _17481_);
  nand (_17485_, _10644_, _07196_);
  or (_17486_, _17249_, _09445_);
  nor (_17487_, _10664_, _07196_);
  or (_17488_, _06854_, \uc8051golden_1.ACC [1]);
  nand (_17489_, _06854_, \uc8051golden_1.ACC [1]);
  nand (_17490_, _17489_, _17488_);
  nor (_17491_, _17490_, _10663_);
  or (_17492_, _17491_, _10654_);
  or (_17493_, _17492_, _17487_);
  and (_17494_, _17493_, _06002_);
  or (_17495_, _17494_, _07212_);
  and (_17496_, _17495_, _07210_);
  and (_17497_, _17496_, _17486_);
  or (_17498_, _07995_, \uc8051golden_1.ACC [1]);
  and (_17499_, _14532_, _07995_);
  not (_17500_, _17499_);
  and (_17501_, _17500_, _17498_);
  and (_17502_, _17501_, _06401_);
  or (_17503_, _17502_, _10677_);
  or (_17504_, _17503_, _17497_);
  nor (_17505_, _10682_, \uc8051golden_1.PSW [6]);
  nor (_17506_, _17505_, \uc8051golden_1.ACC [1]);
  and (_17507_, _17505_, \uc8051golden_1.ACC [1]);
  nor (_17508_, _17507_, _17506_);
  nand (_17509_, _17508_, _10677_);
  and (_17510_, _17509_, _06407_);
  and (_17511_, _17510_, _17504_);
  and (_17512_, _17481_, _06395_);
  and (_17513_, _17477_, _06399_);
  or (_17514_, _17513_, _10644_);
  or (_17515_, _17514_, _17512_);
  or (_17516_, _17515_, _17511_);
  and (_17517_, _17516_, _17485_);
  or (_17518_, _17517_, _07233_);
  or (_17519_, _09445_, _10714_);
  and (_17520_, _17519_, _06414_);
  and (_17521_, _17520_, _17518_);
  nor (_17522_, _08476_, _06414_);
  or (_17523_, _17522_, _10642_);
  or (_17524_, _17523_, _17521_);
  nand (_17525_, _10642_, _10145_);
  and (_17526_, _17525_, _17524_);
  or (_17527_, _17526_, _06393_);
  and (_17528_, _14517_, _08616_);
  or (_17529_, _17528_, _17479_);
  or (_17530_, _17529_, _06844_);
  and (_17531_, _17530_, _07245_);
  and (_17532_, _17531_, _17527_);
  or (_17533_, _17532_, _17484_);
  and (_17534_, _17533_, _09544_);
  nor (_17535_, _09999_, _09998_);
  nor (_17536_, _17535_, _10000_);
  and (_17537_, _17536_, _09538_);
  or (_17538_, _17537_, _17534_);
  and (_17539_, _17538_, _10740_);
  nor (_17540_, _10783_, _06045_);
  or (_17541_, _17540_, _10788_);
  not (_17542_, _17541_);
  nand (_17543_, _17542_, _11142_);
  or (_17544_, _17542_, _11142_);
  and (_17545_, _17544_, _17543_);
  and (_17546_, _17545_, _14157_);
  or (_17547_, _17546_, _12586_);
  or (_17548_, _17547_, _17539_);
  nor (_17549_, _10516_, _06045_);
  or (_17550_, _17549_, _10525_);
  nor (_17551_, _17550_, _11185_);
  and (_17552_, _17550_, _11185_);
  or (_17553_, _17552_, _17551_);
  or (_17554_, _17553_, _12587_);
  and (_17555_, _17554_, _06442_);
  and (_17556_, _17555_, _17548_);
  nor (_17557_, _10574_, _06045_);
  or (_17558_, _17557_, _10620_);
  nand (_17559_, _17558_, _12537_);
  or (_17560_, _17558_, _12537_);
  and (_17561_, _17560_, _06437_);
  and (_17562_, _17561_, _17559_);
  or (_17563_, _17562_, _10572_);
  or (_17564_, _17563_, _17556_);
  and (_17565_, _12243_, \uc8051golden_1.PSW [7]);
  nor (_17566_, _06840_, \uc8051golden_1.ACC [0]);
  nor (_17567_, _17566_, _11260_);
  and (_17568_, _17566_, _11260_);
  nor (_17569_, _17568_, _17567_);
  or (_17570_, _12242_, _10524_);
  and (_17571_, _17570_, _17569_);
  or (_17572_, _17571_, _17565_);
  or (_17573_, _17572_, _10573_);
  and (_17574_, _17573_, _17564_);
  or (_17575_, _17574_, _06022_);
  nand (_17576_, _06228_, _06022_);
  and (_17577_, _17576_, _06446_);
  and (_17578_, _17577_, _17575_);
  or (_17579_, _17479_, _14560_);
  and (_17580_, _17579_, _06300_);
  and (_17581_, _17580_, _17481_);
  or (_17582_, _17581_, _10059_);
  or (_17583_, _17582_, _17578_);
  and (_17584_, _17583_, _17478_);
  or (_17585_, _17584_, _06281_);
  and (_17586_, _07995_, _09445_);
  or (_17587_, _17472_, _06282_);
  or (_17588_, _17587_, _17586_);
  and (_17589_, _17588_, _06279_);
  and (_17590_, _17589_, _17585_);
  or (_17591_, _14615_, _10568_);
  and (_17592_, _17498_, _06015_);
  and (_17593_, _17592_, _17591_);
  or (_17594_, _17593_, _10072_);
  or (_17595_, _17594_, _17590_);
  nand (_17596_, _10329_, _10072_);
  and (_17597_, _17596_, _17595_);
  or (_17598_, _17597_, _05982_);
  nand (_17599_, _06228_, _05982_);
  and (_17600_, _17599_, _06276_);
  and (_17601_, _17600_, _17598_);
  nand (_17602_, _07995_, _07090_);
  and (_17603_, _17498_, _06275_);
  and (_17604_, _17603_, _17602_);
  or (_17605_, _17604_, _10933_);
  or (_17606_, _17605_, _17601_);
  nand (_17607_, _10933_, _06228_);
  nor (_17608_, _10941_, _10565_);
  and (_17609_, _17608_, _17607_);
  and (_17610_, _17609_, _17606_);
  not (_17611_, _17608_);
  and (_17612_, _17611_, _11142_);
  or (_17613_, _17612_, _10950_);
  or (_17614_, _17613_, _17610_);
  or (_17615_, _10951_, _11142_);
  and (_17616_, _17615_, _10959_);
  and (_17617_, _17616_, _17614_);
  and (_17618_, _10953_, _11185_);
  or (_17619_, _17618_, _06580_);
  or (_17620_, _17619_, _17617_);
  and (_17621_, _17620_, _17475_);
  and (_17622_, _10963_, _11260_);
  or (_17623_, _17622_, _17621_);
  and (_17624_, _17623_, _07282_);
  or (_17625_, _14507_, _10568_);
  and (_17626_, _17498_, _06474_);
  and (_17627_, _17626_, _17625_);
  or (_17628_, _17627_, _06582_);
  or (_17629_, _17628_, _17624_);
  and (_17630_, _17629_, _17473_);
  or (_17631_, _17630_, _17471_);
  or (_17632_, _12715_, _11140_);
  and (_17633_, _17632_, _12717_);
  and (_17634_, _17633_, _17631_);
  not (_17635_, _12717_);
  and (_17636_, _17635_, _11140_);
  or (_17637_, _17636_, _10559_);
  or (_17638_, _17637_, _17634_);
  and (_17639_, _17638_, _17470_);
  or (_17640_, _17639_, _06567_);
  or (_17641_, _11222_, _06568_);
  and (_17642_, _17641_, _10990_);
  and (_17643_, _17642_, _17640_);
  and (_17644_, _10989_, _11258_);
  or (_17645_, _17644_, _17643_);
  and (_17646_, _17645_, _07279_);
  or (_17647_, _14505_, _10568_);
  and (_17648_, _17498_, _06478_);
  and (_17649_, _17648_, _17647_);
  or (_17650_, _17649_, _06784_);
  or (_17651_, _17650_, _17646_);
  nor (_17652_, _11141_, _07095_);
  not (_17653_, _07106_);
  nor (_17654_, _07095_, _10552_);
  and (_17655_, _17654_, _17653_);
  or (_17656_, _17655_, _17652_);
  and (_17657_, _17656_, _17651_);
  or (_17658_, _17657_, _17469_);
  and (_17659_, _06285_, _05946_);
  not (_17660_, _17659_);
  and (_17661_, _17660_, _17658_);
  nor (_17662_, _17660_, _11141_);
  or (_17663_, _17662_, _11011_);
  or (_17664_, _17663_, _17661_);
  not (_17665_, _11011_);
  or (_17666_, _17665_, _11183_);
  and (_17667_, _17666_, _06575_);
  and (_17668_, _17667_, _17664_);
  nand (_17669_, _11020_, _11223_);
  and (_17670_, _17669_, _11019_);
  or (_17671_, _17670_, _17668_);
  nand (_17672_, _11017_, _11259_);
  and (_17673_, _17672_, _09043_);
  and (_17674_, _17673_, _17671_);
  or (_17675_, _17602_, _08477_);
  and (_17676_, _17498_, _06479_);
  and (_17677_, _17676_, _17675_);
  or (_17678_, _17677_, _17674_);
  and (_17679_, _17678_, _11028_);
  nor (_17680_, _11039_, _11038_);
  nor (_17681_, _17680_, _11040_);
  and (_17682_, _17681_, _11030_);
  or (_17683_, _17682_, _17463_);
  or (_17684_, _17683_, _17679_);
  and (_17685_, _17684_, _17467_);
  or (_17686_, _17685_, _06984_);
  not (_17687_, _06984_);
  or (_17688_, _17466_, _17687_);
  and (_17689_, _17688_, _06579_);
  and (_17690_, _17689_, _17686_);
  or (_17691_, _17690_, _17462_);
  and (_17692_, _17691_, _11091_);
  or (_17693_, _11100_, _11099_);
  nor (_17694_, _11101_, _11091_);
  and (_17695_, _17694_, _17693_);
  or (_17696_, _17695_, _11089_);
  or (_17697_, _17696_, _17692_);
  nand (_17698_, _11089_, _06045_);
  and (_17699_, _17698_, _11120_);
  and (_17700_, _17699_, _17697_);
  and (_17701_, _07343_, _05970_);
  or (_17702_, _11143_, _11142_);
  nor (_17703_, _11144_, _11120_);
  and (_17704_, _17703_, _17702_);
  or (_17705_, _17704_, _17701_);
  or (_17706_, _17705_, _17700_);
  not (_17707_, _07013_);
  nor (_17708_, _11186_, _11185_);
  nor (_17709_, _17708_, _11187_);
  and (_17710_, _17709_, _17707_);
  or (_17711_, _17710_, _11165_);
  and (_17712_, _17711_, _17706_);
  and (_17713_, _17709_, _07013_);
  or (_17714_, _17713_, _12094_);
  or (_17715_, _17714_, _17712_);
  nor (_17716_, _11225_, _11224_);
  nor (_17717_, _17716_, _11226_);
  or (_17718_, _17717_, _06308_);
  nor (_17719_, _11261_, _11260_);
  nor (_17720_, _17719_, _11262_);
  or (_17721_, _17720_, _14289_);
  and (_17722_, _17721_, _12968_);
  and (_17723_, _17722_, _17718_);
  and (_17724_, _17723_, _17715_);
  and (_17725_, _11243_, \uc8051golden_1.ACC [0]);
  or (_17726_, _17725_, _06606_);
  or (_17727_, _17726_, _17724_);
  or (_17728_, _17501_, _07037_);
  and (_17729_, _17728_, _11286_);
  and (_17730_, _17729_, _17727_);
  nor (_17731_, \uc8051golden_1.ACC [1], \uc8051golden_1.ACC [0]);
  nor (_17732_, _11316_, _17731_);
  nor (_17733_, _17732_, _11286_);
  or (_17734_, _17733_, _17730_);
  or (_17735_, _17734_, _11290_);
  nand (_17736_, _11290_, _10195_);
  and (_17737_, _17736_, _06807_);
  and (_17738_, _17737_, _17735_);
  and (_17739_, _17529_, _06234_);
  or (_17740_, _17739_, _06195_);
  or (_17741_, _17740_, _17738_);
  or (_17742_, _17499_, _17472_);
  or (_17743_, _17742_, _06196_);
  and (_17744_, _17743_, _11309_);
  and (_17745_, _17744_, _17741_);
  and (_17746_, _17732_, _11308_);
  or (_17747_, _17746_, _11315_);
  or (_17748_, _17747_, _17745_);
  nand (_17749_, _11315_, _10195_);
  and (_17750_, _17749_, _01375_);
  and (_17751_, _17750_, _17748_);
  or (_17752_, _17751_, _17459_);
  and (_42898_, _17752_, _42545_);
  nor (_17753_, _01375_, _10195_);
  nand (_17754_, _11243_, _05984_);
  or (_17755_, _11228_, _11221_);
  nor (_17756_, _11229_, _06308_);
  and (_17757_, _17756_, _17755_);
  and (_17758_, _07632_, _05970_);
  nor (_17759_, _10738_, _07009_);
  nor (_17760_, _11146_, _11139_);
  nor (_17761_, _17760_, _11147_);
  and (_17762_, _17761_, _17759_);
  nand (_17763_, _11017_, _11256_);
  and (_17764_, _11002_, _05955_);
  and (_17765_, _17764_, _11137_);
  or (_17766_, _10964_, _11257_);
  nand (_17767_, _06693_, _05982_);
  nor (_17768_, _07995_, _10195_);
  nor (_17769_, _10568_, _07623_);
  or (_17770_, _17769_, _17768_);
  or (_17771_, _17770_, _06293_);
  nor (_17772_, _17567_, _14117_);
  nor (_17773_, _11257_, _17772_);
  and (_17774_, _11257_, _17772_);
  nor (_17775_, _17774_, _17773_);
  nand (_17776_, _17565_, _17775_);
  or (_17777_, _17565_, _17775_);
  and (_17778_, _17777_, _17776_);
  or (_17779_, _17778_, _10573_);
  nand (_17780_, _10644_, _07623_);
  or (_17781_, _17249_, _09444_);
  nor (_17782_, _10664_, _07623_);
  or (_17783_, _06854_, \uc8051golden_1.ACC [2]);
  nand (_17784_, _06854_, \uc8051golden_1.ACC [2]);
  nand (_17785_, _17784_, _17783_);
  nor (_17786_, _17785_, _10663_);
  or (_17787_, _17786_, _10654_);
  or (_17788_, _17787_, _17782_);
  and (_17789_, _17788_, _06002_);
  or (_17790_, _17789_, _07212_);
  and (_17791_, _17790_, _07210_);
  and (_17792_, _17791_, _17781_);
  and (_17793_, _14754_, _07995_);
  or (_17794_, _17793_, _17768_);
  and (_17795_, _17794_, _06401_);
  or (_17796_, _17795_, _10677_);
  or (_17797_, _17796_, _17792_);
  nor (_17798_, _17506_, _10195_);
  and (_17799_, _10681_, \uc8051golden_1.PSW [6]);
  nor (_17800_, _17799_, _17798_);
  nand (_17801_, _17800_, _10677_);
  and (_17802_, _17801_, _06407_);
  and (_17803_, _17802_, _17797_);
  nor (_17804_, _08616_, _10195_);
  and (_17805_, _14751_, _08616_);
  or (_17806_, _17805_, _17804_);
  and (_17807_, _17806_, _06395_);
  and (_17808_, _17770_, _06399_);
  or (_17809_, _17808_, _10644_);
  or (_17810_, _17809_, _17807_);
  or (_17811_, _17810_, _17803_);
  and (_17812_, _17811_, _17780_);
  or (_17813_, _17812_, _07233_);
  or (_17814_, _09444_, _10714_);
  and (_17815_, _17814_, _06414_);
  and (_17816_, _17815_, _17813_);
  nor (_17817_, _08432_, _06414_);
  or (_17818_, _17817_, _10642_);
  or (_17819_, _17818_, _17816_);
  nand (_17820_, _10642_, _10101_);
  and (_17821_, _17820_, _17819_);
  or (_17822_, _17821_, _06393_);
  and (_17823_, _14749_, _08616_);
  or (_17824_, _17823_, _17804_);
  or (_17825_, _17824_, _06844_);
  and (_17826_, _17825_, _07245_);
  and (_17827_, _17826_, _17822_);
  or (_17828_, _17804_, _14778_);
  and (_17829_, _17828_, _06387_);
  and (_17830_, _17829_, _17806_);
  or (_17831_, _17830_, _09538_);
  or (_17832_, _17831_, _17827_);
  nor (_17833_, _10002_, _10000_);
  or (_17834_, _17833_, _10003_);
  nand (_17835_, _17834_, _09538_);
  and (_17836_, _17835_, _10740_);
  and (_17837_, _17836_, _17832_);
  and (_17838_, _07196_, \uc8051golden_1.ACC [1]);
  and (_17839_, _07473_, _06045_);
  nor (_17840_, _17839_, _11142_);
  nor (_17841_, _17840_, _17838_);
  nor (_17842_, _11139_, _17841_);
  and (_17843_, _11139_, _17841_);
  nor (_17844_, _17843_, _17842_);
  nor (_17845_, _17228_, _11142_);
  and (_17846_, _17845_, \uc8051golden_1.PSW [7]);
  or (_17847_, _17846_, _17844_);
  nand (_17848_, _17846_, _17844_);
  and (_17849_, _17848_, _14157_);
  and (_17850_, _17849_, _17847_);
  or (_17851_, _17850_, _12586_);
  or (_17852_, _17851_, _17837_);
  and (_17853_, _09345_, \uc8051golden_1.ACC [1]);
  not (_17854_, _17853_);
  and (_17855_, _09446_, _06045_);
  or (_17856_, _17855_, _11185_);
  and (_17857_, _17856_, _17854_);
  nor (_17858_, _11180_, _17857_);
  and (_17859_, _11180_, _17857_);
  nor (_17860_, _17859_, _17858_);
  nor (_17861_, _17352_, _11185_);
  not (_17862_, _17861_);
  or (_17863_, _17862_, _17860_);
  and (_17864_, _17863_, \uc8051golden_1.PSW [7]);
  nor (_17865_, _17860_, \uc8051golden_1.PSW [7]);
  nor (_17866_, _17865_, _17864_);
  and (_17867_, _17862_, _17860_);
  or (_17868_, _17867_, _12587_);
  or (_17869_, _17868_, _17866_);
  and (_17870_, _17869_, _06442_);
  and (_17871_, _17870_, _17852_);
  and (_17872_, _08476_, \uc8051golden_1.ACC [1]);
  and (_17873_, _08521_, _06045_);
  nor (_17874_, _17873_, _14028_);
  nor (_17875_, _17874_, _17872_);
  nor (_17876_, _17875_, _11221_);
  and (_17877_, _17875_, _11221_);
  nor (_17878_, _17877_, _17876_);
  not (_17879_, _17878_);
  and (_17880_, _12540_, \uc8051golden_1.PSW [7]);
  or (_17881_, _17880_, _17879_);
  nand (_17882_, _17880_, _17879_);
  nand (_17883_, _17882_, _17881_);
  and (_17884_, _17883_, _06437_);
  or (_17885_, _17884_, _10572_);
  or (_17886_, _17885_, _17871_);
  and (_17887_, _17886_, _17779_);
  or (_17888_, _17887_, _06022_);
  nand (_17889_, _06693_, _06022_);
  and (_17890_, _17889_, _06446_);
  and (_17891_, _17890_, _17888_);
  and (_17892_, _14793_, _08616_);
  or (_17893_, _17892_, _17804_);
  and (_17894_, _17893_, _06300_);
  or (_17895_, _17894_, _10059_);
  or (_17896_, _17895_, _17891_);
  and (_17897_, _17896_, _17771_);
  or (_17898_, _17897_, _06281_);
  and (_17899_, _07995_, _09444_);
  or (_17900_, _17768_, _06282_);
  or (_17901_, _17900_, _17899_);
  and (_17902_, _17901_, _06279_);
  and (_17903_, _17902_, _17898_);
  and (_17904_, _14848_, _07995_);
  or (_17905_, _17904_, _17768_);
  and (_17906_, _17905_, _06015_);
  or (_17907_, _17906_, _10072_);
  or (_17908_, _17907_, _17903_);
  or (_17909_, _10264_, _10078_);
  and (_17910_, _17909_, _17908_);
  or (_17911_, _17910_, _05982_);
  and (_17912_, _17911_, _17767_);
  or (_17913_, _17912_, _06275_);
  and (_17914_, _07995_, _08994_);
  or (_17915_, _17914_, _17768_);
  or (_17916_, _17915_, _06276_);
  and (_17917_, _17916_, _10934_);
  and (_17918_, _17917_, _17913_);
  nor (_17919_, _10934_, _06693_);
  or (_17920_, _17919_, _10941_);
  or (_17921_, _17920_, _17918_);
  or (_17922_, _10945_, _11139_);
  and (_17923_, _17922_, _17236_);
  and (_17924_, _17923_, _17921_);
  and (_17925_, _17237_, _11139_);
  or (_17926_, _17925_, _10953_);
  or (_17927_, _17926_, _17924_);
  or (_17928_, _10959_, _11180_);
  and (_17929_, _17928_, _06581_);
  and (_17930_, _17929_, _17927_);
  or (_17931_, _10963_, _11221_);
  and (_17932_, _17931_, _12228_);
  or (_17933_, _17932_, _17930_);
  and (_17934_, _17933_, _17766_);
  or (_17935_, _17934_, _06474_);
  and (_17936_, _14744_, _07995_);
  or (_17937_, _17936_, _17768_);
  or (_17938_, _17937_, _07282_);
  and (_17939_, _17938_, _07284_);
  and (_17940_, _17939_, _17935_);
  and (_17941_, _17768_, _06582_);
  or (_17942_, _17941_, _17471_);
  or (_17943_, _17942_, _17940_);
  nor (_17944_, _12715_, _11137_);
  nor (_17945_, _17944_, _17764_);
  and (_17946_, _17945_, _17943_);
  nor (_17947_, _17946_, _17765_);
  nor (_17948_, _17947_, _06970_);
  and (_17949_, _11137_, _06970_);
  or (_17950_, _17949_, _17948_);
  and (_17951_, _17950_, _10560_);
  and (_17952_, _11178_, _10559_);
  or (_17953_, _17952_, _06567_);
  or (_17954_, _17953_, _17951_);
  or (_17955_, _11219_, _06568_);
  and (_17956_, _17955_, _10990_);
  and (_17957_, _17956_, _17954_);
  and (_17958_, _10989_, _11255_);
  or (_17959_, _17958_, _17957_);
  and (_17960_, _17959_, _07279_);
  nand (_17962_, _17915_, _06478_);
  nor (_17963_, _17962_, _11220_);
  or (_17964_, _17963_, _06784_);
  or (_17965_, _17964_, _17960_);
  nand (_17966_, _11138_, _06784_);
  nor (_17967_, _17659_, _07095_);
  and (_17968_, _17967_, _17966_);
  and (_17969_, _17968_, _17965_);
  nor (_17970_, _17967_, _11138_);
  or (_17971_, _17970_, _11011_);
  or (_17972_, _17971_, _17969_);
  nand (_17973_, _11011_, _11179_);
  and (_17974_, _17973_, _06575_);
  and (_17975_, _17974_, _17972_);
  nand (_17976_, _11020_, _11220_);
  and (_17977_, _17976_, _11019_);
  or (_17978_, _17977_, _17975_);
  and (_17979_, _17978_, _17763_);
  or (_17980_, _17979_, _06479_);
  and (_17981_, _14741_, _07995_);
  or (_17982_, _17768_, _09043_);
  or (_17983_, _17982_, _17981_);
  and (_17984_, _17983_, _11028_);
  and (_17985_, _17984_, _17980_);
  nand (_17986_, _11041_, _10780_);
  nor (_17987_, _11042_, _11028_);
  and (_17988_, _17987_, _17986_);
  or (_17989_, _17988_, _17463_);
  or (_17990_, _17989_, _17985_);
  and (_17991_, _10529_, _10515_);
  nor (_17992_, _17991_, _10530_);
  or (_17993_, _17992_, _17464_);
  and (_17994_, _17993_, _17687_);
  and (_17995_, _17994_, _17990_);
  and (_17996_, _17992_, _06984_);
  or (_17997_, _17996_, _06578_);
  or (_17998_, _17997_, _17995_);
  nand (_17999_, _11072_, _10614_);
  nor (_18000_, _11073_, _11059_);
  and (_18001_, _18000_, _17999_);
  or (_18002_, _18001_, _11060_);
  and (_18003_, _18002_, _17998_);
  and (_18004_, _11102_, _10879_);
  nor (_18005_, _18004_, _11103_);
  and (_18006_, _18005_, _11059_);
  or (_18007_, _18006_, _11089_);
  or (_18008_, _18007_, _18003_);
  and (_18009_, _11089_, _05984_);
  nor (_18010_, _18009_, _17759_);
  and (_18011_, _18010_, _18008_);
  nor (_18012_, _18011_, _17762_);
  nor (_18013_, _18012_, _17758_);
  and (_18014_, _17761_, _17758_);
  nor (_18015_, _18014_, _18013_);
  nor (_18016_, _18015_, _17701_);
  and (_18017_, _11188_, _11181_);
  nor (_18018_, _18017_, _11189_);
  and (_18019_, _18018_, _17701_);
  or (_18020_, _18019_, _07013_);
  or (_18021_, _18020_, _18016_);
  or (_18022_, _18018_, _17707_);
  and (_18023_, _18022_, _06308_);
  and (_18024_, _18023_, _18021_);
  or (_18025_, _18024_, _17757_);
  and (_18026_, _18025_, _14289_);
  or (_18027_, _11264_, _11257_);
  nor (_18028_, _11265_, _14289_);
  and (_18029_, _18028_, _18027_);
  or (_18030_, _18029_, _11243_);
  or (_18031_, _18030_, _18026_);
  and (_18032_, _18031_, _17754_);
  or (_18033_, _18032_, _06606_);
  or (_18034_, _17794_, _07037_);
  and (_18035_, _18034_, _11286_);
  and (_18036_, _18035_, _18033_);
  nor (_18037_, _17731_, _10195_);
  or (_18038_, _18037_, _11291_);
  nor (_18039_, _18038_, _11290_);
  nor (_18040_, _18039_, _12994_);
  or (_18041_, _18040_, _18036_);
  nand (_18042_, _11290_, _10246_);
  and (_18043_, _18042_, _06807_);
  and (_18044_, _18043_, _18041_);
  and (_18045_, _17824_, _06234_);
  or (_18046_, _18045_, _06195_);
  or (_18047_, _18046_, _18044_);
  and (_18048_, _14917_, _07995_);
  or (_18049_, _18048_, _17768_);
  or (_18050_, _18049_, _06196_);
  and (_18051_, _18050_, _11309_);
  and (_18052_, _18051_, _18047_);
  nor (_18053_, _11316_, \uc8051golden_1.ACC [2]);
  nor (_18054_, _18053_, _11317_);
  and (_18055_, _18054_, _11308_);
  or (_18056_, _18055_, _11315_);
  or (_18057_, _18056_, _18052_);
  nand (_18058_, _11315_, _10246_);
  and (_18059_, _18058_, _01375_);
  and (_18060_, _18059_, _18057_);
  or (_18061_, _18060_, _17753_);
  and (_42899_, _18061_, _42545_);
  nor (_18062_, _01375_, _10246_);
  nor (_18063_, _11135_, _11136_);
  nor (_18064_, _11148_, _18063_);
  and (_18065_, _11148_, _18063_);
  or (_18066_, _18065_, _18064_);
  or (_18067_, _18066_, _11120_);
  and (_18068_, _11043_, _10774_);
  nor (_18069_, _18068_, _11044_);
  or (_18070_, _18069_, _11028_);
  nand (_18071_, _11136_, _10556_);
  or (_18072_, _11217_, _06568_);
  and (_18073_, _18072_, _10990_);
  and (_18074_, _10983_, _11135_);
  or (_18075_, _12535_, _06581_);
  and (_18076_, _18075_, _10964_);
  nand (_18077_, _06372_, _05982_);
  nor (_18078_, _07995_, _10246_);
  nor (_18079_, _10568_, _07775_);
  or (_18080_, _18079_, _18078_);
  or (_18081_, _18080_, _06293_);
  and (_18082_, _12244_, \uc8051golden_1.PSW [7]);
  and (_18083_, _06693_, \uc8051golden_1.ACC [2]);
  nor (_18084_, _17773_, _18083_);
  nor (_18085_, _12239_, _18084_);
  and (_18086_, _12239_, _18084_);
  nor (_18087_, _18086_, _18085_);
  not (_18088_, _12243_);
  or (_18089_, _18088_, _17775_);
  or (_18090_, _18089_, _10524_);
  and (_18091_, _18090_, _18087_);
  or (_18092_, _18091_, _10573_);
  or (_18093_, _18092_, _18082_);
  nor (_18094_, _08616_, _10246_);
  and (_18095_, _14951_, _08616_);
  or (_18096_, _18095_, _18094_);
  or (_18097_, _18094_, _14968_);
  and (_18098_, _18097_, _06387_);
  and (_18099_, _18098_, _18096_);
  nand (_18100_, _10644_, _07775_);
  or (_18101_, _18096_, _06396_);
  and (_18102_, _18101_, _07221_);
  and (_18103_, _14947_, _07995_);
  or (_18104_, _18103_, _18078_);
  and (_18105_, _18104_, _06401_);
  nand (_18106_, _10663_, _07775_);
  nor (_18107_, _06854_, _10246_);
  and (_18108_, _06854_, _10246_);
  or (_18109_, _18108_, _18107_);
  or (_18110_, _18109_, _10663_);
  and (_18111_, _18110_, _10655_);
  and (_18112_, _18111_, _18106_);
  and (_18113_, _18112_, _08659_);
  or (_18114_, _18113_, _09443_);
  or (_18115_, _18112_, _10654_);
  and (_18116_, _18115_, _06002_);
  or (_18117_, _18116_, _07212_);
  and (_18118_, _18117_, _07210_);
  and (_18119_, _18118_, _18114_);
  or (_18120_, _18119_, _18105_);
  and (_18121_, _18120_, _10678_);
  not (_18122_, \uc8051golden_1.PSW [6]);
  nor (_18123_, _10681_, _18122_);
  nor (_18124_, _18123_, \uc8051golden_1.ACC [3]);
  nor (_18125_, _18124_, _10682_);
  and (_18126_, _18125_, _10677_);
  or (_18127_, _18126_, _06395_);
  or (_18128_, _18127_, _18121_);
  and (_18129_, _18128_, _18102_);
  and (_18130_, _18080_, _06399_);
  or (_18131_, _18130_, _10644_);
  or (_18132_, _18131_, _18129_);
  and (_18133_, _18132_, _18100_);
  or (_18134_, _18133_, _07233_);
  or (_18135_, _09443_, _10714_);
  and (_18136_, _18135_, _06414_);
  and (_18137_, _18136_, _18134_);
  nor (_18138_, _08388_, _06414_);
  or (_18139_, _18138_, _10642_);
  or (_18140_, _18139_, _18137_);
  nand (_18141_, _10642_, _08651_);
  and (_18142_, _18141_, _18140_);
  or (_18143_, _18142_, _06393_);
  and (_18144_, _14961_, _08616_);
  or (_18145_, _18144_, _18094_);
  or (_18146_, _18145_, _06844_);
  and (_18147_, _18146_, _07245_);
  and (_18148_, _18147_, _18143_);
  or (_18149_, _18148_, _18099_);
  and (_18150_, _18149_, _09544_);
  or (_18151_, _10005_, _10003_);
  nor (_18152_, _10006_, _09544_);
  and (_18153_, _18152_, _18151_);
  or (_18154_, _18153_, _10739_);
  or (_18155_, _18154_, _18150_);
  not (_18156_, _10737_);
  and (_18157_, _07623_, \uc8051golden_1.ACC [2]);
  nor (_18158_, _17842_, _18157_);
  nor (_18159_, _18063_, _18158_);
  and (_18160_, _18063_, _18158_);
  nor (_18161_, _18160_, _18159_);
  and (_18162_, _18161_, \uc8051golden_1.PSW [7]);
  nor (_18163_, _18161_, \uc8051golden_1.PSW [7]);
  nor (_18164_, _18163_, _18162_);
  and (_18165_, _17844_, \uc8051golden_1.PSW [7]);
  nor (_18166_, _17845_, _10524_);
  nor (_18167_, _18166_, _18165_);
  not (_18168_, _18167_);
  and (_18169_, _18168_, _18164_);
  nor (_18170_, _18168_, _18164_);
  nor (_18171_, _18170_, _18169_);
  and (_18172_, _18171_, _18156_);
  or (_18173_, _18172_, _10740_);
  and (_18174_, _18173_, _18155_);
  and (_18175_, _18171_, _10737_);
  or (_18176_, _18175_, _12586_);
  or (_18177_, _18176_, _18174_);
  and (_18178_, _09300_, \uc8051golden_1.ACC [2]);
  nor (_18179_, _17858_, _18178_);
  nor (_18180_, _11176_, _11177_);
  not (_18181_, _18180_);
  nand (_18182_, _18181_, _18179_);
  or (_18183_, _18181_, _18179_);
  and (_18184_, _18183_, _18182_);
  or (_18185_, _18184_, _10524_);
  nand (_18186_, _18184_, _10524_);
  and (_18187_, _18186_, _18185_);
  nand (_18188_, _18187_, _17864_);
  or (_18189_, _18187_, _17864_);
  and (_18190_, _18189_, _18188_);
  or (_18191_, _18190_, _12587_);
  and (_18192_, _18191_, _06442_);
  and (_18193_, _18192_, _18177_);
  and (_18194_, _12541_, \uc8051golden_1.PSW [7]);
  and (_18195_, _08432_, \uc8051golden_1.ACC [2]);
  nor (_18196_, _17876_, _18195_);
  nor (_18197_, _12535_, _18196_);
  and (_18198_, _12535_, _18196_);
  nor (_18199_, _18198_, _18197_);
  and (_18200_, _17882_, _18199_);
  or (_18201_, _18200_, _10572_);
  or (_18202_, _18201_, _18194_);
  and (_18203_, _18202_, _12593_);
  or (_18204_, _18203_, _18193_);
  and (_18205_, _18204_, _18093_);
  or (_18206_, _18205_, _06022_);
  nand (_18207_, _06372_, _06022_);
  and (_18208_, _18207_, _06446_);
  and (_18209_, _18208_, _18206_);
  and (_18210_, _14985_, _08616_);
  or (_18211_, _18210_, _18094_);
  and (_18212_, _18211_, _06300_);
  or (_18213_, _18212_, _10059_);
  or (_18214_, _18213_, _18209_);
  and (_18215_, _18214_, _18081_);
  or (_18216_, _18215_, _06281_);
  and (_18217_, _07995_, _09443_);
  or (_18218_, _18078_, _06282_);
  or (_18219_, _18218_, _18217_);
  and (_18220_, _18219_, _06279_);
  and (_18221_, _18220_, _18216_);
  and (_18222_, _15039_, _07995_);
  or (_18223_, _18222_, _18078_);
  and (_18224_, _18223_, _06015_);
  or (_18225_, _18224_, _10072_);
  or (_18226_, _18225_, _18221_);
  or (_18227_, _10215_, _10078_);
  and (_18228_, _18227_, _18226_);
  or (_18229_, _18228_, _05982_);
  and (_18230_, _18229_, _18077_);
  or (_18231_, _18230_, _06275_);
  and (_18232_, _07995_, _08815_);
  or (_18233_, _18232_, _18078_);
  or (_18234_, _18233_, _06276_);
  and (_18235_, _18234_, _10934_);
  and (_18236_, _18235_, _18231_);
  or (_18237_, _10934_, _06372_);
  not (_18238_, _07104_);
  nor (_18239_, _10941_, _06958_);
  and (_18240_, _18239_, _18238_);
  nand (_18241_, _18240_, _18237_);
  or (_18242_, _18241_, _18236_);
  and (_18243_, _07632_, _05951_);
  not (_18244_, _18243_);
  or (_18245_, _18240_, _18063_);
  and (_18246_, _18245_, _18244_);
  and (_18247_, _18246_, _18242_);
  and (_18248_, _18243_, _18063_);
  or (_18249_, _18248_, _18247_);
  and (_18250_, _18249_, _10959_);
  and (_18251_, _10953_, _18180_);
  or (_18252_, _18251_, _06580_);
  or (_18253_, _18252_, _18250_);
  and (_18254_, _18253_, _18076_);
  and (_18255_, _10963_, _12239_);
  or (_18256_, _18255_, _06474_);
  or (_18257_, _18256_, _18254_);
  and (_18258_, _14934_, _07995_);
  or (_18259_, _18258_, _18078_);
  or (_18260_, _18259_, _07282_);
  and (_18261_, _18260_, _18257_);
  or (_18262_, _18261_, _06582_);
  or (_18263_, _18078_, _07284_);
  and (_18264_, _18263_, _10980_);
  and (_18265_, _18264_, _18262_);
  or (_18266_, _18265_, _18074_);
  and (_18267_, _18266_, _10560_);
  and (_18268_, _11176_, _10559_);
  or (_18269_, _18268_, _06567_);
  or (_18270_, _18269_, _18267_);
  and (_18271_, _18270_, _18073_);
  and (_18272_, _10989_, _11253_);
  or (_18273_, _18272_, _18271_);
  and (_18274_, _18273_, _07279_);
  nand (_18275_, _18233_, _06478_);
  nor (_18276_, _18275_, _11218_);
  or (_18277_, _18276_, _10556_);
  or (_18278_, _18277_, _18274_);
  and (_18279_, _18278_, _18071_);
  or (_18280_, _18279_, _11003_);
  nand (_18281_, _11003_, _11136_);
  and (_18282_, _18281_, _11006_);
  and (_18283_, _18282_, _18280_);
  nor (_18284_, _11136_, _11006_);
  or (_18285_, _18284_, _11011_);
  or (_18286_, _18285_, _18283_);
  nand (_18287_, _11011_, _11177_);
  and (_18288_, _18287_, _06575_);
  and (_18289_, _18288_, _18286_);
  nand (_18290_, _11020_, _11218_);
  and (_18291_, _18290_, _11019_);
  or (_18292_, _18291_, _18289_);
  nand (_18293_, _11017_, _11254_);
  and (_18294_, _18293_, _09043_);
  and (_18295_, _18294_, _18292_);
  and (_18296_, _14931_, _07995_);
  or (_18297_, _18296_, _18078_);
  and (_18298_, _18297_, _06479_);
  or (_18299_, _18298_, _11030_);
  or (_18300_, _18299_, _18295_);
  and (_18301_, _18300_, _18070_);
  or (_18302_, _18301_, _10471_);
  and (_18303_, _10531_, _10508_);
  nor (_18304_, _18303_, _10532_);
  or (_18305_, _18304_, _10472_);
  and (_18306_, _18305_, _06579_);
  and (_18307_, _18306_, _18302_);
  nand (_18308_, _11074_, _10609_);
  nor (_18309_, _11075_, _06579_);
  and (_18310_, _18309_, _18308_);
  or (_18311_, _18310_, _11059_);
  or (_18312_, _18311_, _18307_);
  and (_18313_, _11104_, _10874_);
  nor (_18314_, _18313_, _11105_);
  or (_18315_, _18314_, _11091_);
  and (_18316_, _18315_, _11090_);
  and (_18317_, _18316_, _18312_);
  and (_18318_, _11089_, \uc8051golden_1.ACC [2]);
  or (_18319_, _18318_, _11121_);
  or (_18320_, _18319_, _18317_);
  and (_18321_, _18320_, _18067_);
  or (_18322_, _18321_, _11163_);
  and (_18323_, _11190_, _18180_);
  nor (_18324_, _11190_, _18180_);
  or (_18325_, _18324_, _18323_);
  or (_18326_, _18325_, _11165_);
  and (_18327_, _18326_, _06308_);
  and (_18328_, _18327_, _18322_);
  nor (_18329_, _11230_, _12535_);
  and (_18330_, _11230_, _12535_);
  or (_18331_, _18330_, _18329_);
  and (_18332_, _18331_, _06307_);
  or (_18333_, _18332_, _11203_);
  or (_18334_, _18333_, _18328_);
  and (_18335_, _11266_, _12239_);
  nor (_18336_, _11266_, _12239_);
  or (_18337_, _18336_, _14289_);
  or (_18338_, _18337_, _18335_);
  and (_18339_, _18338_, _12968_);
  and (_18340_, _18339_, _18334_);
  and (_18341_, _11243_, \uc8051golden_1.ACC [2]);
  or (_18342_, _18341_, _06606_);
  or (_18343_, _18342_, _18340_);
  or (_18344_, _18104_, _07037_);
  and (_18345_, _18344_, _11286_);
  and (_18346_, _18345_, _18343_);
  nor (_18347_, _11291_, _10246_);
  or (_18348_, _18347_, _11292_);
  nor (_18349_, _18348_, _11290_);
  nor (_18350_, _18349_, _12994_);
  or (_18351_, _18350_, _18346_);
  nand (_18352_, _11290_, _10119_);
  and (_18353_, _18352_, _06807_);
  and (_18354_, _18353_, _18351_);
  and (_18355_, _18145_, _06234_);
  or (_18356_, _18355_, _06195_);
  or (_18357_, _18356_, _18354_);
  and (_18358_, _15113_, _07995_);
  or (_18359_, _18358_, _18078_);
  or (_18360_, _18359_, _06196_);
  and (_18361_, _18360_, _11309_);
  and (_18362_, _18361_, _18357_);
  nor (_18363_, _11317_, \uc8051golden_1.ACC [3]);
  nor (_18364_, _18363_, _11318_);
  and (_18365_, _18364_, _11308_);
  or (_18366_, _18365_, _11315_);
  or (_18367_, _18366_, _18362_);
  nand (_18368_, _11315_, _10119_);
  and (_18369_, _18368_, _01375_);
  and (_18370_, _18369_, _18367_);
  or (_18371_, _18370_, _18062_);
  and (_42900_, _18371_, _42545_);
  nor (_18372_, _01375_, _10119_);
  nand (_18373_, _11243_, _10246_);
  or (_18374_, _11232_, _11216_);
  and (_18375_, _18374_, _11233_);
  or (_18376_, _18375_, _06308_);
  and (_18377_, _18376_, _14289_);
  or (_18378_, _11076_, _10603_);
  and (_18379_, _18378_, _11077_);
  or (_18380_, _18379_, _06579_);
  and (_18381_, _18380_, _11091_);
  nand (_18382_, _11017_, _11251_);
  and (_18383_, _10983_, _11131_);
  nand (_18384_, _06265_, _05982_);
  nor (_18385_, _07995_, _10119_);
  nor (_18386_, _10568_, _08301_);
  or (_18387_, _18386_, _18385_);
  or (_18388_, _18387_, _06293_);
  nor (_18389_, _12541_, _10524_);
  or (_18390_, _18196_, _14024_);
  and (_18391_, _18390_, _14023_);
  nor (_18392_, _18391_, _11216_);
  and (_18393_, _18391_, _11216_);
  nor (_18394_, _18393_, _18392_);
  and (_18395_, _18394_, \uc8051golden_1.PSW [7]);
  nor (_18396_, _18394_, \uc8051golden_1.PSW [7]);
  nor (_18397_, _18396_, _18395_);
  and (_18398_, _18397_, _18389_);
  nor (_18399_, _18397_, _18389_);
  nor (_18400_, _18399_, _18398_);
  or (_18401_, _18400_, _06442_);
  and (_18402_, _18401_, _10573_);
  or (_18403_, _18169_, _18162_);
  nor (_18404_, _07775_, \uc8051golden_1.ACC [3]);
  nand (_18405_, _07775_, \uc8051golden_1.ACC [3]);
  and (_18406_, _18405_, _18158_);
  or (_18407_, _18406_, _18404_);
  nor (_18408_, _11134_, _18407_);
  and (_18409_, _11134_, _18407_);
  nor (_18410_, _18409_, _18408_);
  and (_18411_, _18410_, \uc8051golden_1.PSW [7]);
  nor (_18412_, _18410_, \uc8051golden_1.PSW [7]);
  nor (_18413_, _18412_, _18411_);
  or (_18414_, _18413_, _18403_);
  and (_18415_, _18413_, _18403_);
  nor (_18416_, _18415_, _10740_);
  and (_18417_, _18416_, _18414_);
  nand (_18418_, _10644_, _08301_);
  nor (_18419_, _08616_, _10119_);
  and (_18420_, _15139_, _08616_);
  or (_18421_, _18420_, _18419_);
  or (_18422_, _18421_, _06396_);
  and (_18423_, _18422_, _07221_);
  and (_18424_, _15130_, _07995_);
  or (_18425_, _18424_, _18385_);
  and (_18426_, _18425_, _06401_);
  or (_18427_, _10655_, _09442_);
  nor (_18428_, _10664_, _08301_);
  or (_18429_, _06854_, \uc8051golden_1.ACC [4]);
  nand (_18430_, _06854_, \uc8051golden_1.ACC [4]);
  nand (_18431_, _18430_, _18429_);
  nor (_18432_, _18431_, _10663_);
  or (_18433_, _18432_, _10654_);
  or (_18434_, _18433_, _18428_);
  and (_18435_, _18434_, _10673_);
  and (_18436_, _18435_, _18427_);
  or (_18437_, _18436_, _18426_);
  and (_18438_, _18437_, _10678_);
  nor (_18439_, _10682_, \uc8051golden_1.ACC [4]);
  nor (_18440_, _18439_, _10683_);
  and (_18441_, _18440_, _10677_);
  or (_18442_, _18441_, _06395_);
  or (_18443_, _18442_, _18438_);
  and (_18444_, _18443_, _18423_);
  and (_18445_, _18387_, _06399_);
  or (_18446_, _18445_, _10644_);
  or (_18447_, _18446_, _18444_);
  and (_18448_, _18447_, _18418_);
  or (_18449_, _18448_, _07233_);
  or (_18450_, _09442_, _10714_);
  and (_18451_, _18450_, _06414_);
  and (_18452_, _18451_, _18449_);
  nor (_18453_, _08344_, _06414_);
  or (_18454_, _18453_, _10642_);
  or (_18455_, _18454_, _18452_);
  nand (_18456_, _10642_, _06045_);
  and (_18457_, _18456_, _18455_);
  or (_18458_, _18457_, _06393_);
  and (_18459_, _15168_, _08616_);
  or (_18460_, _18459_, _18419_);
  or (_18461_, _18460_, _06844_);
  and (_18462_, _18461_, _07245_);
  and (_18463_, _18462_, _18458_);
  or (_18464_, _18419_, _15138_);
  and (_18465_, _18464_, _06387_);
  and (_18466_, _18465_, _18421_);
  or (_18467_, _18466_, _09538_);
  or (_18468_, _18467_, _18463_);
  nor (_18469_, _10008_, _10006_);
  nor (_18470_, _18469_, _10009_);
  or (_18471_, _18470_, _09544_);
  and (_18472_, _18471_, _10740_);
  and (_18473_, _18472_, _18468_);
  or (_18474_, _18473_, _18417_);
  and (_18475_, _18474_, _12587_);
  nand (_18476_, _18188_, _18185_);
  and (_18477_, _09443_, _10246_);
  or (_18478_, _09443_, _10246_);
  and (_18479_, _18478_, _18179_);
  or (_18480_, _18479_, _18477_);
  nor (_18481_, _11175_, _18480_);
  not (_18482_, _18481_);
  nand (_18483_, _11175_, _18480_);
  and (_18484_, _18483_, _18482_);
  nand (_18485_, _18484_, \uc8051golden_1.PSW [7]);
  or (_18486_, _18484_, \uc8051golden_1.PSW [7]);
  and (_18487_, _18486_, _18485_);
  or (_18488_, _18487_, _18476_);
  nand (_18489_, _18487_, _18476_);
  and (_18490_, _12586_, _18489_);
  and (_18491_, _18490_, _18488_);
  or (_18492_, _18491_, _06437_);
  or (_18493_, _18492_, _18475_);
  and (_18494_, _18493_, _18402_);
  nor (_18495_, _12244_, _10524_);
  or (_18496_, _18084_, _14123_);
  and (_18497_, _18496_, _14122_);
  nor (_18498_, _11252_, _18497_);
  and (_18499_, _11252_, _18497_);
  nor (_18500_, _18499_, _18498_);
  and (_18501_, _18500_, \uc8051golden_1.PSW [7]);
  nor (_18502_, _18500_, \uc8051golden_1.PSW [7]);
  nor (_18503_, _18502_, _18501_);
  or (_18504_, _18503_, _18495_);
  and (_18505_, _18503_, _18495_);
  nor (_18506_, _18505_, _10573_);
  and (_18507_, _18506_, _18504_);
  or (_18508_, _18507_, _06022_);
  or (_18509_, _18508_, _18494_);
  nand (_18510_, _06265_, _06022_);
  and (_18511_, _18510_, _06446_);
  and (_18512_, _18511_, _18509_);
  and (_18513_, _15189_, _08616_);
  or (_18514_, _18513_, _18419_);
  and (_18515_, _18514_, _06300_);
  or (_18516_, _18515_, _10059_);
  or (_18517_, _18516_, _18512_);
  and (_18518_, _18517_, _18388_);
  or (_18519_, _18518_, _06281_);
  and (_18520_, _07995_, _09442_);
  or (_18521_, _18385_, _06282_);
  or (_18522_, _18521_, _18520_);
  and (_18523_, _18522_, _06279_);
  and (_18524_, _18523_, _18519_);
  and (_18525_, _15243_, _07995_);
  or (_18526_, _18525_, _18385_);
  and (_18527_, _18526_, _06015_);
  or (_18528_, _18527_, _10072_);
  or (_18529_, _18528_, _18524_);
  or (_18530_, _10163_, _10078_);
  and (_18531_, _18530_, _18529_);
  or (_18532_, _18531_, _05982_);
  and (_18533_, _18532_, _18384_);
  or (_18534_, _18533_, _06275_);
  and (_18535_, _08883_, _07995_);
  or (_18536_, _18535_, _18385_);
  or (_18537_, _18536_, _06276_);
  and (_18538_, _18537_, _10934_);
  and (_18539_, _18538_, _18534_);
  and (_18540_, _06451_, _05951_);
  nor (_18541_, _10934_, _06265_);
  or (_18542_, _18541_, _18540_);
  or (_18543_, _18542_, _18539_);
  not (_18544_, _06958_);
  and (_18545_, _06453_, _05951_);
  nor (_18546_, _18545_, _06961_);
  nand (_18547_, _18546_, _18544_);
  not (_18548_, _18547_);
  and (_18549_, _18548_, _11134_);
  or (_18550_, _18549_, _18239_);
  and (_18551_, _18550_, _18543_);
  and (_18552_, _18547_, _11134_);
  or (_18553_, _18552_, _07104_);
  or (_18554_, _18553_, _18551_);
  or (_18555_, _11134_, _18238_);
  and (_18556_, _18555_, _18244_);
  and (_18557_, _18556_, _18554_);
  and (_18558_, _18243_, _11134_);
  or (_18559_, _18558_, _10953_);
  or (_18560_, _18559_, _18557_);
  or (_18561_, _10959_, _11175_);
  and (_18562_, _18561_, _18560_);
  or (_18563_, _18562_, _06580_);
  or (_18564_, _11216_, _06581_);
  and (_18565_, _18564_, _10964_);
  and (_18566_, _18565_, _18563_);
  and (_18567_, _10963_, _11252_);
  or (_18568_, _18567_, _06474_);
  or (_18569_, _18568_, _18566_);
  and (_18570_, _15135_, _07995_);
  or (_18571_, _18570_, _18385_);
  or (_18572_, _18571_, _07282_);
  and (_18573_, _18572_, _18569_);
  or (_18574_, _18573_, _06582_);
  or (_18575_, _18385_, _07284_);
  and (_18576_, _18575_, _10980_);
  and (_18577_, _18576_, _18574_);
  or (_18578_, _18577_, _18383_);
  and (_18579_, _18578_, _10560_);
  and (_18580_, _11172_, _10559_);
  or (_18581_, _18580_, _06567_);
  or (_18582_, _18581_, _18579_);
  or (_18583_, _11213_, _06568_);
  and (_18584_, _18583_, _10990_);
  and (_18585_, _18584_, _18582_);
  and (_18586_, _10989_, _11249_);
  or (_18587_, _18586_, _18585_);
  and (_18588_, _18587_, _07279_);
  nand (_18589_, _18536_, _06478_);
  nor (_18590_, _18589_, _11215_);
  or (_18591_, _18590_, _06784_);
  or (_18592_, _18591_, _18588_);
  not (_18593_, _06784_);
  or (_18594_, _11133_, _18593_);
  and (_18595_, _18594_, _17468_);
  and (_18596_, _18595_, _18592_);
  and (_18597_, _11133_, _07095_);
  or (_18598_, _18597_, _18596_);
  and (_18599_, _18598_, _17660_);
  and (_18600_, _17659_, _11133_);
  or (_18601_, _18600_, _11011_);
  or (_18602_, _18601_, _18599_);
  or (_18603_, _17665_, _11174_);
  and (_18604_, _18603_, _06575_);
  and (_18605_, _18604_, _18602_);
  nand (_18606_, _11020_, _11215_);
  and (_18607_, _18606_, _11019_);
  or (_18608_, _18607_, _18605_);
  and (_18609_, _18608_, _18382_);
  or (_18610_, _18609_, _06479_);
  and (_18611_, _15134_, _07995_);
  or (_18612_, _18385_, _09043_);
  or (_18613_, _18612_, _18611_);
  and (_18614_, _18613_, _11028_);
  and (_18615_, _18614_, _18610_);
  or (_18616_, _11045_, _10767_);
  and (_18617_, _18616_, _11046_);
  and (_18618_, _18617_, _11030_);
  or (_18619_, _18618_, _17463_);
  or (_18620_, _18619_, _18615_);
  or (_18621_, _10533_, _10501_);
  and (_18622_, _18621_, _10534_);
  or (_18623_, _18622_, _17464_);
  and (_18624_, _18623_, _17687_);
  and (_18625_, _18624_, _18620_);
  and (_18626_, _18622_, _06984_);
  or (_18627_, _18626_, _06578_);
  or (_18628_, _18627_, _18625_);
  and (_18629_, _18628_, _18381_);
  or (_18630_, _11106_, _10868_);
  and (_18631_, _18630_, _11107_);
  and (_18632_, _18631_, _11059_);
  or (_18633_, _18632_, _11089_);
  or (_18634_, _18633_, _18629_);
  nand (_18635_, _11089_, _10246_);
  and (_18636_, _18635_, _11120_);
  and (_18637_, _18636_, _18634_);
  or (_18638_, _11150_, _11134_);
  nor (_18639_, _11151_, _11120_);
  and (_18640_, _18639_, _18638_);
  or (_18641_, _18640_, _17701_);
  or (_18642_, _18641_, _18637_);
  or (_18643_, _11192_, _11175_);
  and (_18644_, _18643_, _11193_);
  and (_18645_, _18644_, _17707_);
  or (_18646_, _18645_, _11165_);
  and (_18647_, _18646_, _18642_);
  and (_18648_, _18644_, _07013_);
  or (_18649_, _18648_, _06307_);
  or (_18650_, _18649_, _18647_);
  and (_18651_, _18650_, _18377_);
  or (_18652_, _11268_, _11252_);
  and (_18653_, _11269_, _11203_);
  and (_18654_, _18653_, _18652_);
  or (_18655_, _18654_, _11243_);
  or (_18656_, _18655_, _18651_);
  and (_18657_, _18656_, _18373_);
  or (_18658_, _18657_, _06606_);
  or (_18659_, _18425_, _07037_);
  and (_18660_, _18659_, _11286_);
  and (_18661_, _18660_, _18658_);
  nor (_18662_, _11292_, _10119_);
  or (_18663_, _18662_, _11293_);
  and (_18664_, _18663_, _11285_);
  or (_18665_, _18664_, _11290_);
  or (_18666_, _18665_, _18661_);
  nand (_18667_, _11290_, _10145_);
  and (_18668_, _18667_, _06807_);
  and (_18669_, _18668_, _18666_);
  and (_18670_, _18460_, _06234_);
  or (_18671_, _18670_, _06195_);
  or (_18672_, _18671_, _18669_);
  and (_18673_, _15315_, _07995_);
  or (_18674_, _18673_, _18385_);
  or (_18675_, _18674_, _06196_);
  and (_18676_, _18675_, _11309_);
  and (_18677_, _18676_, _18672_);
  nor (_18678_, _11318_, \uc8051golden_1.ACC [4]);
  nor (_18679_, _18678_, _11319_);
  and (_18680_, _18679_, _11308_);
  or (_18681_, _18680_, _11315_);
  or (_18682_, _18681_, _18677_);
  nand (_18683_, _11315_, _10145_);
  and (_18684_, _18683_, _01375_);
  and (_18685_, _18684_, _18682_);
  or (_18686_, _18685_, _18372_);
  and (_42901_, _18686_, _42545_);
  nor (_18687_, _01375_, _10145_);
  nor (_18688_, _11153_, _11130_);
  nor (_18689_, _18688_, _11154_);
  or (_18690_, _18689_, _11120_);
  and (_18691_, _11047_, _10760_);
  nor (_18692_, _18691_, _11048_);
  or (_18693_, _18692_, _11028_);
  nand (_18694_, _11129_, _10556_);
  or (_18695_, _11211_, _06568_);
  and (_18696_, _18695_, _10990_);
  nor (_18697_, _12229_, _06958_);
  and (_18698_, _18697_, _18238_);
  and (_18699_, _18546_, _06957_);
  and (_18700_, _18699_, _18698_);
  not (_18701_, _18700_);
  and (_18702_, _18701_, _11130_);
  nand (_18703_, _06650_, _05982_);
  nor (_18704_, _07995_, _10145_);
  nor (_18705_, _10568_, _08207_);
  or (_18706_, _18705_, _18704_);
  or (_18707_, _18706_, _06293_);
  nand (_18708_, _18489_, _18485_);
  and (_18709_, _09210_, \uc8051golden_1.ACC [4]);
  nor (_18710_, _18481_, _18709_);
  nor (_18711_, _11171_, _11170_);
  or (_18712_, _18711_, _18710_);
  nand (_18713_, _18711_, _18710_);
  and (_18714_, _18713_, _18712_);
  and (_18715_, _18714_, \uc8051golden_1.PSW [7]);
  nor (_18716_, _18714_, \uc8051golden_1.PSW [7]);
  nor (_18717_, _18716_, _18715_);
  or (_18718_, _18717_, _18708_);
  nand (_18719_, _18717_, _18708_);
  and (_18720_, _12586_, _18719_);
  and (_18721_, _18720_, _18718_);
  nor (_18722_, _08616_, _10145_);
  and (_18723_, _15341_, _08616_);
  or (_18724_, _18723_, _18722_);
  or (_18725_, _18722_, _15378_);
  and (_18726_, _18725_, _06387_);
  and (_18727_, _18726_, _18724_);
  nand (_18728_, _10644_, _08207_);
  or (_18729_, _10655_, _09441_);
  nor (_18730_, _10664_, _08207_);
  or (_18731_, _06854_, \uc8051golden_1.ACC [5]);
  nand (_18732_, _06854_, \uc8051golden_1.ACC [5]);
  nand (_18733_, _18732_, _18731_);
  nor (_18734_, _18733_, _10663_);
  or (_18735_, _18734_, _10654_);
  or (_18736_, _18735_, _18730_);
  and (_18737_, _18736_, _10673_);
  and (_18738_, _18737_, _18729_);
  and (_18739_, _15348_, _07995_);
  or (_18740_, _18739_, _18704_);
  and (_18741_, _18740_, _06401_);
  or (_18742_, _18741_, _10677_);
  or (_18743_, _18742_, _18738_);
  nor (_18744_, _10699_, _10690_);
  and (_18745_, _10699_, _10690_);
  or (_18746_, _18745_, _18744_);
  or (_18747_, _18746_, _10678_);
  and (_18748_, _18747_, _06407_);
  and (_18750_, _18748_, _18743_);
  and (_18751_, _18724_, _06395_);
  and (_18752_, _18706_, _06399_);
  or (_18753_, _18752_, _10644_);
  or (_18754_, _18753_, _18751_);
  or (_18755_, _18754_, _18750_);
  and (_18756_, _18755_, _18728_);
  or (_18757_, _18756_, _07233_);
  or (_18758_, _09441_, _10714_);
  and (_18759_, _18758_, _06414_);
  and (_18760_, _18759_, _18757_);
  nor (_18761_, _08255_, _06414_);
  or (_18762_, _18761_, _10642_);
  or (_18763_, _18762_, _18760_);
  nand (_18764_, _10642_, _05984_);
  and (_18765_, _18764_, _18763_);
  or (_18766_, _18765_, _06393_);
  and (_18767_, _15345_, _08616_);
  or (_18768_, _18767_, _18722_);
  or (_18769_, _18768_, _06844_);
  and (_18772_, _18769_, _07245_);
  and (_18773_, _18772_, _18766_);
  or (_18774_, _18773_, _18727_);
  and (_18775_, _18774_, _09544_);
  or (_18776_, _10011_, _10009_);
  nor (_18777_, _10012_, _09544_);
  and (_18778_, _18777_, _18776_);
  or (_18779_, _18778_, _14157_);
  or (_18780_, _18779_, _18775_);
  and (_18781_, _08301_, \uc8051golden_1.ACC [4]);
  nor (_18783_, _18408_, _18781_);
  nor (_18784_, _11130_, _18783_);
  and (_18785_, _11130_, _18783_);
  nor (_18786_, _18785_, _18784_);
  and (_18787_, _18786_, \uc8051golden_1.PSW [7]);
  nor (_18788_, _18786_, \uc8051golden_1.PSW [7]);
  nor (_18789_, _18788_, _18787_);
  nor (_18790_, _18415_, _18411_);
  not (_18791_, _18790_);
  and (_18792_, _18791_, _18789_);
  nor (_18794_, _18791_, _18789_);
  nor (_18795_, _18794_, _18792_);
  or (_18796_, _18795_, _10740_);
  and (_18797_, _18796_, _12587_);
  and (_18798_, _18797_, _18780_);
  or (_18799_, _18798_, _06437_);
  or (_18800_, _18799_, _18721_);
  and (_18801_, _08344_, \uc8051golden_1.ACC [4]);
  nor (_18802_, _18392_, _18801_);
  nor (_18803_, _12542_, _18802_);
  and (_18805_, _12542_, _18802_);
  nor (_18806_, _18805_, _18803_);
  and (_18807_, _18806_, \uc8051golden_1.PSW [7]);
  nor (_18808_, _18806_, \uc8051golden_1.PSW [7]);
  nor (_18809_, _18808_, _18807_);
  nor (_18810_, _18398_, _18395_);
  not (_18811_, _18810_);
  and (_18812_, _18811_, _18809_);
  nor (_18813_, _18811_, _18809_);
  nor (_18814_, _18813_, _18812_);
  or (_18816_, _18814_, _06442_);
  and (_18817_, _18816_, _10573_);
  and (_18818_, _18817_, _18800_);
  and (_18819_, _06265_, \uc8051golden_1.ACC [4]);
  nor (_18820_, _18498_, _18819_);
  nor (_18821_, _12245_, _18820_);
  and (_18822_, _12245_, _18820_);
  nor (_18823_, _18822_, _18821_);
  and (_18824_, _18823_, \uc8051golden_1.PSW [7]);
  nor (_18825_, _18823_, \uc8051golden_1.PSW [7]);
  nor (_18827_, _18825_, _18824_);
  nor (_18828_, _18505_, _18501_);
  not (_18829_, _18828_);
  and (_18830_, _18829_, _18827_);
  nor (_18831_, _18829_, _18827_);
  nor (_18832_, _18831_, _18830_);
  and (_18833_, _18832_, _10572_);
  or (_18834_, _18833_, _06022_);
  or (_18835_, _18834_, _18818_);
  nand (_18836_, _06650_, _06022_);
  and (_18838_, _18836_, _06446_);
  and (_18839_, _18838_, _18835_);
  or (_18840_, _18722_, _15342_);
  and (_18841_, _18840_, _06300_);
  and (_18842_, _18841_, _18724_);
  or (_18843_, _18842_, _10059_);
  or (_18844_, _18843_, _18839_);
  and (_18845_, _18844_, _18707_);
  or (_18846_, _18845_, _06281_);
  and (_18847_, _07995_, _09441_);
  or (_18849_, _18704_, _06282_);
  or (_18850_, _18849_, _18847_);
  and (_18851_, _18850_, _06279_);
  and (_18852_, _18851_, _18846_);
  and (_18853_, _15446_, _07995_);
  or (_18854_, _18853_, _18704_);
  and (_18855_, _18854_, _06015_);
  or (_18856_, _18855_, _10072_);
  or (_18857_, _18856_, _18852_);
  or (_18858_, _10133_, _10078_);
  and (_18860_, _18858_, _18857_);
  or (_18861_, _18860_, _05982_);
  and (_18862_, _18861_, _18703_);
  or (_18863_, _18862_, _06275_);
  and (_18864_, _08958_, _07995_);
  or (_18865_, _18864_, _18704_);
  or (_18866_, _18865_, _06276_);
  and (_18867_, _18866_, _10934_);
  and (_18868_, _18867_, _18863_);
  nor (_18869_, _10934_, _06650_);
  or (_18871_, _18869_, _18540_);
  or (_18872_, _18871_, _18868_);
  not (_18873_, _18540_);
  or (_18874_, _11130_, _18873_);
  and (_18875_, _18874_, _18700_);
  and (_18876_, _18875_, _18872_);
  nor (_18877_, _18876_, _18702_);
  nor (_18878_, _18877_, _06959_);
  and (_18879_, _11130_, _06959_);
  or (_18880_, _18879_, _18878_);
  and (_18882_, _18880_, _10959_);
  and (_18883_, _10953_, _18711_);
  or (_18884_, _18883_, _06580_);
  or (_18885_, _18884_, _18882_);
  or (_18886_, _12542_, _06581_);
  and (_18887_, _18886_, _10964_);
  and (_18888_, _18887_, _18885_);
  and (_18889_, _10963_, _12245_);
  or (_18890_, _18889_, _06474_);
  or (_18891_, _18890_, _18888_);
  and (_18893_, _15338_, _07995_);
  or (_18894_, _18893_, _18704_);
  or (_18895_, _18894_, _07282_);
  and (_18896_, _18895_, _18891_);
  or (_18897_, _18896_, _06582_);
  or (_18898_, _06291_, _12714_);
  or (_18899_, _18704_, _07284_);
  and (_18900_, _18899_, _18898_);
  and (_18901_, _18900_, _18897_);
  or (_18902_, _12716_, _11128_);
  and (_18904_, _18902_, _10983_);
  or (_18905_, _18904_, _18901_);
  not (_18906_, _12716_);
  or (_18907_, _18906_, _11128_);
  and (_18908_, _18907_, _10560_);
  and (_18909_, _18908_, _18905_);
  and (_18910_, _11170_, _10559_);
  or (_18911_, _18910_, _06567_);
  or (_18912_, _18911_, _18909_);
  and (_18913_, _18912_, _18696_);
  and (_18915_, _10989_, _11247_);
  or (_18916_, _18915_, _18913_);
  and (_18917_, _18916_, _07279_);
  nand (_18918_, _18865_, _06478_);
  nor (_18919_, _18918_, _11212_);
  or (_18920_, _18919_, _10556_);
  or (_18921_, _18920_, _18917_);
  and (_18922_, _18921_, _18694_);
  or (_18923_, _18922_, _11003_);
  nand (_18924_, _11003_, _11129_);
  and (_18925_, _18924_, _11006_);
  and (_18926_, _18925_, _18923_);
  nor (_18927_, _11129_, _11006_);
  or (_18928_, _18927_, _11011_);
  or (_18929_, _18928_, _18926_);
  nand (_18930_, _11011_, _11171_);
  and (_18931_, _18930_, _06575_);
  and (_18932_, _18931_, _18929_);
  nand (_18933_, _11020_, _11212_);
  and (_18934_, _18933_, _11019_);
  or (_18936_, _18934_, _18932_);
  nand (_18937_, _11017_, _11248_);
  and (_18938_, _18937_, _09043_);
  and (_18939_, _18938_, _18936_);
  and (_18940_, _15335_, _07995_);
  or (_18941_, _18940_, _18704_);
  and (_18942_, _18941_, _06479_);
  or (_18943_, _18942_, _11030_);
  or (_18944_, _18943_, _18939_);
  and (_18945_, _18944_, _18693_);
  or (_18947_, _18945_, _10471_);
  and (_18948_, _10535_, _10494_);
  nor (_18949_, _18948_, _10536_);
  or (_18950_, _18949_, _10472_);
  and (_18951_, _18950_, _06579_);
  and (_18952_, _18951_, _18947_);
  nand (_18953_, _11078_, _10600_);
  nor (_18954_, _11079_, _06579_);
  and (_18955_, _18954_, _18953_);
  or (_18956_, _18955_, _11059_);
  or (_18958_, _18956_, _18952_);
  and (_18959_, _11108_, _10865_);
  nor (_18960_, _18959_, _11109_);
  or (_18961_, _18960_, _11091_);
  and (_18962_, _18961_, _11090_);
  and (_18963_, _18962_, _18958_);
  and (_18964_, _11089_, \uc8051golden_1.ACC [4]);
  or (_18965_, _18964_, _11121_);
  or (_18966_, _18965_, _18963_);
  and (_18967_, _18966_, _18690_);
  or (_18969_, _18967_, _11163_);
  and (_18970_, _11194_, _18711_);
  nor (_18971_, _11194_, _18711_);
  or (_18972_, _18971_, _11165_);
  or (_18973_, _18972_, _18970_);
  and (_18974_, _18973_, _06308_);
  and (_18975_, _18974_, _18969_);
  and (_18976_, _11234_, _12542_);
  nor (_18977_, _11234_, _12542_);
  or (_18978_, _18977_, _11203_);
  or (_18980_, _18978_, _18976_);
  and (_18981_, _18980_, _12094_);
  or (_18982_, _18981_, _18975_);
  and (_18983_, _11270_, _12245_);
  nor (_18984_, _11270_, _12245_);
  or (_18985_, _18984_, _14289_);
  or (_18986_, _18985_, _18983_);
  and (_18987_, _18986_, _12968_);
  and (_18988_, _18987_, _18982_);
  and (_18989_, _11243_, \uc8051golden_1.ACC [4]);
  or (_18991_, _18989_, _06606_);
  or (_18992_, _18991_, _18988_);
  or (_18993_, _18740_, _07037_);
  and (_18994_, _18993_, _11286_);
  and (_18995_, _18994_, _18992_);
  nor (_18996_, _11293_, _10145_);
  or (_18997_, _18996_, _11294_);
  and (_18998_, _18997_, _11285_);
  or (_18999_, _18998_, _11290_);
  or (_19000_, _18999_, _18995_);
  nand (_19002_, _11290_, _10101_);
  and (_19003_, _19002_, _06807_);
  and (_19004_, _19003_, _19000_);
  and (_19005_, _18768_, _06234_);
  or (_19006_, _19005_, _06195_);
  or (_19007_, _19006_, _19004_);
  and (_19008_, _15509_, _07995_);
  or (_19009_, _19008_, _18704_);
  or (_19010_, _19009_, _06196_);
  and (_19011_, _19010_, _11309_);
  and (_19013_, _19011_, _19007_);
  nor (_19014_, _11319_, \uc8051golden_1.ACC [5]);
  nor (_19015_, _19014_, _11320_);
  and (_19016_, _19015_, _11308_);
  or (_19017_, _19016_, _11315_);
  or (_19018_, _19017_, _19013_);
  nand (_19019_, _11315_, _10101_);
  and (_19020_, _19019_, _01375_);
  and (_19021_, _19020_, _19018_);
  or (_19022_, _19021_, _18687_);
  and (_42902_, _19022_, _42545_);
  nor (_19024_, _01375_, _10101_);
  nand (_19025_, _11243_, _10145_);
  or (_19026_, _11236_, _11210_);
  and (_19027_, _19026_, _11237_);
  or (_19028_, _19027_, _06308_);
  and (_19029_, _19028_, _14289_);
  nor (_19030_, _11080_, _10633_);
  nor (_19031_, _19030_, _11081_);
  or (_19032_, _19031_, _06579_);
  and (_19034_, _19032_, _11091_);
  nand (_19035_, _11017_, _11245_);
  and (_19036_, _10983_, _11124_);
  nor (_19037_, _07995_, _10101_);
  and (_19038_, _15639_, _07995_);
  or (_19039_, _19038_, _19037_);
  and (_19040_, _19039_, _06015_);
  nor (_19041_, _10568_, _08118_);
  or (_19042_, _19041_, _19037_);
  or (_19043_, _19042_, _06293_);
  nand (_19045_, _10644_, _08118_);
  or (_19046_, _10655_, _09440_);
  nor (_19047_, _10664_, _08118_);
  or (_19048_, _06854_, \uc8051golden_1.ACC [6]);
  nand (_19049_, _06854_, \uc8051golden_1.ACC [6]);
  nand (_19050_, _19049_, _19048_);
  nor (_19051_, _19050_, _10663_);
  or (_19052_, _19051_, _10654_);
  or (_19053_, _19052_, _19047_);
  and (_19054_, _19053_, _10673_);
  and (_19056_, _19054_, _19046_);
  and (_19057_, _15550_, _07995_);
  or (_19058_, _19057_, _19037_);
  and (_19059_, _19058_, _06401_);
  or (_19060_, _19059_, _10677_);
  or (_19061_, _19060_, _19056_);
  or (_19062_, _18744_, _10693_);
  nand (_19063_, _18744_, _10693_);
  and (_19064_, _19063_, _19062_);
  or (_19065_, _19064_, _10678_);
  and (_19067_, _19065_, _06407_);
  and (_19068_, _19067_, _19061_);
  nor (_19069_, _08616_, _10101_);
  and (_19070_, _15535_, _08616_);
  or (_19071_, _19070_, _19069_);
  and (_19072_, _19071_, _06395_);
  and (_19073_, _19042_, _06399_);
  or (_19074_, _19073_, _10644_);
  or (_19075_, _19074_, _19072_);
  or (_19076_, _19075_, _19068_);
  and (_19078_, _19076_, _19045_);
  or (_19079_, _19078_, _07233_);
  or (_19080_, _09440_, _10714_);
  and (_19081_, _19080_, _06414_);
  and (_19082_, _19081_, _19079_);
  nor (_19083_, _08161_, _06414_);
  or (_19084_, _19083_, _10642_);
  or (_19085_, _19084_, _19082_);
  nand (_19086_, _10642_, _10195_);
  and (_19087_, _19086_, _19085_);
  or (_19089_, _19087_, _06393_);
  and (_19090_, _15561_, _08616_);
  or (_19091_, _19090_, _19069_);
  or (_19092_, _19091_, _06844_);
  and (_19093_, _19092_, _07245_);
  and (_19094_, _19093_, _19089_);
  or (_19095_, _19069_, _15568_);
  and (_19096_, _19071_, _06387_);
  and (_19097_, _19096_, _19095_);
  or (_19098_, _19097_, _09538_);
  or (_19100_, _19098_, _19094_);
  nor (_19101_, _10014_, _10012_);
  nor (_19102_, _19101_, _10015_);
  or (_19103_, _19102_, _09544_);
  and (_19104_, _19103_, _10740_);
  and (_19105_, _19104_, _19100_);
  nand (_19106_, _08207_, \uc8051golden_1.ACC [5]);
  nor (_19107_, _08207_, \uc8051golden_1.ACC [5]);
  or (_19108_, _18783_, _19107_);
  and (_19109_, _19108_, _19106_);
  nor (_19111_, _19109_, _11127_);
  and (_19112_, _19109_, _11127_);
  nor (_19113_, _19112_, _19111_);
  nor (_19114_, _18792_, _18787_);
  and (_19115_, _19114_, \uc8051golden_1.PSW [7]);
  or (_19116_, _19115_, _19113_);
  nand (_19117_, _19115_, _19113_);
  and (_19118_, _19117_, _19116_);
  and (_19119_, _19118_, _14157_);
  or (_19120_, _19119_, _19105_);
  and (_19122_, _19120_, _12587_);
  or (_19123_, _09441_, _10145_);
  and (_19124_, _09441_, _10145_);
  or (_19125_, _18710_, _19124_);
  and (_19126_, _19125_, _19123_);
  nor (_19127_, _19126_, _11169_);
  and (_19128_, _19126_, _11169_);
  nor (_19129_, _19128_, _19127_);
  or (_19130_, _18714_, _10524_);
  nor (_19131_, _18708_, _19130_);
  or (_19133_, _19131_, _19129_);
  nand (_19134_, _19131_, _19129_);
  and (_19135_, _19134_, _12586_);
  and (_19136_, _19135_, _19133_);
  or (_19137_, _19136_, _19122_);
  or (_19138_, _19137_, _06437_);
  or (_19139_, _18802_, _14036_);
  and (_19140_, _19139_, _14035_);
  nor (_19141_, _19140_, _11210_);
  and (_19142_, _19140_, _11210_);
  nor (_19144_, _19142_, _19141_);
  nor (_19145_, _18812_, _18807_);
  and (_19146_, _19145_, \uc8051golden_1.PSW [7]);
  not (_19147_, _19146_);
  nor (_19148_, _19147_, _19144_);
  and (_19149_, _19147_, _19144_);
  or (_19150_, _19149_, _19148_);
  or (_19151_, _19150_, _06442_);
  and (_19152_, _19151_, _10573_);
  and (_19153_, _19152_, _19138_);
  or (_19155_, _18820_, _14130_);
  and (_19156_, _19155_, _14129_);
  nor (_19157_, _19156_, _11246_);
  and (_19158_, _19156_, _11246_);
  nor (_19159_, _19158_, _19157_);
  nor (_19160_, _18830_, _18824_);
  and (_19161_, _19160_, \uc8051golden_1.PSW [7]);
  nand (_19162_, _19161_, _19159_);
  or (_19163_, _19161_, _19159_);
  and (_19164_, _19163_, _10572_);
  and (_19166_, _19164_, _19162_);
  or (_19167_, _19166_, _06022_);
  or (_19168_, _19167_, _19153_);
  nand (_19169_, _06340_, _06022_);
  and (_19170_, _19169_, _06446_);
  and (_19171_, _19170_, _19168_);
  and (_19172_, _15585_, _08616_);
  or (_19173_, _19172_, _19069_);
  and (_19174_, _19173_, _06300_);
  or (_19175_, _19174_, _10059_);
  or (_19177_, _19175_, _19171_);
  and (_19178_, _19177_, _19043_);
  or (_19179_, _19178_, _06281_);
  and (_19180_, _07995_, _09440_);
  or (_19181_, _19037_, _06282_);
  or (_19182_, _19181_, _19180_);
  and (_19183_, _19182_, _06279_);
  and (_19184_, _19183_, _19179_);
  or (_19185_, _19184_, _19040_);
  and (_19186_, _19185_, _12616_);
  nor (_19188_, _06340_, _06021_);
  not (_19189_, _10106_);
  or (_19190_, _19189_, _10102_);
  nor (_19191_, _19190_, _05981_);
  and (_19192_, _19191_, _10072_);
  or (_19193_, _19192_, _19188_);
  or (_19194_, _19193_, _19186_);
  and (_19195_, _19194_, _06276_);
  and (_19196_, _15646_, _07995_);
  nor (_19197_, _19196_, _19037_);
  nor (_19199_, _19197_, _06276_);
  or (_19200_, _19199_, _10933_);
  or (_19201_, _19200_, _19195_);
  and (_19202_, _06742_, _05951_);
  and (_19203_, _10933_, _06340_);
  nor (_19204_, _19203_, _19202_);
  and (_19205_, _19204_, _19201_);
  and (_19206_, _11127_, _19202_);
  or (_19207_, _19206_, _18545_);
  or (_19208_, _19207_, _19205_);
  not (_19210_, _18545_);
  or (_19211_, _11127_, _19210_);
  and (_19212_, _19211_, _10944_);
  and (_19213_, _19212_, _19208_);
  and (_19214_, _11127_, _10565_);
  nor (_19215_, _19214_, _19213_);
  or (_19216_, _19215_, _12229_);
  nand (_19217_, _12229_, _11127_);
  nand (_19218_, _19217_, _19216_);
  or (_19219_, _19218_, _06959_);
  and (_19221_, _10959_, _11127_);
  or (_19222_, _19221_, _12231_);
  and (_19223_, _19222_, _19219_);
  and (_19224_, _10953_, _11169_);
  or (_19225_, _19224_, _06580_);
  or (_19226_, _19225_, _19223_);
  or (_19227_, _11210_, _06581_);
  and (_19228_, _19227_, _10964_);
  and (_19229_, _19228_, _19226_);
  and (_19230_, _10963_, _11246_);
  or (_19232_, _19230_, _06474_);
  or (_19233_, _19232_, _19229_);
  and (_19234_, _15531_, _07995_);
  or (_19235_, _19234_, _19037_);
  or (_19236_, _19235_, _07282_);
  and (_19237_, _19236_, _19233_);
  or (_19238_, _19237_, _06582_);
  or (_19239_, _19037_, _07284_);
  and (_19240_, _19239_, _10980_);
  and (_19241_, _19240_, _19238_);
  or (_19243_, _19241_, _19036_);
  and (_19244_, _19243_, _10560_);
  and (_19245_, _11166_, _10559_);
  or (_19246_, _19245_, _06567_);
  or (_19247_, _19246_, _19244_);
  or (_19248_, _11207_, _06568_);
  and (_19249_, _19248_, _10990_);
  and (_19250_, _19249_, _19247_);
  and (_19251_, _10989_, _11244_);
  or (_19252_, _19251_, _19250_);
  nand (_19254_, _19252_, _07279_);
  or (_19255_, _19197_, _07279_);
  or (_19256_, _19255_, _11209_);
  and (_19257_, _19256_, _19254_);
  nor (_19258_, _19257_, _07106_);
  or (_19259_, _11126_, _17653_);
  nand (_19260_, _19259_, _17654_);
  or (_19261_, _19260_, _19258_);
  not (_19262_, _11126_);
  or (_19263_, _17654_, _19262_);
  and (_19265_, _19263_, _17660_);
  and (_19266_, _19265_, _19261_);
  nor (_19267_, _17660_, _11126_);
  or (_19268_, _19267_, _11011_);
  or (_19269_, _19268_, _19266_);
  or (_19270_, _17665_, _11168_);
  and (_19271_, _19270_, _06575_);
  and (_19272_, _19271_, _19269_);
  nand (_19273_, _11020_, _11209_);
  and (_19274_, _19273_, _11019_);
  or (_19276_, _19274_, _19272_);
  and (_19277_, _19276_, _19035_);
  or (_19278_, _19277_, _06479_);
  and (_19279_, _15528_, _07995_);
  or (_19280_, _19037_, _09043_);
  or (_19281_, _19280_, _19279_);
  and (_19282_, _19281_, _11028_);
  and (_19283_, _19282_, _19278_);
  or (_19284_, _11049_, _10804_);
  nor (_19285_, _11050_, _11028_);
  and (_19287_, _19285_, _19284_);
  or (_19288_, _19287_, _17463_);
  or (_19289_, _19288_, _19283_);
  or (_19290_, _10537_, _10487_);
  and (_19291_, _19290_, _10538_);
  or (_19292_, _19291_, _17464_);
  and (_19293_, _19292_, _17687_);
  and (_19294_, _19293_, _19289_);
  and (_19295_, _19291_, _06984_);
  or (_19296_, _19295_, _06578_);
  or (_19298_, _19296_, _19294_);
  and (_19299_, _19298_, _19034_);
  or (_19300_, _11110_, _10899_);
  and (_19301_, _11111_, _11059_);
  and (_19302_, _19301_, _19300_);
  or (_19303_, _19302_, _11089_);
  or (_19304_, _19303_, _19299_);
  nand (_19305_, _11089_, _10145_);
  and (_19306_, _19305_, _11120_);
  and (_19307_, _19306_, _19304_);
  or (_19309_, _11155_, _11127_);
  and (_19310_, _11156_, _11121_);
  and (_19311_, _19310_, _19309_);
  or (_19312_, _19311_, _17701_);
  or (_19313_, _19312_, _19307_);
  or (_19314_, _11196_, _11169_);
  and (_19315_, _19314_, _11197_);
  and (_19316_, _19315_, _17707_);
  or (_19317_, _19316_, _11165_);
  and (_19318_, _19317_, _19313_);
  and (_19320_, _19315_, _07013_);
  or (_19321_, _19320_, _06307_);
  or (_19322_, _19321_, _19318_);
  and (_19323_, _19322_, _19029_);
  or (_19324_, _11272_, _11246_);
  nor (_19325_, _11273_, _14289_);
  and (_19326_, _19325_, _19324_);
  or (_19327_, _19326_, _11243_);
  or (_19328_, _19327_, _19323_);
  and (_19329_, _19328_, _19025_);
  or (_19331_, _19329_, _06606_);
  or (_19332_, _19058_, _07037_);
  and (_19333_, _19332_, _11286_);
  and (_19334_, _19333_, _19331_);
  nor (_19335_, _11294_, _10101_);
  or (_19336_, _19335_, _11295_);
  and (_19337_, _19336_, _11285_);
  or (_19338_, _19337_, _11290_);
  or (_19339_, _19338_, _19334_);
  nand (_19340_, _11290_, _08651_);
  and (_19342_, _19340_, _06807_);
  and (_19343_, _19342_, _19339_);
  and (_19344_, _19091_, _06234_);
  or (_19345_, _19344_, _06195_);
  or (_19346_, _19345_, _19343_);
  and (_19347_, _15713_, _07995_);
  or (_19348_, _19347_, _19037_);
  or (_19349_, _19348_, _06196_);
  and (_19350_, _19349_, _11309_);
  and (_19351_, _19350_, _19346_);
  nor (_19353_, _11320_, \uc8051golden_1.ACC [6]);
  nor (_19354_, _19353_, _11321_);
  and (_19355_, _19354_, _11308_);
  or (_19356_, _19355_, _11315_);
  or (_19357_, _19356_, _19351_);
  nand (_19358_, _11315_, _08651_);
  and (_19359_, _19358_, _01375_);
  and (_19360_, _19359_, _19357_);
  or (_19361_, _19360_, _19024_);
  and (_42903_, _19361_, _42545_);
  not (_19363_, \uc8051golden_1.PCON [0]);
  nor (_19364_, _01375_, _19363_);
  nand (_19365_, _11225_, _08002_);
  nor (_19366_, _08002_, _19363_);
  nor (_19367_, _19366_, _07276_);
  nand (_19368_, _19367_, _19365_);
  and (_19369_, _08002_, _07473_);
  or (_19370_, _19369_, _19366_);
  or (_19371_, _19370_, _06293_);
  nor (_19372_, _08521_, _11332_);
  or (_19374_, _19372_, _19366_);
  or (_19375_, _19374_, _07210_);
  and (_19376_, _08002_, \uc8051golden_1.ACC [0]);
  or (_19377_, _19376_, _19366_);
  and (_19378_, _19377_, _07199_);
  nor (_19379_, _07199_, _19363_);
  or (_19380_, _19379_, _06401_);
  or (_19381_, _19380_, _19378_);
  and (_19382_, _19381_, _07221_);
  and (_19383_, _19382_, _19375_);
  and (_19385_, _19370_, _06399_);
  or (_19386_, _19385_, _19383_);
  and (_19387_, _19386_, _06414_);
  and (_19388_, _19377_, _06406_);
  or (_19389_, _19388_, _10059_);
  or (_19390_, _19389_, _19387_);
  and (_19391_, _19390_, _19371_);
  or (_19392_, _19391_, _06281_);
  and (_19393_, _08002_, _09446_);
  or (_19394_, _19366_, _06282_);
  or (_19396_, _19394_, _19393_);
  and (_19397_, _19396_, _19392_);
  or (_19398_, _19397_, _06015_);
  and (_19399_, _14426_, _08002_);
  or (_19400_, _19366_, _06279_);
  or (_19401_, _19400_, _19399_);
  and (_19402_, _19401_, _06276_);
  and (_19403_, _19402_, _19398_);
  and (_19404_, _08002_, _08817_);
  or (_19405_, _19404_, _19366_);
  and (_19407_, _19405_, _06275_);
  or (_19408_, _19407_, _06474_);
  or (_19409_, _19408_, _19403_);
  and (_19410_, _14324_, _08002_);
  or (_19411_, _19410_, _19366_);
  or (_19412_, _19411_, _07282_);
  and (_19413_, _19412_, _07284_);
  and (_19414_, _19413_, _19409_);
  nor (_19415_, _12538_, _11332_);
  or (_19416_, _19415_, _19366_);
  and (_19418_, _19365_, _06582_);
  and (_19419_, _19418_, _19416_);
  or (_19420_, _19419_, _19414_);
  and (_19421_, _19420_, _07279_);
  nand (_19422_, _19405_, _06478_);
  nor (_19423_, _19422_, _19372_);
  or (_19424_, _19423_, _06569_);
  or (_19425_, _19424_, _19421_);
  and (_19426_, _19425_, _19368_);
  or (_19427_, _19426_, _06479_);
  and (_19429_, _14320_, _08002_);
  or (_19430_, _19429_, _19366_);
  or (_19431_, _19430_, _09043_);
  and (_19432_, _19431_, _09048_);
  and (_19433_, _19432_, _19427_);
  not (_19434_, _06700_);
  and (_19435_, _19416_, _06572_);
  or (_19436_, _19435_, _19434_);
  or (_19437_, _19436_, _19433_);
  or (_19438_, _19374_, _06700_);
  and (_19440_, _19438_, _01375_);
  and (_19441_, _19440_, _19437_);
  or (_19442_, _19441_, _19364_);
  and (_42905_, _19442_, _42545_);
  not (_19443_, \uc8051golden_1.PCON [1]);
  nor (_19444_, _01375_, _19443_);
  nand (_19445_, _08002_, _07090_);
  or (_19446_, _08002_, \uc8051golden_1.PCON [1]);
  and (_19447_, _19446_, _06275_);
  and (_19448_, _19447_, _19445_);
  and (_19450_, _08002_, _09445_);
  nor (_19451_, _08002_, _19443_);
  or (_19452_, _19451_, _06282_);
  or (_19453_, _19452_, _19450_);
  and (_19454_, _14532_, _08002_);
  not (_19455_, _19454_);
  and (_19456_, _19455_, _19446_);
  or (_19457_, _19456_, _07210_);
  and (_19458_, _08002_, \uc8051golden_1.ACC [1]);
  or (_19459_, _19458_, _19451_);
  and (_19461_, _19459_, _07199_);
  nor (_19462_, _07199_, _19443_);
  or (_19463_, _19462_, _06401_);
  or (_19464_, _19463_, _19461_);
  and (_19465_, _19464_, _07221_);
  and (_19466_, _19465_, _19457_);
  nor (_19467_, _11332_, _07196_);
  or (_19468_, _19467_, _19451_);
  and (_19469_, _19468_, _06399_);
  or (_19470_, _19469_, _19466_);
  and (_19472_, _19470_, _06414_);
  and (_19473_, _19459_, _06406_);
  or (_19474_, _19473_, _10059_);
  or (_19475_, _19474_, _19472_);
  or (_19476_, _19468_, _06293_);
  and (_19477_, _19476_, _19475_);
  or (_19478_, _19477_, _06281_);
  and (_19479_, _19478_, _06279_);
  and (_19480_, _19479_, _19453_);
  or (_19481_, _14615_, _11332_);
  and (_19483_, _19446_, _06015_);
  and (_19484_, _19483_, _19481_);
  or (_19485_, _19484_, _19480_);
  and (_19486_, _19485_, _06276_);
  or (_19487_, _19486_, _19448_);
  and (_19488_, _19487_, _07282_);
  or (_19489_, _14507_, _11332_);
  and (_19490_, _19446_, _06474_);
  and (_19491_, _19490_, _19489_);
  or (_19492_, _19491_, _06582_);
  or (_19494_, _19492_, _19488_);
  nor (_19495_, _11223_, _11332_);
  or (_19496_, _19495_, _19451_);
  nand (_19497_, _11222_, _08002_);
  and (_19498_, _19497_, _19496_);
  or (_19499_, _19498_, _07284_);
  and (_19500_, _19499_, _07279_);
  and (_19501_, _19500_, _19494_);
  or (_19502_, _14505_, _11332_);
  and (_19503_, _19446_, _06478_);
  and (_19505_, _19503_, _19502_);
  or (_19506_, _19505_, _06569_);
  or (_19507_, _19506_, _19501_);
  nor (_19508_, _19451_, _07276_);
  nand (_19509_, _19508_, _19497_);
  and (_19510_, _19509_, _09043_);
  and (_19511_, _19510_, _19507_);
  or (_19512_, _19445_, _08477_);
  and (_19513_, _19446_, _06479_);
  and (_19514_, _19513_, _19512_);
  or (_19516_, _19514_, _06572_);
  or (_19517_, _19516_, _19511_);
  or (_19518_, _19496_, _09048_);
  and (_19519_, _19518_, _07037_);
  and (_19520_, _19519_, _19517_);
  and (_19521_, _19456_, _06606_);
  or (_19522_, _19521_, _06195_);
  or (_19523_, _19522_, _19520_);
  or (_19524_, _19451_, _06196_);
  or (_19525_, _19524_, _19454_);
  and (_19527_, _19525_, _01375_);
  and (_19528_, _19527_, _19523_);
  or (_19529_, _19528_, _19444_);
  and (_42906_, _19529_, _42545_);
  not (_19530_, \uc8051golden_1.PCON [2]);
  nor (_19531_, _01375_, _19530_);
  and (_19532_, _08002_, _09444_);
  nor (_19533_, _08002_, _19530_);
  or (_19534_, _19533_, _06282_);
  or (_19535_, _19534_, _19532_);
  nor (_19537_, _11332_, _07623_);
  or (_19538_, _19537_, _19533_);
  or (_19539_, _19538_, _06293_);
  and (_19540_, _14754_, _08002_);
  or (_19541_, _19540_, _19533_);
  and (_19542_, _19541_, _06401_);
  nor (_19543_, _07199_, _19530_);
  and (_19544_, _08002_, \uc8051golden_1.ACC [2]);
  or (_19545_, _19544_, _19533_);
  and (_19546_, _19545_, _07199_);
  or (_19548_, _19546_, _19543_);
  and (_19549_, _19548_, _07210_);
  or (_19550_, _19549_, _06399_);
  or (_19551_, _19550_, _19542_);
  or (_19552_, _19538_, _07221_);
  and (_19553_, _19552_, _06414_);
  and (_19554_, _19553_, _19551_);
  and (_19555_, _19545_, _06406_);
  or (_19556_, _19555_, _10059_);
  or (_19557_, _19556_, _19554_);
  and (_19559_, _19557_, _19539_);
  or (_19560_, _19559_, _06281_);
  and (_19561_, _19560_, _19535_);
  or (_19562_, _19561_, _06015_);
  and (_19563_, _14848_, _08002_);
  or (_19564_, _19533_, _06279_);
  or (_19565_, _19564_, _19563_);
  and (_19566_, _19565_, _06276_);
  and (_19567_, _19566_, _19562_);
  and (_19568_, _08002_, _08994_);
  or (_19570_, _19568_, _19533_);
  and (_19571_, _19570_, _06275_);
  or (_19572_, _19571_, _06474_);
  or (_19573_, _19572_, _19567_);
  and (_19574_, _14744_, _08002_);
  or (_19575_, _19574_, _19533_);
  or (_19576_, _19575_, _07282_);
  and (_19577_, _19576_, _07284_);
  and (_19578_, _19577_, _19573_);
  and (_19579_, _11221_, _08002_);
  or (_19581_, _19579_, _19533_);
  and (_19582_, _19581_, _06582_);
  or (_19583_, _19582_, _19578_);
  and (_19584_, _19583_, _07279_);
  or (_19585_, _19533_, _08433_);
  and (_19586_, _19570_, _06478_);
  and (_19587_, _19586_, _19585_);
  or (_19588_, _19587_, _19584_);
  and (_19589_, _19588_, _07276_);
  and (_19590_, _19545_, _06569_);
  and (_19592_, _19590_, _19585_);
  or (_19593_, _19592_, _06479_);
  or (_19594_, _19593_, _19589_);
  and (_19595_, _14741_, _08002_);
  or (_19596_, _19533_, _09043_);
  or (_19597_, _19596_, _19595_);
  and (_19598_, _19597_, _09048_);
  and (_19599_, _19598_, _19594_);
  nor (_19600_, _11220_, _11332_);
  or (_19601_, _19600_, _19533_);
  and (_19603_, _19601_, _06572_);
  or (_19604_, _19603_, _19599_);
  and (_19605_, _19604_, _07037_);
  and (_19606_, _19541_, _06606_);
  or (_19607_, _19606_, _06195_);
  or (_19608_, _19607_, _19605_);
  and (_19609_, _14917_, _08002_);
  or (_19610_, _19533_, _06196_);
  or (_19611_, _19610_, _19609_);
  and (_19612_, _19611_, _01375_);
  and (_19614_, _19612_, _19608_);
  or (_19615_, _19614_, _19531_);
  and (_42907_, _19615_, _42545_);
  and (_19616_, _11332_, \uc8051golden_1.PCON [3]);
  and (_19617_, _08002_, _09443_);
  or (_19618_, _19617_, _19616_);
  and (_19619_, _19618_, _06281_);
  and (_19620_, _14947_, _08002_);
  or (_19621_, _19620_, _19616_);
  or (_19622_, _19621_, _07210_);
  and (_19624_, _08002_, \uc8051golden_1.ACC [3]);
  or (_19625_, _19624_, _19616_);
  and (_19626_, _19625_, _07199_);
  and (_19627_, _07200_, \uc8051golden_1.PCON [3]);
  or (_19628_, _19627_, _06401_);
  or (_19629_, _19628_, _19626_);
  and (_19630_, _19629_, _07221_);
  and (_19631_, _19630_, _19622_);
  nor (_19632_, _11332_, _07775_);
  or (_19633_, _19632_, _19616_);
  and (_19635_, _19633_, _06399_);
  or (_19636_, _19635_, _19631_);
  and (_19637_, _19636_, _06414_);
  and (_19638_, _19625_, _06406_);
  or (_19639_, _19638_, _10059_);
  or (_19640_, _19639_, _19637_);
  or (_19641_, _19633_, _06293_);
  and (_19642_, _19641_, _06282_);
  and (_19643_, _19642_, _19640_);
  or (_19644_, _19643_, _06015_);
  or (_19646_, _19644_, _19619_);
  and (_19647_, _15039_, _08002_);
  or (_19648_, _19616_, _06279_);
  or (_19649_, _19648_, _19647_);
  and (_19650_, _19649_, _06276_);
  and (_19651_, _19650_, _19646_);
  and (_19652_, _08002_, _08815_);
  or (_19653_, _19652_, _19616_);
  and (_19654_, _19653_, _06275_);
  or (_19655_, _19654_, _06474_);
  or (_19657_, _19655_, _19651_);
  and (_19658_, _14934_, _08002_);
  or (_19659_, _19658_, _19616_);
  or (_19660_, _19659_, _07282_);
  and (_19661_, _19660_, _07284_);
  and (_19662_, _19661_, _19657_);
  and (_19663_, _12535_, _08002_);
  or (_19664_, _19663_, _19616_);
  and (_19665_, _19664_, _06582_);
  or (_19666_, _19665_, _19662_);
  and (_19668_, _19666_, _07279_);
  or (_19669_, _19616_, _08389_);
  and (_19670_, _19653_, _06478_);
  and (_19671_, _19670_, _19669_);
  or (_19672_, _19671_, _19668_);
  and (_19673_, _19672_, _07276_);
  and (_19674_, _19625_, _06569_);
  and (_19675_, _19674_, _19669_);
  or (_19676_, _19675_, _06479_);
  or (_19677_, _19676_, _19673_);
  and (_19679_, _14931_, _08002_);
  or (_19680_, _19616_, _09043_);
  or (_19681_, _19680_, _19679_);
  and (_19682_, _19681_, _09048_);
  and (_19683_, _19682_, _19677_);
  nor (_19684_, _11218_, _11332_);
  or (_19685_, _19684_, _19616_);
  and (_19686_, _19685_, _06572_);
  or (_19687_, _19686_, _06606_);
  or (_19688_, _19687_, _19683_);
  or (_19690_, _19621_, _07037_);
  and (_19691_, _19690_, _06196_);
  and (_19692_, _19691_, _19688_);
  and (_19693_, _15113_, _08002_);
  or (_19694_, _19693_, _19616_);
  and (_19695_, _19694_, _06195_);
  or (_19696_, _19695_, _01379_);
  or (_19697_, _19696_, _19692_);
  or (_19698_, _01375_, \uc8051golden_1.PCON [3]);
  and (_19699_, _19698_, _42545_);
  and (_42908_, _19699_, _19697_);
  and (_19701_, _11332_, \uc8051golden_1.PCON [4]);
  and (_19702_, _15130_, _08002_);
  or (_19703_, _19702_, _19701_);
  or (_19704_, _19703_, _07210_);
  and (_19705_, _08002_, \uc8051golden_1.ACC [4]);
  or (_19706_, _19705_, _19701_);
  and (_19707_, _19706_, _07199_);
  and (_19708_, _07200_, \uc8051golden_1.PCON [4]);
  or (_19709_, _19708_, _06401_);
  or (_19711_, _19709_, _19707_);
  and (_19712_, _19711_, _07221_);
  and (_19713_, _19712_, _19704_);
  nor (_19714_, _11332_, _08301_);
  or (_19715_, _19714_, _19701_);
  and (_19716_, _19715_, _06399_);
  or (_19717_, _19716_, _19713_);
  and (_19718_, _19717_, _06414_);
  and (_19719_, _19706_, _06406_);
  or (_19720_, _19719_, _10059_);
  or (_19722_, _19720_, _19718_);
  or (_19723_, _19715_, _06293_);
  and (_19724_, _19723_, _19722_);
  or (_19725_, _19724_, _06281_);
  and (_19726_, _08002_, _09442_);
  or (_19727_, _19701_, _06282_);
  or (_19728_, _19727_, _19726_);
  and (_19729_, _19728_, _06279_);
  and (_19730_, _19729_, _19725_);
  and (_19731_, _15243_, _08002_);
  or (_19733_, _19731_, _19701_);
  and (_19734_, _19733_, _06015_);
  or (_19735_, _19734_, _06275_);
  or (_19736_, _19735_, _19730_);
  and (_19737_, _08883_, _08002_);
  or (_19738_, _19737_, _19701_);
  or (_19739_, _19738_, _06276_);
  and (_19740_, _19739_, _19736_);
  or (_19741_, _19740_, _06474_);
  and (_19742_, _15135_, _08002_);
  or (_19744_, _19742_, _19701_);
  or (_19745_, _19744_, _07282_);
  and (_19746_, _19745_, _07284_);
  and (_19747_, _19746_, _19741_);
  and (_19748_, _11216_, _08002_);
  or (_19749_, _19748_, _19701_);
  and (_19750_, _19749_, _06582_);
  or (_19751_, _19750_, _19747_);
  and (_19752_, _19751_, _07279_);
  or (_19753_, _19701_, _08345_);
  and (_19755_, _19738_, _06478_);
  and (_19756_, _19755_, _19753_);
  or (_19757_, _19756_, _19752_);
  and (_19758_, _19757_, _07276_);
  and (_19759_, _19706_, _06569_);
  and (_19760_, _19759_, _19753_);
  or (_19761_, _19760_, _06479_);
  or (_19762_, _19761_, _19758_);
  and (_19763_, _15134_, _08002_);
  or (_19764_, _19701_, _09043_);
  or (_19767_, _19764_, _19763_);
  and (_19768_, _19767_, _09048_);
  and (_19769_, _19768_, _19762_);
  nor (_19770_, _11215_, _11332_);
  or (_19771_, _19770_, _19701_);
  and (_19772_, _19771_, _06572_);
  or (_19773_, _19772_, _06606_);
  or (_19774_, _19773_, _19769_);
  or (_19775_, _19703_, _07037_);
  and (_19776_, _19775_, _06196_);
  and (_19779_, _19776_, _19774_);
  and (_19780_, _15315_, _08002_);
  or (_19781_, _19780_, _19701_);
  and (_19782_, _19781_, _06195_);
  or (_19783_, _19782_, _01379_);
  or (_19784_, _19783_, _19779_);
  or (_19785_, _01375_, \uc8051golden_1.PCON [4]);
  and (_19786_, _19785_, _42545_);
  and (_42909_, _19786_, _19784_);
  and (_19787_, _11332_, \uc8051golden_1.PCON [5]);
  nor (_19790_, _11332_, _08207_);
  or (_19791_, _19790_, _19787_);
  or (_19792_, _19791_, _06293_);
  and (_19793_, _15348_, _08002_);
  or (_19794_, _19793_, _19787_);
  or (_19795_, _19794_, _07210_);
  and (_19796_, _08002_, \uc8051golden_1.ACC [5]);
  or (_19797_, _19796_, _19787_);
  and (_19798_, _19797_, _07199_);
  and (_19799_, _07200_, \uc8051golden_1.PCON [5]);
  or (_19802_, _19799_, _06401_);
  or (_19803_, _19802_, _19798_);
  and (_19804_, _19803_, _07221_);
  and (_19805_, _19804_, _19795_);
  and (_19806_, _19791_, _06399_);
  or (_19807_, _19806_, _19805_);
  and (_19808_, _19807_, _06414_);
  and (_19809_, _19797_, _06406_);
  or (_19810_, _19809_, _10059_);
  or (_19811_, _19810_, _19808_);
  and (_19814_, _19811_, _19792_);
  or (_19815_, _19814_, _06281_);
  and (_19816_, _08002_, _09441_);
  or (_19817_, _19787_, _06282_);
  or (_19818_, _19817_, _19816_);
  and (_19819_, _19818_, _06279_);
  and (_19820_, _19819_, _19815_);
  and (_19821_, _15446_, _08002_);
  or (_19822_, _19821_, _19787_);
  and (_19823_, _19822_, _06015_);
  or (_19826_, _19823_, _06275_);
  or (_19827_, _19826_, _19820_);
  and (_19828_, _08958_, _08002_);
  or (_19829_, _19828_, _19787_);
  or (_19830_, _19829_, _06276_);
  and (_19831_, _19830_, _19827_);
  or (_19832_, _19831_, _06474_);
  and (_19833_, _15338_, _08002_);
  or (_19834_, _19833_, _19787_);
  or (_19835_, _19834_, _07282_);
  and (_19838_, _19835_, _07284_);
  and (_19839_, _19838_, _19832_);
  and (_19840_, _12542_, _08002_);
  or (_19841_, _19840_, _19787_);
  and (_19842_, _19841_, _06582_);
  or (_19843_, _19842_, _19839_);
  and (_19844_, _19843_, _07279_);
  or (_19845_, _19787_, _08256_);
  and (_19846_, _19829_, _06478_);
  and (_19847_, _19846_, _19845_);
  or (_19849_, _19847_, _19844_);
  and (_19850_, _19849_, _07276_);
  and (_19851_, _19797_, _06569_);
  and (_19852_, _19851_, _19845_);
  or (_19853_, _19852_, _06479_);
  or (_19854_, _19853_, _19850_);
  and (_19855_, _15335_, _08002_);
  or (_19856_, _19787_, _09043_);
  or (_19857_, _19856_, _19855_);
  and (_19858_, _19857_, _09048_);
  and (_19860_, _19858_, _19854_);
  nor (_19861_, _11212_, _11332_);
  or (_19862_, _19861_, _19787_);
  and (_19863_, _19862_, _06572_);
  or (_19864_, _19863_, _06606_);
  or (_19865_, _19864_, _19860_);
  or (_19866_, _19794_, _07037_);
  and (_19867_, _19866_, _06196_);
  and (_19868_, _19867_, _19865_);
  and (_19869_, _15509_, _08002_);
  or (_19871_, _19869_, _19787_);
  and (_19872_, _19871_, _06195_);
  or (_19873_, _19872_, _01379_);
  or (_19874_, _19873_, _19868_);
  or (_19875_, _01375_, \uc8051golden_1.PCON [5]);
  and (_19876_, _19875_, _42545_);
  and (_42910_, _19876_, _19874_);
  and (_19877_, _11332_, \uc8051golden_1.PCON [6]);
  nor (_19878_, _11332_, _08118_);
  or (_19879_, _19878_, _19877_);
  or (_19881_, _19879_, _06293_);
  and (_19882_, _15550_, _08002_);
  or (_19883_, _19882_, _19877_);
  or (_19884_, _19883_, _07210_);
  and (_19885_, _08002_, \uc8051golden_1.ACC [6]);
  or (_19886_, _19885_, _19877_);
  and (_19887_, _19886_, _07199_);
  and (_19888_, _07200_, \uc8051golden_1.PCON [6]);
  or (_19889_, _19888_, _06401_);
  or (_19890_, _19889_, _19887_);
  and (_19892_, _19890_, _07221_);
  and (_19893_, _19892_, _19884_);
  and (_19894_, _19879_, _06399_);
  or (_19895_, _19894_, _19893_);
  and (_19896_, _19895_, _06414_);
  and (_19897_, _19886_, _06406_);
  or (_19898_, _19897_, _10059_);
  or (_19899_, _19898_, _19896_);
  and (_19900_, _19899_, _19881_);
  or (_19901_, _19900_, _06281_);
  and (_19903_, _08002_, _09440_);
  or (_19904_, _19877_, _06282_);
  or (_19905_, _19904_, _19903_);
  and (_19906_, _19905_, _06279_);
  and (_19907_, _19906_, _19901_);
  and (_19908_, _15639_, _08002_);
  or (_19909_, _19908_, _19877_);
  and (_19910_, _19909_, _06015_);
  or (_19911_, _19910_, _06275_);
  or (_19912_, _19911_, _19907_);
  and (_19914_, _15646_, _08002_);
  or (_19915_, _19914_, _19877_);
  or (_19916_, _19915_, _06276_);
  and (_19917_, _19916_, _19912_);
  or (_19918_, _19917_, _06474_);
  and (_19919_, _15531_, _08002_);
  or (_19920_, _19919_, _19877_);
  or (_19921_, _19920_, _07282_);
  and (_19922_, _19921_, _07284_);
  and (_19923_, _19922_, _19918_);
  and (_19925_, _11210_, _08002_);
  or (_19926_, _19925_, _19877_);
  and (_19927_, _19926_, _06582_);
  or (_19928_, _19927_, _19923_);
  and (_19929_, _19928_, _07279_);
  or (_19930_, _19877_, _08162_);
  and (_19931_, _19915_, _06478_);
  and (_19932_, _19931_, _19930_);
  or (_19933_, _19932_, _19929_);
  and (_19934_, _19933_, _07276_);
  and (_19936_, _19886_, _06569_);
  and (_19937_, _19936_, _19930_);
  or (_19938_, _19937_, _06479_);
  or (_19939_, _19938_, _19934_);
  and (_19940_, _15528_, _08002_);
  or (_19941_, _19877_, _09043_);
  or (_19942_, _19941_, _19940_);
  and (_19943_, _19942_, _09048_);
  and (_19944_, _19943_, _19939_);
  nor (_19945_, _11209_, _11332_);
  or (_19947_, _19945_, _19877_);
  and (_19948_, _19947_, _06572_);
  or (_19949_, _19948_, _06606_);
  or (_19950_, _19949_, _19944_);
  or (_19951_, _19883_, _07037_);
  and (_19952_, _19951_, _06196_);
  and (_19953_, _19952_, _19950_);
  and (_19954_, _15713_, _08002_);
  or (_19955_, _19954_, _19877_);
  and (_19956_, _19955_, _06195_);
  or (_19958_, _19956_, _01379_);
  or (_19959_, _19958_, _19953_);
  or (_19960_, _01375_, \uc8051golden_1.PCON [6]);
  and (_19961_, _19960_, _42545_);
  and (_42911_, _19961_, _19959_);
  not (_19962_, \uc8051golden_1.TMOD [0]);
  nor (_19963_, _01375_, _19962_);
  nand (_19964_, _11225_, _08006_);
  nor (_19965_, _08006_, _19962_);
  nor (_19966_, _19965_, _07276_);
  nand (_19968_, _19966_, _19964_);
  and (_19969_, _08006_, _07473_);
  or (_19970_, _19969_, _19965_);
  or (_19971_, _19970_, _06293_);
  nor (_19972_, _08521_, _11410_);
  or (_19973_, _19972_, _19965_);
  or (_19974_, _19973_, _07210_);
  and (_19975_, _08006_, \uc8051golden_1.ACC [0]);
  or (_19976_, _19975_, _19965_);
  and (_19977_, _19976_, _07199_);
  nor (_19979_, _07199_, _19962_);
  or (_19980_, _19979_, _06401_);
  or (_19981_, _19980_, _19977_);
  and (_19982_, _19981_, _07221_);
  and (_19983_, _19982_, _19974_);
  and (_19984_, _19970_, _06399_);
  or (_19985_, _19984_, _19983_);
  and (_19986_, _19985_, _06414_);
  and (_19987_, _19976_, _06406_);
  or (_19988_, _19987_, _10059_);
  or (_19990_, _19988_, _19986_);
  and (_19991_, _19990_, _19971_);
  or (_19992_, _19991_, _06281_);
  and (_19993_, _08006_, _09446_);
  or (_19994_, _19965_, _06282_);
  or (_19995_, _19994_, _19993_);
  and (_19996_, _19995_, _19992_);
  or (_19997_, _19996_, _06015_);
  and (_19998_, _14426_, _08006_);
  or (_19999_, _19965_, _06279_);
  or (_20001_, _19999_, _19998_);
  and (_20002_, _20001_, _06276_);
  and (_20003_, _20002_, _19997_);
  and (_20004_, _08006_, _08817_);
  or (_20005_, _20004_, _19965_);
  and (_20006_, _20005_, _06275_);
  or (_20007_, _20006_, _06474_);
  or (_20008_, _20007_, _20003_);
  and (_20009_, _14324_, _08006_);
  or (_20010_, _20009_, _19965_);
  or (_20012_, _20010_, _07282_);
  and (_20013_, _20012_, _07284_);
  and (_20014_, _20013_, _20008_);
  nor (_20015_, _12538_, _11410_);
  or (_20016_, _20015_, _19965_);
  and (_20017_, _19964_, _06582_);
  and (_20018_, _20017_, _20016_);
  or (_20019_, _20018_, _20014_);
  and (_20020_, _20019_, _07279_);
  nand (_20021_, _20005_, _06478_);
  nor (_20023_, _20021_, _19972_);
  or (_20024_, _20023_, _06569_);
  or (_20025_, _20024_, _20020_);
  and (_20026_, _20025_, _19968_);
  or (_20027_, _20026_, _06479_);
  and (_20028_, _14320_, _08006_);
  or (_20029_, _19965_, _09043_);
  or (_20030_, _20029_, _20028_);
  and (_20031_, _20030_, _09048_);
  and (_20032_, _20031_, _20027_);
  and (_20034_, _20016_, _06572_);
  or (_20035_, _20034_, _19434_);
  or (_20036_, _20035_, _20032_);
  or (_20037_, _19973_, _06700_);
  and (_20038_, _20037_, _01375_);
  and (_20039_, _20038_, _20036_);
  or (_20040_, _20039_, _19963_);
  and (_42912_, _20040_, _42545_);
  and (_20041_, _01379_, \uc8051golden_1.TMOD [1]);
  nand (_20042_, _08006_, _07090_);
  or (_20044_, _08006_, \uc8051golden_1.TMOD [1]);
  and (_20045_, _20044_, _06275_);
  and (_20046_, _20045_, _20042_);
  and (_20047_, _08006_, _09445_);
  and (_20048_, _11410_, \uc8051golden_1.TMOD [1]);
  or (_20049_, _20048_, _06282_);
  or (_20050_, _20049_, _20047_);
  nor (_20051_, _11410_, _07196_);
  or (_20052_, _20051_, _20048_);
  or (_20053_, _20052_, _06293_);
  and (_20055_, _14532_, _08006_);
  not (_20056_, _20055_);
  and (_20057_, _20056_, _20044_);
  or (_20058_, _20057_, _07210_);
  and (_20059_, _08006_, \uc8051golden_1.ACC [1]);
  or (_20060_, _20059_, _20048_);
  and (_20061_, _20060_, _07199_);
  and (_20062_, _07200_, \uc8051golden_1.TMOD [1]);
  or (_20063_, _20062_, _06401_);
  or (_20064_, _20063_, _20061_);
  and (_20066_, _20064_, _07221_);
  and (_20067_, _20066_, _20058_);
  and (_20068_, _20052_, _06399_);
  or (_20069_, _20068_, _20067_);
  and (_20070_, _20069_, _06414_);
  and (_20071_, _20060_, _06406_);
  or (_20072_, _20071_, _10059_);
  or (_20073_, _20072_, _20070_);
  and (_20074_, _20073_, _20053_);
  or (_20075_, _20074_, _06281_);
  and (_20077_, _20075_, _06279_);
  and (_20078_, _20077_, _20050_);
  or (_20079_, _14615_, _11410_);
  and (_20080_, _20044_, _06015_);
  and (_20081_, _20080_, _20079_);
  or (_20082_, _20081_, _20078_);
  and (_20083_, _20082_, _06276_);
  or (_20084_, _20083_, _20046_);
  and (_20085_, _20084_, _07282_);
  or (_20086_, _14507_, _11410_);
  and (_20088_, _20044_, _06474_);
  and (_20089_, _20088_, _20086_);
  or (_20090_, _20089_, _06582_);
  or (_20091_, _20090_, _20085_);
  and (_20092_, _11224_, _08006_);
  or (_20093_, _20092_, _20048_);
  or (_20094_, _20093_, _07284_);
  and (_20095_, _20094_, _07279_);
  and (_20096_, _20095_, _20091_);
  or (_20097_, _14505_, _11410_);
  and (_20099_, _20044_, _06478_);
  and (_20100_, _20099_, _20097_);
  or (_20101_, _20100_, _06569_);
  or (_20102_, _20101_, _20096_);
  and (_20103_, _20059_, _08477_);
  or (_20104_, _20048_, _07276_);
  or (_20105_, _20104_, _20103_);
  and (_20106_, _20105_, _09043_);
  and (_20107_, _20106_, _20102_);
  or (_20108_, _20042_, _08477_);
  and (_20110_, _20044_, _06479_);
  and (_20111_, _20110_, _20108_);
  or (_20112_, _20111_, _06572_);
  or (_20113_, _20112_, _20107_);
  nor (_20114_, _11223_, _11410_);
  or (_20115_, _20114_, _20048_);
  or (_20116_, _20115_, _09048_);
  and (_20117_, _20116_, _07037_);
  and (_20118_, _20117_, _20113_);
  and (_20119_, _20057_, _06606_);
  or (_20121_, _20119_, _06195_);
  or (_20122_, _20121_, _20118_);
  or (_20123_, _20048_, _06196_);
  or (_20124_, _20123_, _20055_);
  and (_20125_, _20124_, _01375_);
  and (_20126_, _20125_, _20122_);
  or (_20127_, _20126_, _20041_);
  and (_42913_, _20127_, _42545_);
  and (_20128_, _01379_, \uc8051golden_1.TMOD [2]);
  and (_20129_, _08006_, _09444_);
  and (_20131_, _11410_, \uc8051golden_1.TMOD [2]);
  or (_20132_, _20131_, _06282_);
  or (_20133_, _20132_, _20129_);
  nor (_20134_, _11410_, _07623_);
  or (_20135_, _20134_, _20131_);
  or (_20136_, _20135_, _06293_);
  and (_20137_, _14754_, _08006_);
  or (_20138_, _20137_, _20131_);
  and (_20139_, _20138_, _06401_);
  and (_20140_, _07200_, \uc8051golden_1.TMOD [2]);
  and (_20142_, _08006_, \uc8051golden_1.ACC [2]);
  or (_20143_, _20142_, _20131_);
  and (_20144_, _20143_, _07199_);
  or (_20145_, _20144_, _20140_);
  and (_20146_, _20145_, _07210_);
  or (_20147_, _20146_, _06399_);
  or (_20148_, _20147_, _20139_);
  or (_20149_, _20135_, _07221_);
  and (_20150_, _20149_, _06414_);
  and (_20151_, _20150_, _20148_);
  and (_20153_, _20143_, _06406_);
  or (_20154_, _20153_, _10059_);
  or (_20155_, _20154_, _20151_);
  and (_20156_, _20155_, _20136_);
  or (_20157_, _20156_, _06281_);
  and (_20158_, _20157_, _20133_);
  or (_20159_, _20158_, _06015_);
  and (_20160_, _14848_, _08006_);
  or (_20161_, _20131_, _06279_);
  or (_20162_, _20161_, _20160_);
  and (_20164_, _20162_, _06276_);
  and (_20165_, _20164_, _20159_);
  and (_20166_, _08006_, _08994_);
  or (_20167_, _20166_, _20131_);
  and (_20168_, _20167_, _06275_);
  or (_20169_, _20168_, _06474_);
  or (_20170_, _20169_, _20165_);
  and (_20171_, _14744_, _08006_);
  or (_20172_, _20171_, _20131_);
  or (_20173_, _20172_, _07282_);
  and (_20175_, _20173_, _07284_);
  and (_20176_, _20175_, _20170_);
  and (_20177_, _11221_, _08006_);
  or (_20178_, _20177_, _20131_);
  and (_20179_, _20178_, _06582_);
  or (_20180_, _20179_, _20176_);
  and (_20181_, _20180_, _07279_);
  or (_20182_, _20131_, _08433_);
  and (_20183_, _20167_, _06478_);
  and (_20184_, _20183_, _20182_);
  or (_20186_, _20184_, _20181_);
  and (_20187_, _20186_, _07276_);
  and (_20188_, _20143_, _06569_);
  and (_20189_, _20188_, _20182_);
  or (_20190_, _20189_, _06479_);
  or (_20191_, _20190_, _20187_);
  and (_20192_, _14741_, _08006_);
  or (_20193_, _20131_, _09043_);
  or (_20194_, _20193_, _20192_);
  and (_20195_, _20194_, _09048_);
  and (_20197_, _20195_, _20191_);
  nor (_20198_, _11220_, _11410_);
  or (_20199_, _20198_, _20131_);
  and (_20200_, _20199_, _06572_);
  or (_20201_, _20200_, _20197_);
  and (_20202_, _20201_, _07037_);
  and (_20203_, _20138_, _06606_);
  or (_20204_, _20203_, _06195_);
  or (_20205_, _20204_, _20202_);
  and (_20206_, _14917_, _08006_);
  or (_20208_, _20131_, _06196_);
  or (_20209_, _20208_, _20206_);
  and (_20210_, _20209_, _01375_);
  and (_20211_, _20210_, _20205_);
  or (_20212_, _20211_, _20128_);
  and (_42914_, _20212_, _42545_);
  and (_20213_, _11410_, \uc8051golden_1.TMOD [3]);
  nor (_20214_, _11410_, _07775_);
  or (_20215_, _20214_, _20213_);
  or (_20216_, _20215_, _06293_);
  and (_20218_, _14947_, _08006_);
  or (_20219_, _20218_, _20213_);
  or (_20220_, _20219_, _07210_);
  and (_20221_, _08006_, \uc8051golden_1.ACC [3]);
  or (_20222_, _20221_, _20213_);
  and (_20223_, _20222_, _07199_);
  and (_20224_, _07200_, \uc8051golden_1.TMOD [3]);
  or (_20225_, _20224_, _06401_);
  or (_20226_, _20225_, _20223_);
  and (_20227_, _20226_, _07221_);
  and (_20229_, _20227_, _20220_);
  and (_20230_, _20215_, _06399_);
  or (_20231_, _20230_, _20229_);
  and (_20232_, _20231_, _06414_);
  and (_20233_, _20222_, _06406_);
  or (_20234_, _20233_, _10059_);
  or (_20235_, _20234_, _20232_);
  and (_20236_, _20235_, _20216_);
  or (_20237_, _20236_, _06281_);
  and (_20238_, _08006_, _09443_);
  or (_20240_, _20213_, _06282_);
  or (_20241_, _20240_, _20238_);
  and (_20242_, _20241_, _20237_);
  or (_20243_, _20242_, _06015_);
  and (_20244_, _15039_, _08006_);
  or (_20245_, _20213_, _06279_);
  or (_20246_, _20245_, _20244_);
  and (_20247_, _20246_, _06276_);
  and (_20248_, _20247_, _20243_);
  and (_20249_, _08006_, _08815_);
  or (_20251_, _20249_, _20213_);
  and (_20252_, _20251_, _06275_);
  or (_20253_, _20252_, _06474_);
  or (_20254_, _20253_, _20248_);
  and (_20255_, _14934_, _08006_);
  or (_20256_, _20255_, _20213_);
  or (_20257_, _20256_, _07282_);
  and (_20258_, _20257_, _07284_);
  and (_20259_, _20258_, _20254_);
  and (_20260_, _12535_, _08006_);
  or (_20262_, _20260_, _20213_);
  and (_20263_, _20262_, _06582_);
  or (_20264_, _20263_, _20259_);
  and (_20265_, _20264_, _07279_);
  or (_20266_, _20213_, _08389_);
  and (_20267_, _20251_, _06478_);
  and (_20268_, _20267_, _20266_);
  or (_20269_, _20268_, _20265_);
  and (_20270_, _20269_, _07276_);
  and (_20271_, _20222_, _06569_);
  and (_20273_, _20271_, _20266_);
  or (_20274_, _20273_, _06479_);
  or (_20275_, _20274_, _20270_);
  and (_20276_, _14931_, _08006_);
  or (_20277_, _20213_, _09043_);
  or (_20278_, _20277_, _20276_);
  and (_20279_, _20278_, _09048_);
  and (_20280_, _20279_, _20275_);
  nor (_20281_, _11218_, _11410_);
  or (_20282_, _20281_, _20213_);
  and (_20284_, _20282_, _06572_);
  or (_20285_, _20284_, _06606_);
  or (_20286_, _20285_, _20280_);
  or (_20287_, _20219_, _07037_);
  and (_20288_, _20287_, _06196_);
  and (_20289_, _20288_, _20286_);
  and (_20290_, _15113_, _08006_);
  or (_20291_, _20290_, _20213_);
  and (_20292_, _20291_, _06195_);
  or (_20293_, _20292_, _01379_);
  or (_20295_, _20293_, _20289_);
  or (_20296_, _01375_, \uc8051golden_1.TMOD [3]);
  and (_20297_, _20296_, _42545_);
  and (_42916_, _20297_, _20295_);
  and (_20298_, _11410_, \uc8051golden_1.TMOD [4]);
  and (_20299_, _15130_, _08006_);
  or (_20300_, _20299_, _20298_);
  or (_20301_, _20300_, _07210_);
  and (_20302_, _08006_, \uc8051golden_1.ACC [4]);
  or (_20303_, _20302_, _20298_);
  and (_20305_, _20303_, _07199_);
  and (_20306_, _07200_, \uc8051golden_1.TMOD [4]);
  or (_20307_, _20306_, _06401_);
  or (_20308_, _20307_, _20305_);
  and (_20309_, _20308_, _07221_);
  and (_20310_, _20309_, _20301_);
  nor (_20311_, _11410_, _08301_);
  or (_20312_, _20311_, _20298_);
  and (_20313_, _20312_, _06399_);
  or (_20314_, _20313_, _20310_);
  and (_20316_, _20314_, _06414_);
  and (_20317_, _20303_, _06406_);
  or (_20318_, _20317_, _10059_);
  or (_20319_, _20318_, _20316_);
  or (_20320_, _20312_, _06293_);
  and (_20321_, _20320_, _20319_);
  or (_20322_, _20321_, _06281_);
  and (_20323_, _08006_, _09442_);
  or (_20324_, _20298_, _06282_);
  or (_20325_, _20324_, _20323_);
  and (_20327_, _20325_, _06279_);
  and (_20328_, _20327_, _20322_);
  and (_20329_, _15243_, _08006_);
  or (_20330_, _20329_, _20298_);
  and (_20331_, _20330_, _06015_);
  or (_20332_, _20331_, _06275_);
  or (_20333_, _20332_, _20328_);
  and (_20334_, _08883_, _08006_);
  or (_20335_, _20334_, _20298_);
  or (_20336_, _20335_, _06276_);
  and (_20338_, _20336_, _20333_);
  or (_20339_, _20338_, _06474_);
  and (_20340_, _15135_, _08006_);
  or (_20341_, _20340_, _20298_);
  or (_20342_, _20341_, _07282_);
  and (_20343_, _20342_, _07284_);
  and (_20344_, _20343_, _20339_);
  and (_20345_, _11216_, _08006_);
  or (_20346_, _20345_, _20298_);
  and (_20347_, _20346_, _06582_);
  or (_20349_, _20347_, _20344_);
  and (_20350_, _20349_, _07279_);
  or (_20351_, _20298_, _08345_);
  and (_20352_, _20335_, _06478_);
  and (_20353_, _20352_, _20351_);
  or (_20354_, _20353_, _20350_);
  and (_20355_, _20354_, _07276_);
  and (_20356_, _20303_, _06569_);
  and (_20357_, _20356_, _20351_);
  or (_20358_, _20357_, _06479_);
  or (_20360_, _20358_, _20355_);
  and (_20361_, _15134_, _08006_);
  or (_20362_, _20298_, _09043_);
  or (_20363_, _20362_, _20361_);
  and (_20364_, _20363_, _09048_);
  and (_20365_, _20364_, _20360_);
  nor (_20366_, _11215_, _11410_);
  or (_20367_, _20366_, _20298_);
  and (_20368_, _20367_, _06572_);
  or (_20369_, _20368_, _06606_);
  or (_20371_, _20369_, _20365_);
  or (_20372_, _20300_, _07037_);
  and (_20373_, _20372_, _06196_);
  and (_20374_, _20373_, _20371_);
  and (_20375_, _15315_, _08006_);
  or (_20376_, _20375_, _20298_);
  and (_20377_, _20376_, _06195_);
  or (_20378_, _20377_, _01379_);
  or (_20379_, _20378_, _20374_);
  or (_20380_, _01375_, \uc8051golden_1.TMOD [4]);
  and (_20382_, _20380_, _42545_);
  and (_42917_, _20382_, _20379_);
  and (_20383_, _11410_, \uc8051golden_1.TMOD [5]);
  nor (_20384_, _11410_, _08207_);
  or (_20385_, _20384_, _20383_);
  or (_20386_, _20385_, _06293_);
  and (_20387_, _15348_, _08006_);
  or (_20388_, _20387_, _20383_);
  or (_20389_, _20388_, _07210_);
  and (_20390_, _08006_, \uc8051golden_1.ACC [5]);
  or (_20392_, _20390_, _20383_);
  and (_20393_, _20392_, _07199_);
  and (_20394_, _07200_, \uc8051golden_1.TMOD [5]);
  or (_20395_, _20394_, _06401_);
  or (_20396_, _20395_, _20393_);
  and (_20397_, _20396_, _07221_);
  and (_20398_, _20397_, _20389_);
  and (_20399_, _20385_, _06399_);
  or (_20400_, _20399_, _20398_);
  and (_20401_, _20400_, _06414_);
  and (_20403_, _20392_, _06406_);
  or (_20404_, _20403_, _10059_);
  or (_20405_, _20404_, _20401_);
  and (_20406_, _20405_, _20386_);
  or (_20407_, _20406_, _06281_);
  and (_20408_, _08006_, _09441_);
  or (_20409_, _20383_, _06282_);
  or (_20410_, _20409_, _20408_);
  and (_20411_, _20410_, _06279_);
  and (_20412_, _20411_, _20407_);
  and (_20414_, _15446_, _08006_);
  or (_20415_, _20414_, _20383_);
  and (_20416_, _20415_, _06015_);
  or (_20417_, _20416_, _06275_);
  or (_20418_, _20417_, _20412_);
  and (_20419_, _08958_, _08006_);
  or (_20420_, _20419_, _20383_);
  or (_20421_, _20420_, _06276_);
  and (_20422_, _20421_, _20418_);
  or (_20423_, _20422_, _06474_);
  and (_20425_, _15338_, _08006_);
  or (_20426_, _20425_, _20383_);
  or (_20427_, _20426_, _07282_);
  and (_20428_, _20427_, _07284_);
  and (_20429_, _20428_, _20423_);
  and (_20430_, _12542_, _08006_);
  or (_20431_, _20430_, _20383_);
  and (_20432_, _20431_, _06582_);
  or (_20433_, _20432_, _20429_);
  and (_20434_, _20433_, _07279_);
  or (_20436_, _20383_, _08256_);
  and (_20437_, _20420_, _06478_);
  and (_20438_, _20437_, _20436_);
  or (_20439_, _20438_, _20434_);
  and (_20440_, _20439_, _07276_);
  and (_20441_, _20392_, _06569_);
  and (_20442_, _20441_, _20436_);
  or (_20443_, _20442_, _06479_);
  or (_20444_, _20443_, _20440_);
  and (_20445_, _15335_, _08006_);
  or (_20447_, _20383_, _09043_);
  or (_20448_, _20447_, _20445_);
  and (_20449_, _20448_, _09048_);
  and (_20450_, _20449_, _20444_);
  nor (_20451_, _11212_, _11410_);
  or (_20452_, _20451_, _20383_);
  and (_20453_, _20452_, _06572_);
  or (_20454_, _20453_, _06606_);
  or (_20455_, _20454_, _20450_);
  or (_20456_, _20388_, _07037_);
  and (_20458_, _20456_, _06196_);
  and (_20459_, _20458_, _20455_);
  and (_20460_, _15509_, _08006_);
  or (_20461_, _20460_, _20383_);
  and (_20462_, _20461_, _06195_);
  or (_20463_, _20462_, _01379_);
  or (_20464_, _20463_, _20459_);
  or (_20465_, _01375_, \uc8051golden_1.TMOD [5]);
  and (_20466_, _20465_, _42545_);
  and (_42918_, _20466_, _20464_);
  and (_20468_, _11410_, \uc8051golden_1.TMOD [6]);
  nor (_20469_, _11410_, _08118_);
  or (_20470_, _20469_, _20468_);
  or (_20471_, _20470_, _06293_);
  and (_20472_, _15550_, _08006_);
  or (_20473_, _20472_, _20468_);
  or (_20474_, _20473_, _07210_);
  and (_20475_, _08006_, \uc8051golden_1.ACC [6]);
  or (_20476_, _20475_, _20468_);
  and (_20477_, _20476_, _07199_);
  and (_20479_, _07200_, \uc8051golden_1.TMOD [6]);
  or (_20480_, _20479_, _06401_);
  or (_20481_, _20480_, _20477_);
  and (_20482_, _20481_, _07221_);
  and (_20483_, _20482_, _20474_);
  and (_20484_, _20470_, _06399_);
  or (_20485_, _20484_, _20483_);
  and (_20486_, _20485_, _06414_);
  and (_20487_, _20476_, _06406_);
  or (_20488_, _20487_, _10059_);
  or (_20490_, _20488_, _20486_);
  and (_20491_, _20490_, _20471_);
  or (_20492_, _20491_, _06281_);
  and (_20493_, _08006_, _09440_);
  or (_20494_, _20468_, _06282_);
  or (_20495_, _20494_, _20493_);
  and (_20496_, _20495_, _06279_);
  and (_20497_, _20496_, _20492_);
  and (_20498_, _15639_, _08006_);
  or (_20499_, _20498_, _20468_);
  and (_20501_, _20499_, _06015_);
  or (_20502_, _20501_, _06275_);
  or (_20503_, _20502_, _20497_);
  and (_20504_, _15646_, _08006_);
  or (_20505_, _20504_, _20468_);
  or (_20506_, _20505_, _06276_);
  and (_20507_, _20506_, _20503_);
  or (_20508_, _20507_, _06474_);
  and (_20509_, _15531_, _08006_);
  or (_20510_, _20509_, _20468_);
  or (_20512_, _20510_, _07282_);
  and (_20513_, _20512_, _07284_);
  and (_20514_, _20513_, _20508_);
  and (_20515_, _11210_, _08006_);
  or (_20516_, _20515_, _20468_);
  and (_20517_, _20516_, _06582_);
  or (_20518_, _20517_, _20514_);
  and (_20519_, _20518_, _07279_);
  or (_20520_, _20468_, _08162_);
  and (_20521_, _20505_, _06478_);
  and (_20523_, _20521_, _20520_);
  or (_20524_, _20523_, _20519_);
  and (_20525_, _20524_, _07276_);
  and (_20526_, _20476_, _06569_);
  and (_20527_, _20526_, _20520_);
  or (_20528_, _20527_, _06479_);
  or (_20529_, _20528_, _20525_);
  and (_20530_, _15528_, _08006_);
  or (_20531_, _20468_, _09043_);
  or (_20532_, _20531_, _20530_);
  and (_20534_, _20532_, _09048_);
  and (_20535_, _20534_, _20529_);
  nor (_20536_, _11209_, _11410_);
  or (_20537_, _20536_, _20468_);
  and (_20538_, _20537_, _06572_);
  or (_20539_, _20538_, _06606_);
  or (_20540_, _20539_, _20535_);
  or (_20541_, _20473_, _07037_);
  and (_20542_, _20541_, _06196_);
  and (_20543_, _20542_, _20540_);
  and (_20545_, _15713_, _08006_);
  or (_20546_, _20545_, _20468_);
  and (_20547_, _20546_, _06195_);
  or (_20548_, _20547_, _01379_);
  or (_20549_, _20548_, _20543_);
  or (_20550_, _01375_, \uc8051golden_1.TMOD [6]);
  and (_20551_, _20550_, _42545_);
  and (_42919_, _20551_, _20549_);
  not (_20552_, \uc8051golden_1.DPL [0]);
  nor (_20553_, _01375_, _20552_);
  and (_20555_, _07962_, \uc8051golden_1.ACC [0]);
  and (_20556_, _20555_, _08521_);
  nor (_20557_, _07962_, _20552_);
  or (_20558_, _20557_, _07276_);
  or (_20559_, _20558_, _20556_);
  and (_20560_, _07962_, _07473_);
  or (_20561_, _20560_, _20557_);
  or (_20562_, _20561_, _06293_);
  or (_20563_, _20557_, _20555_);
  or (_20564_, _20563_, _06414_);
  nor (_20566_, _08521_, _11493_);
  or (_20567_, _20566_, _20557_);
  or (_20568_, _20567_, _07210_);
  and (_20569_, _20563_, _07199_);
  nor (_20570_, _07199_, _20552_);
  or (_20571_, _20570_, _06401_);
  or (_20572_, _20571_, _20569_);
  and (_20573_, _20572_, _07221_);
  and (_20574_, _20573_, _20568_);
  and (_20575_, _20561_, _06399_);
  or (_20577_, _20575_, _06406_);
  or (_20578_, _20577_, _20574_);
  and (_20579_, _20578_, _20564_);
  or (_20580_, _20579_, _11511_);
  nand (_20581_, _11511_, \uc8051golden_1.DPL [0]);
  and (_20582_, _20581_, _06473_);
  and (_20583_, _20582_, _20580_);
  nor (_20584_, _06943_, _06473_);
  or (_20585_, _20584_, _10059_);
  or (_20586_, _20585_, _20583_);
  and (_20588_, _20586_, _20562_);
  or (_20589_, _20588_, _06281_);
  and (_20590_, _07962_, _09446_);
  or (_20591_, _20557_, _06282_);
  or (_20592_, _20591_, _20590_);
  and (_20593_, _20592_, _20589_);
  or (_20594_, _20593_, _06015_);
  and (_20595_, _14426_, _07962_);
  or (_20596_, _20557_, _06279_);
  or (_20597_, _20596_, _20595_);
  and (_20599_, _20597_, _06276_);
  and (_20600_, _20599_, _20594_);
  and (_20601_, _07962_, _08817_);
  or (_20602_, _20601_, _20557_);
  and (_20603_, _20602_, _06275_);
  or (_20604_, _20603_, _06474_);
  or (_20605_, _20604_, _20600_);
  and (_20606_, _14324_, _07962_);
  or (_20607_, _20606_, _20557_);
  or (_20608_, _20607_, _07282_);
  and (_20610_, _20608_, _07284_);
  and (_20611_, _20610_, _20605_);
  nor (_20612_, _12538_, _11493_);
  or (_20613_, _20612_, _20557_);
  nor (_20614_, _20556_, _07284_);
  and (_20615_, _20614_, _20613_);
  or (_20616_, _20615_, _20611_);
  and (_20617_, _20616_, _07279_);
  nand (_20618_, _20602_, _06478_);
  nor (_20619_, _20618_, _20566_);
  or (_20621_, _20619_, _06569_);
  or (_20622_, _20621_, _20617_);
  and (_20623_, _20622_, _20559_);
  or (_20624_, _20623_, _06479_);
  and (_20625_, _14320_, _07962_);
  or (_20626_, _20625_, _20557_);
  or (_20627_, _20626_, _09043_);
  and (_20628_, _20627_, _09048_);
  and (_20629_, _20628_, _20624_);
  and (_20630_, _20613_, _06572_);
  or (_20632_, _20630_, _19434_);
  or (_20633_, _20632_, _20629_);
  or (_20634_, _20567_, _06700_);
  and (_20635_, _20634_, _01375_);
  and (_20636_, _20635_, _20633_);
  or (_20637_, _20636_, _20553_);
  and (_42921_, _20637_, _42545_);
  not (_20638_, \uc8051golden_1.DPL [1]);
  nor (_20639_, _01375_, _20638_);
  nor (_20640_, _07962_, _20638_);
  nor (_20642_, _11493_, _07196_);
  or (_20643_, _20642_, _20640_);
  or (_20644_, _20643_, _06293_);
  or (_20645_, _07962_, \uc8051golden_1.DPL [1]);
  and (_20646_, _14532_, _07962_);
  not (_20647_, _20646_);
  and (_20648_, _20647_, _20645_);
  or (_20649_, _20648_, _07210_);
  and (_20650_, _07962_, \uc8051golden_1.ACC [1]);
  or (_20651_, _20650_, _20640_);
  and (_20653_, _20651_, _07199_);
  nor (_20654_, _07199_, _20638_);
  or (_20655_, _20654_, _06401_);
  or (_20656_, _20655_, _20653_);
  and (_20657_, _20656_, _07221_);
  and (_20658_, _20657_, _20649_);
  and (_20659_, _20643_, _06399_);
  or (_20660_, _20659_, _06406_);
  or (_20661_, _20660_, _20658_);
  or (_20662_, _20651_, _06414_);
  and (_20663_, _20662_, _11512_);
  and (_20664_, _20663_, _20661_);
  nor (_20665_, \uc8051golden_1.DPL [1], \uc8051golden_1.DPL [0]);
  nor (_20666_, _20665_, _11516_);
  and (_20667_, _20666_, _11511_);
  or (_20668_, _20667_, _20664_);
  and (_20669_, _20668_, _06473_);
  nor (_20670_, _07090_, _06473_);
  or (_20671_, _20670_, _10059_);
  or (_20672_, _20671_, _20669_);
  and (_20674_, _20672_, _20644_);
  or (_20675_, _20674_, _06281_);
  and (_20676_, _20675_, _06279_);
  and (_20677_, _07962_, _09445_);
  or (_20678_, _20677_, _20640_);
  or (_20679_, _20678_, _06282_);
  and (_20680_, _20679_, _20676_);
  or (_20681_, _14615_, _11493_);
  and (_20682_, _20645_, _06015_);
  and (_20683_, _20682_, _20681_);
  or (_20686_, _20683_, _20680_);
  and (_20687_, _20686_, _06276_);
  nand (_20688_, _07962_, _07090_);
  and (_20689_, _20645_, _06275_);
  and (_20690_, _20689_, _20688_);
  or (_20691_, _20690_, _20687_);
  and (_20692_, _20691_, _07282_);
  or (_20693_, _14507_, _11493_);
  and (_20694_, _20645_, _06474_);
  and (_20695_, _20694_, _20693_);
  or (_20697_, _20695_, _06582_);
  or (_20698_, _20697_, _20692_);
  nor (_20699_, _11223_, _11493_);
  or (_20700_, _20699_, _20640_);
  nand (_20701_, _11222_, _07962_);
  and (_20702_, _20701_, _20700_);
  or (_20703_, _20702_, _07284_);
  and (_20704_, _20703_, _07279_);
  and (_20705_, _20704_, _20698_);
  or (_20706_, _14505_, _11493_);
  and (_20707_, _20645_, _06478_);
  and (_20708_, _20707_, _20706_);
  or (_20709_, _20708_, _06569_);
  or (_20710_, _20709_, _20705_);
  nor (_20711_, _20640_, _07276_);
  nand (_20712_, _20711_, _20701_);
  and (_20713_, _20712_, _09043_);
  and (_20714_, _20713_, _20710_);
  or (_20715_, _20688_, _08477_);
  and (_20716_, _20645_, _06479_);
  and (_20718_, _20716_, _20715_);
  or (_20719_, _20718_, _06572_);
  or (_20720_, _20719_, _20714_);
  or (_20721_, _20700_, _09048_);
  and (_20722_, _20721_, _07037_);
  and (_20723_, _20722_, _20720_);
  and (_20724_, _20648_, _06606_);
  or (_20725_, _20724_, _06195_);
  or (_20726_, _20725_, _20723_);
  or (_20727_, _20640_, _06196_);
  or (_20730_, _20727_, _20646_);
  and (_20731_, _20730_, _01375_);
  and (_20732_, _20731_, _20726_);
  or (_20733_, _20732_, _20639_);
  and (_42922_, _20733_, _42545_);
  not (_20734_, \uc8051golden_1.DPL [2]);
  nor (_20735_, _01375_, _20734_);
  nor (_20736_, _07962_, _20734_);
  nor (_20737_, _11493_, _07623_);
  or (_20738_, _20737_, _20736_);
  or (_20739_, _20738_, _06293_);
  or (_20740_, _20738_, _07221_);
  and (_20741_, _14754_, _07962_);
  or (_20742_, _20741_, _20736_);
  and (_20743_, _20742_, _06401_);
  nor (_20744_, _07199_, _20734_);
  and (_20745_, _07962_, \uc8051golden_1.ACC [2]);
  or (_20746_, _20745_, _20736_);
  and (_20747_, _20746_, _07199_);
  or (_20748_, _20747_, _20744_);
  and (_20750_, _20748_, _07210_);
  or (_20751_, _20750_, _06399_);
  or (_20752_, _20751_, _20743_);
  and (_20753_, _20752_, _20740_);
  or (_20754_, _20753_, _06406_);
  or (_20755_, _20746_, _06414_);
  and (_20756_, _20755_, _11512_);
  and (_20757_, _20756_, _20754_);
  nor (_20758_, _11516_, \uc8051golden_1.DPL [2]);
  nor (_20759_, _20758_, _11517_);
  and (_20762_, _20759_, _11511_);
  or (_20763_, _20762_, _20757_);
  and (_20764_, _20763_, _06473_);
  nor (_20765_, _06736_, _06473_);
  or (_20766_, _20765_, _10059_);
  or (_20767_, _20766_, _20764_);
  and (_20768_, _20767_, _20739_);
  or (_20769_, _20768_, _06281_);
  and (_20770_, _07962_, _09444_);
  or (_20771_, _20736_, _06282_);
  or (_20773_, _20771_, _20770_);
  and (_20774_, _20773_, _06279_);
  and (_20775_, _20774_, _20769_);
  and (_20776_, _14848_, _07962_);
  or (_20777_, _20776_, _20736_);
  and (_20778_, _20777_, _06015_);
  or (_20779_, _20778_, _06275_);
  or (_20780_, _20779_, _20775_);
  and (_20781_, _07962_, _08994_);
  or (_20782_, _20781_, _20736_);
  or (_20784_, _20782_, _06276_);
  and (_20785_, _20784_, _20780_);
  or (_20786_, _20785_, _06474_);
  and (_20787_, _14744_, _07962_);
  or (_20788_, _20787_, _20736_);
  or (_20789_, _20788_, _07282_);
  and (_20790_, _20789_, _07284_);
  and (_20791_, _20790_, _20786_);
  and (_20792_, _11221_, _07962_);
  or (_20793_, _20792_, _20736_);
  and (_20795_, _20793_, _06582_);
  or (_20796_, _20795_, _20791_);
  and (_20797_, _20796_, _07279_);
  or (_20798_, _20736_, _08433_);
  and (_20799_, _20782_, _06478_);
  and (_20800_, _20799_, _20798_);
  or (_20801_, _20800_, _20797_);
  and (_20802_, _20801_, _07276_);
  and (_20803_, _20746_, _06569_);
  and (_20804_, _20803_, _20798_);
  or (_20805_, _20804_, _06479_);
  or (_20806_, _20805_, _20802_);
  and (_20807_, _14741_, _07962_);
  or (_20808_, _20736_, _09043_);
  or (_20809_, _20808_, _20807_);
  and (_20810_, _20809_, _09048_);
  and (_20811_, _20810_, _20806_);
  nor (_20812_, _11220_, _11493_);
  or (_20813_, _20812_, _20736_);
  and (_20814_, _20813_, _06572_);
  or (_20817_, _20814_, _20811_);
  and (_20818_, _20817_, _07037_);
  and (_20819_, _20742_, _06606_);
  or (_20820_, _20819_, _06195_);
  or (_20821_, _20820_, _20818_);
  and (_20822_, _14917_, _07962_);
  or (_20823_, _20736_, _06196_);
  or (_20824_, _20823_, _20822_);
  and (_20825_, _20824_, _01375_);
  and (_20826_, _20825_, _20821_);
  or (_20828_, _20826_, _20735_);
  and (_42923_, _20828_, _42545_);
  and (_20829_, _11493_, \uc8051golden_1.DPL [3]);
  nor (_20830_, _11493_, _07775_);
  or (_20831_, _20830_, _20829_);
  or (_20832_, _20831_, _06293_);
  and (_20833_, _14947_, _07962_);
  or (_20834_, _20833_, _20829_);
  or (_20835_, _20834_, _07210_);
  and (_20836_, _07962_, \uc8051golden_1.ACC [3]);
  or (_20838_, _20836_, _20829_);
  and (_20839_, _20838_, _07199_);
  and (_20840_, _07200_, \uc8051golden_1.DPL [3]);
  or (_20841_, _20840_, _06401_);
  or (_20842_, _20841_, _20839_);
  and (_20843_, _20842_, _07221_);
  and (_20844_, _20843_, _20835_);
  and (_20845_, _20831_, _06399_);
  or (_20846_, _20845_, _06406_);
  or (_20847_, _20846_, _20844_);
  or (_20849_, _20838_, _06414_);
  and (_20850_, _20849_, _11512_);
  and (_20851_, _20850_, _20847_);
  nor (_20852_, _11517_, \uc8051golden_1.DPL [3]);
  nor (_20853_, _20852_, _11518_);
  and (_20854_, _20853_, _11511_);
  or (_20855_, _20854_, _20851_);
  and (_20856_, _20855_, _06473_);
  nor (_20857_, _06562_, _06473_);
  or (_20858_, _20857_, _10059_);
  or (_20860_, _20858_, _20856_);
  and (_20861_, _20860_, _20832_);
  or (_20862_, _20861_, _06281_);
  and (_20863_, _07962_, _09443_);
  or (_20864_, _20829_, _06282_);
  or (_20865_, _20864_, _20863_);
  and (_20866_, _20865_, _06279_);
  and (_20867_, _20866_, _20862_);
  and (_20868_, _15039_, _07962_);
  or (_20869_, _20868_, _20829_);
  and (_20871_, _20869_, _06015_);
  or (_20872_, _20871_, _06275_);
  or (_20873_, _20872_, _20867_);
  and (_20874_, _07962_, _08815_);
  or (_20875_, _20874_, _20829_);
  or (_20876_, _20875_, _06276_);
  and (_20877_, _20876_, _20873_);
  or (_20878_, _20877_, _06474_);
  and (_20879_, _14934_, _07962_);
  or (_20880_, _20879_, _20829_);
  or (_20882_, _20880_, _07282_);
  and (_20883_, _20882_, _07284_);
  and (_20884_, _20883_, _20878_);
  and (_20885_, _12535_, _07962_);
  or (_20886_, _20885_, _20829_);
  and (_20887_, _20886_, _06582_);
  or (_20888_, _20887_, _20884_);
  and (_20889_, _20888_, _07279_);
  or (_20890_, _20829_, _08389_);
  and (_20891_, _20875_, _06478_);
  and (_20893_, _20891_, _20890_);
  or (_20894_, _20893_, _20889_);
  and (_20895_, _20894_, _07276_);
  and (_20896_, _20838_, _06569_);
  and (_20897_, _20896_, _20890_);
  or (_20898_, _20897_, _06479_);
  or (_20899_, _20898_, _20895_);
  and (_20900_, _14931_, _07962_);
  or (_20901_, _20829_, _09043_);
  or (_20902_, _20901_, _20900_);
  and (_20904_, _20902_, _09048_);
  and (_20905_, _20904_, _20899_);
  nor (_20906_, _11218_, _11493_);
  or (_20907_, _20906_, _20829_);
  and (_20908_, _20907_, _06572_);
  or (_20909_, _20908_, _06606_);
  or (_20910_, _20909_, _20905_);
  or (_20911_, _20834_, _07037_);
  and (_20912_, _20911_, _06196_);
  and (_20913_, _20912_, _20910_);
  and (_20915_, _15113_, _07962_);
  or (_20916_, _20915_, _20829_);
  and (_20917_, _20916_, _06195_);
  or (_20918_, _20917_, _01379_);
  or (_20919_, _20918_, _20913_);
  or (_20920_, _01375_, \uc8051golden_1.DPL [3]);
  and (_20921_, _20920_, _42545_);
  and (_42924_, _20921_, _20919_);
  and (_20922_, _11493_, \uc8051golden_1.DPL [4]);
  nor (_20923_, _11493_, _08301_);
  or (_20925_, _20923_, _20922_);
  or (_20926_, _20925_, _06293_);
  and (_20927_, _15130_, _07962_);
  or (_20928_, _20927_, _20922_);
  or (_20929_, _20928_, _07210_);
  and (_20930_, _07962_, \uc8051golden_1.ACC [4]);
  or (_20931_, _20930_, _20922_);
  and (_20932_, _20931_, _07199_);
  and (_20933_, _07200_, \uc8051golden_1.DPL [4]);
  or (_20934_, _20933_, _06401_);
  or (_20935_, _20934_, _20932_);
  and (_20936_, _20935_, _07221_);
  and (_20937_, _20936_, _20929_);
  and (_20938_, _20925_, _06399_);
  or (_20939_, _20938_, _06406_);
  or (_20940_, _20939_, _20937_);
  or (_20941_, _20931_, _06414_);
  and (_20942_, _20941_, _11512_);
  and (_20943_, _20942_, _20940_);
  nor (_20944_, _11518_, \uc8051golden_1.DPL [4]);
  nor (_20947_, _20944_, _11519_);
  and (_20948_, _20947_, _11511_);
  or (_20949_, _20948_, _20943_);
  and (_20950_, _20949_, _06473_);
  nor (_20951_, _08882_, _06473_);
  or (_20952_, _20951_, _10059_);
  or (_20953_, _20952_, _20950_);
  and (_20954_, _20953_, _20926_);
  or (_20955_, _20954_, _06281_);
  and (_20956_, _07962_, _09442_);
  or (_20958_, _20922_, _06282_);
  or (_20959_, _20958_, _20956_);
  and (_20960_, _20959_, _06279_);
  and (_20961_, _20960_, _20955_);
  and (_20962_, _15243_, _07962_);
  or (_20963_, _20962_, _20922_);
  and (_20964_, _20963_, _06015_);
  or (_20965_, _20964_, _06275_);
  or (_20966_, _20965_, _20961_);
  and (_20967_, _08883_, _07962_);
  or (_20969_, _20967_, _20922_);
  or (_20970_, _20969_, _06276_);
  and (_20971_, _20970_, _20966_);
  or (_20972_, _20971_, _06474_);
  and (_20973_, _15135_, _07962_);
  or (_20974_, _20973_, _20922_);
  or (_20975_, _20974_, _07282_);
  and (_20976_, _20975_, _07284_);
  and (_20977_, _20976_, _20972_);
  and (_20978_, _11216_, _07962_);
  or (_20980_, _20978_, _20922_);
  and (_20981_, _20980_, _06582_);
  or (_20982_, _20981_, _20977_);
  and (_20983_, _20982_, _07279_);
  or (_20984_, _20922_, _08345_);
  and (_20985_, _20969_, _06478_);
  and (_20986_, _20985_, _20984_);
  or (_20987_, _20986_, _20983_);
  and (_20988_, _20987_, _07276_);
  and (_20989_, _20931_, _06569_);
  and (_20991_, _20989_, _20984_);
  or (_20992_, _20991_, _06479_);
  or (_20993_, _20992_, _20988_);
  and (_20994_, _15134_, _07962_);
  or (_20995_, _20922_, _09043_);
  or (_20996_, _20995_, _20994_);
  and (_20997_, _20996_, _09048_);
  and (_20998_, _20997_, _20993_);
  nor (_20999_, _11215_, _11493_);
  or (_21000_, _20999_, _20922_);
  and (_21002_, _21000_, _06572_);
  or (_21003_, _21002_, _06606_);
  or (_21004_, _21003_, _20998_);
  or (_21005_, _20928_, _07037_);
  and (_21006_, _21005_, _06196_);
  and (_21007_, _21006_, _21004_);
  and (_21008_, _15315_, _07962_);
  or (_21009_, _21008_, _20922_);
  and (_21010_, _21009_, _06195_);
  or (_21011_, _21010_, _01379_);
  or (_21013_, _21011_, _21007_);
  or (_21014_, _01375_, \uc8051golden_1.DPL [4]);
  and (_21015_, _21014_, _42545_);
  and (_42925_, _21015_, _21013_);
  and (_21016_, _11493_, \uc8051golden_1.DPL [5]);
  nor (_21017_, _11493_, _08207_);
  or (_21018_, _21017_, _21016_);
  or (_21019_, _21018_, _06293_);
  and (_21020_, _15348_, _07962_);
  or (_21021_, _21020_, _21016_);
  or (_21023_, _21021_, _07210_);
  and (_21024_, _07962_, \uc8051golden_1.ACC [5]);
  or (_21025_, _21024_, _21016_);
  and (_21026_, _21025_, _07199_);
  and (_21027_, _07200_, \uc8051golden_1.DPL [5]);
  or (_21028_, _21027_, _06401_);
  or (_21029_, _21028_, _21026_);
  and (_21030_, _21029_, _07221_);
  and (_21031_, _21030_, _21023_);
  and (_21032_, _21018_, _06399_);
  or (_21034_, _21032_, _06406_);
  or (_21035_, _21034_, _21031_);
  or (_21036_, _21025_, _06414_);
  and (_21037_, _21036_, _11512_);
  and (_21038_, _21037_, _21035_);
  nor (_21039_, _11519_, \uc8051golden_1.DPL [5]);
  nor (_21040_, _21039_, _11520_);
  and (_21041_, _21040_, _11511_);
  or (_21042_, _21041_, _21038_);
  and (_21043_, _21042_, _06473_);
  nor (_21045_, _08917_, _06473_);
  or (_21046_, _21045_, _10059_);
  or (_21047_, _21046_, _21043_);
  and (_21048_, _21047_, _21019_);
  or (_21049_, _21048_, _06281_);
  and (_21050_, _07962_, _09441_);
  or (_21051_, _21016_, _06282_);
  or (_21052_, _21051_, _21050_);
  and (_21053_, _21052_, _06279_);
  and (_21054_, _21053_, _21049_);
  and (_21056_, _15446_, _07962_);
  or (_21057_, _21056_, _21016_);
  and (_21058_, _21057_, _06015_);
  or (_21059_, _21058_, _06275_);
  or (_21060_, _21059_, _21054_);
  and (_21061_, _08958_, _07962_);
  or (_21062_, _21061_, _21016_);
  or (_21063_, _21062_, _06276_);
  and (_21064_, _21063_, _21060_);
  or (_21065_, _21064_, _06474_);
  and (_21067_, _15338_, _07962_);
  or (_21068_, _21067_, _21016_);
  or (_21069_, _21068_, _07282_);
  and (_21070_, _21069_, _07284_);
  and (_21071_, _21070_, _21065_);
  and (_21072_, _12542_, _07962_);
  or (_21073_, _21072_, _21016_);
  and (_21074_, _21073_, _06582_);
  or (_21075_, _21074_, _21071_);
  and (_21076_, _21075_, _07279_);
  or (_21078_, _21016_, _08256_);
  and (_21079_, _21062_, _06478_);
  and (_21080_, _21079_, _21078_);
  or (_21081_, _21080_, _21076_);
  and (_21082_, _21081_, _07276_);
  and (_21083_, _21025_, _06569_);
  and (_21084_, _21083_, _21078_);
  or (_21085_, _21084_, _06479_);
  or (_21086_, _21085_, _21082_);
  and (_21087_, _15335_, _07962_);
  or (_21089_, _21016_, _09043_);
  or (_21090_, _21089_, _21087_);
  and (_21091_, _21090_, _09048_);
  and (_21092_, _21091_, _21086_);
  nor (_21093_, _11212_, _11493_);
  or (_21094_, _21093_, _21016_);
  and (_21095_, _21094_, _06572_);
  or (_21096_, _21095_, _06606_);
  or (_21097_, _21096_, _21092_);
  or (_21098_, _21021_, _07037_);
  and (_21100_, _21098_, _06196_);
  and (_21101_, _21100_, _21097_);
  and (_21102_, _15509_, _07962_);
  or (_21103_, _21102_, _21016_);
  and (_21104_, _21103_, _06195_);
  or (_21105_, _21104_, _01379_);
  or (_21106_, _21105_, _21101_);
  or (_21107_, _01375_, \uc8051golden_1.DPL [5]);
  and (_21108_, _21107_, _42545_);
  and (_42926_, _21108_, _21106_);
  and (_21109_, _11493_, \uc8051golden_1.DPL [6]);
  nor (_21110_, _11493_, _08118_);
  or (_21111_, _21110_, _21109_);
  or (_21112_, _21111_, _06293_);
  and (_21113_, _15550_, _07962_);
  or (_21114_, _21113_, _21109_);
  or (_21115_, _21114_, _07210_);
  and (_21116_, _07962_, \uc8051golden_1.ACC [6]);
  or (_21117_, _21116_, _21109_);
  and (_21118_, _21117_, _07199_);
  and (_21121_, _07200_, \uc8051golden_1.DPL [6]);
  or (_21122_, _21121_, _06401_);
  or (_21123_, _21122_, _21118_);
  and (_21124_, _21123_, _07221_);
  and (_21125_, _21124_, _21115_);
  and (_21126_, _21111_, _06399_);
  or (_21127_, _21126_, _06406_);
  or (_21128_, _21127_, _21125_);
  or (_21129_, _21117_, _06414_);
  and (_21130_, _21129_, _11512_);
  and (_21132_, _21130_, _21128_);
  nor (_21133_, _11520_, \uc8051golden_1.DPL [6]);
  nor (_21134_, _21133_, _11521_);
  and (_21135_, _21134_, _11511_);
  or (_21136_, _21135_, _21132_);
  and (_21137_, _21136_, _06473_);
  nor (_21138_, _08850_, _06473_);
  or (_21139_, _21138_, _10059_);
  or (_21140_, _21139_, _21137_);
  and (_21141_, _21140_, _21112_);
  or (_21143_, _21141_, _06281_);
  and (_21144_, _07962_, _09440_);
  or (_21145_, _21109_, _06282_);
  or (_21146_, _21145_, _21144_);
  and (_21147_, _21146_, _06279_);
  and (_21148_, _21147_, _21143_);
  and (_21149_, _15639_, _07962_);
  or (_21150_, _21149_, _21109_);
  and (_21151_, _21150_, _06015_);
  or (_21152_, _21151_, _06275_);
  or (_21154_, _21152_, _21148_);
  and (_21155_, _15646_, _07962_);
  or (_21156_, _21155_, _21109_);
  or (_21157_, _21156_, _06276_);
  and (_21158_, _21157_, _21154_);
  or (_21159_, _21158_, _06474_);
  and (_21160_, _15531_, _07962_);
  or (_21161_, _21160_, _21109_);
  or (_21162_, _21161_, _07282_);
  and (_21163_, _21162_, _07284_);
  and (_21165_, _21163_, _21159_);
  and (_21166_, _11210_, _07962_);
  or (_21167_, _21166_, _21109_);
  and (_21168_, _21167_, _06582_);
  or (_21169_, _21168_, _21165_);
  and (_21170_, _21169_, _07279_);
  or (_21171_, _21109_, _08162_);
  and (_21172_, _21156_, _06478_);
  and (_21173_, _21172_, _21171_);
  or (_21174_, _21173_, _21170_);
  and (_21176_, _21174_, _07276_);
  and (_21177_, _21117_, _06569_);
  and (_21178_, _21177_, _21171_);
  or (_21179_, _21178_, _06479_);
  or (_21180_, _21179_, _21176_);
  and (_21181_, _15528_, _07962_);
  or (_21182_, _21109_, _09043_);
  or (_21183_, _21182_, _21181_);
  and (_21184_, _21183_, _09048_);
  and (_21185_, _21184_, _21180_);
  nor (_21187_, _11209_, _11493_);
  or (_21188_, _21187_, _21109_);
  and (_21189_, _21188_, _06572_);
  or (_21190_, _21189_, _06606_);
  or (_21191_, _21190_, _21185_);
  or (_21192_, _21114_, _07037_);
  and (_21193_, _21192_, _06196_);
  and (_21194_, _21193_, _21191_);
  and (_21195_, _15713_, _07962_);
  or (_21196_, _21195_, _21109_);
  and (_21198_, _21196_, _06195_);
  or (_21199_, _21198_, _01379_);
  or (_21200_, _21199_, _21194_);
  or (_21201_, _01375_, \uc8051golden_1.DPL [6]);
  and (_21202_, _21201_, _42545_);
  and (_42927_, _21202_, _21200_);
  nor (_21203_, _01375_, _12642_);
  nor (_21204_, _07966_, _12642_);
  and (_21205_, _07966_, \uc8051golden_1.ACC [0]);
  and (_21206_, _21205_, _08521_);
  or (_21208_, _21206_, _21204_);
  or (_21209_, _21208_, _07276_);
  and (_21210_, _08249_, _07473_);
  or (_21211_, _21210_, _21204_);
  or (_21212_, _21211_, _06293_);
  or (_21213_, _21211_, _07221_);
  nor (_21214_, _08521_, _11589_);
  or (_21215_, _21214_, _21204_);
  and (_21216_, _21215_, _06401_);
  nor (_21217_, _07199_, _12642_);
  or (_21219_, _21205_, _21204_);
  and (_21220_, _21219_, _07199_);
  or (_21221_, _21220_, _21217_);
  and (_21222_, _21221_, _07210_);
  or (_21223_, _21222_, _06399_);
  or (_21224_, _21223_, _21216_);
  and (_21225_, _21224_, _21213_);
  or (_21226_, _21225_, _06406_);
  or (_21227_, _21219_, _06414_);
  and (_21228_, _21227_, _11512_);
  and (_21230_, _21228_, _21226_);
  nor (_21231_, _11523_, \uc8051golden_1.DPH [0]);
  nor (_21232_, _21231_, _11610_);
  and (_21233_, _21232_, _11511_);
  or (_21234_, _21233_, _21230_);
  and (_21235_, _21234_, _06473_);
  nor (_21236_, _06840_, _06473_);
  or (_21237_, _21236_, _10059_);
  or (_21238_, _21237_, _21235_);
  and (_21239_, _21238_, _21212_);
  or (_21241_, _21239_, _06281_);
  or (_21242_, _21204_, _06282_);
  and (_21243_, _07966_, _09446_);
  or (_21244_, _21243_, _21242_);
  and (_21245_, _21244_, _21241_);
  or (_21246_, _21245_, _06015_);
  and (_21247_, _14426_, _08249_);
  or (_21248_, _21204_, _06279_);
  or (_21249_, _21248_, _21247_);
  and (_21250_, _21249_, _06276_);
  and (_21252_, _21250_, _21246_);
  and (_21253_, _07966_, _08817_);
  or (_21254_, _21253_, _21204_);
  and (_21255_, _21254_, _06275_);
  or (_21256_, _21255_, _06474_);
  or (_21257_, _21256_, _21252_);
  and (_21258_, _14324_, _07966_);
  or (_21259_, _21258_, _21204_);
  or (_21260_, _21259_, _07282_);
  and (_21261_, _21260_, _07284_);
  and (_21263_, _21261_, _21257_);
  nor (_21264_, _12538_, _11589_);
  or (_21265_, _21264_, _21204_);
  nor (_21266_, _21206_, _07284_);
  and (_21267_, _21266_, _21265_);
  or (_21268_, _21267_, _21263_);
  and (_21269_, _21268_, _07279_);
  nand (_21270_, _21254_, _06478_);
  nor (_21271_, _21270_, _21214_);
  or (_21272_, _21271_, _06569_);
  or (_21274_, _21272_, _21269_);
  and (_21275_, _21274_, _21209_);
  or (_21276_, _21275_, _06479_);
  and (_21277_, _14320_, _07966_);
  or (_21278_, _21277_, _21204_);
  or (_21279_, _21278_, _09043_);
  and (_21280_, _21279_, _09048_);
  and (_21281_, _21280_, _21276_);
  and (_21282_, _21265_, _06572_);
  or (_21283_, _21282_, _19434_);
  or (_21285_, _21283_, _21281_);
  or (_21286_, _21215_, _06700_);
  and (_21287_, _21286_, _01375_);
  and (_21288_, _21287_, _21285_);
  or (_21289_, _21288_, _21203_);
  and (_42928_, _21289_, _42545_);
  not (_21290_, \uc8051golden_1.DPH [1]);
  nor (_21291_, _07966_, _21290_);
  nor (_21292_, _11223_, _11589_);
  or (_21293_, _21292_, _21291_);
  or (_21295_, _21293_, _09048_);
  or (_21296_, _07966_, \uc8051golden_1.DPH [1]);
  and (_21297_, _21296_, _06275_);
  nand (_21298_, _08249_, _07090_);
  and (_21299_, _21298_, _21297_);
  nor (_21300_, _11589_, _07196_);
  or (_21301_, _21300_, _21291_);
  or (_21302_, _21301_, _06293_);
  nor (_21303_, _11610_, \uc8051golden_1.DPH [1]);
  nor (_21304_, _21303_, _11611_);
  and (_21305_, _21304_, _11511_);
  and (_21306_, _14532_, _08249_);
  not (_21307_, _21306_);
  and (_21308_, _21307_, _21296_);
  or (_21309_, _21308_, _07210_);
  and (_21310_, _07966_, \uc8051golden_1.ACC [1]);
  or (_21311_, _21310_, _21291_);
  and (_21312_, _21311_, _07199_);
  nor (_21313_, _07199_, _21290_);
  or (_21314_, _21313_, _06401_);
  or (_21317_, _21314_, _21312_);
  and (_21318_, _21317_, _07221_);
  and (_21319_, _21318_, _21309_);
  and (_21320_, _21301_, _06399_);
  or (_21321_, _21320_, _06406_);
  or (_21322_, _21321_, _21319_);
  or (_21323_, _21311_, _06414_);
  and (_21324_, _21323_, _11512_);
  and (_21325_, _21324_, _21322_);
  or (_21326_, _21325_, _21305_);
  and (_21328_, _21326_, _06473_);
  nor (_21329_, _06473_, _06228_);
  or (_21330_, _21329_, _10059_);
  or (_21331_, _21330_, _21328_);
  and (_21332_, _21331_, _21302_);
  or (_21333_, _21332_, _06281_);
  and (_21334_, _21333_, _06279_);
  and (_21335_, _07966_, _09445_);
  or (_21336_, _21335_, _21291_);
  or (_21337_, _21336_, _06282_);
  and (_21339_, _21337_, _21334_);
  and (_21340_, _14615_, _07966_);
  or (_21341_, _21340_, _21291_);
  and (_21342_, _21341_, _06015_);
  or (_21343_, _21342_, _21339_);
  and (_21344_, _21343_, _06276_);
  or (_21345_, _21344_, _21299_);
  and (_21346_, _21345_, _07282_);
  or (_21347_, _14507_, _11589_);
  and (_21348_, _21296_, _06474_);
  and (_21350_, _21348_, _21347_);
  or (_21351_, _21350_, _06582_);
  or (_21352_, _21351_, _21346_);
  nand (_21353_, _11222_, _08249_);
  and (_21354_, _21353_, _21293_);
  or (_21355_, _21354_, _07284_);
  and (_21356_, _21355_, _07279_);
  and (_21357_, _21356_, _21352_);
  or (_21358_, _14505_, _11589_);
  and (_21359_, _21296_, _06478_);
  and (_21361_, _21359_, _21358_);
  or (_21362_, _21361_, _06569_);
  or (_21363_, _21362_, _21357_);
  nor (_21364_, _21291_, _07276_);
  nand (_21365_, _21364_, _21353_);
  and (_21366_, _21365_, _09043_);
  and (_21367_, _21366_, _21363_);
  or (_21368_, _21298_, _08477_);
  and (_21369_, _21296_, _06479_);
  and (_21370_, _21369_, _21368_);
  or (_21372_, _21370_, _06572_);
  or (_21373_, _21372_, _21367_);
  and (_21374_, _21373_, _21295_);
  or (_21375_, _21374_, _06606_);
  or (_21376_, _21308_, _07037_);
  and (_21377_, _21376_, _06196_);
  and (_21378_, _21377_, _21375_);
  or (_21379_, _21306_, _21291_);
  and (_21380_, _21379_, _06195_);
  or (_21381_, _21380_, _01379_);
  or (_21383_, _21381_, _21378_);
  or (_21384_, _01375_, \uc8051golden_1.DPH [1]);
  and (_21385_, _21384_, _42545_);
  and (_42929_, _21385_, _21383_);
  not (_21386_, \uc8051golden_1.DPH [2]);
  nor (_21387_, _01375_, _21386_);
  nor (_21388_, _07966_, _21386_);
  and (_21389_, _07966_, _09444_);
  or (_21390_, _21389_, _21388_);
  and (_21391_, _21390_, _06281_);
  or (_21393_, _11611_, \uc8051golden_1.DPH [2]);
  nor (_21394_, _11612_, _11512_);
  and (_21395_, _21394_, _21393_);
  and (_21396_, _14754_, _08249_);
  or (_21397_, _21396_, _21388_);
  or (_21398_, _21397_, _07210_);
  and (_21399_, _07966_, \uc8051golden_1.ACC [2]);
  or (_21400_, _21399_, _21388_);
  and (_21401_, _21400_, _07199_);
  nor (_21402_, _07199_, _21386_);
  or (_21404_, _21402_, _06401_);
  or (_21405_, _21404_, _21401_);
  and (_21406_, _21405_, _07221_);
  and (_21407_, _21406_, _21398_);
  nor (_21408_, _11589_, _07623_);
  or (_21409_, _21408_, _21388_);
  and (_21410_, _21409_, _06399_);
  or (_21411_, _21410_, _06406_);
  or (_21412_, _21411_, _21407_);
  or (_21413_, _21400_, _06414_);
  and (_21415_, _21413_, _11512_);
  and (_21416_, _21415_, _21412_);
  or (_21417_, _21416_, _21395_);
  and (_21418_, _21417_, _06473_);
  nor (_21419_, _06693_, _06473_);
  or (_21420_, _21419_, _10059_);
  or (_21421_, _21420_, _21418_);
  or (_21422_, _21409_, _06293_);
  and (_21423_, _21422_, _06282_);
  and (_21424_, _21423_, _21421_);
  or (_21426_, _21424_, _06015_);
  or (_21427_, _21426_, _21391_);
  and (_21428_, _14848_, _08249_);
  or (_21429_, _21388_, _06279_);
  or (_21430_, _21429_, _21428_);
  and (_21431_, _21430_, _06276_);
  and (_21432_, _21431_, _21427_);
  and (_21433_, _07966_, _08994_);
  or (_21434_, _21433_, _21388_);
  and (_21435_, _21434_, _06275_);
  or (_21437_, _21435_, _06474_);
  or (_21438_, _21437_, _21432_);
  and (_21439_, _14744_, _07966_);
  or (_21440_, _21439_, _21388_);
  or (_21441_, _21440_, _07282_);
  and (_21442_, _21441_, _07284_);
  and (_21443_, _21442_, _21438_);
  and (_21444_, _11221_, _07966_);
  or (_21445_, _21444_, _21388_);
  and (_21446_, _21445_, _06582_);
  or (_21448_, _21446_, _21443_);
  and (_21449_, _21448_, _07279_);
  or (_21450_, _21388_, _08433_);
  and (_21451_, _21434_, _06478_);
  and (_21452_, _21451_, _21450_);
  or (_21453_, _21452_, _21449_);
  and (_21454_, _21453_, _07276_);
  and (_21455_, _21400_, _06569_);
  and (_21456_, _21455_, _21450_);
  or (_21457_, _21456_, _06479_);
  or (_21459_, _21457_, _21454_);
  and (_21460_, _14741_, _08249_);
  or (_21461_, _21388_, _09043_);
  or (_21462_, _21461_, _21460_);
  and (_21463_, _21462_, _09048_);
  and (_21464_, _21463_, _21459_);
  nor (_21465_, _11220_, _11589_);
  or (_21466_, _21465_, _21388_);
  and (_21467_, _21466_, _06572_);
  or (_21468_, _21467_, _21464_);
  and (_21470_, _21468_, _07037_);
  and (_21471_, _21397_, _06606_);
  or (_21472_, _21471_, _06195_);
  or (_21473_, _21472_, _21470_);
  and (_21474_, _14917_, _08249_);
  or (_21475_, _21388_, _06196_);
  or (_21476_, _21475_, _21474_);
  and (_21477_, _21476_, _01375_);
  and (_21478_, _21477_, _21473_);
  or (_21479_, _21478_, _21387_);
  and (_42930_, _21479_, _42545_);
  and (_21481_, _11589_, \uc8051golden_1.DPH [3]);
  nor (_21482_, _11589_, _07775_);
  or (_21483_, _21482_, _21481_);
  or (_21484_, _21483_, _06293_);
  or (_21485_, _11612_, \uc8051golden_1.DPH [3]);
  nor (_21486_, _11613_, _11512_);
  and (_21487_, _21486_, _21485_);
  and (_21488_, _14947_, _08249_);
  or (_21489_, _21488_, _21481_);
  or (_21491_, _21489_, _07210_);
  and (_21492_, _07966_, \uc8051golden_1.ACC [3]);
  or (_21493_, _21492_, _21481_);
  and (_21494_, _21493_, _07199_);
  and (_21495_, _07200_, \uc8051golden_1.DPH [3]);
  or (_21496_, _21495_, _06401_);
  or (_21497_, _21496_, _21494_);
  and (_21498_, _21497_, _07221_);
  and (_21499_, _21498_, _21491_);
  and (_21500_, _21483_, _06399_);
  or (_21502_, _21500_, _06406_);
  or (_21503_, _21502_, _21499_);
  or (_21504_, _21493_, _06414_);
  and (_21505_, _21504_, _11512_);
  and (_21506_, _21505_, _21503_);
  or (_21507_, _21506_, _21487_);
  and (_21508_, _21507_, _06473_);
  nor (_21509_, _06473_, _06372_);
  or (_21510_, _21509_, _10059_);
  or (_21511_, _21510_, _21508_);
  and (_21513_, _21511_, _21484_);
  or (_21514_, _21513_, _06281_);
  or (_21515_, _21481_, _06282_);
  and (_21516_, _07966_, _09443_);
  or (_21517_, _21516_, _21515_);
  and (_21518_, _21517_, _06279_);
  and (_21519_, _21518_, _21514_);
  and (_21520_, _15039_, _07966_);
  or (_21521_, _21520_, _21481_);
  and (_21522_, _21521_, _06015_);
  or (_21524_, _21522_, _06275_);
  or (_21525_, _21524_, _21519_);
  and (_21526_, _07966_, _08815_);
  or (_21527_, _21526_, _21481_);
  or (_21528_, _21527_, _06276_);
  and (_21529_, _21528_, _21525_);
  or (_21530_, _21529_, _06474_);
  and (_21531_, _14934_, _07966_);
  or (_21532_, _21531_, _21481_);
  or (_21533_, _21532_, _07282_);
  and (_21535_, _21533_, _07284_);
  and (_21536_, _21535_, _21530_);
  and (_21537_, _12535_, _07966_);
  or (_21538_, _21537_, _21481_);
  and (_21539_, _21538_, _06582_);
  or (_21540_, _21539_, _21536_);
  and (_21541_, _21540_, _07279_);
  or (_21542_, _21481_, _08389_);
  and (_21543_, _21527_, _06478_);
  and (_21544_, _21543_, _21542_);
  or (_21546_, _21544_, _21541_);
  and (_21547_, _21546_, _07276_);
  and (_21548_, _21493_, _06569_);
  and (_21549_, _21548_, _21542_);
  or (_21550_, _21549_, _06479_);
  or (_21551_, _21550_, _21547_);
  and (_21552_, _14931_, _08249_);
  or (_21553_, _21481_, _09043_);
  or (_21554_, _21553_, _21552_);
  and (_21555_, _21554_, _09048_);
  and (_21557_, _21555_, _21551_);
  nor (_21558_, _11218_, _11589_);
  or (_21559_, _21558_, _21481_);
  and (_21560_, _21559_, _06572_);
  or (_21561_, _21560_, _06606_);
  or (_21562_, _21561_, _21557_);
  or (_21563_, _21489_, _07037_);
  and (_21564_, _21563_, _06196_);
  and (_21565_, _21564_, _21562_);
  and (_21566_, _15113_, _08249_);
  or (_21568_, _21566_, _21481_);
  and (_21569_, _21568_, _06195_);
  or (_21570_, _21569_, _01379_);
  or (_21571_, _21570_, _21565_);
  or (_21572_, _01375_, \uc8051golden_1.DPH [3]);
  and (_21573_, _21572_, _42545_);
  and (_42931_, _21573_, _21571_);
  not (_21574_, \uc8051golden_1.DPH [4]);
  nor (_21575_, _07966_, _21574_);
  nor (_21576_, _11589_, _08301_);
  or (_21578_, _21576_, _21575_);
  or (_21579_, _21578_, _06293_);
  and (_21580_, _15130_, _08249_);
  or (_21581_, _21580_, _21575_);
  or (_21582_, _21581_, _07210_);
  and (_21583_, _07966_, \uc8051golden_1.ACC [4]);
  or (_21584_, _21583_, _21575_);
  and (_21585_, _21584_, _07199_);
  nor (_21586_, _07199_, _21574_);
  or (_21587_, _21586_, _06401_);
  or (_21589_, _21587_, _21585_);
  and (_21590_, _21589_, _07221_);
  and (_21591_, _21590_, _21582_);
  and (_21592_, _21578_, _06399_);
  or (_21593_, _21592_, _06406_);
  or (_21594_, _21593_, _21591_);
  or (_21595_, _21584_, _06414_);
  and (_21596_, _21595_, _11512_);
  and (_21597_, _21596_, _21594_);
  or (_21598_, _11613_, \uc8051golden_1.DPH [4]);
  nor (_21600_, _11614_, _11512_);
  and (_21601_, _21600_, _21598_);
  or (_21602_, _21601_, _21597_);
  and (_21603_, _21602_, _06473_);
  nor (_21604_, _06473_, _06265_);
  or (_21605_, _21604_, _10059_);
  or (_21606_, _21605_, _21603_);
  and (_21607_, _21606_, _21579_);
  or (_21608_, _21607_, _06281_);
  or (_21609_, _21575_, _06282_);
  and (_21611_, _07966_, _09442_);
  or (_21612_, _21611_, _21609_);
  and (_21613_, _21612_, _06279_);
  and (_21614_, _21613_, _21608_);
  and (_21615_, _15243_, _07966_);
  or (_21616_, _21615_, _21575_);
  and (_21617_, _21616_, _06015_);
  or (_21618_, _21617_, _06275_);
  or (_21619_, _21618_, _21614_);
  and (_21620_, _08883_, _07966_);
  or (_21622_, _21620_, _21575_);
  or (_21623_, _21622_, _06276_);
  and (_21624_, _21623_, _21619_);
  or (_21625_, _21624_, _06474_);
  and (_21626_, _15135_, _07966_);
  or (_21627_, _21626_, _21575_);
  or (_21628_, _21627_, _07282_);
  and (_21629_, _21628_, _07284_);
  and (_21630_, _21629_, _21625_);
  and (_21631_, _11216_, _07966_);
  or (_21633_, _21631_, _21575_);
  and (_21634_, _21633_, _06582_);
  or (_21635_, _21634_, _21630_);
  and (_21636_, _21635_, _07279_);
  or (_21637_, _21575_, _08345_);
  and (_21638_, _21622_, _06478_);
  and (_21639_, _21638_, _21637_);
  or (_21640_, _21639_, _21636_);
  and (_21641_, _21640_, _07276_);
  and (_21642_, _21584_, _06569_);
  and (_21644_, _21642_, _21637_);
  or (_21645_, _21644_, _06479_);
  or (_21646_, _21645_, _21641_);
  and (_21647_, _15134_, _08249_);
  or (_21648_, _21575_, _09043_);
  or (_21649_, _21648_, _21647_);
  and (_21650_, _21649_, _09048_);
  and (_21651_, _21650_, _21646_);
  nor (_21652_, _11215_, _11589_);
  or (_21653_, _21652_, _21575_);
  and (_21654_, _21653_, _06572_);
  or (_21655_, _21654_, _06606_);
  or (_21656_, _21655_, _21651_);
  or (_21657_, _21581_, _07037_);
  and (_21658_, _21657_, _06196_);
  and (_21659_, _21658_, _21656_);
  and (_21660_, _15315_, _08249_);
  or (_21661_, _21660_, _21575_);
  and (_21662_, _21661_, _06195_);
  or (_21663_, _21662_, _01379_);
  or (_21666_, _21663_, _21659_);
  or (_21667_, _01375_, \uc8051golden_1.DPH [4]);
  and (_21668_, _21667_, _42545_);
  and (_42932_, _21668_, _21666_);
  and (_21669_, _11589_, \uc8051golden_1.DPH [5]);
  nor (_21670_, _11589_, _08207_);
  or (_21671_, _21670_, _21669_);
  or (_21672_, _21671_, _06293_);
  and (_21673_, _15348_, _08249_);
  or (_21674_, _21673_, _21669_);
  or (_21676_, _21674_, _07210_);
  and (_21677_, _07966_, \uc8051golden_1.ACC [5]);
  or (_21678_, _21677_, _21669_);
  and (_21679_, _21678_, _07199_);
  and (_21680_, _07200_, \uc8051golden_1.DPH [5]);
  or (_21681_, _21680_, _06401_);
  or (_21682_, _21681_, _21679_);
  and (_21683_, _21682_, _07221_);
  and (_21684_, _21683_, _21676_);
  and (_21685_, _21671_, _06399_);
  or (_21687_, _21685_, _06406_);
  or (_21688_, _21687_, _21684_);
  or (_21689_, _21678_, _06414_);
  and (_21690_, _21689_, _11512_);
  and (_21691_, _21690_, _21688_);
  or (_21692_, _11614_, \uc8051golden_1.DPH [5]);
  nor (_21693_, _11615_, _11512_);
  and (_21694_, _21693_, _21692_);
  or (_21695_, _21694_, _21691_);
  and (_21696_, _21695_, _06473_);
  nor (_21698_, _06650_, _06473_);
  or (_21699_, _21698_, _10059_);
  or (_21700_, _21699_, _21696_);
  and (_21701_, _21700_, _21672_);
  or (_21702_, _21701_, _06281_);
  or (_21703_, _21669_, _06282_);
  and (_21704_, _07966_, _09441_);
  or (_21705_, _21704_, _21703_);
  and (_21706_, _21705_, _06279_);
  and (_21707_, _21706_, _21702_);
  and (_21709_, _15446_, _07966_);
  or (_21710_, _21709_, _21669_);
  and (_21711_, _21710_, _06015_);
  or (_21712_, _21711_, _06275_);
  or (_21713_, _21712_, _21707_);
  and (_21714_, _08958_, _07966_);
  or (_21715_, _21714_, _21669_);
  or (_21716_, _21715_, _06276_);
  and (_21717_, _21716_, _21713_);
  or (_21718_, _21717_, _06474_);
  and (_21720_, _15338_, _07966_);
  or (_21721_, _21720_, _21669_);
  or (_21722_, _21721_, _07282_);
  and (_21723_, _21722_, _07284_);
  and (_21724_, _21723_, _21718_);
  and (_21725_, _12542_, _07966_);
  or (_21726_, _21725_, _21669_);
  and (_21727_, _21726_, _06582_);
  or (_21728_, _21727_, _21724_);
  and (_21729_, _21728_, _07279_);
  or (_21731_, _21669_, _08256_);
  and (_21732_, _21715_, _06478_);
  and (_21733_, _21732_, _21731_);
  or (_21734_, _21733_, _21729_);
  and (_21735_, _21734_, _07276_);
  and (_21736_, _21678_, _06569_);
  and (_21737_, _21736_, _21731_);
  or (_21738_, _21737_, _06479_);
  or (_21739_, _21738_, _21735_);
  and (_21740_, _15335_, _08249_);
  or (_21742_, _21669_, _09043_);
  or (_21743_, _21742_, _21740_);
  and (_21744_, _21743_, _09048_);
  and (_21745_, _21744_, _21739_);
  nor (_21746_, _11212_, _11589_);
  or (_21747_, _21746_, _21669_);
  and (_21748_, _21747_, _06572_);
  or (_21749_, _21748_, _06606_);
  or (_21750_, _21749_, _21745_);
  or (_21751_, _21674_, _07037_);
  and (_21753_, _21751_, _06196_);
  and (_21754_, _21753_, _21750_);
  and (_21755_, _15509_, _08249_);
  or (_21756_, _21755_, _21669_);
  and (_21757_, _21756_, _06195_);
  or (_21758_, _21757_, _01379_);
  or (_21759_, _21758_, _21754_);
  or (_21760_, _01375_, \uc8051golden_1.DPH [5]);
  and (_21761_, _21760_, _42545_);
  and (_42934_, _21761_, _21759_);
  not (_21762_, \uc8051golden_1.DPH [6]);
  nor (_21763_, _07966_, _21762_);
  nor (_21764_, _11589_, _08118_);
  or (_21765_, _21764_, _21763_);
  or (_21766_, _21765_, _06293_);
  and (_21767_, _15550_, _08249_);
  or (_21768_, _21767_, _21763_);
  or (_21769_, _21768_, _07210_);
  and (_21770_, _07966_, \uc8051golden_1.ACC [6]);
  or (_21771_, _21770_, _21763_);
  and (_21774_, _21771_, _07199_);
  nor (_21775_, _07199_, _21762_);
  or (_21776_, _21775_, _06401_);
  or (_21777_, _21776_, _21774_);
  and (_21778_, _21777_, _07221_);
  and (_21779_, _21778_, _21769_);
  and (_21780_, _21765_, _06399_);
  or (_21781_, _21780_, _06406_);
  or (_21782_, _21781_, _21779_);
  or (_21783_, _21771_, _06414_);
  and (_21785_, _21783_, _11512_);
  and (_21786_, _21785_, _21782_);
  or (_21787_, _11615_, \uc8051golden_1.DPH [6]);
  nor (_21788_, _11616_, _11512_);
  and (_21789_, _21788_, _21787_);
  or (_21790_, _21789_, _21786_);
  and (_21791_, _21790_, _06473_);
  nor (_21792_, _06473_, _06340_);
  or (_21793_, _21792_, _10059_);
  or (_21794_, _21793_, _21791_);
  and (_21796_, _21794_, _21766_);
  or (_21797_, _21796_, _06281_);
  or (_21798_, _21763_, _06282_);
  and (_21799_, _07966_, _09440_);
  or (_21800_, _21799_, _21798_);
  and (_21801_, _21800_, _06279_);
  and (_21802_, _21801_, _21797_);
  and (_21803_, _15639_, _07966_);
  or (_21804_, _21803_, _21763_);
  and (_21805_, _21804_, _06015_);
  or (_21807_, _21805_, _06275_);
  or (_21808_, _21807_, _21802_);
  and (_21809_, _15646_, _07966_);
  or (_21810_, _21809_, _21763_);
  or (_21811_, _21810_, _06276_);
  and (_21812_, _21811_, _21808_);
  or (_21813_, _21812_, _06474_);
  and (_21814_, _15531_, _07966_);
  or (_21815_, _21814_, _21763_);
  or (_21816_, _21815_, _07282_);
  and (_21818_, _21816_, _07284_);
  and (_21819_, _21818_, _21813_);
  and (_21820_, _11210_, _07966_);
  or (_21821_, _21820_, _21763_);
  and (_21822_, _21821_, _06582_);
  or (_21823_, _21822_, _21819_);
  and (_21824_, _21823_, _07279_);
  or (_21825_, _21763_, _08162_);
  and (_21826_, _21810_, _06478_);
  and (_21827_, _21826_, _21825_);
  or (_21829_, _21827_, _21824_);
  and (_21830_, _21829_, _07276_);
  and (_21831_, _21771_, _06569_);
  and (_21832_, _21831_, _21825_);
  or (_21833_, _21832_, _06479_);
  or (_21834_, _21833_, _21830_);
  and (_21835_, _15528_, _08249_);
  or (_21836_, _21763_, _09043_);
  or (_21837_, _21836_, _21835_);
  and (_21838_, _21837_, _09048_);
  and (_21840_, _21838_, _21834_);
  nor (_21841_, _11209_, _11589_);
  or (_21842_, _21841_, _21763_);
  and (_21843_, _21842_, _06572_);
  or (_21844_, _21843_, _06606_);
  or (_21845_, _21844_, _21840_);
  or (_21846_, _21768_, _07037_);
  and (_21847_, _21846_, _06196_);
  and (_21848_, _21847_, _21845_);
  and (_21849_, _15713_, _08249_);
  or (_21851_, _21849_, _21763_);
  and (_21852_, _21851_, _06195_);
  or (_21853_, _21852_, _01379_);
  or (_21854_, _21853_, _21848_);
  or (_21855_, _01375_, \uc8051golden_1.DPH [6]);
  and (_21856_, _21855_, _42545_);
  and (_42935_, _21856_, _21854_);
  not (_21857_, \uc8051golden_1.TL1 [0]);
  nor (_21858_, _01375_, _21857_);
  nand (_21859_, _11225_, _07976_);
  nor (_21861_, _07976_, _21857_);
  nor (_21862_, _21861_, _07276_);
  nand (_21863_, _21862_, _21859_);
  and (_21864_, _07976_, _07473_);
  or (_21865_, _21864_, _21861_);
  or (_21866_, _21865_, _06293_);
  nor (_21867_, _08521_, _11679_);
  or (_21868_, _21867_, _21861_);
  or (_21869_, _21868_, _07210_);
  and (_21870_, _07976_, \uc8051golden_1.ACC [0]);
  or (_21872_, _21870_, _21861_);
  and (_21873_, _21872_, _07199_);
  nor (_21874_, _07199_, _21857_);
  or (_21875_, _21874_, _06401_);
  or (_21876_, _21875_, _21873_);
  and (_21877_, _21876_, _07221_);
  and (_21878_, _21877_, _21869_);
  and (_21879_, _21865_, _06399_);
  or (_21880_, _21879_, _21878_);
  and (_21881_, _21880_, _06414_);
  and (_21883_, _21872_, _06406_);
  or (_21884_, _21883_, _10059_);
  or (_21885_, _21884_, _21881_);
  and (_21886_, _21885_, _21866_);
  or (_21887_, _21886_, _06281_);
  and (_21888_, _07976_, _09446_);
  or (_21889_, _21861_, _06282_);
  or (_21890_, _21889_, _21888_);
  and (_21891_, _21890_, _21887_);
  or (_21892_, _21891_, _06015_);
  and (_21894_, _14426_, _07976_);
  or (_21895_, _21861_, _06279_);
  or (_21896_, _21895_, _21894_);
  and (_21897_, _21896_, _06276_);
  and (_21898_, _21897_, _21892_);
  and (_21899_, _07976_, _08817_);
  or (_21900_, _21899_, _21861_);
  and (_21901_, _21900_, _06275_);
  or (_21902_, _21901_, _06474_);
  or (_21903_, _21902_, _21898_);
  and (_21905_, _14324_, _07976_);
  or (_21906_, _21905_, _21861_);
  or (_21907_, _21906_, _07282_);
  and (_21908_, _21907_, _07284_);
  and (_21909_, _21908_, _21903_);
  nor (_21910_, _12538_, _11679_);
  or (_21911_, _21910_, _21861_);
  and (_21912_, _21859_, _06582_);
  and (_21913_, _21912_, _21911_);
  or (_21914_, _21913_, _21909_);
  and (_21916_, _21914_, _07279_);
  nand (_21917_, _21900_, _06478_);
  nor (_21918_, _21917_, _21867_);
  or (_21919_, _21918_, _06569_);
  or (_21920_, _21919_, _21916_);
  and (_21921_, _21920_, _21863_);
  or (_21922_, _21921_, _06479_);
  and (_21923_, _14320_, _07976_);
  or (_21924_, _21923_, _21861_);
  or (_21925_, _21924_, _09043_);
  and (_21927_, _21925_, _09048_);
  and (_21928_, _21927_, _21922_);
  and (_21929_, _21911_, _06572_);
  or (_21930_, _21929_, _19434_);
  or (_21931_, _21930_, _21928_);
  or (_21932_, _21868_, _06700_);
  and (_21933_, _21932_, _01375_);
  and (_21934_, _21933_, _21931_);
  or (_21935_, _21934_, _21858_);
  and (_42936_, _21935_, _42545_);
  and (_21937_, _11679_, \uc8051golden_1.TL1 [1]);
  nor (_21938_, _11223_, _11679_);
  or (_21939_, _21938_, _21937_);
  or (_21940_, _21939_, _09048_);
  and (_21941_, _07976_, _09445_);
  or (_21942_, _21937_, _06282_);
  or (_21943_, _21942_, _21941_);
  or (_21944_, _07976_, \uc8051golden_1.TL1 [1]);
  and (_21945_, _14532_, _07976_);
  not (_21946_, _21945_);
  and (_21948_, _21946_, _21944_);
  or (_21949_, _21948_, _07210_);
  and (_21950_, _07976_, \uc8051golden_1.ACC [1]);
  or (_21951_, _21950_, _21937_);
  and (_21952_, _21951_, _07199_);
  and (_21953_, _07200_, \uc8051golden_1.TL1 [1]);
  or (_21954_, _21953_, _06401_);
  or (_21955_, _21954_, _21952_);
  and (_21956_, _21955_, _07221_);
  and (_21957_, _21956_, _21949_);
  nor (_21959_, _11679_, _07196_);
  or (_21960_, _21959_, _21937_);
  and (_21961_, _21960_, _06399_);
  or (_21962_, _21961_, _21957_);
  and (_21963_, _21962_, _06414_);
  and (_21964_, _21951_, _06406_);
  or (_21965_, _21964_, _10059_);
  or (_21966_, _21965_, _21963_);
  or (_21967_, _21960_, _06293_);
  and (_21968_, _21967_, _21966_);
  or (_21970_, _21968_, _06281_);
  and (_21971_, _21970_, _06279_);
  and (_21972_, _21971_, _21943_);
  or (_21973_, _14615_, _11679_);
  and (_21974_, _21944_, _06015_);
  and (_21975_, _21974_, _21973_);
  or (_21976_, _21975_, _21972_);
  and (_21977_, _21976_, _06276_);
  nand (_21978_, _07976_, _07090_);
  and (_21979_, _21944_, _06275_);
  and (_21981_, _21979_, _21978_);
  or (_21982_, _21981_, _21977_);
  and (_21983_, _21982_, _07282_);
  or (_21984_, _14507_, _11679_);
  and (_21985_, _21944_, _06474_);
  and (_21986_, _21985_, _21984_);
  or (_21987_, _21986_, _06582_);
  or (_21988_, _21987_, _21983_);
  nand (_21989_, _11222_, _07976_);
  and (_21990_, _21989_, _21939_);
  or (_21992_, _21990_, _07284_);
  and (_21993_, _21992_, _07279_);
  and (_21994_, _21993_, _21988_);
  or (_21995_, _14505_, _11679_);
  and (_21996_, _21944_, _06478_);
  and (_21997_, _21996_, _21995_);
  or (_21998_, _21997_, _06569_);
  or (_21999_, _21998_, _21994_);
  nor (_22000_, _21937_, _07276_);
  nand (_22001_, _22000_, _21989_);
  and (_22003_, _22001_, _09043_);
  and (_22004_, _22003_, _21999_);
  or (_22005_, _21978_, _08477_);
  and (_22006_, _21944_, _06479_);
  and (_22007_, _22006_, _22005_);
  or (_22008_, _22007_, _06572_);
  or (_22009_, _22008_, _22004_);
  and (_22010_, _22009_, _21940_);
  or (_22011_, _22010_, _06606_);
  or (_22012_, _21948_, _07037_);
  and (_22014_, _22012_, _06196_);
  and (_22015_, _22014_, _22011_);
  or (_22016_, _21945_, _21937_);
  and (_22017_, _22016_, _06195_);
  or (_22018_, _22017_, _01379_);
  or (_22019_, _22018_, _22015_);
  or (_22020_, _01375_, \uc8051golden_1.TL1 [1]);
  and (_22021_, _22020_, _42545_);
  and (_42938_, _22021_, _22019_);
  and (_22022_, _01379_, \uc8051golden_1.TL1 [2]);
  and (_22024_, _07976_, _09444_);
  and (_22025_, _11679_, \uc8051golden_1.TL1 [2]);
  or (_22026_, _22025_, _06282_);
  or (_22027_, _22026_, _22024_);
  nor (_22028_, _11679_, _07623_);
  or (_22029_, _22028_, _22025_);
  or (_22030_, _22029_, _06293_);
  and (_22031_, _14754_, _07976_);
  or (_22032_, _22031_, _22025_);
  and (_22033_, _22032_, _06401_);
  and (_22035_, _07200_, \uc8051golden_1.TL1 [2]);
  and (_22036_, _07976_, \uc8051golden_1.ACC [2]);
  or (_22037_, _22036_, _22025_);
  and (_22038_, _22037_, _07199_);
  or (_22039_, _22038_, _22035_);
  and (_22040_, _22039_, _07210_);
  or (_22041_, _22040_, _06399_);
  or (_22042_, _22041_, _22033_);
  or (_22043_, _22029_, _07221_);
  and (_22044_, _22043_, _06414_);
  and (_22046_, _22044_, _22042_);
  and (_22047_, _22037_, _06406_);
  or (_22048_, _22047_, _10059_);
  or (_22049_, _22048_, _22046_);
  and (_22050_, _22049_, _22030_);
  or (_22051_, _22050_, _06281_);
  and (_22052_, _22051_, _22027_);
  or (_22053_, _22052_, _06015_);
  and (_22054_, _14848_, _07976_);
  or (_22055_, _22025_, _06279_);
  or (_22057_, _22055_, _22054_);
  and (_22058_, _22057_, _06276_);
  and (_22059_, _22058_, _22053_);
  and (_22060_, _07976_, _08994_);
  or (_22061_, _22060_, _22025_);
  and (_22062_, _22061_, _06275_);
  or (_22063_, _22062_, _06474_);
  or (_22064_, _22063_, _22059_);
  and (_22065_, _14744_, _07976_);
  or (_22066_, _22065_, _22025_);
  or (_22068_, _22066_, _07282_);
  and (_22069_, _22068_, _07284_);
  and (_22070_, _22069_, _22064_);
  and (_22071_, _11221_, _07976_);
  or (_22072_, _22071_, _22025_);
  and (_22073_, _22072_, _06582_);
  or (_22074_, _22073_, _22070_);
  and (_22075_, _22074_, _07279_);
  or (_22076_, _22025_, _08433_);
  and (_22077_, _22061_, _06478_);
  and (_22079_, _22077_, _22076_);
  or (_22080_, _22079_, _22075_);
  and (_22081_, _22080_, _07276_);
  and (_22082_, _22037_, _06569_);
  and (_22083_, _22082_, _22076_);
  or (_22084_, _22083_, _06479_);
  or (_22085_, _22084_, _22081_);
  and (_22086_, _14741_, _07976_);
  or (_22087_, _22025_, _09043_);
  or (_22088_, _22087_, _22086_);
  and (_22090_, _22088_, _09048_);
  and (_22091_, _22090_, _22085_);
  nor (_22092_, _11220_, _11679_);
  or (_22093_, _22092_, _22025_);
  and (_22094_, _22093_, _06572_);
  or (_22095_, _22094_, _22091_);
  and (_22096_, _22095_, _07037_);
  and (_22097_, _22032_, _06606_);
  or (_22098_, _22097_, _06195_);
  or (_22099_, _22098_, _22096_);
  and (_22101_, _14917_, _07976_);
  or (_22102_, _22025_, _06196_);
  or (_22103_, _22102_, _22101_);
  and (_22104_, _22103_, _01375_);
  and (_22105_, _22104_, _22099_);
  or (_22106_, _22105_, _22022_);
  and (_42939_, _22106_, _42545_);
  and (_22107_, _11679_, \uc8051golden_1.TL1 [3]);
  and (_22108_, _07976_, _09443_);
  or (_22109_, _22108_, _22107_);
  and (_22111_, _22109_, _06281_);
  and (_22112_, _14947_, _07976_);
  or (_22113_, _22112_, _22107_);
  or (_22114_, _22113_, _07210_);
  and (_22115_, _07976_, \uc8051golden_1.ACC [3]);
  or (_22116_, _22115_, _22107_);
  and (_22117_, _22116_, _07199_);
  and (_22118_, _07200_, \uc8051golden_1.TL1 [3]);
  or (_22119_, _22118_, _06401_);
  or (_22120_, _22119_, _22117_);
  and (_22123_, _22120_, _07221_);
  and (_22124_, _22123_, _22114_);
  nor (_22125_, _11679_, _07775_);
  or (_22126_, _22125_, _22107_);
  and (_22127_, _22126_, _06399_);
  or (_22128_, _22127_, _22124_);
  and (_22129_, _22128_, _06414_);
  and (_22130_, _22116_, _06406_);
  or (_22131_, _22130_, _10059_);
  or (_22132_, _22131_, _22129_);
  or (_22134_, _22126_, _06293_);
  and (_22135_, _22134_, _06282_);
  and (_22136_, _22135_, _22132_);
  or (_22137_, _22136_, _06015_);
  or (_22138_, _22137_, _22111_);
  and (_22139_, _15039_, _07976_);
  or (_22140_, _22107_, _06279_);
  or (_22141_, _22140_, _22139_);
  and (_22142_, _22141_, _06276_);
  and (_22143_, _22142_, _22138_);
  and (_22145_, _07976_, _08815_);
  or (_22146_, _22145_, _22107_);
  and (_22147_, _22146_, _06275_);
  or (_22148_, _22147_, _06474_);
  or (_22149_, _22148_, _22143_);
  and (_22150_, _14934_, _07976_);
  or (_22151_, _22150_, _22107_);
  or (_22152_, _22151_, _07282_);
  and (_22153_, _22152_, _07284_);
  and (_22154_, _22153_, _22149_);
  and (_22156_, _12535_, _07976_);
  or (_22157_, _22156_, _22107_);
  and (_22158_, _22157_, _06582_);
  or (_22159_, _22158_, _22154_);
  and (_22160_, _22159_, _07279_);
  or (_22161_, _22107_, _08389_);
  and (_22162_, _22146_, _06478_);
  and (_22163_, _22162_, _22161_);
  or (_22164_, _22163_, _22160_);
  and (_22165_, _22164_, _07276_);
  and (_22167_, _22116_, _06569_);
  and (_22168_, _22167_, _22161_);
  or (_22169_, _22168_, _06479_);
  or (_22170_, _22169_, _22165_);
  and (_22171_, _14931_, _07976_);
  or (_22172_, _22107_, _09043_);
  or (_22173_, _22172_, _22171_);
  and (_22174_, _22173_, _09048_);
  and (_22175_, _22174_, _22170_);
  nor (_22176_, _11218_, _11679_);
  or (_22178_, _22176_, _22107_);
  and (_22179_, _22178_, _06572_);
  or (_22180_, _22179_, _06606_);
  or (_22181_, _22180_, _22175_);
  or (_22182_, _22113_, _07037_);
  and (_22183_, _22182_, _06196_);
  and (_22184_, _22183_, _22181_);
  and (_22185_, _15113_, _07976_);
  or (_22186_, _22185_, _22107_);
  and (_22187_, _22186_, _06195_);
  or (_22189_, _22187_, _01379_);
  or (_22190_, _22189_, _22184_);
  or (_22191_, _01375_, \uc8051golden_1.TL1 [3]);
  and (_22192_, _22191_, _42545_);
  and (_42940_, _22192_, _22190_);
  and (_22193_, _11679_, \uc8051golden_1.TL1 [4]);
  and (_22194_, _15130_, _07976_);
  or (_22195_, _22194_, _22193_);
  or (_22196_, _22195_, _07210_);
  and (_22197_, _07976_, \uc8051golden_1.ACC [4]);
  or (_22199_, _22197_, _22193_);
  and (_22200_, _22199_, _07199_);
  and (_22201_, _07200_, \uc8051golden_1.TL1 [4]);
  or (_22202_, _22201_, _06401_);
  or (_22203_, _22202_, _22200_);
  and (_22204_, _22203_, _07221_);
  and (_22205_, _22204_, _22196_);
  nor (_22206_, _11679_, _08301_);
  or (_22207_, _22206_, _22193_);
  and (_22208_, _22207_, _06399_);
  or (_22209_, _22208_, _22205_);
  and (_22210_, _22209_, _06414_);
  and (_22211_, _22199_, _06406_);
  or (_22212_, _22211_, _10059_);
  or (_22213_, _22212_, _22210_);
  or (_22214_, _22207_, _06293_);
  and (_22215_, _22214_, _22213_);
  or (_22216_, _22215_, _06281_);
  and (_22217_, _07976_, _09442_);
  or (_22218_, _22193_, _06282_);
  or (_22221_, _22218_, _22217_);
  and (_22222_, _22221_, _06279_);
  and (_22223_, _22222_, _22216_);
  and (_22224_, _15243_, _07976_);
  or (_22225_, _22224_, _22193_);
  and (_22226_, _22225_, _06015_);
  or (_22227_, _22226_, _06275_);
  or (_22228_, _22227_, _22223_);
  and (_22229_, _08883_, _07976_);
  or (_22230_, _22229_, _22193_);
  or (_22232_, _22230_, _06276_);
  and (_22233_, _22232_, _22228_);
  or (_22234_, _22233_, _06474_);
  and (_22235_, _15135_, _07976_);
  or (_22236_, _22235_, _22193_);
  or (_22237_, _22236_, _07282_);
  and (_22238_, _22237_, _07284_);
  and (_22239_, _22238_, _22234_);
  and (_22240_, _11216_, _07976_);
  or (_22241_, _22240_, _22193_);
  and (_22243_, _22241_, _06582_);
  or (_22244_, _22243_, _22239_);
  and (_22245_, _22244_, _07279_);
  or (_22246_, _22193_, _08345_);
  and (_22247_, _22230_, _06478_);
  and (_22248_, _22247_, _22246_);
  or (_22249_, _22248_, _22245_);
  and (_22250_, _22249_, _07276_);
  and (_22251_, _22199_, _06569_);
  and (_22252_, _22251_, _22246_);
  or (_22254_, _22252_, _06479_);
  or (_22255_, _22254_, _22250_);
  and (_22256_, _15134_, _07976_);
  or (_22257_, _22193_, _09043_);
  or (_22258_, _22257_, _22256_);
  and (_22259_, _22258_, _09048_);
  and (_22260_, _22259_, _22255_);
  nor (_22261_, _11215_, _11679_);
  or (_22262_, _22261_, _22193_);
  and (_22263_, _22262_, _06572_);
  or (_22265_, _22263_, _06606_);
  or (_22266_, _22265_, _22260_);
  or (_22267_, _22195_, _07037_);
  and (_22268_, _22267_, _06196_);
  and (_22269_, _22268_, _22266_);
  and (_22270_, _15315_, _07976_);
  or (_22271_, _22270_, _22193_);
  and (_22272_, _22271_, _06195_);
  or (_22273_, _22272_, _01379_);
  or (_22274_, _22273_, _22269_);
  or (_22276_, _01375_, \uc8051golden_1.TL1 [4]);
  and (_22277_, _22276_, _42545_);
  and (_42941_, _22277_, _22274_);
  and (_22278_, _11679_, \uc8051golden_1.TL1 [5]);
  nor (_22279_, _11679_, _08207_);
  or (_22280_, _22279_, _22278_);
  or (_22281_, _22280_, _06293_);
  and (_22282_, _15348_, _07976_);
  or (_22283_, _22282_, _22278_);
  or (_22284_, _22283_, _07210_);
  and (_22286_, _07976_, \uc8051golden_1.ACC [5]);
  or (_22287_, _22286_, _22278_);
  and (_22288_, _22287_, _07199_);
  and (_22289_, _07200_, \uc8051golden_1.TL1 [5]);
  or (_22290_, _22289_, _06401_);
  or (_22291_, _22290_, _22288_);
  and (_22292_, _22291_, _07221_);
  and (_22293_, _22292_, _22284_);
  and (_22294_, _22280_, _06399_);
  or (_22295_, _22294_, _22293_);
  and (_22297_, _22295_, _06414_);
  and (_22298_, _22287_, _06406_);
  or (_22299_, _22298_, _10059_);
  or (_22300_, _22299_, _22297_);
  and (_22301_, _22300_, _22281_);
  or (_22302_, _22301_, _06281_);
  and (_22303_, _07976_, _09441_);
  or (_22304_, _22278_, _06282_);
  or (_22305_, _22304_, _22303_);
  and (_22306_, _22305_, _06279_);
  and (_22308_, _22306_, _22302_);
  and (_22309_, _15446_, _07976_);
  or (_22310_, _22309_, _22278_);
  and (_22311_, _22310_, _06015_);
  or (_22312_, _22311_, _06275_);
  or (_22313_, _22312_, _22308_);
  and (_22314_, _08958_, _07976_);
  or (_22315_, _22314_, _22278_);
  or (_22316_, _22315_, _06276_);
  and (_22317_, _22316_, _22313_);
  or (_22319_, _22317_, _06474_);
  and (_22320_, _15338_, _07976_);
  or (_22321_, _22320_, _22278_);
  or (_22322_, _22321_, _07282_);
  and (_22323_, _22322_, _07284_);
  and (_22324_, _22323_, _22319_);
  and (_22325_, _12542_, _07976_);
  or (_22326_, _22325_, _22278_);
  and (_22327_, _22326_, _06582_);
  or (_22328_, _22327_, _22324_);
  and (_22330_, _22328_, _07279_);
  or (_22331_, _22278_, _08256_);
  and (_22332_, _22315_, _06478_);
  and (_22333_, _22332_, _22331_);
  or (_22334_, _22333_, _22330_);
  and (_22335_, _22334_, _07276_);
  and (_22336_, _22287_, _06569_);
  and (_22337_, _22336_, _22331_);
  or (_22338_, _22337_, _06479_);
  or (_22339_, _22338_, _22335_);
  and (_22341_, _15335_, _07976_);
  or (_22342_, _22278_, _09043_);
  or (_22343_, _22342_, _22341_);
  and (_22344_, _22343_, _09048_);
  and (_22345_, _22344_, _22339_);
  nor (_22346_, _11212_, _11679_);
  or (_22347_, _22346_, _22278_);
  and (_22348_, _22347_, _06572_);
  or (_22349_, _22348_, _06606_);
  or (_22350_, _22349_, _22345_);
  or (_22352_, _22283_, _07037_);
  and (_22353_, _22352_, _06196_);
  and (_22354_, _22353_, _22350_);
  and (_22355_, _15509_, _07976_);
  or (_22356_, _22355_, _22278_);
  and (_22357_, _22356_, _06195_);
  or (_22358_, _22357_, _01379_);
  or (_22359_, _22358_, _22354_);
  or (_22360_, _01375_, \uc8051golden_1.TL1 [5]);
  and (_22361_, _22360_, _42545_);
  and (_42942_, _22361_, _22359_);
  and (_22363_, _11679_, \uc8051golden_1.TL1 [6]);
  nor (_22364_, _11679_, _08118_);
  or (_22365_, _22364_, _22363_);
  or (_22366_, _22365_, _06293_);
  and (_22367_, _15550_, _07976_);
  or (_22368_, _22367_, _22363_);
  or (_22369_, _22368_, _07210_);
  and (_22370_, _07976_, \uc8051golden_1.ACC [6]);
  or (_22371_, _22370_, _22363_);
  and (_22373_, _22371_, _07199_);
  and (_22374_, _07200_, \uc8051golden_1.TL1 [6]);
  or (_22375_, _22374_, _06401_);
  or (_22376_, _22375_, _22373_);
  and (_22377_, _22376_, _07221_);
  and (_22378_, _22377_, _22369_);
  and (_22379_, _22365_, _06399_);
  or (_22380_, _22379_, _22378_);
  and (_22381_, _22380_, _06414_);
  and (_22382_, _22371_, _06406_);
  or (_22384_, _22382_, _10059_);
  or (_22385_, _22384_, _22381_);
  and (_22386_, _22385_, _22366_);
  or (_22387_, _22386_, _06281_);
  and (_22388_, _07976_, _09440_);
  or (_22389_, _22363_, _06282_);
  or (_22390_, _22389_, _22388_);
  and (_22391_, _22390_, _06279_);
  and (_22392_, _22391_, _22387_);
  and (_22393_, _15639_, _07976_);
  or (_22395_, _22393_, _22363_);
  and (_22396_, _22395_, _06015_);
  or (_22397_, _22396_, _06275_);
  or (_22398_, _22397_, _22392_);
  and (_22399_, _15646_, _07976_);
  or (_22400_, _22399_, _22363_);
  or (_22401_, _22400_, _06276_);
  and (_22402_, _22401_, _22398_);
  or (_22403_, _22402_, _06474_);
  and (_22404_, _15531_, _07976_);
  or (_22406_, _22404_, _22363_);
  or (_22407_, _22406_, _07282_);
  and (_22408_, _22407_, _07284_);
  and (_22409_, _22408_, _22403_);
  and (_22410_, _11210_, _07976_);
  or (_22411_, _22410_, _22363_);
  and (_22412_, _22411_, _06582_);
  or (_22413_, _22412_, _22409_);
  and (_22414_, _22413_, _07279_);
  or (_22415_, _22363_, _08162_);
  and (_22417_, _22400_, _06478_);
  and (_22418_, _22417_, _22415_);
  or (_22419_, _22418_, _22414_);
  and (_22420_, _22419_, _07276_);
  and (_22421_, _22371_, _06569_);
  and (_22422_, _22421_, _22415_);
  or (_22423_, _22422_, _06479_);
  or (_22424_, _22423_, _22420_);
  and (_22425_, _15528_, _07976_);
  or (_22426_, _22363_, _09043_);
  or (_22428_, _22426_, _22425_);
  and (_22429_, _22428_, _09048_);
  and (_22430_, _22429_, _22424_);
  nor (_22431_, _11209_, _11679_);
  or (_22432_, _22431_, _22363_);
  and (_22433_, _22432_, _06572_);
  or (_22434_, _22433_, _06606_);
  or (_22435_, _22434_, _22430_);
  or (_22436_, _22368_, _07037_);
  and (_22437_, _22436_, _06196_);
  and (_22439_, _22437_, _22435_);
  and (_22440_, _15713_, _07976_);
  or (_22441_, _22440_, _22363_);
  and (_22442_, _22441_, _06195_);
  or (_22443_, _22442_, _01379_);
  or (_22444_, _22443_, _22439_);
  or (_22445_, _01375_, \uc8051golden_1.TL1 [6]);
  and (_22446_, _22445_, _42545_);
  and (_42943_, _22446_, _22444_);
  not (_22447_, \uc8051golden_1.TL0 [0]);
  nor (_22449_, _01375_, _22447_);
  nand (_22450_, _11225_, _08010_);
  nor (_22451_, _08010_, _22447_);
  nor (_22452_, _22451_, _07276_);
  nand (_22453_, _22452_, _22450_);
  nor (_22454_, _08521_, _11757_);
  or (_22455_, _22454_, _22451_);
  or (_22456_, _22455_, _07210_);
  and (_22457_, _08010_, \uc8051golden_1.ACC [0]);
  or (_22458_, _22457_, _22451_);
  and (_22460_, _22458_, _07199_);
  nor (_22461_, _07199_, _22447_);
  or (_22462_, _22461_, _06401_);
  or (_22463_, _22462_, _22460_);
  and (_22464_, _22463_, _07221_);
  and (_22465_, _22464_, _22456_);
  and (_22466_, _08010_, _07473_);
  or (_22467_, _22466_, _22451_);
  and (_22468_, _22467_, _06399_);
  or (_22469_, _22468_, _22465_);
  and (_22471_, _22469_, _06414_);
  and (_22472_, _22458_, _06406_);
  or (_22473_, _22472_, _10059_);
  or (_22474_, _22473_, _22471_);
  or (_22475_, _22467_, _06293_);
  and (_22476_, _22475_, _22474_);
  or (_22477_, _22476_, _06281_);
  and (_22478_, _08010_, _09446_);
  or (_22479_, _22451_, _06282_);
  or (_22480_, _22479_, _22478_);
  and (_22482_, _22480_, _22477_);
  or (_22483_, _22482_, _06015_);
  and (_22484_, _14426_, _08010_);
  or (_22485_, _22451_, _06279_);
  or (_22486_, _22485_, _22484_);
  and (_22487_, _22486_, _06276_);
  and (_22488_, _22487_, _22483_);
  and (_22489_, _08010_, _08817_);
  or (_22490_, _22489_, _22451_);
  and (_22491_, _22490_, _06275_);
  or (_22493_, _22491_, _06474_);
  or (_22494_, _22493_, _22488_);
  and (_22495_, _14324_, _08010_);
  or (_22496_, _22495_, _22451_);
  or (_22497_, _22496_, _07282_);
  and (_22498_, _22497_, _07284_);
  and (_22499_, _22498_, _22494_);
  nor (_22500_, _12538_, _11757_);
  or (_22501_, _22500_, _22451_);
  and (_22502_, _22450_, _06582_);
  and (_22503_, _22502_, _22501_);
  or (_22504_, _22503_, _22499_);
  and (_22505_, _22504_, _07279_);
  nand (_22506_, _22490_, _06478_);
  nor (_22507_, _22506_, _22454_);
  or (_22508_, _22507_, _06569_);
  or (_22509_, _22508_, _22505_);
  and (_22510_, _22509_, _22453_);
  or (_22511_, _22510_, _06479_);
  and (_22512_, _14320_, _08010_);
  or (_22515_, _22451_, _09043_);
  or (_22516_, _22515_, _22512_);
  and (_22517_, _22516_, _09048_);
  and (_22518_, _22517_, _22511_);
  and (_22519_, _22501_, _06572_);
  or (_22520_, _22519_, _19434_);
  or (_22521_, _22520_, _22518_);
  or (_22522_, _22455_, _06700_);
  and (_22523_, _22522_, _01375_);
  and (_22524_, _22523_, _22521_);
  or (_22526_, _22524_, _22449_);
  and (_42944_, _22526_, _42545_);
  and (_22527_, _11757_, \uc8051golden_1.TL0 [1]);
  nor (_22528_, _11223_, _11757_);
  or (_22529_, _22528_, _22527_);
  or (_22530_, _22529_, _09048_);
  and (_22531_, _08010_, _09445_);
  or (_22532_, _22527_, _06282_);
  or (_22533_, _22532_, _22531_);
  or (_22534_, _08010_, \uc8051golden_1.TL0 [1]);
  and (_22536_, _14532_, _08010_);
  not (_22537_, _22536_);
  and (_22538_, _22537_, _22534_);
  or (_22539_, _22538_, _07210_);
  and (_22540_, _08010_, \uc8051golden_1.ACC [1]);
  or (_22541_, _22540_, _22527_);
  and (_22542_, _22541_, _07199_);
  and (_22543_, _07200_, \uc8051golden_1.TL0 [1]);
  or (_22544_, _22543_, _06401_);
  or (_22545_, _22544_, _22542_);
  and (_22547_, _22545_, _07221_);
  and (_22548_, _22547_, _22539_);
  nor (_22549_, _11757_, _07196_);
  or (_22550_, _22549_, _22527_);
  and (_22551_, _22550_, _06399_);
  or (_22552_, _22551_, _22548_);
  and (_22553_, _22552_, _06414_);
  and (_22554_, _22541_, _06406_);
  or (_22555_, _22554_, _10059_);
  or (_22556_, _22555_, _22553_);
  or (_22558_, _22550_, _06293_);
  and (_22559_, _22558_, _22556_);
  or (_22560_, _22559_, _06281_);
  and (_22561_, _22560_, _06279_);
  and (_22562_, _22561_, _22533_);
  or (_22563_, _14615_, _11757_);
  and (_22564_, _22534_, _06015_);
  and (_22565_, _22564_, _22563_);
  or (_22566_, _22565_, _22562_);
  and (_22567_, _22566_, _06276_);
  nand (_22569_, _08010_, _07090_);
  and (_22570_, _22534_, _06275_);
  and (_22571_, _22570_, _22569_);
  or (_22572_, _22571_, _22567_);
  and (_22573_, _22572_, _07282_);
  or (_22574_, _14507_, _11757_);
  and (_22575_, _22534_, _06474_);
  and (_22576_, _22575_, _22574_);
  or (_22577_, _22576_, _06582_);
  or (_22578_, _22577_, _22573_);
  nand (_22580_, _11222_, _08010_);
  and (_22581_, _22580_, _22529_);
  or (_22582_, _22581_, _07284_);
  and (_22583_, _22582_, _07279_);
  and (_22584_, _22583_, _22578_);
  or (_22585_, _14505_, _11757_);
  and (_22586_, _22534_, _06478_);
  and (_22587_, _22586_, _22585_);
  or (_22588_, _22587_, _06569_);
  or (_22589_, _22588_, _22584_);
  nor (_22591_, _22527_, _07276_);
  nand (_22592_, _22591_, _22580_);
  and (_22593_, _22592_, _09043_);
  and (_22594_, _22593_, _22589_);
  or (_22595_, _22569_, _08477_);
  and (_22596_, _22534_, _06479_);
  and (_22597_, _22596_, _22595_);
  or (_22598_, _22597_, _06572_);
  or (_22599_, _22598_, _22594_);
  and (_22600_, _22599_, _22530_);
  or (_22602_, _22600_, _06606_);
  or (_22603_, _22538_, _07037_);
  and (_22604_, _22603_, _06196_);
  and (_22605_, _22604_, _22602_);
  or (_22606_, _22536_, _22527_);
  and (_22607_, _22606_, _06195_);
  or (_22608_, _22607_, _01379_);
  or (_22609_, _22608_, _22605_);
  or (_22610_, _01375_, \uc8051golden_1.TL0 [1]);
  and (_22611_, _22610_, _42545_);
  and (_42945_, _22611_, _22609_);
  and (_22612_, _01379_, \uc8051golden_1.TL0 [2]);
  and (_22613_, _08010_, _09444_);
  and (_22614_, _11757_, \uc8051golden_1.TL0 [2]);
  or (_22615_, _22614_, _06282_);
  or (_22616_, _22615_, _22613_);
  nor (_22617_, _11757_, _07623_);
  or (_22618_, _22617_, _22614_);
  or (_22619_, _22618_, _06293_);
  and (_22620_, _14754_, _08010_);
  or (_22623_, _22620_, _22614_);
  and (_22624_, _22623_, _06401_);
  and (_22625_, _07200_, \uc8051golden_1.TL0 [2]);
  and (_22626_, _08010_, \uc8051golden_1.ACC [2]);
  or (_22627_, _22626_, _22614_);
  and (_22628_, _22627_, _07199_);
  or (_22629_, _22628_, _22625_);
  and (_22630_, _22629_, _07210_);
  or (_22631_, _22630_, _06399_);
  or (_22632_, _22631_, _22624_);
  or (_22634_, _22618_, _07221_);
  and (_22635_, _22634_, _06414_);
  and (_22636_, _22635_, _22632_);
  and (_22637_, _22627_, _06406_);
  or (_22638_, _22637_, _10059_);
  or (_22639_, _22638_, _22636_);
  and (_22640_, _22639_, _22619_);
  or (_22641_, _22640_, _06281_);
  and (_22642_, _22641_, _22616_);
  or (_22643_, _22642_, _06015_);
  and (_22645_, _14848_, _08010_);
  or (_22646_, _22614_, _06279_);
  or (_22647_, _22646_, _22645_);
  and (_22648_, _22647_, _06276_);
  and (_22649_, _22648_, _22643_);
  and (_22650_, _08010_, _08994_);
  or (_22651_, _22650_, _22614_);
  and (_22652_, _22651_, _06275_);
  or (_22653_, _22652_, _06474_);
  or (_22654_, _22653_, _22649_);
  and (_22656_, _14744_, _08010_);
  or (_22657_, _22656_, _22614_);
  or (_22658_, _22657_, _07282_);
  and (_22659_, _22658_, _07284_);
  and (_22660_, _22659_, _22654_);
  and (_22661_, _11221_, _08010_);
  or (_22662_, _22661_, _22614_);
  and (_22663_, _22662_, _06582_);
  or (_22664_, _22663_, _22660_);
  and (_22665_, _22664_, _07279_);
  or (_22667_, _22614_, _08433_);
  and (_22668_, _22651_, _06478_);
  and (_22669_, _22668_, _22667_);
  or (_22670_, _22669_, _22665_);
  and (_22671_, _22670_, _07276_);
  and (_22672_, _22627_, _06569_);
  and (_22673_, _22672_, _22667_);
  or (_22674_, _22673_, _06479_);
  or (_22675_, _22674_, _22671_);
  and (_22676_, _14741_, _08010_);
  or (_22678_, _22614_, _09043_);
  or (_22679_, _22678_, _22676_);
  and (_22680_, _22679_, _09048_);
  and (_22681_, _22680_, _22675_);
  nor (_22682_, _11220_, _11757_);
  or (_22683_, _22682_, _22614_);
  and (_22684_, _22683_, _06572_);
  or (_22685_, _22684_, _22681_);
  and (_22686_, _22685_, _07037_);
  and (_22687_, _22623_, _06606_);
  or (_22689_, _22687_, _06195_);
  or (_22690_, _22689_, _22686_);
  and (_22691_, _14917_, _08010_);
  or (_22692_, _22614_, _06196_);
  or (_22693_, _22692_, _22691_);
  and (_22694_, _22693_, _01375_);
  and (_22695_, _22694_, _22690_);
  or (_22696_, _22695_, _22612_);
  and (_42946_, _22696_, _42545_);
  and (_22697_, _11757_, \uc8051golden_1.TL0 [3]);
  and (_22699_, _14947_, _08010_);
  or (_22700_, _22699_, _22697_);
  or (_22701_, _22700_, _07210_);
  and (_22702_, _08010_, \uc8051golden_1.ACC [3]);
  or (_22703_, _22702_, _22697_);
  and (_22704_, _22703_, _07199_);
  and (_22705_, _07200_, \uc8051golden_1.TL0 [3]);
  or (_22706_, _22705_, _06401_);
  or (_22707_, _22706_, _22704_);
  and (_22708_, _22707_, _07221_);
  and (_22710_, _22708_, _22701_);
  nor (_22711_, _11757_, _07775_);
  or (_22712_, _22711_, _22697_);
  and (_22713_, _22712_, _06399_);
  or (_22714_, _22713_, _22710_);
  and (_22715_, _22714_, _06414_);
  and (_22716_, _22703_, _06406_);
  or (_22717_, _22716_, _10059_);
  or (_22718_, _22717_, _22715_);
  or (_22719_, _22712_, _06293_);
  and (_22721_, _22719_, _22718_);
  or (_22722_, _22721_, _06281_);
  and (_22723_, _08010_, _09443_);
  or (_22724_, _22697_, _06282_);
  or (_22725_, _22724_, _22723_);
  and (_22726_, _22725_, _22722_);
  or (_22727_, _22726_, _06015_);
  and (_22728_, _15039_, _08010_);
  or (_22729_, _22697_, _06279_);
  or (_22730_, _22729_, _22728_);
  and (_22732_, _22730_, _06276_);
  and (_22733_, _22732_, _22727_);
  and (_22734_, _08010_, _08815_);
  or (_22735_, _22734_, _22697_);
  and (_22736_, _22735_, _06275_);
  or (_22737_, _22736_, _06474_);
  or (_22738_, _22737_, _22733_);
  and (_22739_, _14934_, _08010_);
  or (_22740_, _22739_, _22697_);
  or (_22741_, _22740_, _07282_);
  and (_22743_, _22741_, _07284_);
  and (_22744_, _22743_, _22738_);
  and (_22745_, _12535_, _08010_);
  or (_22746_, _22745_, _22697_);
  and (_22747_, _22746_, _06582_);
  or (_22748_, _22747_, _22744_);
  and (_22749_, _22748_, _07279_);
  or (_22750_, _22697_, _08389_);
  and (_22751_, _22735_, _06478_);
  and (_22752_, _22751_, _22750_);
  or (_22754_, _22752_, _22749_);
  and (_22755_, _22754_, _07276_);
  and (_22756_, _22703_, _06569_);
  and (_22757_, _22756_, _22750_);
  or (_22758_, _22757_, _06479_);
  or (_22759_, _22758_, _22755_);
  and (_22760_, _14931_, _08010_);
  or (_22761_, _22697_, _09043_);
  or (_22762_, _22761_, _22760_);
  and (_22763_, _22762_, _09048_);
  and (_22765_, _22763_, _22759_);
  nor (_22766_, _11218_, _11757_);
  or (_22767_, _22766_, _22697_);
  and (_22768_, _22767_, _06572_);
  or (_22769_, _22768_, _06606_);
  or (_22770_, _22769_, _22765_);
  or (_22771_, _22700_, _07037_);
  and (_22772_, _22771_, _06196_);
  and (_22773_, _22772_, _22770_);
  and (_22774_, _15113_, _08010_);
  or (_22776_, _22774_, _22697_);
  and (_22777_, _22776_, _06195_);
  or (_22778_, _22777_, _01379_);
  or (_22779_, _22778_, _22773_);
  or (_22780_, _01375_, \uc8051golden_1.TL0 [3]);
  and (_22781_, _22780_, _42545_);
  and (_42947_, _22781_, _22779_);
  and (_22782_, _11757_, \uc8051golden_1.TL0 [4]);
  and (_22783_, _15130_, _08010_);
  or (_22784_, _22783_, _22782_);
  or (_22786_, _22784_, _07210_);
  and (_22787_, _08010_, \uc8051golden_1.ACC [4]);
  or (_22788_, _22787_, _22782_);
  and (_22789_, _22788_, _07199_);
  and (_22790_, _07200_, \uc8051golden_1.TL0 [4]);
  or (_22791_, _22790_, _06401_);
  or (_22792_, _22791_, _22789_);
  and (_22793_, _22792_, _07221_);
  and (_22794_, _22793_, _22786_);
  nor (_22795_, _11757_, _08301_);
  or (_22797_, _22795_, _22782_);
  and (_22798_, _22797_, _06399_);
  or (_22799_, _22798_, _22794_);
  and (_22800_, _22799_, _06414_);
  and (_22801_, _22788_, _06406_);
  or (_22802_, _22801_, _10059_);
  or (_22803_, _22802_, _22800_);
  or (_22804_, _22797_, _06293_);
  and (_22805_, _22804_, _22803_);
  or (_22806_, _22805_, _06281_);
  and (_22808_, _08010_, _09442_);
  or (_22809_, _22782_, _06282_);
  or (_22810_, _22809_, _22808_);
  and (_22811_, _22810_, _06279_);
  and (_22812_, _22811_, _22806_);
  and (_22813_, _15243_, _08010_);
  or (_22814_, _22813_, _22782_);
  and (_22815_, _22814_, _06015_);
  or (_22816_, _22815_, _06275_);
  or (_22817_, _22816_, _22812_);
  and (_22819_, _08883_, _08010_);
  or (_22820_, _22819_, _22782_);
  or (_22821_, _22820_, _06276_);
  and (_22822_, _22821_, _22817_);
  or (_22823_, _22822_, _06474_);
  and (_22824_, _15135_, _08010_);
  or (_22825_, _22824_, _22782_);
  or (_22826_, _22825_, _07282_);
  and (_22827_, _22826_, _07284_);
  and (_22828_, _22827_, _22823_);
  and (_22829_, _11216_, _08010_);
  or (_22830_, _22829_, _22782_);
  and (_22831_, _22830_, _06582_);
  or (_22832_, _22831_, _22828_);
  and (_22833_, _22832_, _07279_);
  or (_22834_, _22782_, _08345_);
  and (_22835_, _22820_, _06478_);
  and (_22836_, _22835_, _22834_);
  or (_22837_, _22836_, _22833_);
  and (_22838_, _22837_, _07276_);
  and (_22841_, _22788_, _06569_);
  and (_22842_, _22841_, _22834_);
  or (_22843_, _22842_, _06479_);
  or (_22844_, _22843_, _22838_);
  and (_22845_, _15134_, _08010_);
  or (_22846_, _22782_, _09043_);
  or (_22847_, _22846_, _22845_);
  and (_22848_, _22847_, _09048_);
  and (_22849_, _22848_, _22844_);
  nor (_22850_, _11215_, _11757_);
  or (_22852_, _22850_, _22782_);
  and (_22853_, _22852_, _06572_);
  or (_22854_, _22853_, _06606_);
  or (_22855_, _22854_, _22849_);
  or (_22856_, _22784_, _07037_);
  and (_22857_, _22856_, _06196_);
  and (_22858_, _22857_, _22855_);
  and (_22859_, _15315_, _08010_);
  or (_22860_, _22859_, _22782_);
  and (_22861_, _22860_, _06195_);
  or (_22863_, _22861_, _01379_);
  or (_22864_, _22863_, _22858_);
  or (_22865_, _01375_, \uc8051golden_1.TL0 [4]);
  and (_22866_, _22865_, _42545_);
  and (_42948_, _22866_, _22864_);
  and (_22867_, _11757_, \uc8051golden_1.TL0 [5]);
  nor (_22868_, _11757_, _08207_);
  or (_22869_, _22868_, _22867_);
  or (_22870_, _22869_, _06293_);
  and (_22871_, _15348_, _08010_);
  or (_22873_, _22871_, _22867_);
  or (_22874_, _22873_, _07210_);
  and (_22875_, _08010_, \uc8051golden_1.ACC [5]);
  or (_22876_, _22875_, _22867_);
  and (_22877_, _22876_, _07199_);
  and (_22878_, _07200_, \uc8051golden_1.TL0 [5]);
  or (_22879_, _22878_, _06401_);
  or (_22880_, _22879_, _22877_);
  and (_22881_, _22880_, _07221_);
  and (_22882_, _22881_, _22874_);
  and (_22884_, _22869_, _06399_);
  or (_22885_, _22884_, _22882_);
  and (_22886_, _22885_, _06414_);
  and (_22887_, _22876_, _06406_);
  or (_22888_, _22887_, _10059_);
  or (_22889_, _22888_, _22886_);
  and (_22890_, _22889_, _22870_);
  or (_22891_, _22890_, _06281_);
  and (_22892_, _08010_, _09441_);
  or (_22893_, _22867_, _06282_);
  or (_22895_, _22893_, _22892_);
  and (_22896_, _22895_, _06279_);
  and (_22897_, _22896_, _22891_);
  and (_22898_, _15446_, _08010_);
  or (_22899_, _22898_, _22867_);
  and (_22900_, _22899_, _06015_);
  or (_22901_, _22900_, _06275_);
  or (_22902_, _22901_, _22897_);
  and (_22903_, _08958_, _08010_);
  or (_22904_, _22903_, _22867_);
  or (_22906_, _22904_, _06276_);
  and (_22907_, _22906_, _22902_);
  or (_22908_, _22907_, _06474_);
  and (_22909_, _15338_, _08010_);
  or (_22910_, _22909_, _22867_);
  or (_22911_, _22910_, _07282_);
  and (_22912_, _22911_, _07284_);
  and (_22913_, _22912_, _22908_);
  and (_22914_, _12542_, _08010_);
  or (_22915_, _22914_, _22867_);
  and (_22917_, _22915_, _06582_);
  or (_22918_, _22917_, _22913_);
  and (_22919_, _22918_, _07279_);
  or (_22920_, _22867_, _08256_);
  and (_22921_, _22904_, _06478_);
  and (_22922_, _22921_, _22920_);
  or (_22923_, _22922_, _22919_);
  and (_22924_, _22923_, _07276_);
  and (_22925_, _22876_, _06569_);
  and (_22926_, _22925_, _22920_);
  or (_22928_, _22926_, _06479_);
  or (_22929_, _22928_, _22924_);
  and (_22930_, _15335_, _08010_);
  or (_22931_, _22867_, _09043_);
  or (_22932_, _22931_, _22930_);
  and (_22933_, _22932_, _09048_);
  and (_22934_, _22933_, _22929_);
  nor (_22935_, _11212_, _11757_);
  or (_22936_, _22935_, _22867_);
  and (_22937_, _22936_, _06572_);
  or (_22939_, _22937_, _06606_);
  or (_22940_, _22939_, _22934_);
  or (_22941_, _22873_, _07037_);
  and (_22942_, _22941_, _06196_);
  and (_22943_, _22942_, _22940_);
  and (_22944_, _15509_, _08010_);
  or (_22945_, _22944_, _22867_);
  and (_22946_, _22945_, _06195_);
  or (_22947_, _22946_, _01379_);
  or (_22948_, _22947_, _22943_);
  or (_22950_, _01375_, \uc8051golden_1.TL0 [5]);
  and (_22951_, _22950_, _42545_);
  and (_42949_, _22951_, _22948_);
  and (_22952_, _11757_, \uc8051golden_1.TL0 [6]);
  nor (_22953_, _11757_, _08118_);
  or (_22954_, _22953_, _22952_);
  or (_22955_, _22954_, _06293_);
  and (_22956_, _15550_, _08010_);
  or (_22957_, _22956_, _22952_);
  or (_22958_, _22957_, _07210_);
  and (_22960_, _08010_, \uc8051golden_1.ACC [6]);
  or (_22961_, _22960_, _22952_);
  and (_22962_, _22961_, _07199_);
  and (_22963_, _07200_, \uc8051golden_1.TL0 [6]);
  or (_22964_, _22963_, _06401_);
  or (_22965_, _22964_, _22962_);
  and (_22966_, _22965_, _07221_);
  and (_22967_, _22966_, _22958_);
  and (_22968_, _22954_, _06399_);
  or (_22969_, _22968_, _22967_);
  and (_22971_, _22969_, _06414_);
  and (_22972_, _22961_, _06406_);
  or (_22973_, _22972_, _10059_);
  or (_22974_, _22973_, _22971_);
  and (_22975_, _22974_, _22955_);
  or (_22976_, _22975_, _06281_);
  and (_22977_, _08010_, _09440_);
  or (_22978_, _22952_, _06282_);
  or (_22979_, _22978_, _22977_);
  and (_22980_, _22979_, _06279_);
  and (_22982_, _22980_, _22976_);
  and (_22983_, _15639_, _08010_);
  or (_22984_, _22983_, _22952_);
  and (_22985_, _22984_, _06015_);
  or (_22986_, _22985_, _06275_);
  or (_22987_, _22986_, _22982_);
  and (_22988_, _15646_, _08010_);
  or (_22989_, _22988_, _22952_);
  or (_22990_, _22989_, _06276_);
  and (_22991_, _22990_, _22987_);
  or (_22993_, _22991_, _06474_);
  and (_22994_, _15531_, _08010_);
  or (_22995_, _22994_, _22952_);
  or (_22996_, _22995_, _07282_);
  and (_22997_, _22996_, _07284_);
  and (_22998_, _22997_, _22993_);
  and (_22999_, _11210_, _08010_);
  or (_23000_, _22999_, _22952_);
  and (_23001_, _23000_, _06582_);
  or (_23002_, _23001_, _22998_);
  and (_23004_, _23002_, _07279_);
  or (_23005_, _22952_, _08162_);
  and (_23006_, _22989_, _06478_);
  and (_23007_, _23006_, _23005_);
  or (_23008_, _23007_, _23004_);
  and (_23009_, _23008_, _07276_);
  and (_23010_, _22961_, _06569_);
  and (_23011_, _23010_, _23005_);
  or (_23012_, _23011_, _06479_);
  or (_23013_, _23012_, _23009_);
  and (_23015_, _15528_, _08010_);
  or (_23016_, _22952_, _09043_);
  or (_23017_, _23016_, _23015_);
  and (_23018_, _23017_, _09048_);
  and (_23019_, _23018_, _23013_);
  nor (_23020_, _11209_, _11757_);
  or (_23021_, _23020_, _22952_);
  and (_23022_, _23021_, _06572_);
  or (_23023_, _23022_, _06606_);
  or (_23024_, _23023_, _23019_);
  or (_23026_, _22957_, _07037_);
  and (_23027_, _23026_, _06196_);
  and (_23028_, _23027_, _23024_);
  and (_23029_, _15713_, _08010_);
  or (_23030_, _23029_, _22952_);
  and (_23031_, _23030_, _06195_);
  or (_23032_, _23031_, _01379_);
  or (_23033_, _23032_, _23028_);
  or (_23034_, _01375_, \uc8051golden_1.TL0 [6]);
  and (_23035_, _23034_, _42545_);
  and (_42950_, _23035_, _23033_);
  not (_23037_, \uc8051golden_1.TCON [0]);
  nor (_23038_, _01375_, _23037_);
  nand (_23039_, _11225_, _08017_);
  nor (_23040_, _08017_, _23037_);
  nor (_23041_, _23040_, _07276_);
  nand (_23042_, _23041_, _23039_);
  nor (_23043_, _08521_, _11836_);
  or (_23044_, _23043_, _23040_);
  and (_23045_, _23044_, _06401_);
  nor (_23047_, _07199_, _23037_);
  and (_23048_, _08017_, \uc8051golden_1.ACC [0]);
  or (_23049_, _23048_, _23040_);
  and (_23050_, _23049_, _07199_);
  or (_23051_, _23050_, _23047_);
  and (_23052_, _23051_, _07210_);
  or (_23053_, _23052_, _06395_);
  or (_23054_, _23053_, _23045_);
  and (_23055_, _14339_, _08623_);
  nor (_23056_, _08623_, _23037_);
  or (_23058_, _23056_, _06396_);
  or (_23059_, _23058_, _23055_);
  and (_23060_, _23059_, _07221_);
  and (_23061_, _23060_, _23054_);
  and (_23062_, _08017_, _07473_);
  or (_23063_, _23062_, _23040_);
  and (_23064_, _23063_, _06399_);
  or (_23065_, _23064_, _06406_);
  or (_23066_, _23065_, _23061_);
  or (_23067_, _23049_, _06414_);
  and (_23069_, _23067_, _06844_);
  and (_23070_, _23069_, _23066_);
  and (_23071_, _23040_, _06393_);
  or (_23072_, _23071_, _06387_);
  or (_23073_, _23072_, _23070_);
  or (_23074_, _23044_, _07245_);
  and (_23075_, _23074_, _06446_);
  and (_23076_, _23075_, _23073_);
  and (_23077_, _14371_, _08623_);
  or (_23078_, _23077_, _23056_);
  and (_23080_, _23078_, _06300_);
  or (_23081_, _23080_, _10059_);
  or (_23082_, _23081_, _23076_);
  or (_23083_, _23063_, _06293_);
  and (_23084_, _23083_, _23082_);
  or (_23085_, _23084_, _06281_);
  and (_23086_, _08017_, _09446_);
  or (_23087_, _23040_, _06282_);
  or (_23088_, _23087_, _23086_);
  and (_23089_, _23088_, _06279_);
  and (_23090_, _23089_, _23085_);
  and (_23091_, _14426_, _08017_);
  or (_23092_, _23091_, _23040_);
  and (_23093_, _23092_, _06015_);
  or (_23094_, _23093_, _06275_);
  or (_23095_, _23094_, _23090_);
  and (_23096_, _08017_, _08817_);
  or (_23097_, _23096_, _23040_);
  or (_23098_, _23097_, _06276_);
  and (_23099_, _23098_, _23095_);
  or (_23102_, _23099_, _06474_);
  and (_23103_, _14324_, _08017_);
  or (_23104_, _23103_, _23040_);
  or (_23105_, _23104_, _07282_);
  and (_23106_, _23105_, _07284_);
  and (_23107_, _23106_, _23102_);
  nor (_23108_, _12538_, _11836_);
  or (_23109_, _23108_, _23040_);
  and (_23110_, _23039_, _06582_);
  and (_23111_, _23110_, _23109_);
  or (_23113_, _23111_, _23107_);
  and (_23114_, _23113_, _07279_);
  nand (_23115_, _23097_, _06478_);
  nor (_23116_, _23115_, _23043_);
  or (_23117_, _23116_, _06569_);
  or (_23118_, _23117_, _23114_);
  and (_23119_, _23118_, _23042_);
  or (_23120_, _23119_, _06479_);
  and (_23121_, _14320_, _08017_);
  or (_23122_, _23040_, _09043_);
  or (_23124_, _23122_, _23121_);
  and (_23125_, _23124_, _09048_);
  and (_23126_, _23125_, _23120_);
  and (_23127_, _23109_, _06572_);
  or (_23128_, _23127_, _06606_);
  or (_23129_, _23128_, _23126_);
  or (_23130_, _23044_, _07037_);
  and (_23131_, _23130_, _23129_);
  or (_23132_, _23131_, _06234_);
  or (_23133_, _23040_, _06807_);
  and (_23135_, _23133_, _23132_);
  or (_23136_, _23135_, _06195_);
  or (_23137_, _23044_, _06196_);
  and (_23138_, _23137_, _01375_);
  and (_23139_, _23138_, _23136_);
  or (_23140_, _23139_, _23038_);
  and (_42952_, _23140_, _42545_);
  not (_23141_, \uc8051golden_1.TCON [1]);
  nor (_23142_, _01375_, _23141_);
  nor (_23143_, _08017_, _23141_);
  nor (_23145_, _11223_, _11836_);
  or (_23146_, _23145_, _23143_);
  or (_23147_, _23146_, _09048_);
  nor (_23148_, _11836_, _07196_);
  or (_23149_, _23148_, _23143_);
  or (_23150_, _23149_, _07221_);
  or (_23151_, _08017_, \uc8051golden_1.TCON [1]);
  and (_23152_, _14532_, _08017_);
  not (_23153_, _23152_);
  and (_23154_, _23153_, _23151_);
  or (_23156_, _23154_, _07210_);
  and (_23157_, _08017_, \uc8051golden_1.ACC [1]);
  or (_23158_, _23157_, _23143_);
  and (_23159_, _23158_, _07199_);
  nor (_23160_, _07199_, _23141_);
  or (_23161_, _23160_, _06401_);
  or (_23162_, _23161_, _23159_);
  and (_23163_, _23162_, _06396_);
  and (_23164_, _23163_, _23156_);
  nor (_23165_, _08623_, _23141_);
  and (_23167_, _14514_, _08623_);
  or (_23168_, _23167_, _23165_);
  and (_23169_, _23168_, _06395_);
  or (_23170_, _23169_, _06399_);
  or (_23171_, _23170_, _23164_);
  and (_23172_, _23171_, _23150_);
  or (_23173_, _23172_, _06406_);
  or (_23174_, _23158_, _06414_);
  and (_23175_, _23174_, _06844_);
  and (_23176_, _23175_, _23173_);
  and (_23178_, _14517_, _08623_);
  or (_23179_, _23178_, _23165_);
  and (_23180_, _23179_, _06393_);
  or (_23181_, _23180_, _06387_);
  or (_23182_, _23181_, _23176_);
  and (_23183_, _23167_, _14513_);
  or (_23184_, _23165_, _07245_);
  or (_23185_, _23184_, _23183_);
  and (_23186_, _23185_, _06446_);
  and (_23187_, _23186_, _23182_);
  or (_23189_, _23165_, _14560_);
  and (_23190_, _23189_, _06300_);
  and (_23191_, _23190_, _23168_);
  or (_23192_, _23191_, _10059_);
  or (_23193_, _23192_, _23187_);
  or (_23194_, _23149_, _06293_);
  and (_23195_, _23194_, _23193_);
  or (_23196_, _23195_, _06281_);
  and (_23197_, _08017_, _09445_);
  or (_23198_, _23143_, _06282_);
  or (_23200_, _23198_, _23197_);
  and (_23201_, _23200_, _06279_);
  and (_23202_, _23201_, _23196_);
  and (_23203_, _14615_, _08017_);
  or (_23204_, _23203_, _23143_);
  and (_23205_, _23204_, _06015_);
  or (_23206_, _23205_, _23202_);
  and (_23207_, _23206_, _06276_);
  nand (_23208_, _08017_, _07090_);
  and (_23209_, _23151_, _06275_);
  and (_23211_, _23209_, _23208_);
  or (_23212_, _23211_, _23207_);
  and (_23213_, _23212_, _07282_);
  or (_23214_, _14507_, _11836_);
  and (_23215_, _23151_, _06474_);
  and (_23216_, _23215_, _23214_);
  or (_23217_, _23216_, _06582_);
  or (_23218_, _23217_, _23213_);
  nand (_23219_, _11222_, _08017_);
  and (_23220_, _23219_, _23146_);
  or (_23222_, _23220_, _07284_);
  and (_23223_, _23222_, _07279_);
  and (_23224_, _23223_, _23218_);
  or (_23225_, _14505_, _11836_);
  and (_23226_, _23151_, _06478_);
  and (_23227_, _23226_, _23225_);
  or (_23228_, _23227_, _06569_);
  or (_23229_, _23228_, _23224_);
  nor (_23230_, _23143_, _07276_);
  nand (_23231_, _23230_, _23219_);
  and (_23233_, _23231_, _09043_);
  and (_23234_, _23233_, _23229_);
  or (_23235_, _23208_, _08477_);
  and (_23236_, _23151_, _06479_);
  and (_23237_, _23236_, _23235_);
  or (_23238_, _23237_, _06572_);
  or (_23239_, _23238_, _23234_);
  and (_23240_, _23239_, _23147_);
  or (_23241_, _23240_, _06606_);
  or (_23242_, _23154_, _07037_);
  and (_23244_, _23242_, _06807_);
  and (_23245_, _23244_, _23241_);
  and (_23246_, _23179_, _06234_);
  or (_23247_, _23246_, _06195_);
  or (_23248_, _23247_, _23245_);
  or (_23249_, _23143_, _06196_);
  or (_23250_, _23249_, _23152_);
  and (_23251_, _23250_, _01375_);
  and (_23252_, _23251_, _23248_);
  or (_23253_, _23252_, _23142_);
  and (_42953_, _23253_, _42545_);
  and (_23255_, _01379_, \uc8051golden_1.TCON [2]);
  and (_23256_, _11836_, \uc8051golden_1.TCON [2]);
  nor (_23257_, _11836_, _07623_);
  or (_23258_, _23257_, _23256_);
  or (_23259_, _23258_, _06293_);
  or (_23260_, _23258_, _07221_);
  and (_23261_, _14754_, _08017_);
  or (_23262_, _23261_, _23256_);
  or (_23263_, _23262_, _07210_);
  and (_23265_, _08017_, \uc8051golden_1.ACC [2]);
  or (_23266_, _23265_, _23256_);
  and (_23267_, _23266_, _07199_);
  and (_23268_, _07200_, \uc8051golden_1.TCON [2]);
  or (_23269_, _23268_, _06401_);
  or (_23270_, _23269_, _23267_);
  and (_23271_, _23270_, _06396_);
  and (_23272_, _23271_, _23263_);
  and (_23273_, _11844_, \uc8051golden_1.TCON [2]);
  and (_23274_, _14751_, _08623_);
  or (_23276_, _23274_, _23273_);
  and (_23277_, _23276_, _06395_);
  or (_23278_, _23277_, _06399_);
  or (_23279_, _23278_, _23272_);
  and (_23280_, _23279_, _23260_);
  or (_23281_, _23280_, _06406_);
  or (_23282_, _23266_, _06414_);
  and (_23283_, _23282_, _06844_);
  and (_23284_, _23283_, _23281_);
  and (_23285_, _14749_, _08623_);
  or (_23287_, _23285_, _23273_);
  and (_23288_, _23287_, _06393_);
  or (_23289_, _23288_, _06387_);
  or (_23290_, _23289_, _23284_);
  and (_23291_, _23274_, _14778_);
  or (_23292_, _23273_, _07245_);
  or (_23293_, _23292_, _23291_);
  and (_23294_, _23293_, _06446_);
  and (_23295_, _23294_, _23290_);
  and (_23296_, _14793_, _08623_);
  or (_23298_, _23296_, _23273_);
  and (_23299_, _23298_, _06300_);
  or (_23300_, _23299_, _10059_);
  or (_23301_, _23300_, _23295_);
  and (_23302_, _23301_, _23259_);
  or (_23303_, _23302_, _06281_);
  and (_23304_, _08017_, _09444_);
  or (_23305_, _23256_, _06282_);
  or (_23306_, _23305_, _23304_);
  and (_23307_, _23306_, _06279_);
  and (_23309_, _23307_, _23303_);
  and (_23310_, _14848_, _08017_);
  or (_23311_, _23310_, _23256_);
  and (_23312_, _23311_, _06015_);
  or (_23313_, _23312_, _06275_);
  or (_23314_, _23313_, _23309_);
  and (_23315_, _08017_, _08994_);
  or (_23316_, _23315_, _23256_);
  or (_23317_, _23316_, _06276_);
  and (_23318_, _23317_, _23314_);
  or (_23320_, _23318_, _06474_);
  and (_23321_, _14744_, _08017_);
  or (_23322_, _23321_, _23256_);
  or (_23323_, _23322_, _07282_);
  and (_23324_, _23323_, _07284_);
  and (_23325_, _23324_, _23320_);
  and (_23326_, _11221_, _08017_);
  or (_23327_, _23326_, _23256_);
  and (_23328_, _23327_, _06582_);
  or (_23329_, _23328_, _23325_);
  and (_23331_, _23329_, _07279_);
  or (_23332_, _23256_, _08433_);
  and (_23333_, _23316_, _06478_);
  and (_23334_, _23333_, _23332_);
  or (_23335_, _23334_, _23331_);
  and (_23336_, _23335_, _07276_);
  and (_23337_, _23266_, _06569_);
  and (_23338_, _23337_, _23332_);
  or (_23339_, _23338_, _06479_);
  or (_23340_, _23339_, _23336_);
  and (_23342_, _14741_, _08017_);
  or (_23343_, _23256_, _09043_);
  or (_23344_, _23343_, _23342_);
  and (_23345_, _23344_, _09048_);
  and (_23346_, _23345_, _23340_);
  nor (_23347_, _11220_, _11836_);
  or (_23348_, _23347_, _23256_);
  and (_23349_, _23348_, _06572_);
  or (_23350_, _23349_, _06606_);
  or (_23351_, _23350_, _23346_);
  or (_23353_, _23262_, _07037_);
  and (_23354_, _23353_, _06807_);
  and (_23355_, _23354_, _23351_);
  and (_23356_, _23287_, _06234_);
  or (_23357_, _23356_, _06195_);
  or (_23358_, _23357_, _23355_);
  and (_23359_, _14917_, _08017_);
  or (_23360_, _23256_, _06196_);
  or (_23361_, _23360_, _23359_);
  and (_23362_, _23361_, _01375_);
  and (_23364_, _23362_, _23358_);
  or (_23365_, _23364_, _23255_);
  and (_42954_, _23365_, _42545_);
  and (_23366_, _01379_, \uc8051golden_1.TCON [3]);
  and (_23367_, _11836_, \uc8051golden_1.TCON [3]);
  nor (_23368_, _11836_, _07775_);
  or (_23369_, _23368_, _23367_);
  or (_23370_, _23369_, _06293_);
  and (_23371_, _14947_, _08017_);
  or (_23372_, _23371_, _23367_);
  or (_23373_, _23372_, _07210_);
  and (_23374_, _08017_, \uc8051golden_1.ACC [3]);
  or (_23375_, _23374_, _23367_);
  and (_23376_, _23375_, _07199_);
  and (_23377_, _07200_, \uc8051golden_1.TCON [3]);
  or (_23378_, _23377_, _06401_);
  or (_23379_, _23378_, _23376_);
  and (_23380_, _23379_, _06396_);
  and (_23381_, _23380_, _23373_);
  and (_23382_, _11844_, \uc8051golden_1.TCON [3]);
  and (_23385_, _14951_, _08623_);
  or (_23386_, _23385_, _23382_);
  and (_23387_, _23386_, _06395_);
  or (_23388_, _23387_, _06399_);
  or (_23389_, _23388_, _23381_);
  or (_23390_, _23369_, _07221_);
  and (_23391_, _23390_, _23389_);
  or (_23392_, _23391_, _06406_);
  or (_23393_, _23375_, _06414_);
  and (_23394_, _23393_, _06844_);
  and (_23396_, _23394_, _23392_);
  and (_23397_, _14961_, _08623_);
  or (_23398_, _23397_, _23382_);
  and (_23399_, _23398_, _06393_);
  or (_23400_, _23399_, _06387_);
  or (_23401_, _23400_, _23396_);
  or (_23402_, _23382_, _14968_);
  and (_23403_, _23402_, _23386_);
  or (_23404_, _23403_, _07245_);
  and (_23405_, _23404_, _06446_);
  and (_23407_, _23405_, _23401_);
  and (_23408_, _14985_, _08623_);
  or (_23409_, _23408_, _23382_);
  and (_23410_, _23409_, _06300_);
  or (_23411_, _23410_, _10059_);
  or (_23412_, _23411_, _23407_);
  and (_23413_, _23412_, _23370_);
  or (_23414_, _23413_, _06281_);
  and (_23415_, _08017_, _09443_);
  or (_23416_, _23367_, _06282_);
  or (_23418_, _23416_, _23415_);
  and (_23419_, _23418_, _06279_);
  and (_23420_, _23419_, _23414_);
  and (_23421_, _15039_, _08017_);
  or (_23422_, _23421_, _23367_);
  and (_23423_, _23422_, _06015_);
  or (_23424_, _23423_, _06275_);
  or (_23425_, _23424_, _23420_);
  and (_23426_, _08017_, _08815_);
  or (_23427_, _23426_, _23367_);
  or (_23429_, _23427_, _06276_);
  and (_23430_, _23429_, _23425_);
  or (_23431_, _23430_, _06474_);
  and (_23432_, _14934_, _08017_);
  or (_23433_, _23432_, _23367_);
  or (_23434_, _23433_, _07282_);
  and (_23435_, _23434_, _07284_);
  and (_23436_, _23435_, _23431_);
  and (_23437_, _12535_, _08017_);
  or (_23438_, _23437_, _23367_);
  and (_23440_, _23438_, _06582_);
  or (_23441_, _23440_, _23436_);
  and (_23442_, _23441_, _07279_);
  or (_23443_, _23367_, _08389_);
  and (_23444_, _23427_, _06478_);
  and (_23445_, _23444_, _23443_);
  or (_23446_, _23445_, _23442_);
  and (_23447_, _23446_, _07276_);
  and (_23448_, _23375_, _06569_);
  and (_23449_, _23448_, _23443_);
  or (_23451_, _23449_, _06479_);
  or (_23452_, _23451_, _23447_);
  and (_23453_, _14931_, _08017_);
  or (_23454_, _23367_, _09043_);
  or (_23455_, _23454_, _23453_);
  and (_23456_, _23455_, _09048_);
  and (_23457_, _23456_, _23452_);
  nor (_23458_, _11218_, _11836_);
  or (_23459_, _23458_, _23367_);
  and (_23460_, _23459_, _06572_);
  or (_23462_, _23460_, _06606_);
  or (_23463_, _23462_, _23457_);
  or (_23464_, _23372_, _07037_);
  and (_23465_, _23464_, _06807_);
  and (_23466_, _23465_, _23463_);
  and (_23467_, _23398_, _06234_);
  or (_23468_, _23467_, _06195_);
  or (_23469_, _23468_, _23466_);
  and (_23470_, _15113_, _08017_);
  or (_23471_, _23367_, _06196_);
  or (_23473_, _23471_, _23470_);
  and (_23474_, _23473_, _01375_);
  and (_23475_, _23474_, _23469_);
  or (_23476_, _23475_, _23366_);
  and (_42956_, _23476_, _42545_);
  and (_23477_, _01379_, \uc8051golden_1.TCON [4]);
  and (_23478_, _11836_, \uc8051golden_1.TCON [4]);
  nor (_23479_, _11836_, _08301_);
  or (_23480_, _23479_, _23478_);
  or (_23481_, _23480_, _06293_);
  and (_23483_, _15130_, _08017_);
  or (_23484_, _23483_, _23478_);
  or (_23485_, _23484_, _07210_);
  and (_23486_, _08017_, \uc8051golden_1.ACC [4]);
  or (_23487_, _23486_, _23478_);
  and (_23488_, _23487_, _07199_);
  and (_23489_, _07200_, \uc8051golden_1.TCON [4]);
  or (_23490_, _23489_, _06401_);
  or (_23491_, _23490_, _23488_);
  and (_23492_, _23491_, _06396_);
  and (_23494_, _23492_, _23485_);
  and (_23495_, _11844_, \uc8051golden_1.TCON [4]);
  and (_23496_, _15139_, _08623_);
  or (_23497_, _23496_, _23495_);
  and (_23498_, _23497_, _06395_);
  or (_23499_, _23498_, _06399_);
  or (_23500_, _23499_, _23494_);
  or (_23501_, _23480_, _07221_);
  and (_23502_, _23501_, _23500_);
  or (_23503_, _23502_, _06406_);
  or (_23505_, _23487_, _06414_);
  and (_23506_, _23505_, _06844_);
  and (_23507_, _23506_, _23503_);
  and (_23508_, _15168_, _08623_);
  or (_23509_, _23508_, _23495_);
  and (_23510_, _23509_, _06393_);
  or (_23511_, _23510_, _06387_);
  or (_23512_, _23511_, _23507_);
  or (_23513_, _23495_, _15138_);
  and (_23514_, _23513_, _23497_);
  or (_23516_, _23514_, _07245_);
  and (_23517_, _23516_, _06446_);
  and (_23518_, _23517_, _23512_);
  and (_23519_, _15189_, _08623_);
  or (_23520_, _23519_, _23495_);
  and (_23521_, _23520_, _06300_);
  or (_23522_, _23521_, _10059_);
  or (_23523_, _23522_, _23518_);
  and (_23524_, _23523_, _23481_);
  or (_23525_, _23524_, _06281_);
  and (_23527_, _08017_, _09442_);
  or (_23528_, _23478_, _06282_);
  or (_23529_, _23528_, _23527_);
  and (_23530_, _23529_, _06279_);
  and (_23531_, _23530_, _23525_);
  and (_23532_, _15243_, _08017_);
  or (_23533_, _23532_, _23478_);
  and (_23534_, _23533_, _06015_);
  or (_23535_, _23534_, _06275_);
  or (_23536_, _23535_, _23531_);
  and (_23538_, _08883_, _08017_);
  or (_23539_, _23538_, _23478_);
  or (_23540_, _23539_, _06276_);
  and (_23541_, _23540_, _23536_);
  or (_23542_, _23541_, _06474_);
  and (_23543_, _15135_, _08017_);
  or (_23544_, _23543_, _23478_);
  or (_23545_, _23544_, _07282_);
  and (_23546_, _23545_, _07284_);
  and (_23547_, _23546_, _23542_);
  and (_23549_, _11216_, _08017_);
  or (_23550_, _23549_, _23478_);
  and (_23551_, _23550_, _06582_);
  or (_23552_, _23551_, _23547_);
  and (_23553_, _23552_, _07279_);
  or (_23554_, _23478_, _08345_);
  and (_23555_, _23539_, _06478_);
  and (_23556_, _23555_, _23554_);
  or (_23557_, _23556_, _23553_);
  and (_23558_, _23557_, _07276_);
  and (_23560_, _23487_, _06569_);
  and (_23561_, _23560_, _23554_);
  or (_23562_, _23561_, _06479_);
  or (_23563_, _23562_, _23558_);
  and (_23564_, _15134_, _08017_);
  or (_23565_, _23478_, _09043_);
  or (_23566_, _23565_, _23564_);
  and (_23567_, _23566_, _09048_);
  and (_23568_, _23567_, _23563_);
  nor (_23569_, _11215_, _11836_);
  or (_23571_, _23569_, _23478_);
  and (_23572_, _23571_, _06572_);
  or (_23573_, _23572_, _06606_);
  or (_23574_, _23573_, _23568_);
  or (_23575_, _23484_, _07037_);
  and (_23576_, _23575_, _06807_);
  and (_23577_, _23576_, _23574_);
  and (_23578_, _23509_, _06234_);
  or (_23579_, _23578_, _06195_);
  or (_23580_, _23579_, _23577_);
  and (_23582_, _15315_, _08017_);
  or (_23583_, _23478_, _06196_);
  or (_23584_, _23583_, _23582_);
  and (_23585_, _23584_, _01375_);
  and (_23586_, _23585_, _23580_);
  or (_23587_, _23586_, _23477_);
  and (_42957_, _23587_, _42545_);
  and (_23588_, _01379_, \uc8051golden_1.TCON [5]);
  and (_23589_, _11836_, \uc8051golden_1.TCON [5]);
  nor (_23590_, _11836_, _08207_);
  or (_23592_, _23590_, _23589_);
  or (_23593_, _23592_, _06293_);
  and (_23594_, _15348_, _08017_);
  or (_23595_, _23594_, _23589_);
  or (_23596_, _23595_, _07210_);
  and (_23597_, _08017_, \uc8051golden_1.ACC [5]);
  or (_23598_, _23597_, _23589_);
  and (_23599_, _23598_, _07199_);
  and (_23600_, _07200_, \uc8051golden_1.TCON [5]);
  or (_23601_, _23600_, _06401_);
  or (_23602_, _23601_, _23599_);
  and (_23603_, _23602_, _06396_);
  and (_23604_, _23603_, _23596_);
  and (_23605_, _11844_, \uc8051golden_1.TCON [5]);
  and (_23606_, _15341_, _08623_);
  or (_23607_, _23606_, _23605_);
  and (_23608_, _23607_, _06395_);
  or (_23609_, _23608_, _06399_);
  or (_23610_, _23609_, _23604_);
  or (_23611_, _23592_, _07221_);
  and (_23613_, _23611_, _23610_);
  or (_23614_, _23613_, _06406_);
  or (_23615_, _23598_, _06414_);
  and (_23616_, _23615_, _06844_);
  and (_23617_, _23616_, _23614_);
  and (_23618_, _15345_, _08623_);
  or (_23619_, _23618_, _23605_);
  and (_23620_, _23619_, _06393_);
  or (_23621_, _23620_, _06387_);
  or (_23622_, _23621_, _23617_);
  or (_23624_, _23605_, _15378_);
  and (_23625_, _23624_, _23607_);
  or (_23626_, _23625_, _07245_);
  and (_23627_, _23626_, _06446_);
  and (_23628_, _23627_, _23622_);
  or (_23629_, _23605_, _15342_);
  and (_23630_, _23629_, _06300_);
  and (_23631_, _23630_, _23607_);
  or (_23632_, _23631_, _10059_);
  or (_23633_, _23632_, _23628_);
  and (_23635_, _23633_, _23593_);
  or (_23636_, _23635_, _06281_);
  and (_23637_, _08017_, _09441_);
  or (_23638_, _23589_, _06282_);
  or (_23639_, _23638_, _23637_);
  and (_23640_, _23639_, _06279_);
  and (_23641_, _23640_, _23636_);
  and (_23642_, _15446_, _08017_);
  or (_23643_, _23642_, _23589_);
  and (_23644_, _23643_, _06015_);
  or (_23645_, _23644_, _06275_);
  or (_23646_, _23645_, _23641_);
  and (_23647_, _08958_, _08017_);
  or (_23648_, _23647_, _23589_);
  or (_23649_, _23648_, _06276_);
  and (_23650_, _23649_, _23646_);
  or (_23651_, _23650_, _06474_);
  and (_23652_, _15338_, _08017_);
  or (_23653_, _23652_, _23589_);
  or (_23654_, _23653_, _07282_);
  and (_23656_, _23654_, _07284_);
  and (_23657_, _23656_, _23651_);
  and (_23658_, _12542_, _08017_);
  or (_23659_, _23658_, _23589_);
  and (_23660_, _23659_, _06582_);
  or (_23661_, _23660_, _23657_);
  and (_23662_, _23661_, _07279_);
  or (_23663_, _23589_, _08256_);
  and (_23664_, _23648_, _06478_);
  and (_23665_, _23664_, _23663_);
  or (_23666_, _23665_, _23662_);
  and (_23667_, _23666_, _07276_);
  and (_23668_, _23598_, _06569_);
  and (_23669_, _23668_, _23663_);
  or (_23670_, _23669_, _06479_);
  or (_23671_, _23670_, _23667_);
  and (_23672_, _15335_, _08017_);
  or (_23673_, _23589_, _09043_);
  or (_23674_, _23673_, _23672_);
  and (_23675_, _23674_, _09048_);
  and (_23677_, _23675_, _23671_);
  nor (_23678_, _11212_, _11836_);
  or (_23679_, _23678_, _23589_);
  and (_23680_, _23679_, _06572_);
  or (_23681_, _23680_, _06606_);
  or (_23682_, _23681_, _23677_);
  or (_23683_, _23595_, _07037_);
  and (_23684_, _23683_, _06807_);
  and (_23685_, _23684_, _23682_);
  and (_23686_, _23619_, _06234_);
  or (_23688_, _23686_, _06195_);
  or (_23689_, _23688_, _23685_);
  and (_23690_, _15509_, _08017_);
  or (_23691_, _23589_, _06196_);
  or (_23692_, _23691_, _23690_);
  and (_23693_, _23692_, _01375_);
  and (_23694_, _23693_, _23689_);
  or (_23695_, _23694_, _23588_);
  and (_42958_, _23695_, _42545_);
  and (_23696_, _01379_, \uc8051golden_1.TCON [6]);
  and (_23697_, _11836_, \uc8051golden_1.TCON [6]);
  nor (_23698_, _11836_, _08118_);
  or (_23699_, _23698_, _23697_);
  or (_23700_, _23699_, _06293_);
  and (_23701_, _15550_, _08017_);
  or (_23702_, _23701_, _23697_);
  or (_23703_, _23702_, _07210_);
  and (_23704_, _08017_, \uc8051golden_1.ACC [6]);
  or (_23705_, _23704_, _23697_);
  and (_23706_, _23705_, _07199_);
  and (_23708_, _07200_, \uc8051golden_1.TCON [6]);
  or (_23709_, _23708_, _06401_);
  or (_23710_, _23709_, _23706_);
  and (_23711_, _23710_, _06396_);
  and (_23712_, _23711_, _23703_);
  and (_23713_, _11844_, \uc8051golden_1.TCON [6]);
  and (_23714_, _15535_, _08623_);
  or (_23715_, _23714_, _23713_);
  and (_23716_, _23715_, _06395_);
  or (_23717_, _23716_, _06399_);
  or (_23719_, _23717_, _23712_);
  or (_23720_, _23699_, _07221_);
  and (_23721_, _23720_, _23719_);
  or (_23722_, _23721_, _06406_);
  or (_23723_, _23705_, _06414_);
  and (_23724_, _23723_, _06844_);
  and (_23725_, _23724_, _23722_);
  and (_23726_, _15561_, _08623_);
  or (_23727_, _23726_, _23713_);
  and (_23728_, _23727_, _06393_);
  or (_23729_, _23728_, _06387_);
  or (_23730_, _23729_, _23725_);
  or (_23731_, _23713_, _15568_);
  and (_23732_, _23731_, _23715_);
  or (_23733_, _23732_, _07245_);
  and (_23734_, _23733_, _06446_);
  and (_23735_, _23734_, _23730_);
  and (_23736_, _15585_, _08623_);
  or (_23737_, _23736_, _23713_);
  and (_23738_, _23737_, _06300_);
  or (_23740_, _23738_, _10059_);
  or (_23741_, _23740_, _23735_);
  and (_23742_, _23741_, _23700_);
  or (_23743_, _23742_, _06281_);
  and (_23744_, _08017_, _09440_);
  or (_23745_, _23697_, _06282_);
  or (_23746_, _23745_, _23744_);
  and (_23747_, _23746_, _06279_);
  and (_23748_, _23747_, _23743_);
  and (_23749_, _15639_, _08017_);
  or (_23751_, _23749_, _23697_);
  and (_23752_, _23751_, _06015_);
  or (_23753_, _23752_, _06275_);
  or (_23754_, _23753_, _23748_);
  and (_23755_, _15646_, _08017_);
  or (_23756_, _23755_, _23697_);
  or (_23757_, _23756_, _06276_);
  and (_23758_, _23757_, _23754_);
  or (_23759_, _23758_, _06474_);
  and (_23760_, _15531_, _08017_);
  or (_23761_, _23760_, _23697_);
  or (_23762_, _23761_, _07282_);
  and (_23763_, _23762_, _07284_);
  and (_23764_, _23763_, _23759_);
  and (_23765_, _11210_, _08017_);
  or (_23766_, _23765_, _23697_);
  and (_23767_, _23766_, _06582_);
  or (_23768_, _23767_, _23764_);
  and (_23769_, _23768_, _07279_);
  or (_23770_, _23697_, _08162_);
  and (_23772_, _23756_, _06478_);
  and (_23773_, _23772_, _23770_);
  or (_23774_, _23773_, _23769_);
  and (_23775_, _23774_, _07276_);
  and (_23776_, _23705_, _06569_);
  and (_23777_, _23776_, _23770_);
  or (_23778_, _23777_, _06479_);
  or (_23779_, _23778_, _23775_);
  and (_23780_, _15528_, _08017_);
  or (_23781_, _23697_, _09043_);
  or (_23783_, _23781_, _23780_);
  and (_23784_, _23783_, _09048_);
  and (_23785_, _23784_, _23779_);
  nor (_23786_, _11209_, _11836_);
  or (_23787_, _23786_, _23697_);
  and (_23788_, _23787_, _06572_);
  or (_23789_, _23788_, _06606_);
  or (_23790_, _23789_, _23785_);
  or (_23791_, _23702_, _07037_);
  and (_23792_, _23791_, _06807_);
  and (_23793_, _23792_, _23790_);
  and (_23794_, _23727_, _06234_);
  or (_23795_, _23794_, _06195_);
  or (_23796_, _23795_, _23793_);
  and (_23797_, _15713_, _08017_);
  or (_23798_, _23697_, _06196_);
  or (_23799_, _23798_, _23797_);
  and (_23800_, _23799_, _01375_);
  and (_23801_, _23800_, _23796_);
  or (_23802_, _23801_, _23696_);
  and (_42959_, _23802_, _42545_);
  not (_23803_, \uc8051golden_1.TH1 [0]);
  nor (_23804_, _01375_, _23803_);
  nand (_23805_, _11225_, _07980_);
  nor (_23806_, _07980_, _23803_);
  nor (_23807_, _23806_, _07276_);
  nand (_23808_, _23807_, _23805_);
  nor (_23809_, _08521_, _11938_);
  or (_23810_, _23809_, _23806_);
  or (_23811_, _23810_, _07210_);
  and (_23814_, _07980_, \uc8051golden_1.ACC [0]);
  or (_23815_, _23814_, _23806_);
  and (_23816_, _23815_, _07199_);
  nor (_23817_, _07199_, _23803_);
  or (_23818_, _23817_, _06401_);
  or (_23819_, _23818_, _23816_);
  and (_23820_, _23819_, _07221_);
  and (_23821_, _23820_, _23811_);
  and (_23822_, _07980_, _07473_);
  or (_23823_, _23822_, _23806_);
  and (_23824_, _23823_, _06399_);
  or (_23825_, _23824_, _23821_);
  and (_23826_, _23825_, _06414_);
  and (_23827_, _23815_, _06406_);
  or (_23828_, _23827_, _10059_);
  or (_23829_, _23828_, _23826_);
  or (_23830_, _23823_, _06293_);
  and (_23831_, _23830_, _23829_);
  or (_23832_, _23831_, _06281_);
  and (_23833_, _07980_, _09446_);
  or (_23835_, _23806_, _06282_);
  or (_23836_, _23835_, _23833_);
  and (_23837_, _23836_, _23832_);
  or (_23838_, _23837_, _06015_);
  and (_23839_, _14426_, _07980_);
  or (_23840_, _23806_, _06279_);
  or (_23841_, _23840_, _23839_);
  and (_23842_, _23841_, _06276_);
  and (_23843_, _23842_, _23838_);
  and (_23844_, _07980_, _08817_);
  or (_23846_, _23844_, _23806_);
  and (_23847_, _23846_, _06275_);
  or (_23848_, _23847_, _06474_);
  or (_23849_, _23848_, _23843_);
  and (_23850_, _14324_, _07980_);
  or (_23851_, _23850_, _23806_);
  or (_23852_, _23851_, _07282_);
  and (_23853_, _23852_, _07284_);
  and (_23854_, _23853_, _23849_);
  nor (_23855_, _12538_, _11938_);
  or (_23856_, _23855_, _23806_);
  and (_23857_, _23805_, _06582_);
  and (_23858_, _23857_, _23856_);
  or (_23859_, _23858_, _23854_);
  and (_23860_, _23859_, _07279_);
  nand (_23861_, _23846_, _06478_);
  nor (_23862_, _23861_, _23809_);
  or (_23863_, _23862_, _06569_);
  or (_23864_, _23863_, _23860_);
  and (_23865_, _23864_, _23808_);
  or (_23867_, _23865_, _06479_);
  and (_23868_, _14320_, _07980_);
  or (_23869_, _23806_, _09043_);
  or (_23870_, _23869_, _23868_);
  and (_23871_, _23870_, _09048_);
  and (_23872_, _23871_, _23867_);
  and (_23873_, _23856_, _06572_);
  or (_23874_, _23873_, _19434_);
  or (_23875_, _23874_, _23872_);
  or (_23876_, _23810_, _06700_);
  and (_23878_, _23876_, _01375_);
  and (_23879_, _23878_, _23875_);
  or (_23880_, _23879_, _23804_);
  and (_42960_, _23880_, _42545_);
  and (_23881_, _01379_, \uc8051golden_1.TH1 [1]);
  nand (_23882_, _07980_, _07090_);
  or (_23883_, _07980_, \uc8051golden_1.TH1 [1]);
  and (_23884_, _23883_, _06275_);
  and (_23885_, _23884_, _23882_);
  and (_23886_, _07980_, _09445_);
  and (_23887_, _11938_, \uc8051golden_1.TH1 [1]);
  or (_23888_, _23887_, _06282_);
  or (_23889_, _23888_, _23886_);
  nor (_23890_, _11938_, _07196_);
  and (_23891_, _06293_, _07221_);
  or (_23892_, _23891_, _23887_);
  or (_23893_, _23892_, _23890_);
  and (_23894_, _07980_, \uc8051golden_1.ACC [1]);
  or (_23895_, _23894_, _23887_);
  and (_23896_, _23895_, _06406_);
  or (_23898_, _23896_, _10059_);
  and (_23899_, _14532_, _07980_);
  not (_23900_, _23899_);
  and (_23901_, _23900_, _23883_);
  and (_23902_, _23901_, _06401_);
  and (_23903_, _07200_, \uc8051golden_1.TH1 [1]);
  and (_23904_, _23895_, _07199_);
  or (_23905_, _23904_, _23903_);
  and (_23906_, _23905_, _07210_);
  or (_23907_, _23906_, _06399_);
  or (_23909_, _23907_, _23902_);
  and (_23910_, _23909_, _06414_);
  or (_23911_, _23910_, _23898_);
  and (_23912_, _23911_, _23893_);
  or (_23913_, _23912_, _06281_);
  and (_23914_, _23913_, _06279_);
  and (_23915_, _23914_, _23889_);
  or (_23916_, _14615_, _11938_);
  and (_23917_, _23883_, _06015_);
  and (_23918_, _23917_, _23916_);
  or (_23919_, _23918_, _23915_);
  and (_23920_, _23919_, _06276_);
  or (_23921_, _23920_, _23885_);
  and (_23922_, _23921_, _07282_);
  or (_23923_, _14507_, _11938_);
  and (_23924_, _23883_, _06474_);
  and (_23925_, _23924_, _23923_);
  or (_23926_, _23925_, _06582_);
  or (_23927_, _23926_, _23922_);
  and (_23928_, _11224_, _07980_);
  or (_23930_, _23928_, _23887_);
  or (_23931_, _23930_, _07284_);
  and (_23932_, _23931_, _07279_);
  and (_23933_, _23932_, _23927_);
  or (_23934_, _14505_, _11938_);
  and (_23935_, _23883_, _06478_);
  and (_23936_, _23935_, _23934_);
  or (_23937_, _23936_, _06569_);
  or (_23938_, _23937_, _23933_);
  and (_23939_, _23894_, _08477_);
  or (_23941_, _23887_, _07276_);
  or (_23942_, _23941_, _23939_);
  and (_23943_, _23942_, _09043_);
  and (_23944_, _23943_, _23938_);
  or (_23945_, _23882_, _08477_);
  and (_23946_, _23883_, _06479_);
  and (_23947_, _23946_, _23945_);
  or (_23948_, _23947_, _06572_);
  or (_23949_, _23948_, _23944_);
  nor (_23950_, _11223_, _11938_);
  or (_23951_, _23950_, _23887_);
  or (_23952_, _23951_, _09048_);
  and (_23953_, _23952_, _07037_);
  and (_23954_, _23953_, _23949_);
  and (_23955_, _23901_, _06606_);
  or (_23956_, _23955_, _06195_);
  or (_23957_, _23956_, _23954_);
  or (_23958_, _23887_, _06196_);
  or (_23959_, _23958_, _23899_);
  and (_23960_, _23959_, _01375_);
  and (_23962_, _23960_, _23957_);
  or (_23963_, _23962_, _23881_);
  and (_42961_, _23963_, _42545_);
  and (_23964_, _01379_, \uc8051golden_1.TH1 [2]);
  and (_23965_, _11938_, \uc8051golden_1.TH1 [2]);
  and (_23966_, _14754_, _07980_);
  or (_23967_, _23966_, _23965_);
  or (_23968_, _23967_, _07210_);
  and (_23969_, _07980_, \uc8051golden_1.ACC [2]);
  or (_23970_, _23969_, _23965_);
  and (_23972_, _23970_, _07199_);
  and (_23973_, _07200_, \uc8051golden_1.TH1 [2]);
  or (_23974_, _23973_, _06401_);
  or (_23975_, _23974_, _23972_);
  and (_23976_, _23975_, _07221_);
  and (_23977_, _23976_, _23968_);
  nor (_23978_, _11938_, _07623_);
  or (_23979_, _23978_, _23965_);
  and (_23980_, _23979_, _06399_);
  or (_23981_, _23980_, _23977_);
  and (_23982_, _23981_, _06414_);
  and (_23983_, _23970_, _06406_);
  or (_23984_, _23983_, _10059_);
  or (_23985_, _23984_, _23982_);
  or (_23986_, _23979_, _06293_);
  and (_23987_, _23986_, _23985_);
  or (_23988_, _23987_, _06281_);
  and (_23989_, _07980_, _09444_);
  or (_23990_, _23965_, _06282_);
  or (_23991_, _23990_, _23989_);
  and (_23993_, _23991_, _23988_);
  or (_23994_, _23993_, _06015_);
  and (_23995_, _14848_, _07980_);
  or (_23996_, _23965_, _06279_);
  or (_23997_, _23996_, _23995_);
  and (_23998_, _23997_, _06276_);
  and (_23999_, _23998_, _23994_);
  and (_24000_, _07980_, _08994_);
  or (_24001_, _24000_, _23965_);
  and (_24002_, _24001_, _06275_);
  or (_24004_, _24002_, _06474_);
  or (_24005_, _24004_, _23999_);
  and (_24006_, _14744_, _07980_);
  or (_24007_, _24006_, _23965_);
  or (_24008_, _24007_, _07282_);
  and (_24009_, _24008_, _07284_);
  and (_24010_, _24009_, _24005_);
  and (_24011_, _11221_, _07980_);
  or (_24012_, _24011_, _23965_);
  and (_24013_, _24012_, _06582_);
  or (_24015_, _24013_, _24010_);
  and (_24016_, _24015_, _07279_);
  or (_24017_, _23965_, _08433_);
  and (_24018_, _24001_, _06478_);
  and (_24019_, _24018_, _24017_);
  or (_24020_, _24019_, _24016_);
  and (_24021_, _24020_, _07276_);
  and (_24022_, _23970_, _06569_);
  and (_24023_, _24022_, _24017_);
  or (_24024_, _24023_, _06479_);
  or (_24025_, _24024_, _24021_);
  and (_24026_, _14741_, _07980_);
  or (_24027_, _23965_, _09043_);
  or (_24028_, _24027_, _24026_);
  and (_24029_, _24028_, _09048_);
  and (_24030_, _24029_, _24025_);
  nor (_24031_, _11220_, _11938_);
  or (_24032_, _24031_, _23965_);
  and (_24033_, _24032_, _06572_);
  or (_24034_, _24033_, _24030_);
  and (_24036_, _24034_, _07037_);
  and (_24037_, _23967_, _06606_);
  or (_24038_, _24037_, _06195_);
  or (_24039_, _24038_, _24036_);
  and (_24040_, _14917_, _07980_);
  or (_24041_, _23965_, _06196_);
  or (_24042_, _24041_, _24040_);
  and (_24043_, _24042_, _01375_);
  and (_24044_, _24043_, _24039_);
  or (_24045_, _24044_, _23964_);
  and (_42962_, _24045_, _42545_);
  and (_24047_, _11938_, \uc8051golden_1.TH1 [3]);
  and (_24048_, _07980_, _09443_);
  or (_24049_, _24048_, _24047_);
  and (_24050_, _24049_, _06281_);
  and (_24051_, _14947_, _07980_);
  or (_24052_, _24051_, _24047_);
  or (_24053_, _24052_, _07210_);
  and (_24054_, _07980_, \uc8051golden_1.ACC [3]);
  or (_24055_, _24054_, _24047_);
  and (_24056_, _24055_, _07199_);
  and (_24057_, _07200_, \uc8051golden_1.TH1 [3]);
  or (_24058_, _24057_, _06401_);
  or (_24059_, _24058_, _24056_);
  and (_24060_, _24059_, _07221_);
  and (_24061_, _24060_, _24053_);
  nor (_24062_, _11938_, _07775_);
  or (_24063_, _24062_, _24047_);
  and (_24064_, _24063_, _06399_);
  or (_24065_, _24064_, _24061_);
  and (_24067_, _24065_, _06414_);
  and (_24068_, _24055_, _06406_);
  or (_24069_, _24068_, _10059_);
  or (_24070_, _24069_, _24067_);
  or (_24071_, _24063_, _06293_);
  and (_24072_, _24071_, _06282_);
  and (_24073_, _24072_, _24070_);
  or (_24074_, _24073_, _06015_);
  or (_24075_, _24074_, _24050_);
  and (_24076_, _15039_, _07980_);
  or (_24078_, _24047_, _06279_);
  or (_24079_, _24078_, _24076_);
  and (_24080_, _24079_, _06276_);
  and (_24081_, _24080_, _24075_);
  and (_24082_, _07980_, _08815_);
  or (_24083_, _24082_, _24047_);
  and (_24084_, _24083_, _06275_);
  or (_24085_, _24084_, _06474_);
  or (_24086_, _24085_, _24081_);
  and (_24087_, _14934_, _07980_);
  or (_24089_, _24087_, _24047_);
  or (_24090_, _24089_, _07282_);
  and (_24091_, _24090_, _07284_);
  and (_24092_, _24091_, _24086_);
  and (_24093_, _12535_, _07980_);
  or (_24094_, _24093_, _24047_);
  and (_24095_, _24094_, _06582_);
  or (_24096_, _24095_, _24092_);
  and (_24097_, _24096_, _07279_);
  or (_24098_, _24047_, _08389_);
  and (_24099_, _24083_, _06478_);
  and (_24100_, _24099_, _24098_);
  or (_24101_, _24100_, _24097_);
  and (_24102_, _24101_, _07276_);
  and (_24103_, _24055_, _06569_);
  and (_24104_, _24103_, _24098_);
  or (_24105_, _24104_, _06479_);
  or (_24106_, _24105_, _24102_);
  and (_24107_, _14931_, _07980_);
  or (_24108_, _24047_, _09043_);
  or (_24110_, _24108_, _24107_);
  and (_24111_, _24110_, _09048_);
  and (_24112_, _24111_, _24106_);
  nor (_24113_, _11218_, _11938_);
  or (_24114_, _24113_, _24047_);
  and (_24115_, _24114_, _06572_);
  or (_24116_, _24115_, _06606_);
  or (_24117_, _24116_, _24112_);
  or (_24118_, _24052_, _07037_);
  and (_24119_, _24118_, _06196_);
  and (_24121_, _24119_, _24117_);
  and (_24122_, _15113_, _07980_);
  or (_24123_, _24122_, _24047_);
  and (_24124_, _24123_, _06195_);
  or (_24125_, _24124_, _01379_);
  or (_24126_, _24125_, _24121_);
  or (_24127_, _01375_, \uc8051golden_1.TH1 [3]);
  and (_24128_, _24127_, _42545_);
  and (_42963_, _24128_, _24126_);
  and (_24129_, _11938_, \uc8051golden_1.TH1 [4]);
  and (_24130_, _15130_, _07980_);
  or (_24131_, _24130_, _24129_);
  or (_24132_, _24131_, _07210_);
  and (_24133_, _07980_, \uc8051golden_1.ACC [4]);
  or (_24134_, _24133_, _24129_);
  and (_24135_, _24134_, _07199_);
  and (_24136_, _07200_, \uc8051golden_1.TH1 [4]);
  or (_24137_, _24136_, _06401_);
  or (_24138_, _24137_, _24135_);
  and (_24139_, _24138_, _07221_);
  and (_24141_, _24139_, _24132_);
  nor (_24142_, _11938_, _08301_);
  or (_24143_, _24142_, _24129_);
  and (_24144_, _24143_, _06399_);
  or (_24145_, _24144_, _24141_);
  and (_24146_, _24145_, _06414_);
  and (_24147_, _24134_, _06406_);
  or (_24148_, _24147_, _10059_);
  or (_24149_, _24148_, _24146_);
  or (_24150_, _24143_, _06293_);
  and (_24152_, _24150_, _24149_);
  or (_24153_, _24152_, _06281_);
  and (_24154_, _07980_, _09442_);
  or (_24155_, _24129_, _06282_);
  or (_24156_, _24155_, _24154_);
  and (_24157_, _24156_, _06279_);
  and (_24158_, _24157_, _24153_);
  and (_24159_, _15243_, _07980_);
  or (_24160_, _24159_, _24129_);
  and (_24161_, _24160_, _06015_);
  or (_24163_, _24161_, _06275_);
  or (_24164_, _24163_, _24158_);
  and (_24165_, _08883_, _07980_);
  or (_24166_, _24165_, _24129_);
  or (_24167_, _24166_, _06276_);
  and (_24168_, _24167_, _24164_);
  or (_24169_, _24168_, _06474_);
  and (_24170_, _15135_, _07980_);
  or (_24171_, _24170_, _24129_);
  or (_24172_, _24171_, _07282_);
  and (_24174_, _24172_, _07284_);
  and (_24175_, _24174_, _24169_);
  and (_24176_, _11216_, _07980_);
  or (_24177_, _24176_, _24129_);
  and (_24178_, _24177_, _06582_);
  or (_24179_, _24178_, _24175_);
  and (_24180_, _24179_, _07279_);
  or (_24181_, _24129_, _08345_);
  and (_24182_, _24166_, _06478_);
  and (_24183_, _24182_, _24181_);
  or (_24185_, _24183_, _24180_);
  and (_24186_, _24185_, _07276_);
  and (_24187_, _24134_, _06569_);
  and (_24188_, _24187_, _24181_);
  or (_24189_, _24188_, _06479_);
  or (_24190_, _24189_, _24186_);
  and (_24191_, _15134_, _07980_);
  or (_24192_, _24129_, _09043_);
  or (_24193_, _24192_, _24191_);
  and (_24194_, _24193_, _09048_);
  and (_24196_, _24194_, _24190_);
  nor (_24197_, _11215_, _11938_);
  or (_24198_, _24197_, _24129_);
  and (_24199_, _24198_, _06572_);
  or (_24200_, _24199_, _06606_);
  or (_24201_, _24200_, _24196_);
  or (_24202_, _24131_, _07037_);
  and (_24203_, _24202_, _06196_);
  and (_24204_, _24203_, _24201_);
  and (_24205_, _15315_, _07980_);
  or (_24207_, _24205_, _24129_);
  and (_24208_, _24207_, _06195_);
  or (_24209_, _24208_, _01379_);
  or (_24210_, _24209_, _24204_);
  or (_24211_, _01375_, \uc8051golden_1.TH1 [4]);
  and (_24212_, _24211_, _42545_);
  and (_42964_, _24212_, _24210_);
  and (_24213_, _11938_, \uc8051golden_1.TH1 [5]);
  nor (_24214_, _11938_, _08207_);
  or (_24215_, _24214_, _24213_);
  or (_24217_, _24215_, _06293_);
  and (_24218_, _15348_, _07980_);
  or (_24219_, _24218_, _24213_);
  or (_24220_, _24219_, _07210_);
  and (_24221_, _07980_, \uc8051golden_1.ACC [5]);
  or (_24222_, _24221_, _24213_);
  and (_24223_, _24222_, _07199_);
  and (_24224_, _07200_, \uc8051golden_1.TH1 [5]);
  or (_24225_, _24224_, _06401_);
  or (_24226_, _24225_, _24223_);
  and (_24228_, _24226_, _07221_);
  and (_24229_, _24228_, _24220_);
  and (_24230_, _24215_, _06399_);
  or (_24231_, _24230_, _24229_);
  and (_24232_, _24231_, _06414_);
  and (_24233_, _24222_, _06406_);
  or (_24234_, _24233_, _10059_);
  or (_24235_, _24234_, _24232_);
  and (_24236_, _24235_, _24217_);
  or (_24237_, _24236_, _06281_);
  and (_24238_, _07980_, _09441_);
  or (_24239_, _24213_, _06282_);
  or (_24240_, _24239_, _24238_);
  and (_24241_, _24240_, _06279_);
  and (_24242_, _24241_, _24237_);
  and (_24243_, _15446_, _07980_);
  or (_24244_, _24243_, _24213_);
  and (_24245_, _24244_, _06015_);
  or (_24246_, _24245_, _06275_);
  or (_24247_, _24246_, _24242_);
  and (_24248_, _08958_, _07980_);
  or (_24249_, _24248_, _24213_);
  or (_24250_, _24249_, _06276_);
  and (_24251_, _24250_, _24247_);
  or (_24252_, _24251_, _06474_);
  and (_24253_, _15338_, _07980_);
  or (_24254_, _24253_, _24213_);
  or (_24255_, _24254_, _07282_);
  and (_24256_, _24255_, _07284_);
  and (_24257_, _24256_, _24252_);
  and (_24259_, _12542_, _07980_);
  or (_24260_, _24259_, _24213_);
  and (_24261_, _24260_, _06582_);
  or (_24262_, _24261_, _24257_);
  and (_24263_, _24262_, _07279_);
  or (_24264_, _24213_, _08256_);
  and (_24265_, _24249_, _06478_);
  and (_24266_, _24265_, _24264_);
  or (_24267_, _24266_, _24263_);
  and (_24268_, _24267_, _07276_);
  and (_24270_, _24222_, _06569_);
  and (_24271_, _24270_, _24264_);
  or (_24272_, _24271_, _06479_);
  or (_24273_, _24272_, _24268_);
  and (_24274_, _15335_, _07980_);
  or (_24275_, _24213_, _09043_);
  or (_24276_, _24275_, _24274_);
  and (_24277_, _24276_, _09048_);
  and (_24278_, _24277_, _24273_);
  nor (_24279_, _11212_, _11938_);
  or (_24282_, _24279_, _24213_);
  and (_24283_, _24282_, _06572_);
  or (_24284_, _24283_, _06606_);
  or (_24285_, _24284_, _24278_);
  or (_24286_, _24219_, _07037_);
  and (_24287_, _24286_, _06196_);
  and (_24288_, _24287_, _24285_);
  and (_24289_, _15509_, _07980_);
  or (_24290_, _24289_, _24213_);
  and (_24291_, _24290_, _06195_);
  or (_24293_, _24291_, _01379_);
  or (_24294_, _24293_, _24288_);
  or (_24295_, _01375_, \uc8051golden_1.TH1 [5]);
  and (_24296_, _24295_, _42545_);
  and (_42965_, _24296_, _24294_);
  and (_24297_, _11938_, \uc8051golden_1.TH1 [6]);
  nor (_24298_, _11938_, _08118_);
  or (_24299_, _24298_, _24297_);
  or (_24300_, _24299_, _06293_);
  and (_24301_, _15550_, _07980_);
  or (_24303_, _24301_, _24297_);
  or (_24304_, _24303_, _07210_);
  and (_24305_, _07980_, \uc8051golden_1.ACC [6]);
  or (_24306_, _24305_, _24297_);
  and (_24307_, _24306_, _07199_);
  and (_24308_, _07200_, \uc8051golden_1.TH1 [6]);
  or (_24309_, _24308_, _06401_);
  or (_24310_, _24309_, _24307_);
  and (_24311_, _24310_, _07221_);
  and (_24312_, _24311_, _24304_);
  and (_24314_, _24299_, _06399_);
  or (_24315_, _24314_, _24312_);
  and (_24316_, _24315_, _06414_);
  and (_24317_, _24306_, _06406_);
  or (_24318_, _24317_, _10059_);
  or (_24319_, _24318_, _24316_);
  and (_24320_, _24319_, _24300_);
  or (_24321_, _24320_, _06281_);
  and (_24322_, _07980_, _09440_);
  or (_24323_, _24297_, _06282_);
  or (_24325_, _24323_, _24322_);
  and (_24326_, _24325_, _06279_);
  and (_24327_, _24326_, _24321_);
  and (_24328_, _15639_, _07980_);
  or (_24329_, _24328_, _24297_);
  and (_24330_, _24329_, _06015_);
  or (_24331_, _24330_, _06275_);
  or (_24332_, _24331_, _24327_);
  and (_24333_, _15646_, _07980_);
  or (_24334_, _24333_, _24297_);
  or (_24336_, _24334_, _06276_);
  and (_24337_, _24336_, _24332_);
  or (_24338_, _24337_, _06474_);
  and (_24339_, _15531_, _07980_);
  or (_24340_, _24339_, _24297_);
  or (_24341_, _24340_, _07282_);
  and (_24342_, _24341_, _07284_);
  and (_24343_, _24342_, _24338_);
  and (_24344_, _11210_, _07980_);
  or (_24345_, _24344_, _24297_);
  and (_24347_, _24345_, _06582_);
  or (_24348_, _24347_, _24343_);
  and (_24349_, _24348_, _07279_);
  or (_24350_, _24297_, _08162_);
  and (_24351_, _24334_, _06478_);
  and (_24352_, _24351_, _24350_);
  or (_24353_, _24352_, _24349_);
  and (_24354_, _24353_, _07276_);
  and (_24355_, _24306_, _06569_);
  and (_24356_, _24355_, _24350_);
  or (_24358_, _24356_, _06479_);
  or (_24359_, _24358_, _24354_);
  and (_24360_, _15528_, _07980_);
  or (_24361_, _24297_, _09043_);
  or (_24362_, _24361_, _24360_);
  and (_24363_, _24362_, _09048_);
  and (_24364_, _24363_, _24359_);
  nor (_24365_, _11209_, _11938_);
  or (_24366_, _24365_, _24297_);
  and (_24367_, _24366_, _06572_);
  or (_24369_, _24367_, _06606_);
  or (_24370_, _24369_, _24364_);
  or (_24371_, _24303_, _07037_);
  and (_24372_, _24371_, _06196_);
  and (_24373_, _24372_, _24370_);
  and (_24374_, _15713_, _07980_);
  or (_24375_, _24374_, _24297_);
  and (_24376_, _24375_, _06195_);
  or (_24377_, _24376_, _01379_);
  or (_24378_, _24377_, _24373_);
  or (_24380_, _01375_, \uc8051golden_1.TH1 [6]);
  and (_24381_, _24380_, _42545_);
  and (_42966_, _24381_, _24378_);
  and (_24382_, _01379_, \uc8051golden_1.TH0 [0]);
  and (_24383_, _08013_, \uc8051golden_1.ACC [0]);
  and (_24384_, _24383_, _08521_);
  and (_24385_, _12016_, \uc8051golden_1.TH0 [0]);
  or (_24386_, _24385_, _07276_);
  or (_24387_, _24386_, _24384_);
  and (_24388_, _08013_, _07473_);
  or (_24390_, _24388_, _24385_);
  or (_24391_, _24390_, _06293_);
  nor (_24392_, _08521_, _12016_);
  or (_24393_, _24392_, _24385_);
  or (_24394_, _24393_, _07210_);
  or (_24395_, _24385_, _24383_);
  and (_24396_, _24395_, _07199_);
  and (_24397_, _07200_, \uc8051golden_1.TH0 [0]);
  or (_24398_, _24397_, _06401_);
  or (_24399_, _24398_, _24396_);
  and (_24401_, _24399_, _07221_);
  and (_24402_, _24401_, _24394_);
  and (_24403_, _24390_, _06399_);
  or (_24404_, _24403_, _24402_);
  and (_24405_, _24404_, _06414_);
  and (_24406_, _24395_, _06406_);
  or (_24407_, _24406_, _10059_);
  or (_24408_, _24407_, _24405_);
  and (_24409_, _24408_, _24391_);
  or (_24410_, _24409_, _06281_);
  and (_24412_, _08013_, _09446_);
  or (_24413_, _24385_, _06282_);
  or (_24414_, _24413_, _24412_);
  and (_24415_, _24414_, _24410_);
  or (_24416_, _24415_, _06015_);
  and (_24417_, _14426_, _08013_);
  or (_24418_, _24385_, _06279_);
  or (_24419_, _24418_, _24417_);
  and (_24420_, _24419_, _06276_);
  and (_24421_, _24420_, _24416_);
  and (_24423_, _08013_, _08817_);
  or (_24424_, _24423_, _24385_);
  and (_24425_, _24424_, _06275_);
  or (_24426_, _24425_, _06474_);
  or (_24427_, _24426_, _24421_);
  and (_24428_, _14324_, _08013_);
  or (_24429_, _24428_, _24385_);
  or (_24430_, _24429_, _07282_);
  and (_24431_, _24430_, _07284_);
  and (_24432_, _24431_, _24427_);
  nor (_24434_, _12538_, _12016_);
  or (_24435_, _24434_, _24385_);
  nor (_24436_, _24384_, _07284_);
  and (_24437_, _24436_, _24435_);
  or (_24438_, _24437_, _24432_);
  and (_24439_, _24438_, _07279_);
  nand (_24440_, _24424_, _06478_);
  nor (_24441_, _24440_, _24392_);
  or (_24442_, _24441_, _06569_);
  or (_24443_, _24442_, _24439_);
  and (_24445_, _24443_, _24387_);
  or (_24446_, _24445_, _06479_);
  and (_24447_, _14320_, _08013_);
  or (_24448_, _24385_, _09043_);
  or (_24449_, _24448_, _24447_);
  and (_24450_, _24449_, _09048_);
  and (_24451_, _24450_, _24446_);
  and (_24452_, _24435_, _06572_);
  or (_24453_, _24452_, _19434_);
  or (_24454_, _24453_, _24451_);
  or (_24456_, _24393_, _06700_);
  and (_24457_, _24456_, _01375_);
  and (_24458_, _24457_, _24454_);
  or (_24459_, _24458_, _24382_);
  and (_42968_, _24459_, _42545_);
  and (_24460_, _12016_, \uc8051golden_1.TH0 [1]);
  nor (_24461_, _11223_, _12016_);
  or (_24462_, _24461_, _24460_);
  or (_24463_, _24462_, _09048_);
  and (_24464_, _08013_, _09445_);
  or (_24466_, _24460_, _06282_);
  or (_24467_, _24466_, _24464_);
  or (_24468_, _08013_, \uc8051golden_1.TH0 [1]);
  and (_24469_, _14532_, _08013_);
  not (_24470_, _24469_);
  and (_24471_, _24470_, _24468_);
  or (_24472_, _24471_, _07210_);
  and (_24473_, _08013_, \uc8051golden_1.ACC [1]);
  or (_24474_, _24473_, _24460_);
  and (_24475_, _24474_, _07199_);
  and (_24477_, _07200_, \uc8051golden_1.TH0 [1]);
  or (_24478_, _24477_, _06401_);
  or (_24479_, _24478_, _24475_);
  and (_24480_, _24479_, _07221_);
  and (_24481_, _24480_, _24472_);
  nor (_24482_, _12016_, _07196_);
  or (_24483_, _24482_, _24460_);
  and (_24484_, _24483_, _06399_);
  or (_24485_, _24484_, _24481_);
  and (_24486_, _24485_, _06414_);
  and (_24488_, _24474_, _06406_);
  or (_24489_, _24488_, _10059_);
  or (_24490_, _24489_, _24486_);
  or (_24491_, _24483_, _06293_);
  and (_24492_, _24491_, _24490_);
  or (_24493_, _24492_, _06281_);
  and (_24494_, _24493_, _06279_);
  and (_24495_, _24494_, _24467_);
  or (_24496_, _14615_, _12016_);
  and (_24497_, _24468_, _06015_);
  and (_24499_, _24497_, _24496_);
  or (_24500_, _24499_, _24495_);
  and (_24501_, _24500_, _06276_);
  nand (_24502_, _08013_, _07090_);
  and (_24503_, _24468_, _06275_);
  and (_24504_, _24503_, _24502_);
  or (_24505_, _24504_, _24501_);
  and (_24506_, _24505_, _07282_);
  or (_24507_, _14507_, _12016_);
  and (_24508_, _24468_, _06474_);
  and (_24509_, _24508_, _24507_);
  or (_24510_, _24509_, _06582_);
  or (_24511_, _24510_, _24506_);
  nand (_24512_, _11222_, _08013_);
  and (_24513_, _24512_, _24462_);
  or (_24514_, _24513_, _07284_);
  and (_24515_, _24514_, _07279_);
  and (_24516_, _24515_, _24511_);
  or (_24517_, _14505_, _12016_);
  and (_24518_, _24468_, _06478_);
  and (_24521_, _24518_, _24517_);
  or (_24522_, _24521_, _06569_);
  or (_24523_, _24522_, _24516_);
  nor (_24524_, _24460_, _07276_);
  nand (_24525_, _24524_, _24512_);
  and (_24526_, _24525_, _09043_);
  and (_24527_, _24526_, _24523_);
  or (_24528_, _24502_, _08477_);
  and (_24529_, _24468_, _06479_);
  and (_24530_, _24529_, _24528_);
  or (_24532_, _24530_, _06572_);
  or (_24533_, _24532_, _24527_);
  and (_24534_, _24533_, _24463_);
  or (_24535_, _24534_, _06606_);
  or (_24536_, _24471_, _07037_);
  and (_24537_, _24536_, _06196_);
  and (_24538_, _24537_, _24535_);
  or (_24539_, _24469_, _24460_);
  and (_24540_, _24539_, _06195_);
  or (_24541_, _24540_, _01379_);
  or (_24543_, _24541_, _24538_);
  or (_24544_, _01375_, \uc8051golden_1.TH0 [1]);
  and (_24545_, _24544_, _42545_);
  and (_42969_, _24545_, _24543_);
  and (_24546_, _01379_, \uc8051golden_1.TH0 [2]);
  and (_24547_, _12016_, \uc8051golden_1.TH0 [2]);
  and (_24548_, _14754_, _08013_);
  or (_24549_, _24548_, _24547_);
  or (_24550_, _24549_, _07210_);
  and (_24551_, _08013_, \uc8051golden_1.ACC [2]);
  or (_24553_, _24551_, _24547_);
  and (_24554_, _24553_, _07199_);
  and (_24555_, _07200_, \uc8051golden_1.TH0 [2]);
  or (_24556_, _24555_, _06401_);
  or (_24557_, _24556_, _24554_);
  and (_24558_, _24557_, _07221_);
  and (_24559_, _24558_, _24550_);
  nor (_24560_, _12016_, _07623_);
  or (_24561_, _24560_, _24547_);
  and (_24562_, _24561_, _06399_);
  or (_24564_, _24562_, _24559_);
  and (_24565_, _24564_, _06414_);
  and (_24566_, _24553_, _06406_);
  or (_24567_, _24566_, _10059_);
  or (_24568_, _24567_, _24565_);
  or (_24569_, _24561_, _06293_);
  and (_24570_, _24569_, _24568_);
  or (_24571_, _24570_, _06281_);
  and (_24572_, _08013_, _09444_);
  or (_24573_, _24547_, _06282_);
  or (_24575_, _24573_, _24572_);
  and (_24576_, _24575_, _24571_);
  or (_24577_, _24576_, _06015_);
  and (_24578_, _14848_, _08013_);
  or (_24579_, _24547_, _06279_);
  or (_24580_, _24579_, _24578_);
  and (_24581_, _24580_, _06276_);
  and (_24582_, _24581_, _24577_);
  and (_24583_, _08013_, _08994_);
  or (_24584_, _24583_, _24547_);
  and (_24586_, _24584_, _06275_);
  or (_24587_, _24586_, _06474_);
  or (_24588_, _24587_, _24582_);
  and (_24589_, _14744_, _08013_);
  or (_24590_, _24589_, _24547_);
  or (_24591_, _24590_, _07282_);
  and (_24592_, _24591_, _07284_);
  and (_24593_, _24592_, _24588_);
  and (_24594_, _11221_, _08013_);
  or (_24595_, _24594_, _24547_);
  and (_24597_, _24595_, _06582_);
  or (_24598_, _24597_, _24593_);
  and (_24599_, _24598_, _07279_);
  or (_24600_, _24547_, _08433_);
  and (_24601_, _24584_, _06478_);
  and (_24602_, _24601_, _24600_);
  or (_24603_, _24602_, _24599_);
  and (_24604_, _24603_, _07276_);
  and (_24605_, _24553_, _06569_);
  and (_24606_, _24605_, _24600_);
  or (_24608_, _24606_, _06479_);
  or (_24609_, _24608_, _24604_);
  and (_24610_, _14741_, _08013_);
  or (_24611_, _24547_, _09043_);
  or (_24612_, _24611_, _24610_);
  and (_24613_, _24612_, _09048_);
  and (_24614_, _24613_, _24609_);
  nor (_24615_, _11220_, _12016_);
  or (_24616_, _24615_, _24547_);
  and (_24617_, _24616_, _06572_);
  or (_24619_, _24617_, _24614_);
  and (_24620_, _24619_, _07037_);
  and (_24621_, _24549_, _06606_);
  or (_24622_, _24621_, _06195_);
  or (_24623_, _24622_, _24620_);
  and (_24624_, _14917_, _08013_);
  or (_24625_, _24547_, _06196_);
  or (_24626_, _24625_, _24624_);
  and (_24627_, _24626_, _01375_);
  and (_24628_, _24627_, _24623_);
  or (_24630_, _24628_, _24546_);
  and (_42970_, _24630_, _42545_);
  and (_24631_, _12016_, \uc8051golden_1.TH0 [3]);
  and (_24632_, _14947_, _08013_);
  or (_24633_, _24632_, _24631_);
  or (_24634_, _24633_, _07210_);
  and (_24635_, _08013_, \uc8051golden_1.ACC [3]);
  or (_24636_, _24635_, _24631_);
  and (_24637_, _24636_, _07199_);
  and (_24638_, _07200_, \uc8051golden_1.TH0 [3]);
  or (_24640_, _24638_, _06401_);
  or (_24641_, _24640_, _24637_);
  and (_24642_, _24641_, _07221_);
  and (_24643_, _24642_, _24634_);
  nor (_24644_, _12016_, _07775_);
  or (_24645_, _24644_, _24631_);
  and (_24646_, _24645_, _06399_);
  or (_24647_, _24646_, _24643_);
  and (_24648_, _24647_, _06414_);
  and (_24649_, _24636_, _06406_);
  or (_24651_, _24649_, _10059_);
  or (_24652_, _24651_, _24648_);
  or (_24653_, _24645_, _06293_);
  and (_24654_, _24653_, _24652_);
  or (_24655_, _24654_, _06281_);
  and (_24656_, _08013_, _09443_);
  or (_24657_, _24631_, _06282_);
  or (_24658_, _24657_, _24656_);
  and (_24659_, _24658_, _24655_);
  or (_24660_, _24659_, _06015_);
  and (_24662_, _15039_, _08013_);
  or (_24663_, _24631_, _06279_);
  or (_24664_, _24663_, _24662_);
  and (_24665_, _24664_, _06276_);
  and (_24666_, _24665_, _24660_);
  and (_24667_, _08013_, _08815_);
  or (_24668_, _24667_, _24631_);
  and (_24669_, _24668_, _06275_);
  or (_24670_, _24669_, _06474_);
  or (_24671_, _24670_, _24666_);
  and (_24673_, _14934_, _08013_);
  or (_24674_, _24673_, _24631_);
  or (_24675_, _24674_, _07282_);
  and (_24676_, _24675_, _07284_);
  and (_24677_, _24676_, _24671_);
  and (_24678_, _12535_, _08013_);
  or (_24679_, _24678_, _24631_);
  and (_24680_, _24679_, _06582_);
  or (_24681_, _24680_, _24677_);
  and (_24682_, _24681_, _07279_);
  or (_24684_, _24631_, _08389_);
  and (_24685_, _24668_, _06478_);
  and (_24686_, _24685_, _24684_);
  or (_24687_, _24686_, _24682_);
  and (_24688_, _24687_, _07276_);
  and (_24689_, _24636_, _06569_);
  and (_24690_, _24689_, _24684_);
  or (_24691_, _24690_, _06479_);
  or (_24692_, _24691_, _24688_);
  and (_24693_, _14931_, _08013_);
  or (_24695_, _24631_, _09043_);
  or (_24696_, _24695_, _24693_);
  and (_24697_, _24696_, _09048_);
  and (_24698_, _24697_, _24692_);
  nor (_24699_, _11218_, _12016_);
  or (_24700_, _24699_, _24631_);
  and (_24701_, _24700_, _06572_);
  or (_24702_, _24701_, _06606_);
  or (_24703_, _24702_, _24698_);
  or (_24704_, _24633_, _07037_);
  and (_24706_, _24704_, _06196_);
  and (_24707_, _24706_, _24703_);
  and (_24708_, _15113_, _08013_);
  or (_24709_, _24708_, _24631_);
  and (_24710_, _24709_, _06195_);
  or (_24711_, _24710_, _01379_);
  or (_24712_, _24711_, _24707_);
  or (_24713_, _01375_, \uc8051golden_1.TH0 [3]);
  and (_24714_, _24713_, _42545_);
  and (_42971_, _24714_, _24712_);
  and (_24716_, _12016_, \uc8051golden_1.TH0 [4]);
  and (_24717_, _15130_, _08013_);
  or (_24718_, _24717_, _24716_);
  or (_24719_, _24718_, _07210_);
  and (_24720_, _08013_, \uc8051golden_1.ACC [4]);
  or (_24721_, _24720_, _24716_);
  and (_24722_, _24721_, _07199_);
  and (_24723_, _07200_, \uc8051golden_1.TH0 [4]);
  or (_24724_, _24723_, _06401_);
  or (_24725_, _24724_, _24722_);
  and (_24727_, _24725_, _07221_);
  and (_24728_, _24727_, _24719_);
  nor (_24729_, _12016_, _08301_);
  or (_24730_, _24729_, _24716_);
  and (_24731_, _24730_, _06399_);
  or (_24732_, _24731_, _24728_);
  and (_24733_, _24732_, _06414_);
  and (_24734_, _24721_, _06406_);
  or (_24735_, _24734_, _10059_);
  or (_24736_, _24735_, _24733_);
  or (_24738_, _24730_, _06293_);
  and (_24739_, _24738_, _24736_);
  or (_24740_, _24739_, _06281_);
  and (_24741_, _08013_, _09442_);
  or (_24742_, _24716_, _06282_);
  or (_24743_, _24742_, _24741_);
  and (_24744_, _24743_, _06279_);
  and (_24745_, _24744_, _24740_);
  and (_24746_, _15243_, _08013_);
  or (_24747_, _24746_, _24716_);
  and (_24749_, _24747_, _06015_);
  or (_24750_, _24749_, _06275_);
  or (_24751_, _24750_, _24745_);
  and (_24752_, _08883_, _08013_);
  or (_24753_, _24752_, _24716_);
  or (_24754_, _24753_, _06276_);
  and (_24755_, _24754_, _24751_);
  or (_24756_, _24755_, _06474_);
  and (_24757_, _15135_, _08013_);
  or (_24758_, _24757_, _24716_);
  or (_24760_, _24758_, _07282_);
  and (_24761_, _24760_, _07284_);
  and (_24762_, _24761_, _24756_);
  and (_24763_, _11216_, _08013_);
  or (_24764_, _24763_, _24716_);
  and (_24765_, _24764_, _06582_);
  or (_24766_, _24765_, _24762_);
  and (_24767_, _24766_, _07279_);
  or (_24768_, _24716_, _08345_);
  and (_24769_, _24753_, _06478_);
  and (_24771_, _24769_, _24768_);
  or (_24772_, _24771_, _24767_);
  and (_24773_, _24772_, _07276_);
  and (_24774_, _24721_, _06569_);
  and (_24775_, _24774_, _24768_);
  or (_24776_, _24775_, _06479_);
  or (_24777_, _24776_, _24773_);
  and (_24778_, _15134_, _08013_);
  or (_24779_, _24716_, _09043_);
  or (_24780_, _24779_, _24778_);
  and (_24782_, _24780_, _09048_);
  and (_24783_, _24782_, _24777_);
  nor (_24784_, _11215_, _12016_);
  or (_24785_, _24784_, _24716_);
  and (_24786_, _24785_, _06572_);
  or (_24787_, _24786_, _06606_);
  or (_24788_, _24787_, _24783_);
  or (_24789_, _24718_, _07037_);
  and (_24790_, _24789_, _06196_);
  and (_24791_, _24790_, _24788_);
  and (_24793_, _15315_, _08013_);
  or (_24794_, _24793_, _24716_);
  and (_24795_, _24794_, _06195_);
  or (_24796_, _24795_, _01379_);
  or (_24797_, _24796_, _24791_);
  or (_24798_, _01375_, \uc8051golden_1.TH0 [4]);
  and (_24799_, _24798_, _42545_);
  and (_42972_, _24799_, _24797_);
  and (_24800_, _12016_, \uc8051golden_1.TH0 [5]);
  nor (_24801_, _12016_, _08207_);
  or (_24803_, _24801_, _24800_);
  or (_24804_, _24803_, _06293_);
  and (_24805_, _15348_, _08013_);
  or (_24806_, _24805_, _24800_);
  or (_24807_, _24806_, _07210_);
  and (_24808_, _08013_, \uc8051golden_1.ACC [5]);
  or (_24809_, _24808_, _24800_);
  and (_24810_, _24809_, _07199_);
  and (_24811_, _07200_, \uc8051golden_1.TH0 [5]);
  or (_24812_, _24811_, _06401_);
  or (_24814_, _24812_, _24810_);
  and (_24815_, _24814_, _07221_);
  and (_24816_, _24815_, _24807_);
  and (_24817_, _24803_, _06399_);
  or (_24818_, _24817_, _24816_);
  and (_24819_, _24818_, _06414_);
  and (_24820_, _24809_, _06406_);
  or (_24821_, _24820_, _10059_);
  or (_24822_, _24821_, _24819_);
  and (_24823_, _24822_, _24804_);
  or (_24825_, _24823_, _06281_);
  and (_24826_, _08013_, _09441_);
  or (_24827_, _24800_, _06282_);
  or (_24828_, _24827_, _24826_);
  and (_24829_, _24828_, _06279_);
  and (_24830_, _24829_, _24825_);
  and (_24831_, _15446_, _08013_);
  or (_24832_, _24831_, _24800_);
  and (_24833_, _24832_, _06015_);
  or (_24834_, _24833_, _06275_);
  or (_24836_, _24834_, _24830_);
  and (_24837_, _08958_, _08013_);
  or (_24838_, _24837_, _24800_);
  or (_24839_, _24838_, _06276_);
  and (_24840_, _24839_, _24836_);
  or (_24841_, _24840_, _06474_);
  and (_24842_, _15338_, _08013_);
  or (_24843_, _24842_, _24800_);
  or (_24844_, _24843_, _07282_);
  and (_24845_, _24844_, _07284_);
  and (_24847_, _24845_, _24841_);
  and (_24848_, _12542_, _08013_);
  or (_24849_, _24848_, _24800_);
  and (_24850_, _24849_, _06582_);
  or (_24851_, _24850_, _24847_);
  and (_24852_, _24851_, _07279_);
  or (_24853_, _24800_, _08256_);
  and (_24854_, _24838_, _06478_);
  and (_24855_, _24854_, _24853_);
  or (_24856_, _24855_, _24852_);
  and (_24858_, _24856_, _07276_);
  and (_24859_, _24809_, _06569_);
  and (_24860_, _24859_, _24853_);
  or (_24861_, _24860_, _06479_);
  or (_24862_, _24861_, _24858_);
  and (_24863_, _15335_, _08013_);
  or (_24864_, _24800_, _09043_);
  or (_24865_, _24864_, _24863_);
  and (_24866_, _24865_, _09048_);
  and (_24867_, _24866_, _24862_);
  nor (_24869_, _11212_, _12016_);
  or (_24870_, _24869_, _24800_);
  and (_24871_, _24870_, _06572_);
  or (_24872_, _24871_, _06606_);
  or (_24873_, _24872_, _24867_);
  or (_24874_, _24806_, _07037_);
  and (_24875_, _24874_, _06196_);
  and (_24876_, _24875_, _24873_);
  and (_24877_, _15509_, _08013_);
  or (_24878_, _24877_, _24800_);
  and (_24880_, _24878_, _06195_);
  or (_24881_, _24880_, _01379_);
  or (_24882_, _24881_, _24876_);
  or (_24883_, _01375_, \uc8051golden_1.TH0 [5]);
  and (_24884_, _24883_, _42545_);
  and (_42974_, _24884_, _24882_);
  and (_24885_, _12016_, \uc8051golden_1.TH0 [6]);
  and (_24886_, _15550_, _08013_);
  or (_24887_, _24886_, _24885_);
  or (_24888_, _24887_, _07210_);
  and (_24890_, _08013_, \uc8051golden_1.ACC [6]);
  or (_24891_, _24890_, _24885_);
  and (_24892_, _24891_, _07199_);
  and (_24893_, _07200_, \uc8051golden_1.TH0 [6]);
  or (_24894_, _24893_, _06401_);
  or (_24895_, _24894_, _24892_);
  and (_24896_, _24895_, _07221_);
  and (_24897_, _24896_, _24888_);
  nor (_24898_, _12016_, _08118_);
  or (_24899_, _24898_, _24885_);
  and (_24901_, _24899_, _06399_);
  or (_24902_, _24901_, _24897_);
  and (_24903_, _24902_, _06414_);
  and (_24904_, _24891_, _06406_);
  or (_24905_, _24904_, _10059_);
  or (_24906_, _24905_, _24903_);
  or (_24907_, _24899_, _06293_);
  and (_24908_, _24907_, _24906_);
  or (_24909_, _24908_, _06281_);
  and (_24910_, _08013_, _09440_);
  or (_24912_, _24885_, _06282_);
  or (_24913_, _24912_, _24910_);
  and (_24914_, _24913_, _06279_);
  and (_24915_, _24914_, _24909_);
  and (_24916_, _15639_, _08013_);
  or (_24917_, _24916_, _24885_);
  and (_24918_, _24917_, _06015_);
  or (_24919_, _24918_, _06275_);
  or (_24920_, _24919_, _24915_);
  and (_24921_, _15646_, _08013_);
  or (_24923_, _24921_, _24885_);
  or (_24924_, _24923_, _06276_);
  and (_24925_, _24924_, _24920_);
  or (_24926_, _24925_, _06474_);
  and (_24927_, _15531_, _08013_);
  or (_24928_, _24927_, _24885_);
  or (_24929_, _24928_, _07282_);
  and (_24930_, _24929_, _07284_);
  and (_24931_, _24930_, _24926_);
  and (_24932_, _11210_, _08013_);
  or (_24934_, _24932_, _24885_);
  and (_24935_, _24934_, _06582_);
  or (_24936_, _24935_, _24931_);
  and (_24937_, _24936_, _07279_);
  or (_24938_, _24885_, _08162_);
  and (_24939_, _24923_, _06478_);
  and (_24940_, _24939_, _24938_);
  or (_24941_, _24940_, _24937_);
  and (_24942_, _24941_, _07276_);
  and (_24943_, _24891_, _06569_);
  and (_24945_, _24943_, _24938_);
  or (_24946_, _24945_, _06479_);
  or (_24947_, _24946_, _24942_);
  and (_24948_, _15528_, _08013_);
  or (_24949_, _24885_, _09043_);
  or (_24950_, _24949_, _24948_);
  and (_24951_, _24950_, _09048_);
  and (_24952_, _24951_, _24947_);
  nor (_24953_, _11209_, _12016_);
  or (_24954_, _24953_, _24885_);
  and (_24956_, _24954_, _06572_);
  or (_24957_, _24956_, _06606_);
  or (_24958_, _24957_, _24952_);
  or (_24959_, _24887_, _07037_);
  and (_24960_, _24959_, _06196_);
  and (_24961_, _24960_, _24958_);
  and (_24962_, _15713_, _08013_);
  or (_24963_, _24962_, _24885_);
  and (_24964_, _24963_, _06195_);
  or (_24965_, _24964_, _01379_);
  or (_24967_, _24965_, _24961_);
  or (_24968_, _01375_, \uc8051golden_1.TH0 [6]);
  and (_24969_, _24968_, _42545_);
  and (_42975_, _24969_, _24967_);
  and (_24970_, _13030_, _05685_);
  nor (_24971_, _06475_, _05963_);
  not (_24972_, _24971_);
  and (_24973_, _24972_, _06943_);
  and (_24974_, _12958_, \uc8051golden_1.PC [0]);
  and (_24975_, _06943_, \uc8051golden_1.PC [0]);
  nor (_24977_, _24975_, _12317_);
  nor (_24978_, _24977_, _12958_);
  nor (_24979_, _24978_, _24974_);
  and (_24980_, _24979_, _06234_);
  and (_24981_, _12987_, _12994_);
  nor (_24982_, _24981_, _05685_);
  and (_24983_, _12108_, _12968_);
  nor (_24984_, _24983_, _05685_);
  and (_24985_, _10881_, \uc8051golden_1.PC [0]);
  nor (_24986_, _10881_, \uc8051golden_1.PC [0]);
  nor (_24988_, _24986_, _24985_);
  and (_24989_, _24988_, _12217_);
  nor (_24990_, _12224_, _06479_);
  nor (_24991_, _24990_, _05685_);
  not (_24992_, _05956_);
  and (_24993_, _12719_, _07279_);
  nor (_24994_, _24993_, _05685_);
  not (_24995_, _05952_);
  and (_24996_, _12233_, _07282_);
  nor (_24997_, _24996_, _05685_);
  and (_24999_, _06275_, _05685_);
  nor (_25000_, _06943_, _06007_);
  and (_25001_, _12546_, _05685_);
  not (_25002_, _24977_);
  nor (_25003_, _25002_, _12546_);
  nor (_25004_, _25003_, _25001_);
  nor (_25005_, _25004_, _06842_);
  and (_25006_, _12405_, _05685_);
  and (_25007_, _24977_, _12407_);
  or (_25008_, _25007_, _12411_);
  nor (_25010_, _25008_, _25006_);
  nor (_25011_, _06943_, _06000_);
  and (_25012_, _12517_, _12509_);
  nor (_25013_, _25012_, _05685_);
  and (_25014_, _06943_, _06790_);
  and (_25015_, _12481_, \uc8051golden_1.PC [0]);
  nor (_25016_, _12492_, _05685_);
  and (_25017_, _12492_, _05685_);
  nor (_25018_, _25017_, _25016_);
  nor (_25019_, _12481_, _06790_);
  not (_25021_, _25019_);
  nor (_25022_, _25021_, _25018_);
  nor (_25023_, _25022_, _25015_);
  not (_25024_, _25023_);
  nor (_25025_, _25024_, _25014_);
  nor (_25026_, _25025_, _08643_);
  and (_25027_, _12476_, \uc8051golden_1.PC [0]);
  and (_25028_, _06840_, _05685_);
  nor (_25029_, _25028_, _12163_);
  and (_25030_, _25029_, _12474_);
  or (_25032_, _25030_, _25027_);
  nor (_25033_, _25032_, _08644_);
  nor (_25034_, _25033_, _25026_);
  nor (_25035_, _25034_, _07212_);
  and (_25036_, _07212_, \uc8051golden_1.PC [0]);
  nor (_25037_, _25036_, _06401_);
  not (_25038_, _25037_);
  nor (_25039_, _25038_, _25035_);
  not (_25040_, _25039_);
  not (_25041_, _12458_);
  and (_25043_, _25002_, _12464_);
  and (_25044_, _12466_, \uc8051golden_1.PC [0]);
  or (_25045_, _25044_, _07210_);
  nor (_25046_, _25045_, _25043_);
  nor (_25047_, _25046_, _25041_);
  and (_25048_, _25047_, _25040_);
  nor (_25049_, _12458_, _05685_);
  nor (_25050_, _25049_, _07351_);
  not (_25051_, _25050_);
  nor (_25052_, _25051_, _25048_);
  nor (_25053_, _06943_, _05997_);
  not (_25054_, _25012_);
  nor (_25055_, _25054_, _25053_);
  not (_25056_, _25055_);
  nor (_25057_, _25056_, _25052_);
  or (_25058_, _25057_, _12521_);
  nor (_25059_, _25058_, _25013_);
  nor (_25060_, _25059_, _25011_);
  or (_25061_, _25060_, _12450_);
  and (_25062_, _12444_, \uc8051golden_1.PC [0]);
  nor (_25065_, _24977_, _12444_);
  or (_25066_, _25065_, _12449_);
  or (_25067_, _25066_, _25062_);
  and (_25068_, _25067_, _12411_);
  and (_25069_, _25068_, _25061_);
  nor (_25070_, _25069_, _06420_);
  not (_25071_, _25070_);
  nor (_25072_, _25071_, _25010_);
  nor (_25073_, _25072_, _25005_);
  nor (_25074_, _25073_, _06482_);
  and (_25076_, _12249_, _05685_);
  nor (_25077_, _25002_, _12249_);
  or (_25078_, _25077_, _25076_);
  and (_25079_, _25078_, _06482_);
  or (_25080_, _25079_, _25074_);
  and (_25081_, _25080_, _12238_);
  and (_25082_, _12237_, _05685_);
  or (_25083_, _25082_, _25081_);
  and (_25084_, _25083_, _05994_);
  nor (_25085_, _06943_, _05994_);
  nor (_25087_, _25085_, _12580_);
  not (_25088_, _25087_);
  nor (_25089_, _25088_, _25084_);
  not (_25090_, _06007_);
  nor (_25091_, _12576_, _05685_);
  nor (_25092_, _25091_, _25090_);
  not (_25093_, _25092_);
  nor (_25094_, _25093_, _25089_);
  and (_25095_, _12588_, _06023_);
  not (_25096_, _25095_);
  or (_25098_, _25096_, _25094_);
  nor (_25099_, _25098_, _25000_);
  nor (_25100_, _25095_, _05685_);
  nor (_25101_, _25100_, _06017_);
  not (_25102_, _25101_);
  nor (_25103_, _25102_, _25099_);
  nor (_25104_, _06943_, _07846_);
  nor (_25105_, _06472_, _06015_);
  and (_25106_, _25105_, _12616_);
  not (_25107_, _25106_);
  nor (_25109_, _25107_, _25104_);
  not (_25110_, _25109_);
  nor (_25111_, _25110_, _25103_);
  nor (_25112_, _25106_, _05685_);
  nor (_25113_, _25112_, _05936_);
  not (_25114_, _25113_);
  nor (_25115_, _25114_, _25111_);
  not (_25116_, _05936_);
  nor (_25117_, _06943_, _25116_);
  or (_25118_, _25117_, _12624_);
  nor (_25120_, _25118_, _25115_);
  nor (_25121_, _25029_, _12625_);
  nor (_25122_, _25121_, _25120_);
  and (_25123_, _25122_, _06276_);
  or (_25124_, _25123_, _24999_);
  and (_25125_, _25124_, _12640_);
  and (_25126_, _12639_, _06053_);
  or (_25127_, _25126_, _25125_);
  and (_25128_, _25127_, _13854_);
  nor (_25129_, _06943_, _13854_);
  or (_25131_, _25129_, _25128_);
  and (_25132_, _25131_, _12681_);
  not (_25133_, _24996_);
  nor (_25134_, _25029_, _11297_);
  and (_25135_, _11297_, _05685_);
  nor (_25136_, _25135_, _12681_);
  not (_25137_, _25136_);
  nor (_25138_, _25137_, _25134_);
  nor (_25139_, _25138_, _25133_);
  not (_25140_, _25139_);
  nor (_25142_, _25140_, _25132_);
  nor (_25143_, _25142_, _24997_);
  and (_25144_, _25143_, _24995_);
  nor (_25145_, _06943_, _24995_);
  or (_25146_, _25145_, _25144_);
  and (_25147_, _25146_, _12705_);
  not (_25148_, _24993_);
  nor (_25149_, _11297_, _05685_);
  and (_25150_, _25029_, _11297_);
  or (_25151_, _25150_, _25149_);
  and (_25153_, _25151_, _12704_);
  nor (_25154_, _25153_, _25148_);
  not (_25155_, _25154_);
  nor (_25156_, _25155_, _25147_);
  nor (_25157_, _25156_, _24994_);
  and (_25158_, _25157_, _24992_);
  nor (_25159_, _06943_, _24992_);
  or (_25160_, _25159_, _25158_);
  and (_25161_, _25160_, _12736_);
  not (_25162_, _24990_);
  and (_25164_, \uc8051golden_1.PSW [7], \uc8051golden_1.PC [0]);
  and (_25165_, _25029_, _10524_);
  or (_25166_, _25165_, _25164_);
  and (_25167_, _25166_, _12735_);
  nor (_25168_, _25167_, _25162_);
  not (_25169_, _25168_);
  nor (_25170_, _25169_, _25161_);
  nor (_25171_, _25170_, _24991_);
  and (_25172_, _25171_, _05948_);
  nor (_25173_, _06943_, _05948_);
  or (_25175_, _25173_, _25172_);
  and (_25176_, _25175_, _12756_);
  and (_25177_, _12761_, _11090_);
  not (_25178_, _25177_);
  or (_25179_, _25178_, _25176_);
  nor (_25180_, _25179_, _24989_);
  nor (_25181_, _25177_, _05685_);
  nor (_25182_, _25181_, _06588_);
  not (_25183_, _25182_);
  nor (_25184_, _25183_, _25180_);
  and (_25186_, _09446_, _06588_);
  or (_25187_, _25186_, _25184_);
  and (_25188_, _25187_, _05967_);
  nor (_25189_, _06943_, _05967_);
  or (_25190_, _25189_, _25188_);
  and (_25191_, _25190_, _06596_);
  and (_25192_, _25002_, _12958_);
  nor (_25193_, _12958_, _05685_);
  or (_25194_, _25193_, _06596_);
  or (_25195_, _25194_, _25192_);
  and (_25197_, _25195_, _24983_);
  not (_25198_, _25197_);
  nor (_25199_, _25198_, _25191_);
  nor (_25200_, _25199_, _24984_);
  and (_25201_, _25200_, _06306_);
  and (_25202_, _09446_, _06305_);
  or (_25203_, _25202_, _25201_);
  and (_25204_, _25203_, _12979_);
  nor (_25205_, _06943_, _12979_);
  nor (_25206_, _25205_, _25204_);
  nor (_25208_, _25206_, _06487_);
  not (_25209_, _24981_);
  and (_25210_, _24979_, _06487_);
  nor (_25211_, _25210_, _25209_);
  not (_25212_, _25211_);
  nor (_25213_, _25212_, _25208_);
  nor (_25214_, _25213_, _24982_);
  nor (_25215_, _25214_, _07887_);
  and (_25216_, _07887_, _06943_);
  nor (_25217_, _25216_, _06234_);
  not (_25219_, _25217_);
  nor (_25220_, _25219_, _25215_);
  nor (_25221_, _25220_, _24980_);
  and (_25222_, _13019_, _13011_);
  not (_25223_, _25222_);
  nor (_25224_, _25223_, _25221_);
  nor (_25225_, _25222_, \uc8051golden_1.PC [0]);
  nor (_25226_, _25225_, _24972_);
  not (_25227_, _25226_);
  nor (_25228_, _25227_, _25224_);
  or (_25230_, _25228_, _13030_);
  nor (_25231_, _25230_, _24973_);
  nor (_25232_, _25231_, _24970_);
  nand (_25233_, _25232_, _01375_);
  or (_25234_, _01375_, \uc8051golden_1.PC [0]);
  and (_25235_, _25234_, _42545_);
  and (_42976_, _25235_, _25233_);
  nor (_25236_, _13019_, _06024_);
  nor (_25237_, _12994_, _06024_);
  nand (_25238_, _07694_, _06011_);
  and (_25240_, _25238_, _09061_);
  nor (_25241_, _25240_, _06024_);
  nor (_25242_, _12108_, _06024_);
  nor (_25243_, _06291_, _06988_);
  and (_25244_, _25243_, _05985_);
  nor (_25245_, _12721_, _05653_);
  nor (_25246_, _12715_, _06024_);
  nor (_25247_, _12233_, _06024_);
  nor (_25248_, _09012_, _05653_);
  nand (_25249_, _12444_, _05985_);
  nor (_25251_, _12319_, _12317_);
  or (_25252_, _25251_, _12320_);
  or (_25253_, _25252_, _12444_);
  and (_25254_, _25253_, _25249_);
  and (_25255_, _25254_, _12450_);
  nor (_25256_, _12165_, _12163_);
  or (_25257_, _25256_, _12166_);
  or (_25258_, _25257_, _12476_);
  or (_25259_, _12474_, \uc8051golden_1.PC [1]);
  and (_25260_, _25259_, _25258_);
  and (_25262_, _25260_, _08643_);
  and (_25263_, _07090_, _06790_);
  and (_25264_, _12481_, _05985_);
  and (_25265_, _07332_, \uc8051golden_1.PC [0]);
  and (_25266_, _06854_, _05685_);
  nor (_25267_, _25266_, _12484_);
  nor (_25268_, _25267_, _25265_);
  nor (_25269_, _25268_, _05653_);
  and (_25270_, _25268_, _05653_);
  or (_25271_, _25270_, _25269_);
  and (_25273_, _25271_, _25019_);
  or (_25274_, _25273_, _25264_);
  or (_25275_, _25274_, _25263_);
  and (_25276_, _25275_, _08644_);
  or (_25277_, _25276_, _07212_);
  or (_25278_, _25277_, _25262_);
  nand (_25279_, _07212_, _06024_);
  and (_25280_, _25279_, _07210_);
  and (_25281_, _25280_, _25278_);
  or (_25282_, _25252_, _12466_);
  or (_25284_, _12464_, _06024_);
  and (_25285_, _25284_, _06401_);
  and (_25286_, _25285_, _25282_);
  or (_25287_, _25286_, _25281_);
  and (_25288_, _25287_, _12458_);
  nor (_25289_, _12458_, _06024_);
  or (_25290_, _25289_, _06395_);
  or (_25291_, _25290_, _25288_);
  nand (_25292_, _06395_, _05653_);
  and (_25293_, _25292_, _05997_);
  and (_25295_, _25293_, _25291_);
  and (_25296_, _07090_, _07351_);
  or (_25297_, _25296_, _06399_);
  or (_25298_, _25297_, _25295_);
  nand (_25299_, _06399_, _05653_);
  and (_25300_, _25299_, _12509_);
  and (_25301_, _25300_, _25298_);
  nor (_25302_, _12509_, _06024_);
  or (_25303_, _25302_, _06406_);
  or (_25304_, _25303_, _25301_);
  nand (_25306_, _06406_, _05653_);
  and (_25307_, _25306_, _12517_);
  and (_25308_, _25307_, _25304_);
  nor (_25309_, _12517_, _06024_);
  or (_25310_, _25309_, _06393_);
  or (_25311_, _25310_, _25308_);
  nand (_25312_, _06393_, _05653_);
  and (_25313_, _25312_, _06000_);
  and (_25314_, _25313_, _25311_);
  and (_25315_, _07090_, _12521_);
  or (_25316_, _25315_, _06419_);
  or (_25317_, _25316_, _25314_);
  nand (_25318_, _06419_, _05653_);
  and (_25319_, _25318_, _12449_);
  and (_25320_, _25319_, _25317_);
  or (_25321_, _25320_, _25255_);
  and (_25322_, _25321_, _12411_);
  or (_25323_, _12407_, _06024_);
  or (_25324_, _25252_, _12405_);
  and (_25325_, _25324_, _25323_);
  and (_25328_, _25325_, _06457_);
  or (_25329_, _25328_, _06420_);
  or (_25330_, _25329_, _25322_);
  or (_25331_, _25252_, _12546_);
  nand (_25332_, _12546_, _05985_);
  and (_25333_, _25332_, _25331_);
  or (_25334_, _25333_, _06842_);
  and (_25335_, _25334_, _25330_);
  or (_25336_, _25335_, _06482_);
  nand (_25337_, _12249_, _05985_);
  or (_25339_, _25252_, _12249_);
  and (_25340_, _25339_, _25337_);
  or (_25341_, _25340_, _12534_);
  and (_25342_, _25341_, _12238_);
  and (_25343_, _25342_, _25336_);
  nand (_25344_, _12237_, _05985_);
  nand (_25345_, _25344_, _12557_);
  or (_25346_, _25345_, _25343_);
  or (_25347_, _07090_, _05994_);
  nand (_25348_, _06387_, _05653_);
  and (_25350_, _25348_, _12569_);
  and (_25351_, _25350_, _25347_);
  and (_25352_, _25351_, _25346_);
  nor (_25353_, _12569_, _05653_);
  or (_25354_, _25353_, _12573_);
  or (_25355_, _25354_, _25352_);
  nand (_25356_, _12573_, _06024_);
  and (_25357_, _25356_, _12575_);
  and (_25358_, _25357_, _25355_);
  nor (_25359_, _12575_, _06024_);
  or (_25361_, _25359_, _06433_);
  or (_25362_, _25361_, _25358_);
  nand (_25363_, _06433_, _05653_);
  and (_25364_, _25363_, _06007_);
  and (_25365_, _25364_, _25362_);
  and (_25366_, _07090_, _25090_);
  or (_25367_, _25366_, _06432_);
  or (_25368_, _25367_, _25365_);
  not (_25369_, _10738_);
  or (_25370_, _25369_, _11002_);
  and (_25372_, _25370_, _06016_);
  and (_25373_, _06452_, _06016_);
  nor (_25374_, _12586_, _25373_);
  nand (_25375_, _06432_, _05653_);
  nand (_25376_, _25375_, _25374_);
  nor (_25377_, _25376_, _25372_);
  and (_25378_, _25377_, _25368_);
  nor (_25379_, _12588_, _06024_);
  or (_25380_, _25379_, _25378_);
  and (_25381_, _25380_, _12592_);
  nor (_25383_, _12592_, _05653_);
  or (_25384_, _25383_, _06022_);
  or (_25385_, _25384_, _25381_);
  nand (_25386_, _06022_, _06024_);
  and (_25387_, _25386_, _06446_);
  and (_25388_, _25387_, _25385_);
  and (_25389_, _06300_, \uc8051golden_1.PC [1]);
  or (_25390_, _25389_, _25388_);
  and (_25391_, _25390_, _07846_);
  and (_25392_, _07090_, _06017_);
  or (_25394_, _25392_, _06472_);
  or (_25395_, _25394_, _25391_);
  nand (_25396_, _06472_, _05985_);
  and (_25397_, _25396_, _06294_);
  and (_25398_, _25397_, _25395_);
  nor (_25399_, _06294_, _05653_);
  or (_25400_, _25399_, _06015_);
  or (_25401_, _25400_, _25398_);
  nand (_25402_, _06015_, _05985_);
  and (_25403_, _25402_, _12616_);
  and (_25405_, _25403_, _25401_);
  nor (_25406_, _12616_, _06024_);
  or (_25407_, _25406_, _06376_);
  or (_25408_, _25407_, _25405_);
  nand (_25409_, _06376_, _05653_);
  and (_25410_, _25409_, _25116_);
  and (_25411_, _25410_, _25408_);
  and (_25412_, _07090_, _05936_);
  or (_25413_, _25412_, _12624_);
  or (_25414_, _25413_, _25411_);
  or (_25416_, _25257_, _12625_);
  and (_25417_, _25416_, _09012_);
  and (_25418_, _25417_, _25414_);
  or (_25419_, _25418_, _25248_);
  and (_25420_, _25419_, _06276_);
  and (_25421_, _06275_, _06024_);
  or (_25422_, _25421_, _10933_);
  or (_25423_, _25422_, _25420_);
  nand (_25424_, _10933_, _05653_);
  and (_25425_, _25424_, _12640_);
  and (_25427_, _25425_, _25423_);
  nor (_25428_, _12640_, _06034_);
  or (_25429_, _25428_, _06375_);
  or (_25430_, _25429_, _25427_);
  nand (_25431_, _06375_, _05653_);
  and (_25432_, _25431_, _13854_);
  and (_25433_, _25432_, _25430_);
  and (_25434_, _07090_, _05943_);
  or (_25435_, _25434_, _12680_);
  or (_25436_, _25435_, _25433_);
  and (_25438_, _25257_, _12687_);
  nand (_25439_, _11297_, \uc8051golden_1.PC [1]);
  nand (_25440_, _25439_, _12680_);
  or (_25441_, _25440_, _25438_);
  and (_25442_, _25441_, _12233_);
  and (_25443_, _25442_, _25436_);
  or (_25444_, _25443_, _25247_);
  and (_25445_, _25444_, _12227_);
  nor (_25446_, _12227_, _05653_);
  or (_25447_, _25446_, _06474_);
  or (_25449_, _25447_, _25445_);
  nand (_25450_, _06474_, _05985_);
  and (_25451_, _25450_, _07284_);
  and (_25452_, _25451_, _25449_);
  and (_25453_, _06582_, \uc8051golden_1.PC [1]);
  or (_25454_, _25453_, _25452_);
  and (_25455_, _25454_, _24995_);
  and (_25456_, _07090_, _05952_);
  or (_25457_, _25456_, _12704_);
  or (_25458_, _25457_, _25455_);
  and (_25460_, _25257_, _11297_);
  or (_25461_, _11297_, _05653_);
  nand (_25462_, _25461_, _12704_);
  or (_25463_, _25462_, _25460_);
  and (_25464_, _25463_, _12715_);
  and (_25465_, _25464_, _25458_);
  or (_25466_, _25465_, _25246_);
  nand (_25467_, _10559_, _05979_);
  and (_25468_, _25467_, _12717_);
  and (_25469_, _25468_, _25466_);
  nor (_25471_, _25468_, _06024_);
  or (_25472_, _25471_, _06969_);
  or (_25473_, _25472_, _25469_);
  nand (_25474_, _06969_, _06024_);
  and (_25475_, _25474_, _12721_);
  and (_25476_, _25475_, _25473_);
  or (_25477_, _25476_, _25245_);
  and (_25478_, _25477_, _07279_);
  and (_25479_, _06478_, _06024_);
  or (_25480_, _25479_, _06569_);
  or (_25482_, _25480_, _25478_);
  nand (_25483_, _06569_, _05653_);
  and (_25484_, _25483_, _24992_);
  and (_25485_, _25484_, _25482_);
  and (_25486_, _07090_, _05956_);
  or (_25487_, _25486_, _12735_);
  or (_25488_, _25487_, _25485_);
  and (_25489_, _25257_, _10524_);
  nand (_25490_, \uc8051golden_1.PSW [7], \uc8051golden_1.PC [1]);
  nand (_25491_, _25490_, _12735_);
  or (_25493_, _25491_, _25489_);
  and (_25494_, _25493_, _12225_);
  and (_25495_, _25494_, _25488_);
  and (_25496_, _12224_, _05985_);
  or (_25497_, _25496_, _25495_);
  and (_25498_, _25497_, _11018_);
  nor (_25499_, _11018_, _05653_);
  or (_25500_, _25499_, _06479_);
  or (_25501_, _25500_, _25498_);
  nand (_25502_, _06479_, _05985_);
  and (_25504_, _25502_, _09048_);
  and (_25505_, _25504_, _25501_);
  and (_25506_, _06572_, \uc8051golden_1.PC [1]);
  or (_25507_, _25506_, _25505_);
  and (_25508_, _25507_, _05948_);
  and (_25509_, _07090_, _05947_);
  or (_25510_, _25509_, _12217_);
  or (_25511_, _25510_, _25508_);
  and (_25512_, _25257_, \uc8051golden_1.PSW [7]);
  or (_25513_, \uc8051golden_1.PSW [7], _05653_);
  nand (_25515_, _25513_, _12217_);
  nor (_25516_, _25515_, _25512_);
  nor (_25517_, _25516_, _25243_);
  and (_25518_, _25517_, _25511_);
  or (_25519_, _25518_, _25244_);
  and (_25520_, _06285_, _05965_);
  nor (_25521_, _17463_, _25520_);
  and (_25522_, _25521_, _25519_);
  nor (_25523_, _25521_, _06024_);
  or (_25524_, _25523_, _06984_);
  or (_25526_, _25524_, _25522_);
  nand (_25527_, _06984_, _06024_);
  and (_25528_, _25527_, _11060_);
  and (_25529_, _25528_, _25526_);
  nor (_25530_, _11060_, _05653_);
  or (_25531_, _25530_, _11089_);
  or (_25532_, _25531_, _25529_);
  nand (_25533_, _11089_, _06024_);
  and (_25534_, _25533_, _13881_);
  and (_25535_, _25534_, _25532_);
  and (_25537_, _09345_, _06588_);
  or (_25538_, _25537_, _25535_);
  and (_25539_, _25538_, _05967_);
  and (_25540_, _07090_, _05966_);
  or (_25541_, _25540_, _06460_);
  or (_25542_, _25541_, _25539_);
  and (_25543_, _25252_, _12958_);
  nor (_25544_, _12958_, _05985_);
  or (_25545_, _25544_, _06596_);
  or (_25546_, _25545_, _25543_);
  and (_25548_, _25546_, _12108_);
  and (_25549_, _25548_, _25542_);
  or (_25550_, _25549_, _25242_);
  and (_25551_, _25550_, _11204_);
  nor (_25552_, _11204_, _05653_);
  or (_25553_, _25552_, _11243_);
  or (_25554_, _25553_, _25551_);
  nand (_25555_, _11243_, _06024_);
  and (_25556_, _25555_, _06306_);
  and (_25557_, _25556_, _25554_);
  and (_25559_, _09345_, _06305_);
  or (_25560_, _25559_, _25557_);
  and (_25561_, _25560_, _12979_);
  and (_25562_, _07090_, _05971_);
  or (_25563_, _25562_, _06487_);
  or (_25564_, _25563_, _25561_);
  nand (_25565_, _12958_, _05985_);
  or (_25566_, _25252_, _12958_);
  and (_25567_, _25566_, _25565_);
  or (_25568_, _25567_, _12978_);
  and (_25570_, _25568_, _25240_);
  and (_25571_, _25570_, _25564_);
  or (_25572_, _25571_, _25241_);
  nor (_25573_, _07305_, _09066_);
  and (_25574_, _25573_, _25572_);
  nor (_25575_, _25573_, _06024_);
  or (_25576_, _25575_, _06606_);
  or (_25577_, _25576_, _25574_);
  nand (_25578_, _06606_, _05653_);
  and (_25579_, _25578_, _12994_);
  and (_25581_, _25579_, _25577_);
  or (_25582_, _25581_, _25237_);
  and (_25583_, _25582_, _07312_);
  and (_25584_, _07887_, _07090_);
  or (_25585_, _25584_, _06234_);
  or (_25586_, _25585_, _25583_);
  or (_25587_, _25567_, _06807_);
  and (_25588_, _25587_, _14683_);
  and (_25589_, _25588_, _25586_);
  nor (_25590_, _14683_, _06024_);
  or (_25592_, _25590_, _25589_);
  nor (_25593_, _07320_, _07048_);
  and (_25594_, _25593_, _25592_);
  nor (_25595_, _25593_, _06024_);
  or (_25596_, _25595_, _06195_);
  or (_25597_, _25596_, _25594_);
  nand (_25598_, _06195_, _05653_);
  and (_25599_, _25598_, _13019_);
  and (_25600_, _25599_, _25597_);
  or (_25601_, _25600_, _25236_);
  nand (_25603_, _25601_, _24971_);
  and (_25604_, _24972_, _07090_);
  nor (_25605_, _25604_, _13030_);
  and (_25606_, _25605_, _25603_);
  and (_25607_, _13030_, _06024_);
  or (_25608_, _25607_, _25606_);
  or (_25609_, _25608_, _01379_);
  or (_25610_, _01375_, \uc8051golden_1.PC [1]);
  and (_25611_, _25610_, _42545_);
  and (_42977_, _25611_, _25609_);
  and (_25613_, _13030_, _06071_);
  and (_25614_, _06195_, _06065_);
  and (_25615_, _06606_, _06065_);
  nor (_25616_, _12108_, _06071_);
  nor (_25617_, _12761_, _06071_);
  not (_25618_, _06071_);
  and (_25619_, _12224_, _25618_);
  nor (_25620_, _12719_, _06071_);
  nor (_25621_, _12233_, _06071_);
  nor (_25622_, _12569_, _06065_);
  and (_25623_, _12237_, _25618_);
  and (_25624_, _12324_, _12321_);
  nor (_25625_, _25624_, _12325_);
  not (_25626_, _25625_);
  or (_25627_, _25626_, _12405_);
  or (_25628_, _12407_, _12314_);
  nand (_25629_, _25628_, _25627_);
  nand (_25630_, _25629_, _06457_);
  or (_25631_, _25625_, _12466_);
  or (_25632_, _12464_, _12313_);
  and (_25635_, _25632_, _25631_);
  or (_25636_, _25635_, _07210_);
  and (_25637_, _12476_, _06065_);
  and (_25638_, _12170_, _12167_);
  nor (_25639_, _25638_, _12171_);
  and (_25640_, _25639_, _12474_);
  nor (_25641_, _25640_, _25637_);
  nand (_25642_, _25641_, _08643_);
  or (_25643_, _07366_, _06736_);
  and (_25644_, _07199_, _06500_);
  or (_25646_, _25644_, _06854_);
  or (_25647_, _07332_, _05663_);
  and (_25648_, _25647_, _07200_);
  or (_25649_, _25648_, _25646_);
  or (_25650_, _12492_, _25618_);
  and (_25651_, _25650_, _12491_);
  and (_25652_, _25651_, _25649_);
  or (_25653_, _25652_, _06790_);
  and (_25654_, _25653_, _25643_);
  and (_25655_, _12481_, _25618_);
  or (_25657_, _25655_, _25654_);
  and (_25658_, _25657_, _08644_);
  nor (_25659_, _25658_, _07212_);
  and (_25660_, _25659_, _25642_);
  and (_25661_, _07212_, _06071_);
  or (_25662_, _25661_, _06401_);
  or (_25663_, _25662_, _25660_);
  nand (_25664_, _25663_, _25636_);
  nand (_25665_, _25664_, _12458_);
  nor (_25666_, _12458_, _06071_);
  nor (_25668_, _25666_, _06395_);
  nand (_25669_, _25668_, _25665_);
  and (_25670_, _06395_, _06065_);
  nor (_25671_, _25670_, _07351_);
  nand (_25672_, _25671_, _25669_);
  and (_25673_, _06736_, _07351_);
  nor (_25674_, _25673_, _06399_);
  nand (_25675_, _25674_, _25672_);
  and (_25676_, _06399_, _06065_);
  nor (_25677_, _25676_, _12510_);
  nand (_25679_, _25677_, _25675_);
  nor (_25680_, _12509_, _06071_);
  nor (_25681_, _25680_, _06406_);
  nand (_25682_, _25681_, _25679_);
  and (_25683_, _06406_, _06065_);
  nor (_25684_, _25683_, _12519_);
  nand (_25685_, _25684_, _25682_);
  nor (_25686_, _12517_, _06071_);
  nor (_25687_, _25686_, _06393_);
  nand (_25688_, _25687_, _25685_);
  and (_25690_, _06393_, _06065_);
  nor (_25691_, _25690_, _12521_);
  nand (_25692_, _25691_, _25688_);
  and (_25693_, _06736_, _12521_);
  nor (_25694_, _25693_, _06419_);
  nand (_25695_, _25694_, _25692_);
  and (_25696_, _06419_, _06065_);
  nor (_25697_, _25696_, _12450_);
  nand (_25698_, _25697_, _25695_);
  and (_25699_, _12444_, _12313_);
  nor (_25701_, _25626_, _12444_);
  or (_25702_, _25701_, _12449_);
  nor (_25703_, _25702_, _25699_);
  nor (_25704_, _25703_, _06457_);
  nand (_25705_, _25704_, _25698_);
  and (_25706_, _25705_, _25630_);
  or (_25707_, _25706_, _06420_);
  nor (_25708_, _25626_, _12546_);
  and (_25709_, _12546_, _12313_);
  nor (_25710_, _25709_, _25708_);
  or (_25712_, _25710_, _06842_);
  and (_25713_, _25712_, _25707_);
  or (_25714_, _25713_, _06482_);
  and (_25715_, _12314_, _12249_);
  nor (_25716_, _25625_, _12249_);
  or (_25717_, _25716_, _12534_);
  or (_25718_, _25717_, _25715_);
  and (_25719_, _25718_, _12238_);
  and (_25720_, _25719_, _25714_);
  or (_25721_, _25720_, _25623_);
  nand (_25723_, _25721_, _07245_);
  and (_25724_, _06387_, _06500_);
  nor (_25725_, _25724_, _07349_);
  nand (_25726_, _25725_, _25723_);
  not (_25727_, _12569_);
  nor (_25728_, _06736_, _05994_);
  nor (_25729_, _25728_, _25727_);
  and (_25730_, _25729_, _25726_);
  or (_25731_, _25730_, _25622_);
  nand (_25732_, _25731_, _12576_);
  nor (_25734_, _12576_, _06071_);
  nor (_25735_, _25734_, _06433_);
  nand (_25736_, _25735_, _25732_);
  and (_25737_, _06433_, _06065_);
  nor (_25738_, _25737_, _25090_);
  nand (_25739_, _25738_, _25736_);
  and (_25740_, _06736_, _25090_);
  nor (_25741_, _25740_, _06432_);
  nand (_25742_, _25741_, _25739_);
  and (_25743_, _06432_, _06065_);
  nor (_25745_, _25743_, _12594_);
  and (_25746_, _25745_, _25742_);
  nor (_25747_, _12588_, _06071_);
  or (_25748_, _25747_, _25746_);
  nand (_25749_, _25748_, _12592_);
  nor (_25750_, _12592_, _06065_);
  nor (_25751_, _25750_, _06022_);
  nand (_25752_, _25751_, _25749_);
  and (_25753_, _06071_, _06022_);
  nor (_25754_, _25753_, _06300_);
  and (_25756_, _25754_, _25752_);
  and (_25757_, _06300_, _06500_);
  or (_25758_, _25757_, _25756_);
  nand (_25759_, _25758_, _07846_);
  and (_25760_, _06736_, _06017_);
  nor (_25761_, _25760_, _06472_);
  nand (_25762_, _25761_, _25759_);
  and (_25763_, _06849_, _05935_);
  not (_25764_, _25763_);
  and (_25765_, _07343_, _05935_);
  nor (_25767_, _25765_, _06286_);
  and (_25768_, _25767_, _25764_);
  and (_25769_, _12313_, _06472_);
  nor (_25770_, _25769_, _06292_);
  and (_25771_, _25770_, _25768_);
  nand (_25772_, _25771_, _25762_);
  nor (_25773_, _06294_, _06065_);
  nor (_25774_, _25773_, _06015_);
  nand (_25775_, _25774_, _25772_);
  and (_25776_, _12313_, _06015_);
  nor (_25778_, _25776_, _12620_);
  nand (_25779_, _25778_, _25775_);
  nor (_25780_, _12616_, _06071_);
  nor (_25781_, _25780_, _06376_);
  and (_25782_, _25781_, _25779_);
  and (_25783_, _06376_, _06065_);
  or (_25784_, _25783_, _05936_);
  nor (_25785_, _25784_, _25782_);
  and (_25786_, _06736_, _05936_);
  or (_25787_, _25786_, _25785_);
  nand (_25789_, _25787_, _12625_);
  nor (_25790_, _25639_, _12625_);
  nor (_25791_, _25790_, _09011_);
  and (_25792_, _25791_, _25789_);
  nor (_25793_, _07268_, _06065_);
  nor (_25794_, _25793_, _09012_);
  or (_25795_, _25794_, _25792_);
  and (_25796_, _07268_, _06500_);
  nor (_25797_, _25796_, _06275_);
  nand (_25798_, _25797_, _25795_);
  and (_25800_, _12313_, _06275_);
  nor (_25801_, _25800_, _10933_);
  and (_25802_, _25801_, _25798_);
  and (_25803_, _10933_, _06500_);
  or (_25804_, _25803_, _25802_);
  nand (_25805_, _25804_, _12640_);
  nor (_25806_, _12640_, _06088_);
  nor (_25807_, _25806_, _06375_);
  nand (_25808_, _25807_, _25805_);
  and (_25809_, _06375_, _06065_);
  nor (_25811_, _25809_, _05943_);
  nand (_25812_, _25811_, _25808_);
  and (_25813_, _06736_, _05943_);
  nor (_25814_, _25813_, _12680_);
  nand (_25815_, _25814_, _25812_);
  nor (_25816_, _25639_, _11297_);
  and (_25817_, _11297_, _06500_);
  nor (_25818_, _25817_, _12681_);
  not (_25819_, _25818_);
  nor (_25820_, _25819_, _25816_);
  nor (_25822_, _25820_, _12685_);
  and (_25823_, _25822_, _25815_);
  or (_25824_, _25823_, _25621_);
  nand (_25825_, _25824_, _12227_);
  nor (_25826_, _12227_, _06065_);
  nor (_25827_, _25826_, _06474_);
  nand (_25828_, _25827_, _25825_);
  and (_25829_, _12313_, _06474_);
  nor (_25830_, _25829_, _06582_);
  and (_25831_, _25830_, _25828_);
  and (_25833_, _06582_, _06500_);
  or (_25834_, _25833_, _25831_);
  nand (_25835_, _25834_, _24995_);
  and (_25836_, _06736_, _05952_);
  nor (_25837_, _25836_, _12704_);
  nand (_25838_, _25837_, _25835_);
  nor (_25839_, _11297_, _06500_);
  and (_25840_, _25639_, _11297_);
  or (_25841_, _25840_, _25839_);
  and (_25842_, _25841_, _12704_);
  nor (_25844_, _25842_, _12723_);
  and (_25845_, _25844_, _25838_);
  or (_25846_, _25845_, _25620_);
  nand (_25847_, _25846_, _12721_);
  nor (_25848_, _12721_, _06065_);
  nor (_25849_, _25848_, _06478_);
  nand (_25850_, _25849_, _25847_);
  and (_25851_, _12313_, _06478_);
  nor (_25852_, _25851_, _06569_);
  and (_25853_, _25852_, _25850_);
  and (_25855_, _06569_, _06500_);
  or (_25856_, _25855_, _25853_);
  nand (_25857_, _25856_, _24992_);
  and (_25858_, _06736_, _05956_);
  nor (_25859_, _25858_, _12735_);
  nand (_25860_, _25859_, _25857_);
  nor (_25861_, _25639_, \uc8051golden_1.PSW [7]);
  nor (_25862_, _06065_, _10524_);
  nor (_25863_, _25862_, _12736_);
  not (_25864_, _25863_);
  nor (_25866_, _25864_, _25861_);
  nor (_25867_, _25866_, _12224_);
  and (_25868_, _25867_, _25860_);
  or (_25869_, _25868_, _25619_);
  nand (_25870_, _25869_, _11018_);
  nor (_25871_, _11018_, _06065_);
  nor (_25872_, _25871_, _06479_);
  nand (_25873_, _25872_, _25870_);
  and (_25874_, _12313_, _06479_);
  nor (_25875_, _25874_, _06572_);
  and (_25877_, _25875_, _25873_);
  and (_25878_, _06572_, _06500_);
  or (_25879_, _25878_, _25877_);
  nand (_25880_, _25879_, _05948_);
  and (_25881_, _06736_, _05947_);
  nor (_25882_, _25881_, _12217_);
  nand (_25883_, _25882_, _25880_);
  nor (_25884_, _25639_, _10524_);
  nor (_25885_, _06065_, \uc8051golden_1.PSW [7]);
  nor (_25886_, _25885_, _12756_);
  not (_25888_, _25886_);
  nor (_25889_, _25888_, _25884_);
  nor (_25890_, _25889_, _12763_);
  and (_25891_, _25890_, _25883_);
  or (_25892_, _25891_, _25617_);
  nand (_25893_, _25892_, _11060_);
  nor (_25894_, _11060_, _06065_);
  nor (_25895_, _25894_, _11089_);
  nand (_25896_, _25895_, _25893_);
  and (_25897_, _11089_, _06071_);
  nor (_25899_, _25897_, _06588_);
  and (_25900_, _25899_, _25896_);
  and (_25901_, _09300_, _06588_);
  or (_25902_, _25901_, _25900_);
  nand (_25903_, _25902_, _05967_);
  and (_25904_, _06736_, _05966_);
  nor (_25905_, _25904_, _06460_);
  nand (_25906_, _25905_, _25903_);
  nor (_25907_, _12313_, _12958_);
  and (_25908_, _25626_, _12958_);
  or (_25910_, _25908_, _06596_);
  nor (_25911_, _25910_, _25907_);
  nor (_25912_, _25911_, _12779_);
  and (_25913_, _25912_, _25906_);
  or (_25914_, _25913_, _25616_);
  nand (_25915_, _25914_, _11204_);
  nor (_25916_, _11204_, _06065_);
  nor (_25917_, _25916_, _11243_);
  nand (_25918_, _25917_, _25915_);
  and (_25919_, _11243_, _06071_);
  nor (_25921_, _25919_, _06305_);
  and (_25922_, _25921_, _25918_);
  and (_25923_, _09300_, _06305_);
  or (_25924_, _25923_, _25922_);
  nand (_25925_, _25924_, _12979_);
  and (_25926_, _06736_, _05971_);
  nor (_25927_, _25926_, _06487_);
  nand (_25928_, _25927_, _25925_);
  nor (_25929_, _25625_, _12958_);
  and (_25930_, _12314_, _12958_);
  nor (_25932_, _25930_, _25929_);
  and (_25933_, _25932_, _06487_);
  nor (_25934_, _25933_, _12988_);
  nand (_25935_, _25934_, _25928_);
  nor (_25936_, _12987_, _06071_);
  nor (_25937_, _25936_, _06606_);
  and (_25938_, _25937_, _25935_);
  or (_25939_, _25938_, _25615_);
  nand (_25940_, _25939_, _12994_);
  nor (_25941_, _12994_, _25618_);
  nor (_25943_, _25941_, _07887_);
  nand (_25944_, _25943_, _25940_);
  and (_25945_, _07887_, _06736_);
  nor (_25946_, _25945_, _06234_);
  nand (_25947_, _25946_, _25944_);
  and (_25948_, _25932_, _06234_);
  nor (_25949_, _25948_, _13012_);
  nand (_25950_, _25949_, _25947_);
  nor (_25951_, _13011_, _06071_);
  nor (_25952_, _25951_, _06195_);
  and (_25953_, _25952_, _25950_);
  or (_25954_, _25953_, _25614_);
  nand (_25955_, _25954_, _13019_);
  nor (_25956_, _13019_, _25618_);
  nor (_25957_, _25956_, _24972_);
  nand (_25958_, _25957_, _25955_);
  and (_25959_, _24972_, _06736_);
  nor (_25960_, _25959_, _13030_);
  and (_25961_, _25960_, _25958_);
  or (_25962_, _25961_, _25613_);
  or (_25965_, _25962_, _01379_);
  or (_25966_, _01375_, \uc8051golden_1.PC [2]);
  and (_25967_, _25966_, _42545_);
  and (_42978_, _25967_, _25965_);
  and (_25968_, _06195_, _06124_);
  nor (_25969_, _12994_, _06120_);
  nor (_25970_, _12108_, _06120_);
  nor (_25971_, _12761_, _06120_);
  and (_25972_, _12224_, _06102_);
  nor (_25973_, _12719_, _06120_);
  nor (_25975_, _12233_, _06120_);
  nor (_25976_, _09012_, _06124_);
  nor (_25977_, _12569_, _06124_);
  and (_25978_, _12237_, _06102_);
  or (_25979_, _12311_, _12310_);
  and (_25980_, _25979_, _12326_);
  nor (_25981_, _25979_, _12326_);
  nor (_25982_, _25981_, _25980_);
  not (_25983_, _25982_);
  or (_25984_, _25983_, _12405_);
  or (_25986_, _12407_, _12309_);
  nand (_25987_, _25986_, _25984_);
  nand (_25988_, _25987_, _06457_);
  or (_25989_, _12464_, _12308_);
  or (_25990_, _25982_, _12466_);
  and (_25991_, _25990_, _25989_);
  or (_25992_, _25991_, _07210_);
  and (_25993_, _12476_, _06124_);
  or (_25994_, _12160_, _12159_);
  and (_25995_, _25994_, _12172_);
  nor (_25997_, _25994_, _12172_);
  nor (_25998_, _25997_, _25995_);
  and (_25999_, _25998_, _12474_);
  nor (_26000_, _25999_, _25993_);
  nand (_26001_, _26000_, _08643_);
  or (_26002_, _07366_, _06562_);
  and (_26003_, _07199_, _06134_);
  or (_26004_, _26003_, _06854_);
  or (_26005_, _07332_, _05655_);
  and (_26006_, _26005_, _07200_);
  or (_26008_, _26006_, _26004_);
  or (_26009_, _12492_, _06102_);
  and (_26010_, _26009_, _12491_);
  and (_26011_, _26010_, _26008_);
  or (_26012_, _26011_, _06790_);
  and (_26013_, _26012_, _26002_);
  and (_26014_, _12481_, _06102_);
  or (_26015_, _26014_, _26013_);
  and (_26016_, _26015_, _08644_);
  nor (_26017_, _26016_, _07212_);
  and (_26019_, _26017_, _26001_);
  and (_26020_, _07212_, _06120_);
  or (_26021_, _26020_, _06401_);
  or (_26022_, _26021_, _26019_);
  nand (_26023_, _26022_, _25992_);
  nand (_26024_, _26023_, _12458_);
  nor (_26025_, _12458_, _06120_);
  nor (_26026_, _26025_, _06395_);
  nand (_26027_, _26026_, _26024_);
  and (_26028_, _06395_, _06124_);
  nor (_26030_, _26028_, _07351_);
  nand (_26031_, _26030_, _26027_);
  and (_26032_, _06562_, _07351_);
  nor (_26033_, _26032_, _06399_);
  nand (_26034_, _26033_, _26031_);
  and (_26035_, _06399_, _06124_);
  nor (_26036_, _26035_, _12510_);
  nand (_26037_, _26036_, _26034_);
  nor (_26038_, _12509_, _06120_);
  nor (_26039_, _26038_, _06406_);
  nand (_26041_, _26039_, _26037_);
  and (_26042_, _06406_, _06124_);
  nor (_26043_, _26042_, _12519_);
  nand (_26044_, _26043_, _26041_);
  nor (_26045_, _12517_, _06120_);
  nor (_26046_, _26045_, _06393_);
  nand (_26047_, _26046_, _26044_);
  and (_26048_, _06393_, _06124_);
  nor (_26049_, _26048_, _12521_);
  nand (_26050_, _26049_, _26047_);
  and (_26052_, _06562_, _12521_);
  nor (_26053_, _26052_, _06419_);
  nand (_26054_, _26053_, _26050_);
  and (_26055_, _06419_, _06124_);
  nor (_26056_, _26055_, _12450_);
  nand (_26057_, _26056_, _26054_);
  and (_26058_, _12444_, _12308_);
  nor (_26059_, _25983_, _12444_);
  or (_26060_, _26059_, _26058_);
  nor (_26061_, _26060_, _12449_);
  nor (_26063_, _26061_, _06457_);
  nand (_26064_, _26063_, _26057_);
  and (_26065_, _26064_, _06842_);
  nand (_26066_, _26065_, _25988_);
  nor (_26067_, _25983_, _12546_);
  not (_26068_, _26067_);
  and (_26069_, _12546_, _12308_);
  nor (_26070_, _26069_, _06842_);
  and (_26071_, _26070_, _26068_);
  nor (_26072_, _26071_, _06482_);
  nand (_26074_, _26072_, _26066_);
  nor (_26075_, _25982_, _12249_);
  and (_26076_, _12309_, _12249_);
  or (_26077_, _26076_, _12534_);
  nor (_26078_, _26077_, _26075_);
  nor (_26079_, _26078_, _12237_);
  and (_26080_, _26079_, _26074_);
  or (_26081_, _26080_, _25978_);
  nand (_26082_, _26081_, _07245_);
  and (_26083_, _06387_, _06134_);
  nor (_26085_, _26083_, _07349_);
  nand (_26086_, _26085_, _26082_);
  nor (_26087_, _06562_, _05994_);
  nor (_26088_, _26087_, _25727_);
  and (_26089_, _26088_, _26086_);
  or (_26090_, _26089_, _25977_);
  nand (_26091_, _26090_, _12576_);
  nor (_26092_, _12576_, _06120_);
  nor (_26093_, _26092_, _06433_);
  nand (_26094_, _26093_, _26091_);
  and (_26096_, _06433_, _06124_);
  nor (_26097_, _26096_, _25090_);
  nand (_26098_, _26097_, _26094_);
  and (_26099_, _06562_, _25090_);
  nor (_26100_, _26099_, _06432_);
  nand (_26101_, _26100_, _26098_);
  and (_26102_, _06432_, _06124_);
  nor (_26103_, _26102_, _12594_);
  and (_26104_, _26103_, _26101_);
  nor (_26105_, _12588_, _06120_);
  or (_26107_, _26105_, _26104_);
  nand (_26108_, _26107_, _12592_);
  nor (_26109_, _12592_, _06124_);
  nor (_26110_, _26109_, _06022_);
  nand (_26111_, _26110_, _26108_);
  and (_26112_, _06022_, _06120_);
  nor (_26113_, _26112_, _06300_);
  and (_26114_, _26113_, _26111_);
  and (_26115_, _06300_, _06134_);
  or (_26116_, _26115_, _26114_);
  nand (_26118_, _26116_, _07846_);
  and (_26119_, _06562_, _06017_);
  nor (_26120_, _26119_, _06472_);
  nand (_26121_, _26120_, _26118_);
  and (_26122_, _12308_, _06472_);
  nor (_26123_, _26122_, _13788_);
  nand (_26124_, _26123_, _26121_);
  nor (_26125_, _06294_, _06124_);
  nor (_26126_, _26125_, _06015_);
  nand (_26127_, _26126_, _26124_);
  and (_26129_, _12308_, _06015_);
  nor (_26130_, _26129_, _12620_);
  nand (_26131_, _26130_, _26127_);
  nor (_26132_, _12616_, _06120_);
  nor (_26133_, _26132_, _06376_);
  nand (_26134_, _26133_, _26131_);
  and (_26135_, _06376_, _06124_);
  nor (_26136_, _26135_, _05936_);
  nand (_26137_, _26136_, _26134_);
  and (_26138_, _06562_, _05936_);
  nor (_26140_, _26138_, _12624_);
  nand (_26141_, _26140_, _26137_);
  and (_26142_, _25998_, _12624_);
  nor (_26143_, _26142_, _09013_);
  and (_26144_, _26143_, _26141_);
  or (_26145_, _26144_, _25976_);
  nand (_26146_, _26145_, _06276_);
  and (_26147_, _12309_, _06275_);
  nor (_26148_, _26147_, _10933_);
  nand (_26149_, _26148_, _26146_);
  and (_26151_, _10933_, _06124_);
  nor (_26152_, _26151_, _12639_);
  nand (_26153_, _26152_, _26149_);
  nor (_26154_, _12640_, _06117_);
  nor (_26155_, _26154_, _06375_);
  nand (_26156_, _26155_, _26153_);
  and (_26157_, _06375_, _06124_);
  nor (_26158_, _26157_, _05943_);
  nand (_26159_, _26158_, _26156_);
  and (_26160_, _06562_, _05943_);
  nor (_26162_, _26160_, _12680_);
  nand (_26163_, _26162_, _26159_);
  and (_26164_, _11297_, _06124_);
  and (_26165_, _25998_, _12687_);
  or (_26166_, _26165_, _26164_);
  and (_26167_, _26166_, _12680_);
  nor (_26168_, _26167_, _12685_);
  and (_26169_, _26168_, _26163_);
  or (_26170_, _26169_, _25975_);
  nand (_26171_, _26170_, _12227_);
  nor (_26173_, _12227_, _06124_);
  nor (_26174_, _26173_, _06474_);
  nand (_26175_, _26174_, _26171_);
  and (_26176_, _12308_, _06474_);
  nor (_26177_, _26176_, _06582_);
  and (_26178_, _26177_, _26175_);
  and (_26179_, _06582_, _06134_);
  or (_26180_, _26179_, _26178_);
  nand (_26181_, _26180_, _24995_);
  and (_26182_, _06562_, _05952_);
  nor (_26184_, _26182_, _12704_);
  nand (_26185_, _26184_, _26181_);
  nor (_26186_, _11297_, _06134_);
  and (_26187_, _25998_, _11297_);
  or (_26188_, _26187_, _26186_);
  and (_26189_, _26188_, _12704_);
  nor (_26190_, _26189_, _12723_);
  and (_26191_, _26190_, _26185_);
  or (_26192_, _26191_, _25973_);
  nand (_26193_, _26192_, _12721_);
  nor (_26195_, _12721_, _06124_);
  nor (_26196_, _26195_, _06478_);
  nand (_26197_, _26196_, _26193_);
  and (_26198_, _12308_, _06478_);
  nor (_26199_, _26198_, _06569_);
  and (_26200_, _26199_, _26197_);
  and (_26201_, _06569_, _06134_);
  or (_26202_, _26201_, _26200_);
  nand (_26203_, _26202_, _24992_);
  and (_26204_, _06562_, _05956_);
  nor (_26206_, _26204_, _12735_);
  nand (_26207_, _26206_, _26203_);
  nor (_26208_, _25998_, \uc8051golden_1.PSW [7]);
  nor (_26209_, _06124_, _10524_);
  nor (_26210_, _26209_, _12736_);
  not (_26211_, _26210_);
  nor (_26212_, _26211_, _26208_);
  nor (_26213_, _26212_, _12224_);
  and (_26214_, _26213_, _26207_);
  or (_26215_, _26214_, _25972_);
  nand (_26217_, _26215_, _11018_);
  nor (_26218_, _11018_, _06124_);
  nor (_26219_, _26218_, _06479_);
  and (_26220_, _26219_, _26217_);
  and (_26221_, _12308_, _06479_);
  or (_26222_, _26221_, _06572_);
  nor (_26223_, _26222_, _26220_);
  and (_26224_, _06572_, _06134_);
  or (_26225_, _26224_, _26223_);
  nand (_26226_, _26225_, _05948_);
  and (_26228_, _06562_, _05947_);
  nor (_26229_, _26228_, _12217_);
  nand (_26230_, _26229_, _26226_);
  and (_26231_, _06124_, _10524_);
  and (_26232_, _25998_, \uc8051golden_1.PSW [7]);
  or (_26233_, _26232_, _26231_);
  and (_26234_, _26233_, _12217_);
  nor (_26235_, _26234_, _12763_);
  and (_26236_, _26235_, _26230_);
  or (_26237_, _26236_, _25971_);
  nand (_26239_, _26237_, _11060_);
  nor (_26240_, _11060_, _06124_);
  nor (_26241_, _26240_, _11089_);
  nand (_26242_, _26241_, _26239_);
  and (_26243_, _11089_, _06120_);
  nor (_26244_, _26243_, _06588_);
  and (_26245_, _26244_, _26242_);
  and (_26246_, _09255_, _06588_);
  or (_26247_, _26246_, _26245_);
  nand (_26248_, _26247_, _05967_);
  and (_26250_, _06562_, _05966_);
  nor (_26251_, _26250_, _06460_);
  nand (_26252_, _26251_, _26248_);
  and (_26253_, _25983_, _12958_);
  nor (_26254_, _12308_, _12958_);
  or (_26255_, _26254_, _06596_);
  or (_26256_, _26255_, _26253_);
  and (_26257_, _26256_, _12108_);
  and (_26258_, _26257_, _26252_);
  or (_26259_, _26258_, _25970_);
  nand (_26261_, _26259_, _11204_);
  nor (_26262_, _11204_, _06124_);
  nor (_26263_, _26262_, _11243_);
  nand (_26264_, _26263_, _26261_);
  and (_26265_, _11243_, _06120_);
  nor (_26266_, _26265_, _06305_);
  and (_26267_, _26266_, _26264_);
  and (_26268_, _09255_, _06305_);
  or (_26269_, _26268_, _26267_);
  nand (_26270_, _26269_, _12979_);
  and (_26272_, _06562_, _05971_);
  nor (_26273_, _26272_, _06487_);
  nand (_26274_, _26273_, _26270_);
  nor (_26275_, _25982_, _12958_);
  and (_26276_, _12309_, _12958_);
  nor (_26277_, _26276_, _26275_);
  and (_26278_, _26277_, _06487_);
  nor (_26279_, _26278_, _12988_);
  nand (_26280_, _26279_, _26274_);
  nor (_26281_, _12987_, _06120_);
  nor (_26283_, _26281_, _06606_);
  nand (_26284_, _26283_, _26280_);
  and (_26285_, _06606_, _06124_);
  nor (_26286_, _26285_, _12995_);
  and (_26287_, _26286_, _26284_);
  or (_26288_, _26287_, _25969_);
  nand (_26289_, _26288_, _07312_);
  and (_26290_, _07887_, _06562_);
  nor (_26291_, _26290_, _06234_);
  nand (_26292_, _26291_, _26289_);
  and (_26294_, _26277_, _06234_);
  nor (_26295_, _26294_, _13012_);
  nand (_26296_, _26295_, _26292_);
  nor (_26297_, _13011_, _06120_);
  nor (_26298_, _26297_, _06195_);
  and (_26299_, _26298_, _26296_);
  or (_26300_, _26299_, _25968_);
  nand (_26301_, _26300_, _13019_);
  nor (_26302_, _13019_, _06102_);
  nor (_26303_, _26302_, _24972_);
  nand (_26305_, _26303_, _26301_);
  and (_26306_, _24972_, _06562_);
  nor (_26307_, _26306_, _13030_);
  and (_26308_, _26307_, _26305_);
  and (_26309_, _13030_, _06120_);
  or (_26310_, _26309_, _26308_);
  or (_26311_, _26310_, _01379_);
  or (_26312_, _01375_, \uc8051golden_1.PC [3]);
  and (_26313_, _26312_, _42545_);
  and (_42980_, _26313_, _26311_);
  not (_26315_, \uc8051golden_1.PC [4]);
  nor (_26316_, _05672_, _26315_);
  and (_26317_, _05672_, _26315_);
  nor (_26318_, _26317_, _26316_);
  and (_26319_, _26318_, _13030_);
  nor (_26320_, _26318_, _13011_);
  nor (_26321_, _12157_, _11297_);
  and (_26322_, _12177_, _12174_);
  nor (_26323_, _26322_, _12178_);
  and (_26324_, _26323_, _11297_);
  or (_26326_, _26324_, _26321_);
  and (_26327_, _26326_, _12704_);
  nor (_26328_, _12156_, _09012_);
  nor (_26329_, _12569_, _12156_);
  not (_26330_, _26318_);
  and (_26331_, _26330_, _12237_);
  and (_26332_, _12546_, _12304_);
  and (_26333_, _12331_, _12328_);
  nor (_26334_, _26333_, _12332_);
  not (_26335_, _26334_);
  nor (_26337_, _26335_, _12546_);
  nor (_26338_, _26337_, _26332_);
  or (_26339_, _26338_, _06842_);
  and (_26340_, _12405_, _12304_);
  and (_26341_, _26334_, _12407_);
  nor (_26342_, _26341_, _26340_);
  nand (_26343_, _26342_, _06457_);
  and (_26344_, _26334_, _12464_);
  and (_26345_, _12466_, _12304_);
  or (_26346_, _26345_, _26344_);
  and (_26348_, _26346_, _06401_);
  or (_26349_, _26323_, _12476_);
  or (_26350_, _12474_, _12156_);
  nand (_26351_, _26350_, _26349_);
  nand (_26352_, _26351_, _08643_);
  and (_26353_, _08882_, _06790_);
  and (_26354_, _12157_, _07199_);
  nor (_26355_, _26354_, _06854_);
  nor (_26356_, _07332_, _26315_);
  or (_26357_, _26356_, _07199_);
  and (_26359_, _26357_, _26355_);
  nor (_26360_, _26330_, _12492_);
  or (_26361_, _26360_, _06790_);
  nor (_26362_, _26361_, _26359_);
  nor (_26363_, _26362_, _12481_);
  not (_26364_, _26363_);
  nor (_26365_, _26364_, _26353_);
  and (_26366_, _26318_, _12481_);
  nor (_26367_, _26366_, _08643_);
  not (_26368_, _26367_);
  nor (_26370_, _26368_, _26365_);
  not (_26371_, _26370_);
  and (_26372_, _26371_, _12497_);
  and (_26373_, _26372_, _26352_);
  or (_26374_, _26373_, _26348_);
  and (_26375_, _26374_, _12458_);
  nor (_26376_, _26330_, _12503_);
  or (_26377_, _26376_, _06395_);
  or (_26378_, _26377_, _26375_);
  and (_26379_, _12157_, _06395_);
  nor (_26381_, _26379_, _07351_);
  nand (_26382_, _26381_, _26378_);
  nor (_26383_, _08882_, _05997_);
  nor (_26384_, _26383_, _06399_);
  nand (_26385_, _26384_, _26382_);
  and (_26386_, _12157_, _06399_);
  nor (_26387_, _26386_, _12510_);
  nand (_26388_, _26387_, _26385_);
  nor (_26389_, _26330_, _12509_);
  nor (_26390_, _26389_, _06406_);
  nand (_26392_, _26390_, _26388_);
  and (_26393_, _12157_, _06406_);
  nor (_26394_, _26393_, _12519_);
  nand (_26395_, _26394_, _26392_);
  nor (_26396_, _26330_, _12517_);
  nor (_26397_, _26396_, _06393_);
  and (_26398_, _26397_, _26395_);
  and (_26399_, _12157_, _06393_);
  or (_26400_, _26399_, _26398_);
  nand (_26401_, _26400_, _06000_);
  and (_26403_, _08882_, _12521_);
  nor (_26404_, _26403_, _06419_);
  nand (_26405_, _26404_, _26401_);
  and (_26406_, _12156_, _06419_);
  nor (_26407_, _26406_, _12450_);
  and (_26408_, _26407_, _26405_);
  and (_26409_, _12444_, _12304_);
  nor (_26410_, _26335_, _12444_);
  or (_26411_, _26410_, _26409_);
  nor (_26412_, _26411_, _12449_);
  or (_26414_, _26412_, _26408_);
  nand (_26415_, _26414_, _12411_);
  nand (_26416_, _26415_, _26343_);
  or (_26417_, _26416_, _06420_);
  and (_26418_, _26417_, _26339_);
  or (_26419_, _26418_, _06482_);
  and (_26420_, _12304_, _12249_);
  not (_26421_, _12249_);
  and (_26422_, _26334_, _26421_);
  or (_26423_, _26422_, _26420_);
  and (_26425_, _26423_, _06482_);
  nor (_26426_, _26425_, _12237_);
  and (_26427_, _26426_, _26419_);
  or (_26428_, _26427_, _26331_);
  nand (_26429_, _26428_, _07245_);
  and (_26430_, _12157_, _06387_);
  nor (_26431_, _26430_, _07349_);
  nand (_26432_, _26431_, _26429_);
  nor (_26433_, _08882_, _05994_);
  nor (_26434_, _26433_, _25727_);
  and (_26435_, _26434_, _26432_);
  or (_26436_, _26435_, _26329_);
  nand (_26437_, _26436_, _12576_);
  nor (_26438_, _26318_, _12576_);
  nor (_26439_, _26438_, _06433_);
  nand (_26440_, _26439_, _26437_);
  and (_26441_, _12156_, _06433_);
  nor (_26442_, _26441_, _25090_);
  nand (_26443_, _26442_, _26440_);
  and (_26444_, _08882_, _25090_);
  nor (_26447_, _26444_, _06432_);
  and (_26448_, _26447_, _26443_);
  and (_26449_, _12156_, _06432_);
  or (_26450_, _26449_, _26448_);
  nand (_26451_, _26450_, _12588_);
  nor (_26452_, _26330_, _12588_);
  nor (_26453_, _26452_, _12593_);
  nand (_26454_, _26453_, _26451_);
  nor (_26455_, _12156_, _12592_);
  nor (_26456_, _26455_, _06022_);
  nand (_26457_, _26456_, _26454_);
  and (_26458_, _26318_, _06022_);
  nor (_26459_, _26458_, _06300_);
  and (_26460_, _26459_, _26457_);
  and (_26461_, _12157_, _06300_);
  or (_26462_, _26461_, _26460_);
  nand (_26463_, _26462_, _07846_);
  and (_26464_, _08882_, _06017_);
  nor (_26465_, _26464_, _06472_);
  nand (_26466_, _26465_, _26463_);
  and (_26468_, _12304_, _06472_);
  nor (_26469_, _26468_, _13788_);
  and (_26470_, _26469_, _26466_);
  nor (_26471_, _12156_, _06294_);
  or (_26472_, _26471_, _26470_);
  nand (_26473_, _26472_, _06279_);
  and (_26474_, _12305_, _06015_);
  nor (_26475_, _26474_, _12620_);
  nand (_26476_, _26475_, _26473_);
  nor (_26477_, _26330_, _12616_);
  nor (_26479_, _26477_, _06376_);
  nand (_26480_, _26479_, _26476_);
  and (_26481_, _12157_, _06376_);
  nor (_26482_, _26481_, _05936_);
  and (_26483_, _26482_, _26480_);
  nor (_26484_, _08882_, _25116_);
  or (_26485_, _26484_, _26483_);
  nand (_26486_, _26485_, _12625_);
  and (_26487_, _26323_, _12624_);
  nor (_26488_, _26487_, _09013_);
  and (_26489_, _26488_, _26486_);
  or (_26490_, _26489_, _26328_);
  nand (_26491_, _26490_, _06276_);
  and (_26492_, _12305_, _06275_);
  nor (_26493_, _26492_, _10933_);
  nand (_26494_, _26493_, _26491_);
  and (_26495_, _12156_, _10933_);
  nor (_26496_, _26495_, _12639_);
  nand (_26497_, _26496_, _26494_);
  and (_26498_, _12654_, _12651_);
  nor (_26499_, _26498_, _12655_);
  nor (_26500_, _26499_, _12640_);
  nor (_26501_, _26500_, _06375_);
  nand (_26502_, _26501_, _26497_);
  and (_26503_, _12156_, _06375_);
  nor (_26504_, _26503_, _05943_);
  nand (_26505_, _26504_, _26502_);
  and (_26506_, _08882_, _05943_);
  nor (_26507_, _26506_, _12680_);
  and (_26508_, _26507_, _26505_);
  and (_26509_, _12156_, _11297_);
  and (_26510_, _26323_, _12687_);
  or (_26511_, _26510_, _26509_);
  and (_26512_, _26511_, _12680_);
  or (_26513_, _26512_, _26508_);
  nand (_26514_, _26513_, _12233_);
  nor (_26515_, _26330_, _12233_);
  nor (_26516_, _26515_, _12228_);
  nand (_26517_, _26516_, _26514_);
  nor (_26518_, _12156_, _12227_);
  nor (_26519_, _26518_, _06474_);
  nand (_26520_, _26519_, _26517_);
  and (_26521_, _12304_, _06474_);
  nor (_26522_, _26521_, _06582_);
  and (_26523_, _26522_, _26520_);
  and (_26524_, _12157_, _06582_);
  or (_26525_, _26524_, _26523_);
  nand (_26526_, _26525_, _24995_);
  and (_26527_, _08882_, _05952_);
  nor (_26528_, _26527_, _12704_);
  and (_26529_, _26528_, _26526_);
  or (_26530_, _26529_, _26327_);
  nand (_26531_, _26530_, _12719_);
  nor (_26532_, _26330_, _12719_);
  nor (_26533_, _26532_, _12722_);
  nand (_26534_, _26533_, _26531_);
  nor (_26535_, _12156_, _12721_);
  nor (_26536_, _26535_, _06478_);
  nand (_26537_, _26536_, _26534_);
  and (_26538_, _12304_, _06478_);
  nor (_26540_, _26538_, _06569_);
  and (_26541_, _26540_, _26537_);
  and (_26542_, _12157_, _06569_);
  or (_26543_, _26542_, _26541_);
  nand (_26544_, _26543_, _24992_);
  and (_26545_, _08882_, _05956_);
  nor (_26546_, _26545_, _12735_);
  and (_26547_, _26546_, _26544_);
  and (_26548_, _12156_, \uc8051golden_1.PSW [7]);
  and (_26549_, _26323_, _10524_);
  or (_26551_, _26549_, _26548_);
  and (_26552_, _26551_, _12735_);
  or (_26553_, _26552_, _26547_);
  nand (_26554_, _26553_, _12225_);
  and (_26555_, _26318_, _12224_);
  nor (_26556_, _26555_, _11019_);
  nand (_26557_, _26556_, _26554_);
  nor (_26558_, _12156_, _11018_);
  nor (_26559_, _26558_, _06479_);
  nand (_26560_, _26559_, _26557_);
  and (_26561_, _12304_, _06479_);
  nor (_26562_, _26561_, _06572_);
  and (_26563_, _26562_, _26560_);
  and (_26564_, _12157_, _06572_);
  or (_26565_, _26564_, _26563_);
  nand (_26566_, _26565_, _05948_);
  and (_26567_, _08882_, _05947_);
  nor (_26568_, _26567_, _12217_);
  and (_26569_, _26568_, _26566_);
  and (_26570_, _12156_, _10524_);
  and (_26572_, _26323_, \uc8051golden_1.PSW [7]);
  or (_26573_, _26572_, _26570_);
  and (_26574_, _26573_, _12217_);
  or (_26575_, _26574_, _26569_);
  nand (_26576_, _26575_, _12761_);
  nor (_26577_, _26330_, _12761_);
  nor (_26578_, _26577_, _11061_);
  nand (_26579_, _26578_, _26576_);
  nor (_26580_, _12156_, _11060_);
  nor (_26581_, _26580_, _11089_);
  nand (_26583_, _26581_, _26579_);
  and (_26584_, _26318_, _11089_);
  nor (_26585_, _26584_, _06588_);
  and (_26586_, _26585_, _26583_);
  and (_26587_, _09210_, _06588_);
  or (_26588_, _26587_, _26586_);
  nand (_26589_, _26588_, _05967_);
  and (_26590_, _08882_, _05966_);
  nor (_26591_, _26590_, _06460_);
  and (_26592_, _26591_, _26589_);
  nor (_26594_, _12305_, _12958_);
  and (_26595_, _26334_, _12958_);
  nor (_26596_, _26595_, _26594_);
  nor (_26597_, _26596_, _06596_);
  or (_26598_, _26597_, _26592_);
  nand (_26599_, _26598_, _12108_);
  nor (_26600_, _26330_, _12108_);
  nor (_26601_, _26600_, _12094_);
  nand (_26602_, _26601_, _26599_);
  nor (_26603_, _12156_, _11204_);
  nor (_26605_, _26603_, _11243_);
  nand (_26606_, _26605_, _26602_);
  and (_26607_, _26318_, _11243_);
  nor (_26608_, _26607_, _06305_);
  nand (_26609_, _26608_, _26606_);
  and (_26610_, _09210_, _06305_);
  nor (_26611_, _26610_, _05971_);
  nand (_26612_, _26611_, _26609_);
  nor (_26613_, _08882_, _12979_);
  nor (_26614_, _26613_, _06487_);
  nand (_26616_, _26614_, _26612_);
  nor (_26617_, _26334_, _12958_);
  and (_26618_, _12305_, _12958_);
  nor (_26619_, _26618_, _26617_);
  nor (_26620_, _26619_, _12978_);
  nor (_26621_, _26620_, _12988_);
  nand (_26622_, _26621_, _26616_);
  nor (_26623_, _26330_, _12987_);
  nor (_26624_, _26623_, _06606_);
  nand (_26625_, _26624_, _26622_);
  and (_26626_, _12157_, _06606_);
  nor (_26627_, _26626_, _12995_);
  nand (_26628_, _26627_, _26625_);
  nor (_26629_, _26330_, _12994_);
  nor (_26630_, _26629_, _07887_);
  nand (_26631_, _26630_, _26628_);
  and (_26632_, _08882_, _07887_);
  nor (_26633_, _26632_, _06234_);
  nand (_26634_, _26633_, _26631_);
  and (_26635_, _26619_, _06234_);
  nor (_26637_, _26635_, _13012_);
  and (_26638_, _26637_, _26634_);
  or (_26639_, _26638_, _26320_);
  nand (_26640_, _26639_, _06196_);
  and (_26641_, _12157_, _06195_);
  nor (_26642_, _26641_, _13020_);
  nand (_26643_, _26642_, _26640_);
  nor (_26644_, _26330_, _13019_);
  nor (_26645_, _26644_, _24972_);
  nand (_26646_, _26645_, _26643_);
  and (_26648_, _24972_, _08882_);
  nor (_26649_, _26648_, _13030_);
  and (_26650_, _26649_, _26646_);
  or (_26651_, _26650_, _26319_);
  or (_26652_, _26651_, _01379_);
  or (_26653_, _01375_, \uc8051golden_1.PC [4]);
  and (_26654_, _26653_, _42545_);
  and (_42981_, _26654_, _26652_);
  nor (_26655_, \uc8051golden_1.PC [5], \uc8051golden_1.PC [0]);
  nor (_26656_, _12151_, _05685_);
  nor (_26657_, _26656_, _26655_);
  and (_26658_, _26657_, _13030_);
  and (_26659_, _12151_, _06195_);
  and (_26660_, _12151_, _06606_);
  nor (_26661_, _26657_, _12108_);
  and (_26662_, _09165_, _06588_);
  nor (_26663_, _26657_, _12761_);
  not (_26664_, _26657_);
  and (_26665_, _26664_, _12224_);
  nor (_26666_, _26657_, _12719_);
  nor (_26669_, _26657_, _12233_);
  nor (_26670_, _12151_, _09012_);
  nor (_26671_, _12569_, _12151_);
  and (_26672_, _26664_, _12237_);
  or (_26673_, _12301_, _12302_);
  and (_26674_, _26673_, _12333_);
  nor (_26675_, _26673_, _12333_);
  nor (_26676_, _26675_, _26674_);
  not (_26677_, _26676_);
  or (_26678_, _26677_, _12405_);
  or (_26680_, _12407_, _12300_);
  nand (_26681_, _26680_, _26678_);
  nand (_26682_, _26681_, _06457_);
  or (_26683_, _12464_, _12299_);
  or (_26684_, _26676_, _12466_);
  and (_26685_, _26684_, _26683_);
  or (_26686_, _26685_, _07210_);
  and (_26687_, _12476_, _12151_);
  or (_26688_, _12154_, _12153_);
  not (_26689_, _26688_);
  nor (_26690_, _26689_, _12179_);
  and (_26691_, _26689_, _12179_);
  nor (_26692_, _26691_, _26690_);
  nor (_26693_, _26692_, _12476_);
  nor (_26694_, _26693_, _26687_);
  nand (_26695_, _26694_, _08643_);
  or (_26696_, _08917_, _07366_);
  and (_26697_, _12152_, _07199_);
  or (_26698_, _26697_, _06854_);
  nand (_26699_, _07333_, \uc8051golden_1.PC [5]);
  and (_26701_, _26699_, _07200_);
  or (_26702_, _26701_, _26698_);
  or (_26703_, _26664_, _12492_);
  and (_26704_, _26703_, _12491_);
  and (_26705_, _26704_, _26702_);
  or (_26706_, _26705_, _06790_);
  and (_26707_, _26706_, _26696_);
  and (_26708_, _26664_, _12481_);
  or (_26709_, _26708_, _26707_);
  and (_26710_, _26709_, _08644_);
  nor (_26712_, _26710_, _07212_);
  and (_26713_, _26712_, _26695_);
  and (_26714_, _26657_, _07212_);
  or (_26715_, _26714_, _06401_);
  or (_26716_, _26715_, _26713_);
  nand (_26717_, _26716_, _26686_);
  nand (_26718_, _26717_, _12458_);
  nor (_26719_, _26657_, _12458_);
  nor (_26720_, _26719_, _06395_);
  nand (_26721_, _26720_, _26718_);
  and (_26723_, _12151_, _06395_);
  nor (_26724_, _26723_, _07351_);
  nand (_26725_, _26724_, _26721_);
  and (_26726_, _08917_, _07351_);
  nor (_26727_, _26726_, _06399_);
  nand (_26728_, _26727_, _26725_);
  and (_26729_, _12151_, _06399_);
  nor (_26730_, _26729_, _12510_);
  nand (_26731_, _26730_, _26728_);
  nor (_26732_, _26657_, _12509_);
  nor (_26734_, _26732_, _06406_);
  nand (_26735_, _26734_, _26731_);
  and (_26736_, _12151_, _06406_);
  nor (_26737_, _26736_, _12519_);
  nand (_26738_, _26737_, _26735_);
  nor (_26739_, _26657_, _12517_);
  nor (_26740_, _26739_, _06393_);
  nand (_26741_, _26740_, _26738_);
  and (_26742_, _12151_, _06393_);
  nor (_26743_, _26742_, _12521_);
  nand (_26745_, _26743_, _26741_);
  and (_26746_, _08917_, _12521_);
  nor (_26747_, _26746_, _06419_);
  nand (_26748_, _26747_, _26745_);
  and (_26749_, _12151_, _06419_);
  nor (_26750_, _26749_, _12450_);
  nand (_26751_, _26750_, _26748_);
  and (_26752_, _12444_, _12299_);
  nor (_26753_, _26677_, _12444_);
  or (_26754_, _26753_, _26752_);
  nor (_26755_, _26754_, _12449_);
  nor (_26756_, _26755_, _06457_);
  nand (_26757_, _26756_, _26751_);
  and (_26758_, _26757_, _06842_);
  nand (_26759_, _26758_, _26682_);
  and (_26760_, _12546_, _12299_);
  not (_26761_, _26760_);
  nor (_26762_, _26677_, _12546_);
  nor (_26763_, _26762_, _06842_);
  and (_26764_, _26763_, _26761_);
  nor (_26766_, _26764_, _06482_);
  nand (_26767_, _26766_, _26759_);
  and (_26768_, _12299_, _12249_);
  and (_26769_, _26676_, _26421_);
  or (_26770_, _26769_, _26768_);
  and (_26771_, _26770_, _06482_);
  nor (_26772_, _26771_, _12237_);
  and (_26773_, _26772_, _26767_);
  or (_26774_, _26773_, _26672_);
  nand (_26775_, _26774_, _07245_);
  and (_26777_, _12152_, _06387_);
  nor (_26778_, _26777_, _07349_);
  nand (_26779_, _26778_, _26775_);
  nor (_26780_, _08917_, _05994_);
  nor (_26781_, _26780_, _25727_);
  and (_26782_, _26781_, _26779_);
  or (_26783_, _26782_, _26671_);
  nand (_26784_, _26783_, _12576_);
  nor (_26785_, _26657_, _12576_);
  nor (_26786_, _26785_, _06433_);
  nand (_26788_, _26786_, _26784_);
  and (_26789_, _12151_, _06433_);
  nor (_26790_, _26789_, _25090_);
  nand (_26791_, _26790_, _26788_);
  and (_26792_, _08917_, _25090_);
  nor (_26793_, _26792_, _06432_);
  nand (_26794_, _26793_, _26791_);
  and (_26795_, _12151_, _06432_);
  nor (_26796_, _26795_, _12594_);
  and (_26797_, _26796_, _26794_);
  nor (_26799_, _26657_, _12588_);
  or (_26800_, _26799_, _26797_);
  nand (_26801_, _26800_, _12592_);
  nor (_26802_, _12151_, _12592_);
  nor (_26803_, _26802_, _06022_);
  nand (_26804_, _26803_, _26801_);
  and (_26805_, _26657_, _06022_);
  nor (_26806_, _26805_, _06300_);
  and (_26807_, _26806_, _26804_);
  and (_26808_, _12152_, _06300_);
  or (_26810_, _26808_, _26807_);
  nand (_26811_, _26810_, _07846_);
  and (_26812_, _08917_, _06017_);
  nor (_26813_, _26812_, _06472_);
  nand (_26814_, _26813_, _26811_);
  and (_26815_, _12299_, _06472_);
  nor (_26816_, _26815_, _13788_);
  nand (_26817_, _26816_, _26814_);
  nor (_26818_, _12151_, _06294_);
  nor (_26819_, _26818_, _06015_);
  nand (_26820_, _26819_, _26817_);
  and (_26821_, _12299_, _06015_);
  nor (_26822_, _26821_, _12620_);
  nand (_26823_, _26822_, _26820_);
  nor (_26824_, _26657_, _12616_);
  nor (_26825_, _26824_, _06376_);
  nand (_26826_, _26825_, _26823_);
  and (_26827_, _12151_, _06376_);
  nor (_26828_, _26827_, _05936_);
  nand (_26829_, _26828_, _26826_);
  and (_26831_, _08917_, _05936_);
  nor (_26832_, _26831_, _12624_);
  nand (_26833_, _26832_, _26829_);
  nor (_26834_, _26692_, _12625_);
  nor (_26835_, _26834_, _09013_);
  and (_26836_, _26835_, _26833_);
  or (_26837_, _26836_, _26670_);
  nand (_26838_, _26837_, _06276_);
  and (_26839_, _12300_, _06275_);
  nor (_26840_, _26839_, _10933_);
  nand (_26842_, _26840_, _26838_);
  and (_26843_, _12151_, _10933_);
  nor (_26844_, _26843_, _12639_);
  and (_26845_, _26844_, _26842_);
  or (_26846_, _12649_, _12648_);
  nand (_26847_, _26846_, _12656_);
  or (_26848_, _26846_, _12656_);
  and (_26849_, _26848_, _26847_);
  nor (_26850_, _26849_, _12640_);
  nor (_26851_, _26850_, _26845_);
  nand (_26853_, _26851_, _06952_);
  and (_26854_, _12151_, _06375_);
  nor (_26855_, _26854_, _05943_);
  nand (_26856_, _26855_, _26853_);
  and (_26857_, _08917_, _05943_);
  nor (_26858_, _26857_, _12680_);
  nand (_26859_, _26858_, _26856_);
  and (_26860_, _12151_, _11297_);
  nor (_26861_, _26692_, _11297_);
  or (_26862_, _26861_, _26860_);
  and (_26864_, _26862_, _12680_);
  nor (_26865_, _26864_, _12685_);
  and (_26866_, _26865_, _26859_);
  or (_26867_, _26866_, _26669_);
  nand (_26868_, _26867_, _12227_);
  nor (_26869_, _12151_, _12227_);
  nor (_26870_, _26869_, _06474_);
  nand (_26871_, _26870_, _26868_);
  and (_26872_, _12299_, _06474_);
  nor (_26873_, _26872_, _06582_);
  and (_26875_, _26873_, _26871_);
  and (_26876_, _12152_, _06582_);
  or (_26877_, _26876_, _26875_);
  nand (_26878_, _26877_, _24995_);
  and (_26879_, _08917_, _05952_);
  nor (_26880_, _26879_, _12704_);
  nand (_26881_, _26880_, _26878_);
  nor (_26882_, _12152_, _11297_);
  nor (_26883_, _26692_, _12687_);
  or (_26884_, _26883_, _26882_);
  and (_26885_, _26884_, _12704_);
  nor (_26886_, _26885_, _12723_);
  and (_26887_, _26886_, _26881_);
  or (_26888_, _26887_, _26666_);
  nand (_26889_, _26888_, _12721_);
  nor (_26890_, _12151_, _12721_);
  nor (_26891_, _26890_, _06478_);
  nand (_26892_, _26891_, _26889_);
  and (_26893_, _12299_, _06478_);
  nor (_26894_, _26893_, _06569_);
  and (_26896_, _26894_, _26892_);
  and (_26897_, _12152_, _06569_);
  or (_26898_, _26897_, _26896_);
  nand (_26899_, _26898_, _24992_);
  and (_26900_, _08917_, _05956_);
  nor (_26901_, _26900_, _12735_);
  nand (_26902_, _26901_, _26899_);
  and (_26903_, _26692_, _10524_);
  nor (_26904_, _12151_, _10524_);
  nor (_26905_, _26904_, _12736_);
  not (_26907_, _26905_);
  nor (_26908_, _26907_, _26903_);
  nor (_26909_, _26908_, _12224_);
  and (_26910_, _26909_, _26902_);
  or (_26911_, _26910_, _26665_);
  nand (_26912_, _26911_, _11018_);
  nor (_26913_, _12151_, _11018_);
  nor (_26914_, _26913_, _06479_);
  nand (_26915_, _26914_, _26912_);
  and (_26916_, _12299_, _06479_);
  nor (_26918_, _26916_, _06572_);
  and (_26919_, _26918_, _26915_);
  and (_26920_, _12152_, _06572_);
  or (_26921_, _26920_, _26919_);
  nand (_26922_, _26921_, _05948_);
  and (_26923_, _08917_, _05947_);
  nor (_26924_, _26923_, _12217_);
  nand (_26925_, _26924_, _26922_);
  and (_26926_, _12151_, _10524_);
  nor (_26927_, _26692_, _10524_);
  or (_26929_, _26927_, _26926_);
  and (_26930_, _26929_, _12217_);
  nor (_26931_, _26930_, _12763_);
  and (_26932_, _26931_, _26925_);
  or (_26933_, _26932_, _26663_);
  nand (_26934_, _26933_, _11060_);
  nor (_26935_, _12151_, _11060_);
  nor (_26936_, _26935_, _11089_);
  nand (_26937_, _26936_, _26934_);
  and (_26938_, _26657_, _11089_);
  nor (_26940_, _26938_, _06588_);
  and (_26941_, _26940_, _26937_);
  or (_26942_, _26941_, _26662_);
  nand (_26943_, _26942_, _05967_);
  and (_26944_, _08917_, _05966_);
  nor (_26945_, _26944_, _06460_);
  nand (_26946_, _26945_, _26943_);
  and (_26947_, _26677_, _12958_);
  nor (_26948_, _12299_, _12958_);
  or (_26949_, _26948_, _06596_);
  or (_26951_, _26949_, _26947_);
  and (_26952_, _26951_, _12108_);
  and (_26953_, _26952_, _26946_);
  or (_26954_, _26953_, _26661_);
  nand (_26955_, _26954_, _11204_);
  nor (_26956_, _12151_, _11204_);
  nor (_26957_, _26956_, _11243_);
  nand (_26958_, _26957_, _26955_);
  and (_26959_, _26657_, _11243_);
  nor (_26960_, _26959_, _06305_);
  and (_26962_, _26960_, _26958_);
  and (_26963_, _09165_, _06305_);
  or (_26964_, _26963_, _26962_);
  nand (_26965_, _26964_, _12979_);
  and (_26966_, _08917_, _05971_);
  nor (_26967_, _26966_, _06487_);
  nand (_26968_, _26967_, _26965_);
  and (_26969_, _12300_, _12958_);
  nor (_26970_, _26676_, _12958_);
  nor (_26971_, _26970_, _26969_);
  and (_26972_, _26971_, _06487_);
  nor (_26973_, _26972_, _12988_);
  nand (_26974_, _26973_, _26968_);
  nor (_26975_, _26657_, _12987_);
  nor (_26976_, _26975_, _06606_);
  and (_26977_, _26976_, _26974_);
  or (_26978_, _26977_, _26660_);
  nand (_26979_, _26978_, _12994_);
  nor (_26980_, _26664_, _12994_);
  nor (_26981_, _26980_, _07887_);
  nand (_26983_, _26981_, _26979_);
  and (_26984_, _08917_, _07887_);
  nor (_26985_, _26984_, _06234_);
  nand (_26986_, _26985_, _26983_);
  and (_26987_, _26971_, _06234_);
  nor (_26988_, _26987_, _13012_);
  nand (_26989_, _26988_, _26986_);
  nor (_26990_, _26657_, _13011_);
  nor (_26991_, _26990_, _06195_);
  and (_26992_, _26991_, _26989_);
  or (_26994_, _26992_, _26659_);
  nand (_26995_, _26994_, _13019_);
  nor (_26996_, _26664_, _13019_);
  nor (_26997_, _26996_, _24972_);
  nand (_26998_, _26997_, _26995_);
  and (_26999_, _24972_, _08917_);
  nor (_27000_, _26999_, _13030_);
  and (_27001_, _27000_, _26998_);
  or (_27002_, _27001_, _26658_);
  or (_27003_, _27002_, _01379_);
  or (_27005_, _01375_, \uc8051golden_1.PC [5]);
  and (_27006_, _27005_, _42545_);
  and (_42982_, _27006_, _27003_);
  nand (_27007_, _08850_, _07887_);
  and (_27008_, _08532_, _12095_);
  nor (_27009_, _27008_, \uc8051golden_1.PC [6]);
  nor (_27010_, _27009_, _12096_);
  not (_27011_, _27010_);
  nand (_27012_, _27011_, _11243_);
  nand (_27013_, _12293_, _06479_);
  nand (_27015_, _12293_, _06478_);
  nand (_27016_, _12293_, _06474_);
  nand (_27017_, _27011_, _12237_);
  nor (_27018_, _12335_, _12296_);
  nor (_27019_, _27018_, _12336_);
  or (_27020_, _27019_, _12405_);
  or (_27021_, _12407_, _12292_);
  and (_27022_, _27021_, _27020_);
  or (_27023_, _27022_, _12411_);
  or (_27024_, _27010_, _12503_);
  and (_27026_, _12466_, _12292_);
  and (_27027_, _27019_, _12464_);
  or (_27028_, _27027_, _07210_);
  or (_27029_, _27028_, _27026_);
  nand (_27030_, _08850_, _06790_);
  nand (_27031_, _12145_, _07199_);
  and (_27032_, _27031_, _06855_);
  and (_27033_, _07333_, \uc8051golden_1.PC [6]);
  or (_27034_, _27033_, _07199_);
  and (_27035_, _27034_, _27032_);
  nor (_27036_, _27011_, _12492_);
  or (_27037_, _27036_, _06790_);
  or (_27038_, _27037_, _27035_);
  and (_27039_, _27038_, _12491_);
  and (_27040_, _27039_, _27030_);
  and (_27041_, _27010_, _12481_);
  or (_27042_, _27041_, _08643_);
  or (_27043_, _27042_, _27040_);
  nor (_27044_, _12182_, _12148_);
  nor (_27045_, _27044_, _12183_);
  and (_27047_, _27045_, _12474_);
  and (_27048_, _12476_, _12144_);
  or (_27049_, _27048_, _08644_);
  or (_27050_, _27049_, _27047_);
  nand (_27051_, _27050_, _27043_);
  nand (_27052_, _27051_, _12497_);
  and (_27053_, _27052_, _27029_);
  or (_27054_, _27053_, _25041_);
  and (_27055_, _27054_, _27024_);
  or (_27056_, _27055_, _06395_);
  nand (_27058_, _12145_, _06395_);
  and (_27059_, _27058_, _05997_);
  and (_27060_, _27059_, _27056_);
  nor (_27061_, _08850_, _05997_);
  or (_27062_, _27061_, _06399_);
  or (_27063_, _27062_, _27060_);
  nand (_27064_, _12145_, _06399_);
  and (_27065_, _27064_, _12509_);
  and (_27066_, _27065_, _27063_);
  nor (_27067_, _27011_, _12509_);
  or (_27069_, _27067_, _06406_);
  or (_27070_, _27069_, _27066_);
  nand (_27071_, _12145_, _06406_);
  and (_27072_, _27071_, _12517_);
  and (_27073_, _27072_, _27070_);
  nor (_27074_, _27011_, _12517_);
  or (_27075_, _27074_, _06393_);
  or (_27076_, _27075_, _27073_);
  nand (_27077_, _12145_, _06393_);
  and (_27078_, _27077_, _27076_);
  or (_27080_, _27078_, _12521_);
  nand (_27081_, _08850_, _12521_);
  and (_27082_, _27081_, _07785_);
  and (_27083_, _27082_, _27080_);
  nand (_27084_, _12144_, _06419_);
  nand (_27085_, _27084_, _12449_);
  or (_27086_, _27085_, _27083_);
  not (_27087_, _27019_);
  nor (_27088_, _27087_, _12444_);
  and (_27089_, _12444_, _12292_);
  or (_27091_, _27089_, _12449_);
  or (_27092_, _27091_, _27088_);
  and (_27093_, _27092_, _27086_);
  or (_27094_, _27093_, _06457_);
  and (_27095_, _27094_, _27023_);
  or (_27096_, _27095_, _06420_);
  nor (_27097_, _27087_, _12546_);
  and (_27098_, _12546_, _12292_);
  or (_27099_, _27098_, _06842_);
  or (_27100_, _27099_, _27097_);
  and (_27102_, _27100_, _12534_);
  and (_27103_, _27102_, _27096_);
  or (_27104_, _27019_, _12249_);
  nand (_27105_, _12293_, _12249_);
  and (_27106_, _27105_, _06482_);
  and (_27107_, _27106_, _27104_);
  or (_27108_, _27107_, _12237_);
  or (_27109_, _27108_, _27103_);
  and (_27110_, _27109_, _27017_);
  or (_27111_, _27110_, _06387_);
  nand (_27113_, _12145_, _06387_);
  and (_27114_, _27113_, _05994_);
  and (_27115_, _27114_, _27111_);
  nor (_27116_, _08850_, _05994_);
  or (_27117_, _27116_, _25727_);
  or (_27118_, _27117_, _27115_);
  or (_27119_, _12569_, _12144_);
  and (_27120_, _27119_, _27118_);
  or (_27121_, _27120_, _12580_);
  or (_27122_, _27010_, _12576_);
  and (_27124_, _27122_, _14016_);
  and (_27125_, _27124_, _27121_);
  and (_27126_, _12144_, _06433_);
  or (_27127_, _27126_, _25090_);
  or (_27128_, _27127_, _27125_);
  nand (_27129_, _08850_, _25090_);
  and (_27130_, _27129_, _14015_);
  and (_27131_, _27130_, _27128_);
  nand (_27132_, _12144_, _06432_);
  nand (_27133_, _27132_, _12588_);
  or (_27135_, _27133_, _27131_);
  or (_27136_, _27010_, _12588_);
  and (_27137_, _27136_, _12592_);
  and (_27138_, _27137_, _27135_);
  nor (_27139_, _12145_, _12592_);
  or (_27140_, _27139_, _06022_);
  or (_27141_, _27140_, _27138_);
  nand (_27142_, _27011_, _06022_);
  and (_27143_, _27142_, _27141_);
  or (_27144_, _27143_, _06300_);
  nand (_27146_, _12145_, _06300_);
  and (_27147_, _27146_, _07846_);
  and (_27148_, _27147_, _27144_);
  nor (_27149_, _08850_, _07846_);
  or (_27150_, _27149_, _06472_);
  or (_27151_, _27150_, _27148_);
  nand (_27152_, _12293_, _06472_);
  and (_27153_, _27152_, _06294_);
  and (_27154_, _27153_, _27151_);
  nor (_27155_, _12145_, _06294_);
  or (_27157_, _27155_, _06015_);
  or (_27158_, _27157_, _27154_);
  nand (_27159_, _12293_, _06015_);
  and (_27160_, _27159_, _12616_);
  and (_27161_, _27160_, _27158_);
  nor (_27162_, _27011_, _12616_);
  or (_27163_, _27162_, _06376_);
  or (_27164_, _27163_, _27161_);
  nand (_27165_, _12145_, _06376_);
  and (_27166_, _27165_, _25116_);
  and (_27168_, _27166_, _27164_);
  nor (_27169_, _08850_, _25116_);
  or (_27170_, _27169_, _12624_);
  or (_27171_, _27170_, _27168_);
  or (_27172_, _27045_, _12625_);
  and (_27173_, _27172_, _09012_);
  and (_27174_, _27173_, _27171_);
  nor (_27175_, _12145_, _09012_);
  or (_27176_, _27175_, _06275_);
  or (_27177_, _27176_, _27174_);
  nand (_27179_, _12293_, _06275_);
  and (_27180_, _27179_, _10934_);
  and (_27181_, _27180_, _27177_);
  and (_27182_, _12144_, _10933_);
  or (_27183_, _27182_, _12639_);
  or (_27184_, _27183_, _27181_);
  nor (_27185_, _12659_, _12647_);
  nor (_27186_, _27185_, _12660_);
  or (_27187_, _27186_, _12640_);
  and (_27188_, _27187_, _06952_);
  and (_27190_, _27188_, _27184_);
  and (_27191_, _12144_, _06375_);
  or (_27192_, _27191_, _05943_);
  or (_27193_, _27192_, _27190_);
  nand (_27194_, _08850_, _05943_);
  and (_27195_, _27194_, _12681_);
  and (_27196_, _27195_, _27193_);
  or (_27197_, _27045_, _11297_);
  nand (_27198_, _12145_, _11297_);
  and (_27199_, _27198_, _12680_);
  and (_27201_, _27199_, _27197_);
  or (_27202_, _27201_, _12685_);
  or (_27203_, _27202_, _27196_);
  or (_27204_, _27010_, _12233_);
  and (_27205_, _27204_, _12227_);
  and (_27206_, _27205_, _27203_);
  nor (_27207_, _12145_, _12227_);
  or (_27208_, _27207_, _06474_);
  or (_27209_, _27208_, _27206_);
  and (_27210_, _27209_, _27016_);
  or (_27212_, _27210_, _06582_);
  nand (_27213_, _12145_, _06582_);
  and (_27214_, _27213_, _24995_);
  and (_27215_, _27214_, _27212_);
  nor (_27216_, _08850_, _24995_);
  or (_27217_, _27216_, _27215_);
  and (_27218_, _27217_, _12705_);
  or (_27219_, _27045_, _12687_);
  or (_27220_, _12144_, _11297_);
  and (_27221_, _27220_, _12704_);
  and (_27223_, _27221_, _27219_);
  or (_27224_, _27223_, _12723_);
  or (_27225_, _27224_, _27218_);
  or (_27226_, _27010_, _12719_);
  and (_27227_, _27226_, _12721_);
  and (_27228_, _27227_, _27225_);
  nor (_27229_, _12145_, _12721_);
  or (_27230_, _27229_, _06478_);
  or (_27231_, _27230_, _27228_);
  and (_27232_, _27231_, _27015_);
  or (_27233_, _27232_, _06569_);
  nand (_27234_, _12145_, _06569_);
  and (_27235_, _27234_, _24992_);
  and (_27236_, _27235_, _27233_);
  nor (_27237_, _08850_, _24992_);
  or (_27238_, _27237_, _27236_);
  and (_27239_, _27238_, _12736_);
  or (_27240_, _27045_, \uc8051golden_1.PSW [7]);
  or (_27241_, _12144_, _10524_);
  and (_27242_, _27241_, _12735_);
  and (_27245_, _27242_, _27240_);
  or (_27246_, _27245_, _12224_);
  or (_27247_, _27246_, _27239_);
  nand (_27248_, _27011_, _12224_);
  and (_27249_, _27248_, _11018_);
  and (_27250_, _27249_, _27247_);
  nor (_27251_, _12145_, _11018_);
  or (_27252_, _27251_, _06479_);
  or (_27253_, _27252_, _27250_);
  and (_27254_, _27253_, _27013_);
  or (_27256_, _27254_, _06572_);
  nand (_27257_, _12145_, _06572_);
  and (_27258_, _27257_, _05948_);
  and (_27259_, _27258_, _27256_);
  nor (_27260_, _08850_, _05948_);
  or (_27261_, _27260_, _27259_);
  and (_27262_, _27261_, _12756_);
  or (_27263_, _27045_, _10524_);
  or (_27264_, _12144_, \uc8051golden_1.PSW [7]);
  and (_27265_, _27264_, _12217_);
  and (_27267_, _27265_, _27263_);
  or (_27268_, _27267_, _12763_);
  or (_27269_, _27268_, _27262_);
  or (_27270_, _27010_, _12761_);
  and (_27271_, _27270_, _11060_);
  and (_27272_, _27271_, _27269_);
  nor (_27273_, _12145_, _11060_);
  or (_27274_, _27273_, _11089_);
  or (_27275_, _27274_, _27272_);
  nand (_27276_, _27011_, _11089_);
  and (_27278_, _27276_, _13881_);
  and (_27279_, _27278_, _27275_);
  and (_27280_, _09440_, _06588_);
  or (_27281_, _27280_, _05966_);
  or (_27282_, _27281_, _27279_);
  nand (_27283_, _08850_, _05966_);
  and (_27284_, _27283_, _06596_);
  and (_27285_, _27284_, _27282_);
  nand (_27286_, _27087_, _12958_);
  or (_27287_, _12292_, _12958_);
  and (_27289_, _27287_, _06460_);
  and (_27290_, _27289_, _27286_);
  or (_27291_, _27290_, _12779_);
  or (_27292_, _27291_, _27285_);
  or (_27293_, _27010_, _12108_);
  and (_27294_, _27293_, _11204_);
  and (_27295_, _27294_, _27292_);
  nor (_27296_, _12145_, _11204_);
  or (_27297_, _27296_, _11243_);
  or (_27298_, _27297_, _27295_);
  and (_27300_, _27298_, _27012_);
  or (_27301_, _27300_, _06305_);
  or (_27302_, _09440_, _06306_);
  and (_27303_, _27302_, _12979_);
  and (_27304_, _27303_, _27301_);
  nor (_27305_, _08850_, _12979_);
  or (_27306_, _27305_, _06487_);
  or (_27307_, _27306_, _27304_);
  nor (_27308_, _27019_, _12958_);
  and (_27309_, _12293_, _12958_);
  nor (_27311_, _27309_, _27308_);
  or (_27312_, _27311_, _12978_);
  and (_27313_, _27312_, _27307_);
  or (_27314_, _27313_, _12988_);
  or (_27315_, _27010_, _12987_);
  and (_27316_, _27315_, _27314_);
  or (_27317_, _27316_, _06606_);
  nand (_27318_, _12145_, _06606_);
  and (_27319_, _27318_, _12994_);
  and (_27320_, _27319_, _27317_);
  nor (_27322_, _27011_, _12994_);
  or (_27323_, _27322_, _07887_);
  or (_27324_, _27323_, _27320_);
  and (_27325_, _27324_, _27007_);
  or (_27326_, _27325_, _06234_);
  nor (_27327_, _27311_, _06807_);
  nor (_27328_, _27327_, _13012_);
  nand (_27329_, _27328_, _27326_);
  nor (_27330_, _27011_, _13011_);
  nor (_27331_, _27330_, _06195_);
  nand (_27333_, _27331_, _27329_);
  and (_27334_, _12145_, _06195_);
  nor (_27335_, _27334_, _13020_);
  nand (_27336_, _27335_, _27333_);
  nor (_27337_, _27011_, _13019_);
  nor (_27338_, _27337_, _24972_);
  nand (_27339_, _27338_, _27336_);
  and (_27340_, _24972_, _08850_);
  nor (_27341_, _27340_, _13030_);
  and (_27342_, _27341_, _27339_);
  and (_27344_, _27010_, _13030_);
  nor (_27345_, _27344_, _27342_);
  nand (_27346_, _27345_, _01375_);
  or (_27347_, _01375_, \uc8051golden_1.PC [6]);
  and (_27348_, _27347_, _42545_);
  and (_42983_, _27348_, _27346_);
  nor (_27349_, _12096_, \uc8051golden_1.PC [7]);
  nor (_27350_, _27349_, _12097_);
  and (_27351_, _27350_, _13030_);
  and (_27352_, _08649_, _06195_);
  nor (_27354_, _27350_, _12108_);
  nor (_27355_, _27350_, _12761_);
  not (_27356_, _27350_);
  and (_27357_, _27356_, _12224_);
  nor (_27358_, _27350_, _12719_);
  nor (_27359_, _27350_, _12233_);
  nor (_27360_, _09012_, _08649_);
  nor (_27361_, _12569_, _08649_);
  and (_27362_, _27356_, _12237_);
  and (_27363_, _12337_, _12289_);
  nor (_27365_, _27363_, _12338_);
  not (_27366_, _27365_);
  or (_27367_, _27366_, _12405_);
  or (_27368_, _12407_, _08540_);
  nand (_27369_, _27368_, _27367_);
  nand (_27370_, _27369_, _06457_);
  or (_27371_, _12464_, _08539_);
  or (_27372_, _27365_, _12466_);
  and (_27373_, _27372_, _27371_);
  or (_27374_, _27373_, _07210_);
  and (_27376_, _12476_, _08649_);
  or (_27377_, _12140_, _12141_);
  and (_27378_, _27377_, _12184_);
  nor (_27379_, _27377_, _12184_);
  nor (_27380_, _27379_, _27378_);
  and (_27381_, _27380_, _12474_);
  nor (_27382_, _27381_, _27376_);
  nand (_27383_, _27382_, _08643_);
  or (_27384_, _08590_, _07366_);
  and (_27385_, _08781_, _07199_);
  or (_27387_, _27385_, _06854_);
  nand (_27388_, _07333_, \uc8051golden_1.PC [7]);
  and (_27389_, _27388_, _07200_);
  or (_27390_, _27389_, _27387_);
  or (_27391_, _27356_, _12492_);
  and (_27392_, _27391_, _12491_);
  and (_27393_, _27392_, _27390_);
  or (_27394_, _27393_, _06790_);
  and (_27395_, _27394_, _27384_);
  and (_27396_, _27356_, _12481_);
  or (_27398_, _27396_, _27395_);
  and (_27399_, _27398_, _08644_);
  nor (_27400_, _27399_, _07212_);
  and (_27401_, _27400_, _27383_);
  and (_27402_, _27350_, _07212_);
  or (_27403_, _27402_, _06401_);
  or (_27404_, _27403_, _27401_);
  nand (_27405_, _27404_, _27374_);
  nand (_27406_, _27405_, _12458_);
  nor (_27407_, _27350_, _12458_);
  nor (_27409_, _27407_, _06395_);
  nand (_27410_, _27409_, _27406_);
  and (_27411_, _08649_, _06395_);
  nor (_27412_, _27411_, _07351_);
  nand (_27413_, _27412_, _27410_);
  and (_27414_, _08590_, _07351_);
  nor (_27415_, _27414_, _06399_);
  nand (_27416_, _27415_, _27413_);
  and (_27417_, _08649_, _06399_);
  nor (_27418_, _27417_, _12510_);
  nand (_27420_, _27418_, _27416_);
  nor (_27421_, _27350_, _12509_);
  nor (_27422_, _27421_, _06406_);
  nand (_27423_, _27422_, _27420_);
  and (_27424_, _08649_, _06406_);
  nor (_27425_, _27424_, _12519_);
  nand (_27426_, _27425_, _27423_);
  nor (_27427_, _27350_, _12517_);
  nor (_27428_, _27427_, _06393_);
  nand (_27429_, _27428_, _27426_);
  and (_27431_, _08649_, _06393_);
  nor (_27432_, _27431_, _12521_);
  nand (_27433_, _27432_, _27429_);
  and (_27434_, _08590_, _12521_);
  nor (_27435_, _27434_, _06419_);
  nand (_27436_, _27435_, _27433_);
  and (_27437_, _08649_, _06419_);
  nor (_27438_, _27437_, _12450_);
  nand (_27439_, _27438_, _27436_);
  and (_27440_, _12444_, _08539_);
  nor (_27442_, _27366_, _12444_);
  or (_27443_, _27442_, _12449_);
  nor (_27444_, _27443_, _27440_);
  nor (_27445_, _27444_, _06457_);
  nand (_27446_, _27445_, _27439_);
  and (_27447_, _27446_, _27370_);
  or (_27448_, _27447_, _06420_);
  and (_27449_, _12546_, _08539_);
  nor (_27450_, _27366_, _12546_);
  nor (_27451_, _27450_, _27449_);
  or (_27453_, _27451_, _06842_);
  and (_27454_, _27453_, _27448_);
  or (_27455_, _27454_, _06482_);
  nor (_27456_, _27365_, _12249_);
  and (_27457_, _12249_, _08540_);
  or (_27458_, _27457_, _12534_);
  or (_27459_, _27458_, _27456_);
  and (_27460_, _27459_, _12238_);
  and (_27461_, _27460_, _27455_);
  or (_27462_, _27461_, _27362_);
  nand (_27464_, _27462_, _07245_);
  and (_27465_, _08781_, _06387_);
  nor (_27466_, _27465_, _07349_);
  nand (_27467_, _27466_, _27464_);
  nor (_27468_, _08590_, _05994_);
  nor (_27469_, _27468_, _25727_);
  and (_27470_, _27469_, _27467_);
  or (_27471_, _27470_, _27361_);
  nand (_27472_, _27471_, _12576_);
  nor (_27473_, _27350_, _12576_);
  nor (_27475_, _27473_, _06433_);
  nand (_27476_, _27475_, _27472_);
  and (_27477_, _08649_, _06433_);
  nor (_27478_, _27477_, _25090_);
  nand (_27479_, _27478_, _27476_);
  and (_27480_, _08590_, _25090_);
  nor (_27481_, _27480_, _06432_);
  nand (_27482_, _27481_, _27479_);
  and (_27483_, _08649_, _06432_);
  nor (_27484_, _27483_, _12594_);
  and (_27486_, _27484_, _27482_);
  nor (_27487_, _27350_, _12588_);
  or (_27488_, _27487_, _27486_);
  nand (_27489_, _27488_, _12592_);
  nor (_27490_, _12592_, _08649_);
  nor (_27491_, _27490_, _06022_);
  nand (_27492_, _27491_, _27489_);
  and (_27493_, _27350_, _06022_);
  nor (_27494_, _27493_, _06300_);
  and (_27495_, _27494_, _27492_);
  and (_27497_, _08781_, _06300_);
  or (_27498_, _27497_, _27495_);
  nand (_27499_, _27498_, _07846_);
  and (_27500_, _08590_, _06017_);
  nor (_27501_, _27500_, _06472_);
  nand (_27502_, _27501_, _27499_);
  and (_27503_, _08539_, _06472_);
  nor (_27504_, _27503_, _13788_);
  nand (_27505_, _27504_, _27502_);
  nor (_27506_, _08649_, _06294_);
  nor (_27508_, _27506_, _06015_);
  nand (_27509_, _27508_, _27505_);
  and (_27510_, _08539_, _06015_);
  nor (_27511_, _27510_, _12620_);
  nand (_27512_, _27511_, _27509_);
  nor (_27513_, _27350_, _12616_);
  nor (_27514_, _27513_, _06376_);
  nand (_27515_, _27514_, _27512_);
  and (_27516_, _08649_, _06376_);
  nor (_27517_, _27516_, _05936_);
  nand (_27519_, _27517_, _27515_);
  and (_27520_, _08590_, _05936_);
  nor (_27521_, _27520_, _12624_);
  nand (_27522_, _27521_, _27519_);
  and (_27523_, _27380_, _12624_);
  nor (_27524_, _27523_, _09013_);
  and (_27525_, _27524_, _27522_);
  or (_27526_, _27525_, _27360_);
  nand (_27527_, _27526_, _06276_);
  and (_27528_, _08540_, _06275_);
  nor (_27530_, _27528_, _10933_);
  and (_27531_, _27530_, _27527_);
  and (_27532_, _10933_, _08649_);
  or (_27533_, _27532_, _27531_);
  nand (_27534_, _27533_, _12640_);
  or (_27535_, _12644_, _12643_);
  nor (_27536_, _27535_, _12661_);
  and (_27537_, _27535_, _12661_);
  or (_27538_, _27537_, _12640_);
  or (_27539_, _27538_, _27536_);
  and (_27541_, _27539_, _06952_);
  and (_27542_, _27541_, _27534_);
  and (_27543_, _08781_, _06375_);
  or (_27544_, _27543_, _27542_);
  nand (_27545_, _27544_, _13854_);
  and (_27546_, _08590_, _05943_);
  nor (_27547_, _27546_, _12680_);
  nand (_27548_, _27547_, _27545_);
  and (_27549_, _11297_, _08649_);
  and (_27550_, _27380_, _12687_);
  or (_27552_, _27550_, _27549_);
  and (_27553_, _27552_, _12680_);
  nor (_27554_, _27553_, _12685_);
  and (_27555_, _27554_, _27548_);
  or (_27556_, _27555_, _27359_);
  nand (_27557_, _27556_, _12227_);
  nor (_27558_, _12227_, _08649_);
  nor (_27559_, _27558_, _06474_);
  nand (_27560_, _27559_, _27557_);
  and (_27561_, _08539_, _06474_);
  nor (_27563_, _27561_, _06582_);
  and (_27564_, _27563_, _27560_);
  and (_27565_, _08781_, _06582_);
  or (_27566_, _27565_, _27564_);
  nand (_27567_, _27566_, _24995_);
  and (_27568_, _08590_, _05952_);
  nor (_27569_, _27568_, _12704_);
  nand (_27570_, _27569_, _27567_);
  nor (_27571_, _11297_, _08781_);
  and (_27572_, _27380_, _11297_);
  or (_27574_, _27572_, _27571_);
  and (_27575_, _27574_, _12704_);
  nor (_27576_, _27575_, _12723_);
  and (_27577_, _27576_, _27570_);
  or (_27578_, _27577_, _27358_);
  nand (_27579_, _27578_, _12721_);
  nor (_27580_, _12721_, _08649_);
  nor (_27581_, _27580_, _06478_);
  nand (_27582_, _27581_, _27579_);
  and (_27583_, _08539_, _06478_);
  nor (_27585_, _27583_, _06569_);
  and (_27586_, _27585_, _27582_);
  and (_27587_, _08781_, _06569_);
  or (_27588_, _27587_, _27586_);
  nand (_27589_, _27588_, _24992_);
  and (_27590_, _08590_, _05956_);
  nor (_27591_, _27590_, _12735_);
  nand (_27592_, _27591_, _27589_);
  nor (_27593_, _27380_, \uc8051golden_1.PSW [7]);
  nor (_27594_, _08649_, _10524_);
  nor (_27596_, _27594_, _12736_);
  not (_27597_, _27596_);
  nor (_27598_, _27597_, _27593_);
  nor (_27599_, _27598_, _12224_);
  and (_27600_, _27599_, _27592_);
  or (_27601_, _27600_, _27357_);
  nand (_27602_, _27601_, _11018_);
  nor (_27603_, _11018_, _08649_);
  nor (_27604_, _27603_, _06479_);
  nand (_27605_, _27604_, _27602_);
  and (_27607_, _08539_, _06479_);
  nor (_27608_, _27607_, _06572_);
  and (_27609_, _27608_, _27605_);
  and (_27610_, _08781_, _06572_);
  or (_27611_, _27610_, _27609_);
  nand (_27612_, _27611_, _05948_);
  and (_27613_, _08590_, _05947_);
  nor (_27614_, _27613_, _12217_);
  nand (_27615_, _27614_, _27612_);
  and (_27616_, _08649_, _10524_);
  and (_27618_, _27380_, \uc8051golden_1.PSW [7]);
  or (_27619_, _27618_, _27616_);
  and (_27620_, _27619_, _12217_);
  nor (_27621_, _27620_, _12763_);
  and (_27622_, _27621_, _27615_);
  or (_27623_, _27622_, _27355_);
  nand (_27624_, _27623_, _11060_);
  nor (_27625_, _11060_, _08649_);
  nor (_27626_, _27625_, _11089_);
  nand (_27627_, _27626_, _27624_);
  and (_27629_, _27350_, _11089_);
  nor (_27630_, _27629_, _06588_);
  and (_27631_, _27630_, _27627_);
  and (_27632_, _09075_, _06588_);
  or (_27633_, _27632_, _27631_);
  nand (_27634_, _27633_, _05967_);
  and (_27635_, _08590_, _05966_);
  nor (_27636_, _27635_, _06460_);
  nand (_27637_, _27636_, _27634_);
  and (_27638_, _27366_, _12958_);
  nor (_27640_, _12958_, _08539_);
  or (_27641_, _27640_, _06596_);
  or (_27642_, _27641_, _27638_);
  and (_27643_, _27642_, _12108_);
  and (_27644_, _27643_, _27637_);
  or (_27645_, _27644_, _27354_);
  nand (_27646_, _27645_, _11204_);
  nor (_27647_, _11204_, _08649_);
  nor (_27648_, _27647_, _11243_);
  nand (_27649_, _27648_, _27646_);
  and (_27651_, _27350_, _11243_);
  nor (_27652_, _27651_, _06305_);
  and (_27653_, _27652_, _27649_);
  and (_27654_, _09075_, _06305_);
  or (_27655_, _27654_, _27653_);
  nand (_27656_, _27655_, _12979_);
  and (_27657_, _08590_, _05971_);
  nor (_27658_, _27657_, _06487_);
  nand (_27659_, _27658_, _27656_);
  and (_27660_, _12958_, _08540_);
  nor (_27662_, _27365_, _12958_);
  nor (_27663_, _27662_, _27660_);
  and (_27664_, _27663_, _06487_);
  nor (_27665_, _27664_, _12988_);
  nand (_27666_, _27665_, _27659_);
  nor (_27667_, _27350_, _12987_);
  nor (_27668_, _27667_, _06606_);
  nand (_27669_, _27668_, _27666_);
  and (_27670_, _08649_, _06606_);
  nor (_27671_, _27670_, _12995_);
  and (_27673_, _27671_, _27669_);
  nor (_27674_, _27350_, _12994_);
  or (_27675_, _27674_, _27673_);
  nand (_27676_, _27675_, _07312_);
  and (_27677_, _08590_, _07887_);
  nor (_27678_, _27677_, _06234_);
  nand (_27679_, _27678_, _27676_);
  and (_27680_, _27663_, _06234_);
  nor (_27681_, _27680_, _13012_);
  nand (_27682_, _27681_, _27679_);
  nor (_27684_, _27350_, _13011_);
  nor (_27685_, _27684_, _06195_);
  and (_27686_, _27685_, _27682_);
  or (_27687_, _27686_, _27352_);
  nand (_27688_, _27687_, _13019_);
  nor (_27689_, _27356_, _13019_);
  nor (_27690_, _27689_, _24972_);
  nand (_27691_, _27690_, _27688_);
  and (_27692_, _24972_, _08590_);
  nor (_27693_, _27692_, _13030_);
  and (_27695_, _27693_, _27691_);
  or (_27696_, _27695_, _27351_);
  or (_27697_, _27696_, _01379_);
  or (_27698_, _01375_, \uc8051golden_1.PC [7]);
  and (_27699_, _27698_, _42545_);
  and (_42984_, _27699_, _27697_);
  nor (_27700_, _06840_, _13023_);
  nor (_27701_, _06840_, _09463_);
  nor (_27702_, _12097_, \uc8051golden_1.PC [8]);
  nor (_27703_, _27702_, _12098_);
  and (_27705_, _27703_, _11243_);
  nor (_27706_, _27703_, _12108_);
  and (_27707_, _27703_, _11089_);
  nor (_27708_, _27703_, _12761_);
  not (_27709_, _27703_);
  and (_27710_, _27709_, _12224_);
  nor (_27711_, _27703_, _12719_);
  and (_27712_, _12341_, _06474_);
  nor (_27713_, _27703_, _12233_);
  nor (_27714_, _12188_, _09012_);
  nor (_27716_, _12624_, _05936_);
  nor (_27717_, _12569_, _12188_);
  and (_27718_, _12346_, _12339_);
  nor (_27719_, _27718_, _12347_);
  and (_27720_, _27719_, _12407_);
  and (_27721_, _12405_, _12341_);
  nor (_27722_, _27721_, _27720_);
  nor (_27723_, _27722_, _12411_);
  and (_27724_, _12188_, _06393_);
  nor (_27725_, _06399_, _07351_);
  and (_27727_, _12188_, _06395_);
  not (_27728_, _27719_);
  and (_27729_, _27728_, _12464_);
  and (_27730_, _12466_, _12342_);
  nor (_27731_, _27730_, _27729_);
  or (_27732_, _27731_, _07210_);
  and (_27733_, _12476_, _12188_);
  nor (_27734_, _12191_, _12186_);
  nor (_27735_, _27734_, _12192_);
  and (_27736_, _27735_, _12474_);
  nor (_27738_, _27736_, _27733_);
  nand (_27739_, _27738_, _08643_);
  or (_27740_, _12481_, _07332_);
  and (_27741_, _27740_, _27709_);
  and (_27742_, _14497_, _07199_);
  or (_27743_, _27742_, _06854_);
  or (_27744_, _07199_, \uc8051golden_1.PC [8]);
  nor (_27745_, _27744_, _07332_);
  or (_27746_, _27745_, _27743_);
  and (_27747_, _27746_, _25019_);
  or (_27749_, _27747_, _27741_);
  nand (_27750_, _27703_, _06854_);
  and (_27751_, _27750_, _08644_);
  and (_27752_, _27751_, _27749_);
  nor (_27753_, _27752_, _07212_);
  and (_27754_, _27753_, _27739_);
  and (_27755_, _27703_, _07212_);
  or (_27756_, _27755_, _06401_);
  or (_27757_, _27756_, _27754_);
  nand (_27758_, _27757_, _27732_);
  nand (_27760_, _27758_, _12458_);
  nor (_27761_, _27703_, _12458_);
  nor (_27762_, _27761_, _06395_);
  and (_27763_, _27762_, _27760_);
  or (_27764_, _27763_, _27727_);
  nand (_27765_, _27764_, _27725_);
  and (_27766_, _12188_, _06399_);
  nor (_27767_, _27766_, _12510_);
  nand (_27768_, _27767_, _27765_);
  nor (_27769_, _27703_, _12509_);
  nor (_27771_, _27769_, _06406_);
  nand (_27772_, _27771_, _27768_);
  and (_27773_, _12188_, _06406_);
  nor (_27774_, _27773_, _12519_);
  nand (_27775_, _27774_, _27772_);
  nor (_27776_, _27703_, _12517_);
  nor (_27777_, _27776_, _06393_);
  and (_27778_, _27777_, _27775_);
  or (_27779_, _27778_, _27724_);
  nand (_27780_, _27779_, _12522_);
  and (_27782_, _12188_, _06419_);
  nor (_27783_, _27782_, _12450_);
  nand (_27784_, _27783_, _27780_);
  and (_27785_, _12444_, _12341_);
  nor (_27786_, _27728_, _12444_);
  or (_27787_, _27786_, _27785_);
  nor (_27788_, _27787_, _12449_);
  nor (_27789_, _27788_, _06457_);
  nand (_27790_, _27789_, _27784_);
  nand (_27791_, _27790_, _06842_);
  or (_27793_, _27791_, _27723_);
  and (_27794_, _12546_, _12341_);
  not (_27795_, _27794_);
  nor (_27796_, _27728_, _12546_);
  nor (_27797_, _27796_, _06842_);
  and (_27798_, _27797_, _27795_);
  nor (_27799_, _27798_, _06482_);
  nand (_27800_, _27799_, _27793_);
  and (_27801_, _12341_, _12249_);
  and (_27802_, _27719_, _26421_);
  or (_27804_, _27802_, _27801_);
  and (_27805_, _27804_, _06482_);
  nor (_27806_, _27805_, _12237_);
  nand (_27807_, _27806_, _27800_);
  and (_27808_, _27709_, _12237_);
  nor (_27809_, _27808_, _06387_);
  nand (_27810_, _27809_, _27807_);
  and (_27811_, _12569_, _05994_);
  and (_27812_, _12188_, _06387_);
  not (_27813_, _27812_);
  and (_27815_, _27813_, _27811_);
  and (_27816_, _27815_, _27810_);
  or (_27817_, _27816_, _27717_);
  nand (_27818_, _27817_, _12576_);
  nor (_27819_, _27703_, _12576_);
  nor (_27820_, _27819_, _06433_);
  nand (_27821_, _27820_, _27818_);
  and (_27822_, _12188_, _06433_);
  nor (_27823_, _27822_, _25090_);
  nand (_27824_, _27823_, _27821_);
  nand (_27826_, _27824_, _14015_);
  and (_27827_, _12188_, _06432_);
  nor (_27828_, _27827_, _12594_);
  and (_27829_, _27828_, _27826_);
  nor (_27830_, _27703_, _12588_);
  or (_27831_, _27830_, _27829_);
  nand (_27832_, _27831_, _12592_);
  nor (_27833_, _12188_, _12592_);
  nor (_27834_, _27833_, _06022_);
  nand (_27835_, _27834_, _27832_);
  and (_27837_, _27703_, _06022_);
  nor (_27838_, _27837_, _06300_);
  nand (_27839_, _27838_, _27835_);
  nor (_27840_, _06472_, _06017_);
  not (_27841_, _27840_);
  and (_27842_, _14497_, _06300_);
  nor (_27843_, _27842_, _27841_);
  nand (_27844_, _27843_, _27839_);
  and (_27845_, _12341_, _06472_);
  nor (_27846_, _27845_, _13788_);
  nand (_27848_, _27846_, _27844_);
  nor (_27849_, _12188_, _06294_);
  nor (_27850_, _27849_, _06015_);
  nand (_27851_, _27850_, _27848_);
  and (_27852_, _12341_, _06015_);
  nor (_27853_, _27852_, _12620_);
  nand (_27854_, _27853_, _27851_);
  nor (_27855_, _27703_, _12616_);
  nor (_27856_, _27855_, _06376_);
  and (_27857_, _27856_, _27854_);
  and (_27859_, _12188_, _06376_);
  or (_27860_, _27859_, _27857_);
  nand (_27861_, _27860_, _27716_);
  and (_27862_, _27735_, _12624_);
  nor (_27863_, _27862_, _09013_);
  and (_27864_, _27863_, _27861_);
  or (_27865_, _27864_, _27714_);
  nand (_27866_, _27865_, _06276_);
  and (_27867_, _12342_, _06275_);
  nor (_27868_, _27867_, _10933_);
  nand (_27869_, _27868_, _27866_);
  and (_27870_, _12188_, _10933_);
  nor (_27871_, _27870_, _12639_);
  nand (_27872_, _27871_, _27869_);
  and (_27873_, _12663_, _12642_);
  nor (_27874_, _27873_, _12664_);
  nor (_27875_, _27874_, _12640_);
  nor (_27876_, _27875_, _06375_);
  nand (_27877_, _27876_, _27872_);
  and (_27878_, _12188_, _06375_);
  nor (_27881_, _27878_, _05943_);
  nand (_27882_, _27881_, _27877_);
  nand (_27883_, _27882_, _12681_);
  and (_27884_, _12188_, _11297_);
  and (_27885_, _27735_, _12687_);
  or (_27886_, _27885_, _27884_);
  and (_27887_, _27886_, _12680_);
  nor (_27888_, _27887_, _12685_);
  and (_27889_, _27888_, _27883_);
  or (_27890_, _27889_, _27713_);
  nand (_27892_, _27890_, _12227_);
  nor (_27893_, _12188_, _12227_);
  nor (_27894_, _27893_, _06474_);
  and (_27895_, _27894_, _27892_);
  or (_27896_, _27895_, _27712_);
  nand (_27897_, _27896_, _07284_);
  and (_27898_, _12188_, _06582_);
  nor (_27899_, _27898_, _05952_);
  nand (_27900_, _27899_, _27897_);
  nand (_27901_, _27900_, _12705_);
  nor (_27903_, _14497_, _11297_);
  and (_27904_, _27735_, _11297_);
  or (_27905_, _27904_, _27903_);
  and (_27906_, _27905_, _12704_);
  nor (_27907_, _27906_, _12723_);
  and (_27908_, _27907_, _27901_);
  or (_27909_, _27908_, _27711_);
  nand (_27910_, _27909_, _12721_);
  nor (_27911_, _12188_, _12721_);
  nor (_27912_, _27911_, _06478_);
  nand (_27914_, _27912_, _27910_);
  and (_27915_, _12341_, _06478_);
  nor (_27916_, _27915_, _06569_);
  nand (_27917_, _27916_, _27914_);
  nor (_27918_, _12735_, _05956_);
  not (_27919_, _27918_);
  and (_27920_, _14497_, _06569_);
  nor (_27921_, _27920_, _27919_);
  nand (_27922_, _27921_, _27917_);
  nor (_27923_, _27735_, \uc8051golden_1.PSW [7]);
  nor (_27925_, _12188_, _10524_);
  nor (_27926_, _27925_, _12736_);
  not (_27927_, _27926_);
  nor (_27928_, _27927_, _27923_);
  nor (_27929_, _27928_, _12224_);
  and (_27930_, _27929_, _27922_);
  or (_27931_, _27930_, _27710_);
  nand (_27932_, _27931_, _11018_);
  nor (_27933_, _12188_, _11018_);
  nor (_27934_, _27933_, _06479_);
  nand (_27936_, _27934_, _27932_);
  and (_27937_, _12341_, _06479_);
  nor (_27938_, _27937_, _06572_);
  nand (_27939_, _27938_, _27936_);
  nor (_27940_, _12217_, _05947_);
  not (_27941_, _27940_);
  and (_27942_, _14497_, _06572_);
  nor (_27943_, _27942_, _27941_);
  nand (_27944_, _27943_, _27939_);
  and (_27945_, _12188_, _10524_);
  and (_27947_, _27735_, \uc8051golden_1.PSW [7]);
  or (_27948_, _27947_, _27945_);
  and (_27949_, _27948_, _12217_);
  nor (_27950_, _27949_, _12763_);
  and (_27951_, _27950_, _27944_);
  or (_27952_, _27951_, _27708_);
  nand (_27953_, _27952_, _11060_);
  nor (_27954_, _12188_, _11060_);
  nor (_27955_, _27954_, _11089_);
  and (_27956_, _27955_, _27953_);
  or (_27958_, _27956_, _27707_);
  nand (_27959_, _27958_, _13881_);
  and (_27960_, _07473_, _06588_);
  nor (_27961_, _27960_, _05966_);
  nand (_27962_, _27961_, _27959_);
  nand (_27963_, _27962_, _06596_);
  nor (_27964_, _12341_, _12958_);
  and (_27965_, _27728_, _12958_);
  or (_27966_, _27965_, _06596_);
  or (_27967_, _27966_, _27964_);
  and (_27969_, _27967_, _12108_);
  and (_27970_, _27969_, _27963_);
  or (_27971_, _27970_, _27706_);
  nand (_27972_, _27971_, _11204_);
  nor (_27973_, _12188_, _11204_);
  nor (_27974_, _27973_, _11243_);
  and (_27975_, _27974_, _27972_);
  or (_27976_, _27975_, _27705_);
  nand (_27977_, _27976_, _06306_);
  and (_27978_, _07473_, _06305_);
  nor (_27980_, _27978_, _05971_);
  nand (_27981_, _27980_, _27977_);
  nand (_27982_, _27981_, _12978_);
  nor (_27983_, _27719_, _12958_);
  and (_27984_, _12342_, _12958_);
  nor (_27985_, _27984_, _27983_);
  and (_27986_, _27985_, _06487_);
  nor (_27987_, _27986_, _12988_);
  nand (_27988_, _27987_, _27982_);
  nor (_27989_, _27703_, _12987_);
  nor (_27991_, _27989_, _06606_);
  nand (_27992_, _27991_, _27988_);
  and (_27993_, _12188_, _06606_);
  nor (_27994_, _27993_, _12995_);
  nand (_27995_, _27994_, _27992_);
  nor (_27996_, _27703_, _12994_);
  nor (_27997_, _27996_, _06465_);
  and (_27998_, _27997_, _27995_);
  or (_27999_, _27998_, _27701_);
  nor (_28000_, _06234_, _05969_);
  nand (_28002_, _28000_, _27999_);
  and (_28003_, _27985_, _06234_);
  nor (_28004_, _28003_, _13012_);
  nand (_28005_, _28004_, _28002_);
  nor (_28006_, _27703_, _13011_);
  nor (_28007_, _28006_, _06195_);
  nand (_28008_, _28007_, _28005_);
  and (_28009_, _12188_, _06195_);
  nor (_28010_, _28009_, _13020_);
  nand (_28011_, _28010_, _28008_);
  nor (_28013_, _27703_, _13019_);
  nor (_28014_, _28013_, _06475_);
  and (_28015_, _28014_, _28011_);
  or (_28016_, _28015_, _27700_);
  nor (_28017_, _13030_, _05963_);
  and (_28018_, _28017_, _28016_);
  and (_28019_, _27703_, _13030_);
  or (_28020_, _28019_, _28018_);
  or (_28021_, _28020_, _01379_);
  or (_28022_, _01375_, \uc8051golden_1.PC [8]);
  and (_28024_, _28022_, _42545_);
  and (_42985_, _28024_, _28021_);
  nor (_28025_, _13023_, _06228_);
  nor (_28026_, _09463_, _06228_);
  nor (_28027_, _12098_, \uc8051golden_1.PC [9]);
  nor (_28028_, _28027_, _12099_);
  nor (_28029_, _28028_, _12108_);
  nor (_28030_, _28028_, _12761_);
  and (_28031_, _12281_, _06479_);
  not (_28032_, _28028_);
  and (_28034_, _28032_, _12224_);
  and (_28035_, _12281_, _06478_);
  nor (_28036_, _28028_, _12719_);
  and (_28037_, _12281_, _06474_);
  nor (_28038_, _28028_, _12233_);
  nor (_28039_, _12136_, _09012_);
  and (_28040_, _12136_, _06376_);
  and (_28041_, _12136_, _06432_);
  nor (_28042_, _28028_, _12576_);
  and (_28043_, _28032_, _12237_);
  nor (_28045_, _12347_, _12343_);
  and (_28046_, _28045_, _12285_);
  nor (_28047_, _28045_, _12285_);
  nor (_28048_, _28047_, _28046_);
  and (_28049_, _28048_, _12407_);
  and (_28050_, _12405_, _12282_);
  nor (_28051_, _28050_, _28049_);
  nor (_28052_, _28051_, _12411_);
  and (_28053_, _28028_, _06854_);
  nand (_28054_, _28032_, _27740_);
  and (_28056_, _14726_, _07199_);
  nor (_28057_, _28056_, _06854_);
  or (_28058_, _07199_, \uc8051golden_1.PC [9]);
  or (_28059_, _28058_, _07332_);
  nand (_28060_, _28059_, _28057_);
  nand (_28061_, _28060_, _25019_);
  and (_28062_, _28061_, _28054_);
  or (_28063_, _28062_, _08643_);
  nor (_28064_, _28063_, _28053_);
  and (_28065_, _12476_, _12136_);
  nor (_28067_, _12192_, _12189_);
  and (_28068_, _28067_, _12139_);
  nor (_28069_, _28067_, _12139_);
  nor (_28070_, _28069_, _28068_);
  nor (_28071_, _28070_, _12476_);
  nor (_28072_, _28071_, _28065_);
  and (_28073_, _28072_, _08643_);
  or (_28074_, _28073_, _28064_);
  nand (_28075_, _28074_, _08659_);
  and (_28076_, _28032_, _07212_);
  nor (_28078_, _28076_, _06401_);
  and (_28079_, _28078_, _28075_);
  or (_28080_, _12464_, _12281_);
  not (_28081_, _28048_);
  or (_28082_, _28081_, _12466_);
  and (_28083_, _28082_, _06401_);
  and (_28084_, _28083_, _28080_);
  or (_28085_, _28084_, _25041_);
  or (_28086_, _28085_, _28079_);
  nor (_28087_, _28028_, _12458_);
  nor (_28089_, _28087_, _06395_);
  nand (_28090_, _28089_, _28086_);
  and (_28091_, _12136_, _06395_);
  nor (_28092_, _28091_, _07351_);
  nand (_28093_, _28092_, _28090_);
  nand (_28094_, _28093_, _07221_);
  and (_28095_, _12136_, _06399_);
  nor (_28096_, _28095_, _12510_);
  nand (_28097_, _28096_, _28094_);
  nor (_28098_, _28028_, _12509_);
  nor (_28100_, _28098_, _06406_);
  nand (_28101_, _28100_, _28097_);
  and (_28102_, _12136_, _06406_);
  nor (_28103_, _28102_, _12519_);
  nand (_28104_, _28103_, _28101_);
  nor (_28105_, _28028_, _12517_);
  nor (_28106_, _28105_, _06393_);
  nand (_28107_, _28106_, _28104_);
  and (_28108_, _12136_, _06393_);
  nor (_28109_, _28108_, _12521_);
  nand (_28111_, _28109_, _28107_);
  nand (_28112_, _28111_, _07785_);
  and (_28113_, _12136_, _06419_);
  nor (_28114_, _28113_, _12450_);
  and (_28115_, _28114_, _28112_);
  and (_28116_, _12444_, _12281_);
  nor (_28117_, _28048_, _12444_);
  or (_28118_, _28117_, _12449_);
  nor (_28119_, _28118_, _28116_);
  or (_28120_, _28119_, _28115_);
  and (_28122_, _28120_, _12411_);
  or (_28123_, _28122_, _28052_);
  or (_28124_, _28123_, _06420_);
  and (_28125_, _12546_, _12281_);
  nor (_28126_, _28048_, _12546_);
  nor (_28127_, _28126_, _28125_);
  or (_28128_, _28127_, _06842_);
  and (_28129_, _28128_, _28124_);
  or (_28130_, _28129_, _06482_);
  and (_28131_, _12281_, _12249_);
  nor (_28133_, _28048_, _12249_);
  or (_28134_, _28133_, _28131_);
  and (_28135_, _28134_, _06482_);
  nor (_28136_, _28135_, _12237_);
  and (_28137_, _28136_, _28130_);
  or (_28138_, _28137_, _28043_);
  nand (_28139_, _28138_, _07245_);
  and (_28140_, _14726_, _06387_);
  not (_28141_, _28140_);
  and (_28142_, _28141_, _27811_);
  nand (_28144_, _28142_, _28139_);
  nor (_28145_, _12569_, _14726_);
  nor (_28146_, _28145_, _12580_);
  and (_28147_, _28146_, _28144_);
  nor (_28148_, _28147_, _28042_);
  or (_28149_, _28148_, _06433_);
  nor (_28150_, _06432_, _25090_);
  nand (_28151_, _14726_, _06433_);
  and (_28152_, _28151_, _28150_);
  and (_28153_, _28152_, _28149_);
  or (_28155_, _28153_, _28041_);
  nand (_28156_, _28155_, _12588_);
  nor (_28157_, _28032_, _12588_);
  nor (_28158_, _28157_, _12593_);
  nand (_28159_, _28158_, _28156_);
  nor (_28160_, _12136_, _12592_);
  nor (_28161_, _28160_, _06022_);
  nand (_28162_, _28161_, _28159_);
  and (_28163_, _28028_, _06022_);
  nor (_28164_, _28163_, _06300_);
  nand (_28166_, _28164_, _28162_);
  and (_28167_, _14726_, _06300_);
  nor (_28168_, _28167_, _27841_);
  nand (_28169_, _28168_, _28166_);
  and (_28170_, _12281_, _06472_);
  nor (_28171_, _28170_, _13788_);
  nand (_28172_, _28171_, _28169_);
  nor (_28173_, _12136_, _06294_);
  nor (_28174_, _28173_, _06015_);
  nand (_28175_, _28174_, _28172_);
  and (_28176_, _12281_, _06015_);
  nor (_28177_, _28176_, _12620_);
  nand (_28178_, _28177_, _28175_);
  nor (_28179_, _28028_, _12616_);
  nor (_28180_, _28179_, _06376_);
  and (_28181_, _28180_, _28178_);
  or (_28182_, _28181_, _28040_);
  nand (_28183_, _28182_, _27716_);
  nor (_28184_, _28070_, _12625_);
  nor (_28185_, _28184_, _09013_);
  and (_28188_, _28185_, _28183_);
  or (_28189_, _28188_, _28039_);
  nand (_28190_, _28189_, _06276_);
  and (_28191_, _12282_, _06275_);
  nor (_28192_, _28191_, _10933_);
  nand (_28193_, _28192_, _28190_);
  and (_28194_, _12136_, _10933_);
  nor (_28195_, _28194_, _12639_);
  nand (_28196_, _28195_, _28193_);
  nor (_28197_, _12664_, \uc8051golden_1.DPH [1]);
  nor (_28199_, _28197_, _12665_);
  nor (_28200_, _28199_, _12640_);
  nor (_28201_, _28200_, _06375_);
  nand (_28202_, _28201_, _28196_);
  and (_28203_, _12136_, _06375_);
  nor (_28204_, _28203_, _05943_);
  nand (_28205_, _28204_, _28202_);
  nand (_28206_, _28205_, _12681_);
  and (_28207_, _12136_, _11297_);
  nor (_28208_, _28070_, _11297_);
  or (_28210_, _28208_, _28207_);
  and (_28211_, _28210_, _12680_);
  nor (_28212_, _28211_, _12685_);
  and (_28213_, _28212_, _28206_);
  or (_28214_, _28213_, _28038_);
  nand (_28215_, _28214_, _12227_);
  nor (_28216_, _12136_, _12227_);
  nor (_28217_, _28216_, _06474_);
  and (_28218_, _28217_, _28215_);
  or (_28219_, _28218_, _28037_);
  nand (_28221_, _28219_, _07284_);
  and (_28222_, _12136_, _06582_);
  nor (_28223_, _28222_, _05952_);
  nand (_28224_, _28223_, _28221_);
  nand (_28225_, _28224_, _12705_);
  and (_28226_, _28070_, _11297_);
  nor (_28227_, _12136_, _11297_);
  nor (_28228_, _28227_, _12705_);
  not (_28229_, _28228_);
  nor (_28230_, _28229_, _28226_);
  nor (_28232_, _28230_, _12723_);
  and (_28233_, _28232_, _28225_);
  or (_28234_, _28233_, _28036_);
  nand (_28235_, _28234_, _12721_);
  nor (_28236_, _12136_, _12721_);
  nor (_28237_, _28236_, _06478_);
  and (_28238_, _28237_, _28235_);
  or (_28239_, _28238_, _28035_);
  nand (_28240_, _28239_, _07276_);
  and (_28241_, _12136_, _06569_);
  nor (_28243_, _28241_, _05956_);
  nand (_28244_, _28243_, _28240_);
  nand (_28245_, _28244_, _12736_);
  and (_28246_, _12136_, \uc8051golden_1.PSW [7]);
  nor (_28247_, _28070_, \uc8051golden_1.PSW [7]);
  or (_28248_, _28247_, _28246_);
  and (_28249_, _28248_, _12735_);
  nor (_28250_, _28249_, _12224_);
  and (_28251_, _28250_, _28245_);
  or (_28252_, _28251_, _28034_);
  nand (_28254_, _28252_, _11018_);
  nor (_28255_, _12136_, _11018_);
  nor (_28256_, _28255_, _06479_);
  and (_28257_, _28256_, _28254_);
  or (_28258_, _28257_, _28031_);
  nand (_28259_, _28258_, _09048_);
  and (_28260_, _12136_, _06572_);
  nor (_28261_, _28260_, _05947_);
  nand (_28262_, _28261_, _28259_);
  nand (_28263_, _28262_, _12756_);
  and (_28265_, _12136_, _10524_);
  nor (_28266_, _28070_, _10524_);
  or (_28267_, _28266_, _28265_);
  and (_28268_, _28267_, _12217_);
  nor (_28269_, _28268_, _12763_);
  and (_28270_, _28269_, _28263_);
  or (_28271_, _28270_, _28030_);
  nand (_28272_, _28271_, _11060_);
  nor (_28273_, _12136_, _11060_);
  nor (_28274_, _28273_, _11089_);
  nand (_28276_, _28274_, _28272_);
  and (_28277_, _28028_, _11089_);
  nor (_28278_, _28277_, _06588_);
  nand (_28279_, _28278_, _28276_);
  nor (_28280_, _06460_, _05966_);
  not (_28281_, _28280_);
  and (_28282_, _07196_, _06588_);
  nor (_28283_, _28282_, _28281_);
  nand (_28284_, _28283_, _28279_);
  and (_28285_, _28048_, _12958_);
  nor (_28287_, _12281_, _12958_);
  or (_28288_, _28287_, _06596_);
  or (_28289_, _28288_, _28285_);
  and (_28290_, _28289_, _12108_);
  and (_28291_, _28290_, _28284_);
  or (_28292_, _28291_, _28029_);
  nand (_28293_, _28292_, _11204_);
  nor (_28294_, _12136_, _11204_);
  nor (_28295_, _28294_, _11243_);
  nand (_28296_, _28295_, _28293_);
  and (_28298_, _28028_, _11243_);
  nor (_28299_, _28298_, _06305_);
  nand (_28300_, _28299_, _28296_);
  nor (_28301_, _06487_, _05971_);
  not (_28302_, _28301_);
  and (_28303_, _07196_, _06305_);
  nor (_28304_, _28303_, _28302_);
  nand (_28305_, _28304_, _28300_);
  and (_28306_, _12282_, _12958_);
  nor (_28307_, _28081_, _12958_);
  nor (_28309_, _28307_, _28306_);
  and (_28310_, _28309_, _06487_);
  nor (_28311_, _28310_, _12988_);
  nand (_28312_, _28311_, _28305_);
  nor (_28313_, _28028_, _12987_);
  nor (_28314_, _28313_, _06606_);
  nand (_28315_, _28314_, _28312_);
  and (_28316_, _12136_, _06606_);
  nor (_28317_, _28316_, _12995_);
  nand (_28318_, _28317_, _28315_);
  nor (_28320_, _28028_, _12994_);
  nor (_28321_, _28320_, _06465_);
  and (_28322_, _28321_, _28318_);
  or (_28323_, _28322_, _28026_);
  nand (_28324_, _28323_, _28000_);
  and (_28325_, _28309_, _06234_);
  nor (_28326_, _28325_, _13012_);
  nand (_28327_, _28326_, _28324_);
  nor (_28328_, _28028_, _13011_);
  nor (_28329_, _28328_, _06195_);
  nand (_28331_, _28329_, _28327_);
  and (_28332_, _12136_, _06195_);
  nor (_28333_, _28332_, _13020_);
  nand (_28334_, _28333_, _28331_);
  nor (_28335_, _28028_, _13019_);
  nor (_28336_, _28335_, _06475_);
  and (_28337_, _28336_, _28334_);
  or (_28338_, _28337_, _28025_);
  and (_28339_, _28338_, _28017_);
  and (_28340_, _28028_, _13030_);
  or (_28342_, _28340_, _28339_);
  or (_28343_, _28342_, _01379_);
  or (_28344_, _01375_, \uc8051golden_1.PC [9]);
  and (_28345_, _28344_, _42545_);
  and (_42986_, _28345_, _28343_);
  and (_28346_, _06693_, _06465_);
  nor (_28347_, _12680_, _05943_);
  nor (_28348_, _12569_, _12124_);
  nor (_28349_, _12099_, \uc8051golden_1.PC [10]);
  nor (_28350_, _28349_, _12100_);
  nor (_28352_, _28350_, _12509_);
  not (_28353_, _12278_);
  nor (_28354_, _12351_, _12348_);
  nor (_28355_, _28354_, _28353_);
  and (_28356_, _28354_, _28353_);
  nor (_28357_, _28356_, _28355_);
  or (_28358_, _28357_, _12466_);
  or (_28359_, _12464_, _12274_);
  and (_28360_, _28359_, _28358_);
  or (_28361_, _28360_, _07210_);
  not (_28363_, _12133_);
  nor (_28364_, _12196_, _12193_);
  nor (_28365_, _28364_, _28363_);
  and (_28366_, _28364_, _28363_);
  nor (_28367_, _28366_, _28365_);
  or (_28368_, _28367_, _12476_);
  or (_28369_, _12474_, _12124_);
  nand (_28370_, _28369_, _28368_);
  nand (_28371_, _28370_, _08643_);
  nand (_28372_, _12124_, _07199_);
  nand (_28374_, _07200_, \uc8051golden_1.PC [10]);
  or (_28375_, _28374_, _07332_);
  and (_28376_, _28375_, _28372_);
  or (_28377_, _28376_, _06854_);
  and (_28378_, _28377_, _07366_);
  or (_28379_, _28378_, _12481_);
  not (_28380_, _28350_);
  or (_28381_, _28380_, _12493_);
  and (_28382_, _28381_, _08644_);
  and (_28383_, _28382_, _28379_);
  nor (_28385_, _28383_, _07212_);
  and (_28386_, _28385_, _28371_);
  and (_28387_, _28350_, _07212_);
  or (_28388_, _28387_, _06401_);
  or (_28389_, _28388_, _28386_);
  nand (_28390_, _28389_, _28361_);
  nand (_28391_, _28390_, _12458_);
  nor (_28392_, _28350_, _12458_);
  nor (_28393_, _28392_, _06395_);
  nand (_28394_, _28393_, _28391_);
  nand (_28396_, _28394_, _05997_);
  nand (_28397_, _28396_, _07221_);
  nor (_28398_, _14927_, _06407_);
  nor (_28399_, _28398_, _12510_);
  and (_28400_, _28399_, _28397_);
  or (_28401_, _28400_, _28352_);
  nand (_28402_, _28401_, _06414_);
  and (_28403_, _14927_, _06406_);
  nor (_28404_, _28403_, _12519_);
  and (_28405_, _28404_, _28402_);
  nor (_28407_, _28380_, _12517_);
  or (_28408_, _28407_, _28405_);
  nand (_28409_, _28408_, _06844_);
  and (_28410_, _12124_, _06393_);
  nor (_28411_, _28410_, _12521_);
  nand (_28412_, _28411_, _28409_);
  nand (_28413_, _28412_, _07785_);
  and (_28414_, _12124_, _06419_);
  nor (_28415_, _28414_, _12450_);
  and (_28416_, _28415_, _28413_);
  and (_28418_, _12444_, _12274_);
  not (_28419_, _28357_);
  nor (_28420_, _28419_, _12444_);
  or (_28421_, _28420_, _28418_);
  nor (_28422_, _28421_, _12449_);
  or (_28423_, _28422_, _28416_);
  nand (_28424_, _28423_, _12411_);
  and (_28425_, _12405_, _12274_);
  and (_28426_, _28357_, _12407_);
  or (_28427_, _28426_, _28425_);
  nor (_28429_, _28427_, _12411_);
  nor (_28430_, _28429_, _06420_);
  nand (_28431_, _28430_, _28424_);
  and (_28432_, _12546_, _12275_);
  nor (_28433_, _28357_, _12546_);
  or (_28434_, _28433_, _06842_);
  or (_28435_, _28434_, _28432_);
  nand (_28436_, _28435_, _28431_);
  nand (_28437_, _28436_, _12534_);
  nand (_28438_, _12274_, _12249_);
  nand (_28440_, _28357_, _26421_);
  and (_28441_, _28440_, _28438_);
  or (_28442_, _28441_, _12534_);
  and (_28443_, _28442_, _28437_);
  or (_28444_, _28443_, _12237_);
  nand (_28445_, _28350_, _12237_);
  and (_28446_, _28445_, _28444_);
  nor (_28447_, _28446_, _06387_);
  and (_28448_, _12124_, _06387_);
  nor (_28449_, _28448_, _28447_);
  and (_28451_, _28449_, _27811_);
  or (_28452_, _28451_, _28348_);
  nand (_28453_, _28452_, _12576_);
  nor (_28454_, _28350_, _12576_);
  nor (_28455_, _28454_, _06433_);
  nand (_28456_, _28455_, _28453_);
  nand (_28457_, _28456_, _06007_);
  nand (_28458_, _28457_, _14015_);
  nor (_28459_, _14927_, _06434_);
  nor (_28460_, _28459_, _12594_);
  nand (_28462_, _28460_, _28458_);
  nor (_28463_, _28350_, _12588_);
  nor (_28464_, _28463_, _12593_);
  nand (_28465_, _28464_, _28462_);
  nor (_28466_, _14927_, _12592_);
  nor (_28467_, _28466_, _06022_);
  nand (_28468_, _28467_, _28465_);
  and (_28469_, _28380_, _06022_);
  nor (_28470_, _28469_, _06300_);
  and (_28471_, _28470_, _28468_);
  and (_28473_, _12124_, _06300_);
  nor (_28474_, _28473_, _28471_);
  and (_28475_, _28474_, _27840_);
  and (_28476_, _12275_, _06472_);
  or (_28477_, _28476_, _28475_);
  and (_28478_, _28477_, _06294_);
  nor (_28479_, _12124_, _06294_);
  or (_28480_, _28479_, _28478_);
  nand (_28481_, _28480_, _06279_);
  and (_28482_, _12275_, _06015_);
  nor (_28484_, _28482_, _12620_);
  and (_28485_, _28484_, _28481_);
  nor (_28486_, _28380_, _12616_);
  nor (_28487_, _28486_, _28485_);
  or (_28488_, _28487_, _06376_);
  and (_28489_, _12124_, _06376_);
  not (_28490_, _28489_);
  and (_28491_, _28490_, _27716_);
  nand (_28492_, _28491_, _28488_);
  nor (_28493_, _28367_, _12625_);
  nor (_28495_, _28493_, _09013_);
  and (_28496_, _28495_, _28492_);
  nor (_28497_, _14927_, _09012_);
  or (_28498_, _28497_, _06275_);
  or (_28499_, _28498_, _28496_);
  and (_28500_, _12275_, _06275_);
  nor (_28501_, _28500_, _10933_);
  nand (_28502_, _28501_, _28499_);
  and (_28503_, _12124_, _10933_);
  nor (_28504_, _28503_, _12639_);
  nand (_28506_, _28504_, _28502_);
  nor (_28507_, _12665_, \uc8051golden_1.DPH [2]);
  nor (_28508_, _28507_, _12666_);
  nor (_28509_, _28508_, _12640_);
  nor (_28510_, _28509_, _06375_);
  and (_28511_, _28510_, _28506_);
  and (_28512_, _12124_, _06375_);
  or (_28513_, _28512_, _28511_);
  nand (_28514_, _28513_, _28347_);
  and (_28515_, _12124_, _11297_);
  and (_28517_, _28367_, _12687_);
  or (_28518_, _28517_, _28515_);
  and (_28519_, _28518_, _12680_);
  nor (_28520_, _28519_, _12685_);
  nand (_28521_, _28520_, _28514_);
  nor (_28522_, _28350_, _12233_);
  nor (_28523_, _28522_, _12228_);
  nand (_28524_, _28523_, _28521_);
  nor (_28525_, _14927_, _12227_);
  nor (_28526_, _28525_, _06474_);
  and (_28527_, _28526_, _28524_);
  and (_28528_, _12275_, _06474_);
  or (_28529_, _28528_, _28527_);
  or (_28530_, _28529_, _06582_);
  nand (_28531_, _12124_, _06582_);
  and (_28532_, _28531_, _28530_);
  or (_28533_, _28532_, _05952_);
  or (_28534_, _28533_, _12704_);
  and (_28535_, _12124_, _12687_);
  and (_28536_, _28367_, _11297_);
  or (_28539_, _28536_, _28535_);
  and (_28540_, _28539_, _12704_);
  nor (_28541_, _28540_, _12723_);
  nand (_28542_, _28541_, _28534_);
  nor (_28543_, _28350_, _12719_);
  nor (_28544_, _28543_, _12722_);
  nand (_28545_, _28544_, _28542_);
  nor (_28546_, _14927_, _12721_);
  nor (_28547_, _28546_, _06478_);
  and (_28548_, _28547_, _28545_);
  and (_28550_, _12275_, _06478_);
  or (_28551_, _28550_, _28548_);
  nand (_28552_, _28551_, _07276_);
  and (_28553_, _14927_, _06569_);
  nor (_28554_, _28553_, _27919_);
  nand (_28555_, _28554_, _28552_);
  nor (_28556_, _28367_, \uc8051golden_1.PSW [7]);
  nor (_28557_, _12124_, _10524_);
  nor (_28558_, _28557_, _12736_);
  not (_28559_, _28558_);
  nor (_28561_, _28559_, _28556_);
  nor (_28562_, _28561_, _12224_);
  nand (_28563_, _28562_, _28555_);
  and (_28564_, _28380_, _12224_);
  nor (_28565_, _28564_, _11019_);
  nand (_28566_, _28565_, _28563_);
  nor (_28567_, _14927_, _11018_);
  nor (_28568_, _28567_, _06479_);
  and (_28569_, _28568_, _28566_);
  and (_28570_, _12275_, _06479_);
  or (_28572_, _28570_, _28569_);
  nand (_28573_, _28572_, _09048_);
  and (_28574_, _14927_, _06572_);
  nor (_28575_, _28574_, _27941_);
  nand (_28576_, _28575_, _28573_);
  and (_28577_, _12124_, _10524_);
  and (_28578_, _28367_, \uc8051golden_1.PSW [7]);
  or (_28579_, _28578_, _28577_);
  and (_28580_, _28579_, _12217_);
  nor (_28581_, _28580_, _12763_);
  nand (_28583_, _28581_, _28576_);
  nor (_28584_, _28350_, _12761_);
  nor (_28585_, _28584_, _11061_);
  nand (_28586_, _28585_, _28583_);
  nor (_28587_, _14927_, _11060_);
  nor (_28588_, _28587_, _11089_);
  and (_28589_, _28588_, _28586_);
  and (_28590_, _28380_, _11089_);
  or (_28591_, _28590_, _28589_);
  nand (_28592_, _28591_, _13881_);
  and (_28594_, _07623_, _06588_);
  nor (_28595_, _28594_, _28281_);
  nand (_28596_, _28595_, _28592_);
  and (_28597_, _28419_, _12958_);
  nor (_28598_, _12274_, _12958_);
  or (_28599_, _28598_, _06596_);
  or (_28600_, _28599_, _28597_);
  and (_28601_, _28600_, _12108_);
  nand (_28602_, _28601_, _28596_);
  nor (_28603_, _28350_, _12108_);
  nor (_28605_, _28603_, _12094_);
  nand (_28606_, _28605_, _28602_);
  nor (_28607_, _14927_, _11204_);
  nor (_28608_, _28607_, _11243_);
  and (_28609_, _28608_, _28606_);
  and (_28610_, _28380_, _11243_);
  or (_28611_, _28610_, _28609_);
  nand (_28612_, _28611_, _06306_);
  and (_28613_, _07623_, _06305_);
  nor (_28614_, _28613_, _28302_);
  nand (_28616_, _28614_, _28612_);
  nor (_28617_, _28357_, _12958_);
  and (_28618_, _12275_, _12958_);
  nor (_28619_, _28618_, _28617_);
  and (_28620_, _28619_, _06487_);
  nor (_28621_, _28620_, _12988_);
  and (_28622_, _28621_, _28616_);
  nor (_28623_, _28350_, _12987_);
  or (_28624_, _28623_, _28622_);
  nand (_28625_, _28624_, _07037_);
  and (_28627_, _14927_, _06606_);
  nor (_28628_, _28627_, _12995_);
  nand (_28629_, _28628_, _28625_);
  nor (_28630_, _28380_, _12994_);
  nor (_28631_, _28630_, _06465_);
  nand (_28632_, _28631_, _28629_);
  nand (_28633_, _28632_, _28000_);
  or (_28634_, _28633_, _28346_);
  and (_28635_, _28619_, _06234_);
  nor (_28636_, _28635_, _13012_);
  and (_28638_, _28636_, _28634_);
  nor (_28639_, _28350_, _13011_);
  or (_28640_, _28639_, _28638_);
  nand (_28641_, _28640_, _06196_);
  and (_28642_, _14927_, _06195_);
  nor (_28643_, _28642_, _13020_);
  nand (_28644_, _28643_, _28641_);
  nor (_28645_, _28380_, _13019_);
  nor (_28646_, _28645_, _06475_);
  nand (_28647_, _28646_, _28644_);
  not (_28649_, _28017_);
  and (_28650_, _06693_, _06475_);
  nor (_28651_, _28650_, _28649_);
  and (_28652_, _28651_, _28647_);
  and (_28653_, _28350_, _13030_);
  or (_28654_, _28653_, _28652_);
  or (_28655_, _28654_, _01379_);
  or (_28656_, _01375_, \uc8051golden_1.PC [10]);
  and (_28657_, _28656_, _42545_);
  and (_42987_, _28657_, _28655_);
  nor (_28659_, _12100_, \uc8051golden_1.PC [11]);
  nor (_28660_, _28659_, _12101_);
  or (_28661_, _28660_, _12108_);
  or (_28662_, _28660_, _12761_);
  or (_28663_, _28660_, _12225_);
  or (_28664_, _28660_, _12719_);
  or (_28665_, _28660_, _12233_);
  or (_28666_, _12128_, _09012_);
  and (_28667_, _12268_, _06015_);
  or (_28668_, _28660_, _12509_);
  or (_28670_, _28660_, _12503_);
  nor (_28671_, _28355_, _12276_);
  and (_28672_, _28671_, _12272_);
  nor (_28673_, _28671_, _12272_);
  or (_28674_, _28673_, _28672_);
  or (_28675_, _28674_, _12466_);
  or (_28676_, _12464_, _12268_);
  and (_28677_, _28676_, _28675_);
  or (_28678_, _28677_, _07210_);
  nor (_28679_, _28365_, _12125_);
  nor (_28681_, _28679_, _12131_);
  and (_28682_, _28679_, _12131_);
  or (_28683_, _28682_, _28681_);
  or (_28684_, _28683_, _12476_);
  or (_28685_, _12474_, _12128_);
  and (_28686_, _28685_, _08643_);
  and (_28687_, _28686_, _28684_);
  nor (_28688_, _28660_, _12493_);
  or (_28689_, _12128_, _07200_);
  or (_28690_, _07199_, \uc8051golden_1.PC [11]);
  or (_28692_, _28690_, _07332_);
  nand (_28693_, _28692_, _28689_);
  and (_28694_, _25019_, _06855_);
  and (_28695_, _28694_, _28693_);
  nor (_28696_, _12128_, _07366_);
  or (_28697_, _28696_, _08643_);
  or (_28698_, _28697_, _28695_);
  or (_28699_, _28698_, _28688_);
  nand (_28700_, _28699_, _12497_);
  or (_28701_, _28700_, _28687_);
  and (_28703_, _28701_, _28678_);
  nand (_28704_, _12509_, _12458_);
  or (_28705_, _28704_, _28703_);
  and (_28706_, _28705_, _28670_);
  or (_28707_, _28706_, _12502_);
  and (_28708_, _28707_, _28668_);
  or (_28709_, _28708_, _06406_);
  and (_28710_, _12455_, _06414_);
  or (_28711_, _28710_, _12128_);
  and (_28712_, _28711_, _12517_);
  and (_28714_, _28712_, _28709_);
  and (_28715_, _28660_, _12519_);
  or (_28716_, _28715_, _12524_);
  or (_28717_, _28716_, _28714_);
  or (_28718_, _12523_, _12128_);
  and (_28719_, _28718_, _28717_);
  or (_28720_, _28719_, _12450_);
  or (_28721_, _28674_, _12444_);
  nand (_28722_, _12444_, _12269_);
  and (_28723_, _28722_, _28721_);
  or (_28725_, _28723_, _12449_);
  and (_28726_, _28725_, _28720_);
  or (_28727_, _28726_, _06457_);
  and (_28728_, _12405_, _12268_);
  and (_28729_, _28674_, _12407_);
  or (_28730_, _28729_, _12411_);
  or (_28731_, _28730_, _28728_);
  and (_28732_, _28731_, _06842_);
  and (_28733_, _28732_, _28727_);
  and (_28734_, _12546_, _12268_);
  and (_28736_, _28674_, _12548_);
  or (_28737_, _28736_, _28734_);
  and (_28738_, _28737_, _06420_);
  or (_28739_, _28738_, _28733_);
  and (_28740_, _28739_, _12534_);
  or (_28741_, _28674_, _12249_);
  nand (_28742_, _12269_, _12249_);
  and (_28743_, _28742_, _06482_);
  and (_28744_, _28743_, _28741_);
  or (_28745_, _28744_, _28740_);
  and (_28747_, _28745_, _12238_);
  nand (_28748_, _28660_, _12237_);
  nand (_28749_, _28748_, _12570_);
  or (_28750_, _28749_, _28747_);
  or (_28751_, _12570_, _12128_);
  and (_28752_, _28751_, _12576_);
  and (_28753_, _28752_, _28750_);
  and (_28754_, _28660_, _12580_);
  or (_28755_, _28754_, _12583_);
  or (_28756_, _28755_, _28753_);
  or (_28758_, _12582_, _12128_);
  and (_28759_, _28758_, _12588_);
  and (_28760_, _28759_, _28756_);
  and (_28761_, _28660_, _12594_);
  or (_28762_, _28761_, _12593_);
  or (_28763_, _28762_, _28760_);
  or (_28764_, _12128_, _12592_);
  and (_28765_, _28764_, _06023_);
  and (_28766_, _28765_, _28763_);
  nand (_28767_, _28660_, _06022_);
  nand (_28769_, _28767_, _12602_);
  or (_28770_, _28769_, _28766_);
  or (_28771_, _12602_, _12128_);
  and (_28772_, _28771_, _06473_);
  and (_28773_, _28772_, _28770_);
  nand (_28774_, _12268_, _06472_);
  nand (_28775_, _28774_, _06294_);
  or (_28776_, _28775_, _28773_);
  or (_28777_, _12128_, _06294_);
  and (_28778_, _28777_, _06279_);
  and (_28780_, _28778_, _28776_);
  or (_28781_, _28780_, _28667_);
  and (_28782_, _28781_, _12616_);
  and (_28783_, _28660_, _12620_);
  or (_28784_, _28783_, _12619_);
  or (_28785_, _28784_, _28782_);
  or (_28786_, _12618_, _12128_);
  and (_28787_, _28786_, _12625_);
  and (_28788_, _28787_, _28785_);
  and (_28789_, _28683_, _12624_);
  or (_28791_, _28789_, _09013_);
  or (_28792_, _28791_, _28788_);
  and (_28793_, _28792_, _28666_);
  or (_28794_, _28793_, _06275_);
  nand (_28795_, _12269_, _06275_);
  and (_28796_, _28795_, _10934_);
  and (_28797_, _28796_, _28794_);
  and (_28798_, _12128_, _10933_);
  or (_28799_, _28798_, _28797_);
  and (_28800_, _28799_, _12640_);
  or (_28802_, _12666_, \uc8051golden_1.DPH [3]);
  nor (_28803_, _12667_, _12640_);
  and (_28804_, _28803_, _28802_);
  or (_28805_, _28804_, _12677_);
  or (_28806_, _28805_, _28800_);
  or (_28807_, _12676_, _12128_);
  and (_28808_, _28807_, _12681_);
  and (_28809_, _28808_, _28806_);
  or (_28810_, _28683_, _11297_);
  or (_28811_, _12128_, _12687_);
  and (_28813_, _28811_, _12680_);
  and (_28814_, _28813_, _28810_);
  or (_28815_, _28814_, _12685_);
  or (_28816_, _28815_, _28809_);
  and (_28817_, _28816_, _28665_);
  or (_28818_, _28817_, _12228_);
  or (_28819_, _12128_, _12227_);
  and (_28820_, _28819_, _07282_);
  and (_28821_, _28820_, _28818_);
  nand (_28822_, _12268_, _06474_);
  nand (_28824_, _28822_, _12700_);
  or (_28825_, _28824_, _28821_);
  or (_28826_, _12700_, _12128_);
  and (_28827_, _28826_, _12705_);
  and (_28828_, _28827_, _28825_);
  or (_28829_, _28683_, _12687_);
  or (_28830_, _12128_, _11297_);
  and (_28831_, _28830_, _12704_);
  and (_28832_, _28831_, _28829_);
  or (_28833_, _28832_, _12723_);
  or (_28835_, _28833_, _28828_);
  and (_28836_, _28835_, _28664_);
  or (_28837_, _28836_, _12722_);
  or (_28838_, _12128_, _12721_);
  and (_28839_, _28838_, _07279_);
  and (_28840_, _28839_, _28837_);
  nand (_28841_, _12268_, _06478_);
  nand (_28842_, _28841_, _12731_);
  or (_28843_, _28842_, _28840_);
  or (_28844_, _12731_, _12128_);
  and (_28846_, _28844_, _12736_);
  and (_28847_, _28846_, _28843_);
  or (_28848_, _28683_, \uc8051golden_1.PSW [7]);
  or (_28849_, _12128_, _10524_);
  and (_28850_, _28849_, _12735_);
  and (_28851_, _28850_, _28848_);
  or (_28852_, _28851_, _12224_);
  or (_28853_, _28852_, _28847_);
  and (_28854_, _28853_, _28663_);
  or (_28855_, _28854_, _11019_);
  or (_28857_, _12128_, _11018_);
  and (_28858_, _28857_, _09043_);
  and (_28859_, _28858_, _28855_);
  nand (_28860_, _12268_, _06479_);
  nand (_28861_, _28860_, _12752_);
  or (_28862_, _28861_, _28859_);
  or (_28863_, _12752_, _12128_);
  and (_28864_, _28863_, _12756_);
  and (_28865_, _28864_, _28862_);
  or (_28866_, _28683_, _10524_);
  or (_28868_, _12128_, \uc8051golden_1.PSW [7]);
  and (_28869_, _28868_, _12217_);
  and (_28870_, _28869_, _28866_);
  or (_28871_, _28870_, _12763_);
  or (_28872_, _28871_, _28865_);
  and (_28873_, _28872_, _28662_);
  or (_28874_, _28873_, _11061_);
  or (_28875_, _12128_, _11060_);
  and (_28876_, _28875_, _11090_);
  and (_28877_, _28876_, _28874_);
  and (_28879_, _28660_, _11089_);
  or (_28880_, _28879_, _06588_);
  or (_28881_, _28880_, _28877_);
  nand (_28882_, _07775_, _06588_);
  and (_28883_, _28882_, _28881_);
  or (_28884_, _28883_, _05966_);
  or (_28885_, _12128_, _05967_);
  and (_28886_, _28885_, _06596_);
  and (_28887_, _28886_, _28884_);
  or (_28888_, _28674_, _12959_);
  or (_28890_, _12268_, _12958_);
  and (_28891_, _28890_, _06460_);
  and (_28892_, _28891_, _28888_);
  or (_28893_, _28892_, _12779_);
  or (_28894_, _28893_, _28887_);
  and (_28895_, _28894_, _28661_);
  or (_28896_, _28895_, _12094_);
  or (_28897_, _12128_, _11204_);
  and (_28898_, _28897_, _12968_);
  and (_28899_, _28898_, _28896_);
  and (_28900_, _28660_, _11243_);
  or (_28901_, _28900_, _06305_);
  or (_28902_, _28901_, _28899_);
  nand (_28903_, _07775_, _06305_);
  and (_28904_, _28903_, _28902_);
  or (_28905_, _28904_, _05971_);
  or (_28906_, _12128_, _12979_);
  and (_28907_, _28906_, _12978_);
  and (_28908_, _28907_, _28905_);
  or (_28909_, _28674_, _12958_);
  nand (_28912_, _12269_, _12958_);
  and (_28913_, _28912_, _28909_);
  and (_28914_, _28913_, _06487_);
  or (_28915_, _28914_, _12988_);
  or (_28916_, _28915_, _28908_);
  or (_28917_, _28660_, _12987_);
  and (_28918_, _28917_, _07037_);
  and (_28919_, _28918_, _28916_);
  nand (_28920_, _12128_, _06606_);
  nand (_28921_, _28920_, _12994_);
  or (_28923_, _28921_, _28919_);
  or (_28924_, _28660_, _12994_);
  and (_28925_, _28924_, _09463_);
  and (_28926_, _28925_, _28923_);
  nor (_28927_, _09463_, _06372_);
  or (_28928_, _28927_, _05969_);
  or (_28929_, _28928_, _28926_);
  or (_28930_, _12128_, _13005_);
  and (_28931_, _28930_, _06807_);
  and (_28932_, _28931_, _28929_);
  and (_28934_, _28913_, _06234_);
  or (_28935_, _28934_, _13012_);
  or (_28936_, _28935_, _28932_);
  or (_28937_, _28660_, _13011_);
  and (_28938_, _28937_, _06196_);
  and (_28939_, _28938_, _28936_);
  nand (_28940_, _12128_, _06195_);
  nand (_28941_, _28940_, _13019_);
  or (_28942_, _28941_, _28939_);
  or (_28943_, _28660_, _13019_);
  and (_28945_, _28943_, _13023_);
  and (_28946_, _28945_, _28942_);
  nor (_28947_, _13023_, _06372_);
  or (_28948_, _28947_, _05963_);
  or (_28949_, _28948_, _28946_);
  or (_28950_, _12128_, _05964_);
  and (_28951_, _28950_, _13031_);
  and (_28952_, _28951_, _28949_);
  and (_28953_, _28660_, _13030_);
  or (_28954_, _28953_, _28952_);
  or (_28956_, _28954_, _01379_);
  or (_28957_, _01375_, \uc8051golden_1.PC [11]);
  and (_28958_, _28957_, _42545_);
  and (_42988_, _28958_, _28956_);
  and (_28959_, _12097_, _09465_);
  and (_28960_, _28959_, \uc8051golden_1.PC [11]);
  and (_28961_, _28960_, \uc8051golden_1.PC [12]);
  nor (_28962_, _28960_, \uc8051golden_1.PC [12]);
  nor (_28963_, _28962_, _28961_);
  not (_28964_, _28963_);
  and (_28966_, _28964_, _11243_);
  nor (_28967_, _12752_, _15323_);
  nor (_28968_, _12731_, _15323_);
  nor (_28969_, _12700_, _15323_);
  and (_28970_, _12405_, _12262_);
  and (_28971_, _12358_, _12355_);
  nor (_28972_, _28971_, _12359_);
  and (_28973_, _28972_, _12407_);
  nor (_28974_, _28973_, _28970_);
  nand (_28975_, _28974_, _06457_);
  nor (_28977_, _28964_, _12517_);
  nor (_28978_, _28963_, _12509_);
  nand (_28979_, _12466_, _12262_);
  not (_28980_, _28972_);
  or (_28981_, _28980_, _12466_);
  and (_28982_, _28981_, _06401_);
  and (_28983_, _28982_, _28979_);
  and (_28984_, _12203_, _12200_);
  nor (_28985_, _28984_, _12204_);
  nand (_28986_, _28985_, _12474_);
  or (_28988_, _12474_, _15323_);
  and (_28989_, _28988_, _08643_);
  nand (_28990_, _28989_, _28986_);
  and (_28991_, _28964_, _12481_);
  nor (_28992_, _12481_, _12121_);
  nor (_28993_, _28992_, _28991_);
  nor (_28994_, _28993_, _25019_);
  nor (_28995_, _28964_, _12493_);
  not (_28996_, _28995_);
  and (_28997_, _15323_, _07199_);
  nor (_28999_, _28997_, _06854_);
  not (_29000_, _28999_);
  and (_29001_, _07333_, \uc8051golden_1.PC [12]);
  nor (_29002_, _29001_, _07199_);
  nor (_29003_, _29002_, _29000_);
  nor (_29004_, _29003_, _06790_);
  and (_29005_, _29004_, _28996_);
  nor (_29006_, _29005_, _28994_);
  nor (_29007_, _29006_, _08643_);
  nor (_29008_, _29007_, _07212_);
  nand (_29010_, _29008_, _28990_);
  and (_29011_, _28963_, _07212_);
  nor (_29012_, _29011_, _06401_);
  and (_29013_, _29012_, _29010_);
  or (_29014_, _29013_, _28983_);
  nand (_29015_, _29014_, _12458_);
  nor (_29016_, _28963_, _12458_);
  nor (_29017_, _29016_, _12502_);
  nand (_29018_, _29017_, _29015_);
  nor (_29019_, _12455_, _15323_);
  nor (_29021_, _29019_, _12510_);
  and (_29022_, _29021_, _29018_);
  or (_29023_, _29022_, _28978_);
  nand (_29024_, _29023_, _06414_);
  and (_29025_, _15323_, _06406_);
  nor (_29026_, _29025_, _12519_);
  and (_29027_, _29026_, _29024_);
  or (_29028_, _29027_, _28977_);
  nand (_29029_, _29028_, _12523_);
  nor (_29030_, _12523_, _15323_);
  nor (_29032_, _29030_, _12450_);
  and (_29033_, _29032_, _29029_);
  and (_29034_, _12444_, _12262_);
  nor (_29035_, _28980_, _12444_);
  or (_29036_, _29035_, _29034_);
  nor (_29037_, _29036_, _12449_);
  or (_29038_, _29037_, _29033_);
  nand (_29039_, _29038_, _12411_);
  and (_29040_, _29039_, _28975_);
  or (_29041_, _29040_, _06420_);
  nor (_29043_, _28980_, _12546_);
  and (_29044_, _12546_, _12262_);
  or (_29045_, _29044_, _06842_);
  or (_29046_, _29045_, _29043_);
  and (_29047_, _29046_, _12534_);
  nand (_29048_, _29047_, _29041_);
  and (_29049_, _12262_, _12249_);
  and (_29050_, _28972_, _26421_);
  or (_29051_, _29050_, _29049_);
  and (_29052_, _29051_, _06482_);
  nor (_29054_, _29052_, _12237_);
  and (_29055_, _29054_, _29048_);
  and (_29056_, _28964_, _12237_);
  or (_29057_, _29056_, _29055_);
  and (_29058_, _29057_, _12570_);
  nor (_29059_, _12570_, _12121_);
  or (_29060_, _29059_, _29058_);
  nand (_29061_, _29060_, _12576_);
  nor (_29062_, _28963_, _12576_);
  nor (_29063_, _29062_, _12583_);
  nand (_29065_, _29063_, _29061_);
  nor (_29066_, _12582_, _15323_);
  nor (_29067_, _29066_, _12594_);
  nand (_29068_, _29067_, _29065_);
  nor (_29069_, _28963_, _12588_);
  nor (_29070_, _29069_, _12593_);
  nand (_29071_, _29070_, _29068_);
  nor (_29072_, _15323_, _12592_);
  nor (_29073_, _29072_, _06022_);
  nand (_29074_, _29073_, _29071_);
  and (_29076_, _28964_, _06022_);
  nor (_29077_, _29076_, _12603_);
  nand (_29078_, _29077_, _29074_);
  nor (_29079_, _12602_, _15323_);
  nor (_29080_, _29079_, _06472_);
  nand (_29081_, _29080_, _29078_);
  and (_29082_, _12263_, _06472_);
  nor (_29083_, _29082_, _13788_);
  nand (_29084_, _29083_, _29081_);
  nor (_29085_, _15323_, _06294_);
  nor (_29087_, _29085_, _06015_);
  nand (_29088_, _29087_, _29084_);
  and (_29089_, _12263_, _06015_);
  nor (_29090_, _29089_, _12620_);
  nand (_29091_, _29090_, _29088_);
  nor (_29092_, _28964_, _12616_);
  nor (_29093_, _29092_, _12619_);
  nand (_29094_, _29093_, _29091_);
  nor (_29095_, _12618_, _12121_);
  nor (_29096_, _29095_, _12624_);
  and (_29098_, _29096_, _29094_);
  and (_29099_, _28985_, _12624_);
  nor (_29100_, _29099_, _29098_);
  or (_29101_, _29100_, _09013_);
  or (_29102_, _15323_, _09012_);
  and (_29103_, _29102_, _06276_);
  nand (_29104_, _29103_, _29101_);
  and (_29105_, _12263_, _06275_);
  nor (_29106_, _29105_, _10933_);
  nand (_29107_, _29106_, _29104_);
  and (_29109_, _12121_, _10933_);
  nor (_29110_, _29109_, _12639_);
  and (_29111_, _29110_, _29107_);
  nor (_29112_, _12667_, \uc8051golden_1.DPH [4]);
  nor (_29113_, _29112_, _12668_);
  nor (_29114_, _29113_, _12640_);
  or (_29115_, _29114_, _29111_);
  nand (_29116_, _29115_, _12676_);
  nor (_29117_, _12676_, _12121_);
  nor (_29118_, _29117_, _12680_);
  nand (_29120_, _29118_, _29116_);
  nor (_29121_, _12121_, _12687_);
  nor (_29122_, _28985_, _11297_);
  or (_29123_, _29122_, _12681_);
  or (_29124_, _29123_, _29121_);
  and (_29125_, _29124_, _12233_);
  nand (_29126_, _29125_, _29120_);
  nor (_29127_, _28963_, _12233_);
  nor (_29128_, _29127_, _12228_);
  nand (_29129_, _29128_, _29126_);
  nor (_29131_, _15323_, _12227_);
  nor (_29132_, _29131_, _06474_);
  nand (_29133_, _29132_, _29129_);
  and (_29134_, _12263_, _06474_);
  nor (_29135_, _29134_, _12701_);
  and (_29136_, _29135_, _29133_);
  or (_29137_, _29136_, _28969_);
  nand (_29138_, _29137_, _12705_);
  and (_29139_, _12121_, _12687_);
  and (_29140_, _28985_, _11297_);
  or (_29142_, _29140_, _29139_);
  and (_29143_, _29142_, _12704_);
  nor (_29144_, _29143_, _12723_);
  nand (_29145_, _29144_, _29138_);
  nor (_29146_, _28963_, _12719_);
  nor (_29147_, _29146_, _12722_);
  nand (_29148_, _29147_, _29145_);
  nor (_29149_, _15323_, _12721_);
  nor (_29150_, _29149_, _06478_);
  nand (_29151_, _29150_, _29148_);
  and (_29153_, _12263_, _06478_);
  nor (_29154_, _29153_, _12732_);
  and (_29155_, _29154_, _29151_);
  or (_29156_, _29155_, _28968_);
  nand (_29157_, _29156_, _12736_);
  and (_29158_, _12121_, \uc8051golden_1.PSW [7]);
  and (_29159_, _28985_, _10524_);
  or (_29160_, _29159_, _29158_);
  and (_29161_, _29160_, _12735_);
  nor (_29162_, _29161_, _12224_);
  nand (_29164_, _29162_, _29157_);
  and (_29165_, _28964_, _12224_);
  nor (_29166_, _29165_, _11019_);
  nand (_29167_, _29166_, _29164_);
  nor (_29168_, _15323_, _11018_);
  nor (_29169_, _29168_, _06479_);
  nand (_29170_, _29169_, _29167_);
  and (_29171_, _12263_, _06479_);
  nor (_29172_, _29171_, _12753_);
  and (_29173_, _29172_, _29170_);
  or (_29175_, _29173_, _28967_);
  nand (_29176_, _29175_, _12756_);
  and (_29177_, _12121_, _10524_);
  and (_29178_, _28985_, \uc8051golden_1.PSW [7]);
  or (_29179_, _29178_, _29177_);
  and (_29180_, _29179_, _12217_);
  nor (_29181_, _29180_, _12763_);
  nand (_29182_, _29181_, _29176_);
  nor (_29183_, _28963_, _12761_);
  nor (_29184_, _29183_, _11061_);
  nand (_29186_, _29184_, _29182_);
  nor (_29187_, _15323_, _11060_);
  nor (_29188_, _29187_, _11089_);
  nand (_29189_, _29188_, _29186_);
  and (_29190_, _28964_, _11089_);
  nor (_29191_, _29190_, _06588_);
  and (_29192_, _29191_, _29189_);
  nor (_29193_, _08301_, _13881_);
  or (_29194_, _29193_, _05966_);
  or (_29195_, _29194_, _29192_);
  and (_29197_, _15323_, _05966_);
  nor (_29198_, _29197_, _06460_);
  nand (_29199_, _29198_, _29195_);
  nor (_29200_, _12262_, _12958_);
  and (_29201_, _28980_, _12958_);
  or (_29202_, _29201_, _06596_);
  or (_29203_, _29202_, _29200_);
  and (_29204_, _29203_, _12108_);
  nand (_29205_, _29204_, _29199_);
  nor (_29206_, _28963_, _12108_);
  nor (_29208_, _29206_, _12094_);
  nand (_29209_, _29208_, _29205_);
  nor (_29210_, _15323_, _11204_);
  nor (_29211_, _29210_, _11243_);
  and (_29212_, _29211_, _29209_);
  or (_29213_, _29212_, _28966_);
  nand (_29214_, _29213_, _06306_);
  and (_29215_, _08301_, _06305_);
  nor (_29216_, _29215_, _05971_);
  nand (_29217_, _29216_, _29214_);
  and (_29219_, _12121_, _05971_);
  nor (_29220_, _29219_, _06487_);
  and (_29221_, _29220_, _29217_);
  nor (_29222_, _28972_, _12958_);
  and (_29223_, _12263_, _12958_);
  nor (_29224_, _29223_, _29222_);
  nor (_29225_, _29224_, _12978_);
  or (_29226_, _29225_, _29221_);
  and (_29227_, _29226_, _12987_);
  nor (_29228_, _28963_, _12987_);
  or (_29230_, _29228_, _29227_);
  nand (_29231_, _29230_, _07037_);
  nand (_29232_, _15323_, _06606_);
  and (_29233_, _29232_, _12994_);
  nand (_29234_, _29233_, _29231_);
  nor (_29235_, _28964_, _12994_);
  nor (_29236_, _29235_, _06465_);
  nand (_29237_, _29236_, _29234_);
  and (_29238_, _06465_, _06265_);
  nor (_29239_, _29238_, _05969_);
  nand (_29241_, _29239_, _29237_);
  and (_29242_, _12121_, _05969_);
  nor (_29243_, _29242_, _06234_);
  nand (_29244_, _29243_, _29241_);
  nor (_29245_, _29224_, _06807_);
  nor (_29246_, _29245_, _13012_);
  nand (_29247_, _29246_, _29244_);
  nor (_29248_, _28964_, _13011_);
  nor (_29249_, _29248_, _06195_);
  nand (_29250_, _29249_, _29247_);
  and (_29252_, _15323_, _06195_);
  nor (_29253_, _29252_, _13020_);
  nand (_29254_, _29253_, _29250_);
  nor (_29255_, _28964_, _13019_);
  nor (_29256_, _29255_, _06475_);
  and (_29257_, _29256_, _29254_);
  and (_29258_, _06475_, _06265_);
  or (_29259_, _29258_, _05963_);
  nor (_29260_, _29259_, _29257_);
  and (_29261_, _12121_, _05963_);
  or (_29263_, _29261_, _13030_);
  nor (_29264_, _29263_, _29260_);
  and (_29265_, _28964_, _13030_);
  nor (_29266_, _29265_, _29264_);
  or (_29267_, _29266_, _01379_);
  or (_29268_, _01375_, \uc8051golden_1.PC [12]);
  and (_29269_, _29268_, _42545_);
  and (_42989_, _29269_, _29267_);
  and (_29270_, _28961_, \uc8051golden_1.PC [13]);
  nor (_29271_, _28961_, \uc8051golden_1.PC [13]);
  nor (_29273_, _29271_, _29270_);
  and (_29274_, _29273_, _13030_);
  or (_29275_, _29273_, _12108_);
  or (_29276_, _29273_, _12761_);
  not (_29277_, _29273_);
  nand (_29278_, _29277_, _12224_);
  or (_29279_, _12119_, _12118_);
  not (_29280_, _29279_);
  nor (_29281_, _29280_, _12205_);
  and (_29282_, _29280_, _12205_);
  or (_29284_, _29282_, _29281_);
  or (_29285_, _29284_, _12687_);
  or (_29286_, _12117_, _11297_);
  and (_29287_, _29286_, _12704_);
  and (_29288_, _29287_, _29285_);
  or (_29289_, _29273_, _12233_);
  or (_29290_, _12117_, _09012_);
  and (_29291_, _12258_, _06015_);
  or (_29292_, _29273_, _12588_);
  nor (_29293_, _29277_, _12576_);
  or (_29295_, _12407_, _12258_);
  or (_29296_, _12260_, _12259_);
  not (_29297_, _29296_);
  nor (_29298_, _29297_, _12360_);
  and (_29299_, _29297_, _12360_);
  or (_29300_, _29299_, _29298_);
  or (_29301_, _29300_, _12405_);
  and (_29302_, _29301_, _06457_);
  and (_29303_, _29302_, _29295_);
  or (_29304_, _14077_, _12258_);
  or (_29306_, _29300_, _12444_);
  and (_29307_, _29306_, _12450_);
  and (_29308_, _29307_, _29304_);
  and (_29309_, _12117_, _06406_);
  or (_29310_, _12455_, _12117_);
  or (_29311_, _12464_, _12258_);
  or (_29312_, _29300_, _12466_);
  and (_29313_, _29312_, _06401_);
  and (_29314_, _29313_, _29311_);
  and (_29315_, _12476_, _12117_);
  and (_29317_, _29284_, _12474_);
  or (_29318_, _29317_, _08644_);
  or (_29319_, _29318_, _29315_);
  or (_29320_, _12482_, _12117_);
  or (_29321_, _06790_, \uc8051golden_1.PC [13]);
  or (_29322_, _29321_, _12485_);
  or (_29323_, _29322_, _07332_);
  and (_29324_, _29323_, _29320_);
  or (_29325_, _29324_, _12481_);
  or (_29326_, _29273_, _12493_);
  and (_29328_, _29326_, _29325_);
  or (_29329_, _29328_, _08643_);
  and (_29330_, _29329_, _12497_);
  and (_29331_, _29330_, _29319_);
  or (_29332_, _29331_, _29314_);
  and (_29333_, _29332_, _12458_);
  nor (_29334_, _29277_, _12503_);
  or (_29335_, _29334_, _12502_);
  or (_29336_, _29335_, _29333_);
  and (_29337_, _29336_, _29310_);
  or (_29339_, _29337_, _12510_);
  or (_29340_, _29273_, _12509_);
  and (_29341_, _29340_, _06414_);
  and (_29342_, _29341_, _29339_);
  or (_29343_, _29342_, _29309_);
  and (_29344_, _29343_, _12517_);
  or (_29345_, _29277_, _12517_);
  nand (_29346_, _29345_, _12523_);
  or (_29347_, _29346_, _29344_);
  or (_29348_, _12523_, _12117_);
  and (_29350_, _29348_, _12449_);
  and (_29351_, _29350_, _29347_);
  or (_29352_, _29351_, _29308_);
  and (_29353_, _29352_, _12411_);
  or (_29354_, _29353_, _06420_);
  or (_29355_, _29354_, _29303_);
  and (_29356_, _12546_, _12258_);
  and (_29357_, _29300_, _12548_);
  or (_29358_, _29357_, _06842_);
  or (_29359_, _29358_, _29356_);
  and (_29361_, _29359_, _12534_);
  and (_29362_, _29361_, _29355_);
  or (_29363_, _29300_, _12249_);
  or (_29364_, _12258_, _26421_);
  and (_29365_, _29364_, _06482_);
  and (_29366_, _29365_, _29363_);
  or (_29367_, _29366_, _29362_);
  and (_29368_, _29367_, _12238_);
  nand (_29369_, _29273_, _12237_);
  nand (_29370_, _29369_, _12570_);
  or (_29372_, _29370_, _29368_);
  or (_29373_, _12570_, _12117_);
  and (_29374_, _29373_, _12576_);
  and (_29375_, _29374_, _29372_);
  or (_29376_, _29375_, _29293_);
  and (_29377_, _29376_, _12582_);
  or (_29378_, _12582_, _15518_);
  nand (_29379_, _29378_, _12588_);
  or (_29380_, _29379_, _29377_);
  and (_29381_, _29380_, _29292_);
  or (_29383_, _29381_, _12593_);
  or (_29384_, _12117_, _12592_);
  and (_29385_, _29384_, _06023_);
  and (_29386_, _29385_, _29383_);
  nand (_29387_, _29273_, _06022_);
  nand (_29388_, _29387_, _12602_);
  or (_29389_, _29388_, _29386_);
  or (_29390_, _12602_, _12117_);
  and (_29391_, _29390_, _06473_);
  and (_29392_, _29391_, _29389_);
  nand (_29394_, _12258_, _06472_);
  nand (_29395_, _29394_, _06294_);
  or (_29396_, _29395_, _29392_);
  or (_29397_, _12117_, _06294_);
  and (_29398_, _29397_, _06279_);
  and (_29399_, _29398_, _29396_);
  or (_29400_, _29399_, _29291_);
  and (_29401_, _29400_, _12616_);
  nor (_29402_, _29277_, _12616_);
  or (_29403_, _29402_, _12619_);
  or (_29405_, _29403_, _29401_);
  or (_29406_, _12618_, _12117_);
  and (_29407_, _29406_, _12625_);
  and (_29408_, _29407_, _29405_);
  and (_29409_, _29284_, _12624_);
  or (_29410_, _29409_, _09013_);
  or (_29411_, _29410_, _29408_);
  and (_29412_, _29411_, _29290_);
  or (_29413_, _29412_, _06275_);
  or (_29414_, _12258_, _06276_);
  and (_29416_, _29414_, _10934_);
  and (_29417_, _29416_, _29413_);
  and (_29418_, _12117_, _10933_);
  or (_29419_, _29418_, _29417_);
  and (_29420_, _29419_, _12640_);
  or (_29421_, _12668_, \uc8051golden_1.DPH [5]);
  nor (_29422_, _12669_, _12640_);
  and (_29423_, _29422_, _29421_);
  or (_29424_, _29423_, _12677_);
  or (_29425_, _29424_, _29420_);
  or (_29426_, _12676_, _12117_);
  and (_29427_, _29426_, _12681_);
  and (_29428_, _29427_, _29425_);
  or (_29429_, _29284_, _11297_);
  or (_29430_, _12117_, _12687_);
  and (_29431_, _29430_, _12680_);
  and (_29432_, _29431_, _29429_);
  or (_29433_, _29432_, _12685_);
  or (_29434_, _29433_, _29428_);
  and (_29435_, _29434_, _29289_);
  or (_29438_, _29435_, _12228_);
  or (_29439_, _12117_, _12227_);
  and (_29440_, _29439_, _07282_);
  and (_29441_, _29440_, _29438_);
  nand (_29442_, _12258_, _06474_);
  nand (_29443_, _29442_, _12700_);
  or (_29444_, _29443_, _29441_);
  or (_29445_, _12700_, _12117_);
  and (_29446_, _29445_, _12705_);
  and (_29447_, _29446_, _29444_);
  or (_29449_, _29447_, _29288_);
  and (_29450_, _29449_, _12719_);
  nor (_29451_, _29277_, _12719_);
  or (_29452_, _29451_, _12722_);
  or (_29453_, _29452_, _29450_);
  or (_29454_, _12117_, _12721_);
  and (_29455_, _29454_, _07279_);
  and (_29456_, _29455_, _29453_);
  nand (_29457_, _12258_, _06478_);
  nand (_29458_, _29457_, _12731_);
  or (_29460_, _29458_, _29456_);
  or (_29461_, _12731_, _12117_);
  and (_29462_, _29461_, _12736_);
  and (_29463_, _29462_, _29460_);
  or (_29464_, _29284_, \uc8051golden_1.PSW [7]);
  or (_29465_, _12117_, _10524_);
  and (_29466_, _29465_, _12735_);
  and (_29467_, _29466_, _29464_);
  or (_29468_, _29467_, _12224_);
  or (_29469_, _29468_, _29463_);
  and (_29471_, _29469_, _29278_);
  or (_29472_, _29471_, _11019_);
  or (_29473_, _12117_, _11018_);
  and (_29474_, _29473_, _09043_);
  and (_29475_, _29474_, _29472_);
  nand (_29476_, _12258_, _06479_);
  nand (_29477_, _29476_, _12752_);
  or (_29478_, _29477_, _29475_);
  or (_29479_, _12752_, _12117_);
  and (_29480_, _29479_, _12756_);
  and (_29482_, _29480_, _29478_);
  or (_29483_, _29284_, _10524_);
  or (_29484_, _12117_, \uc8051golden_1.PSW [7]);
  and (_29485_, _29484_, _12217_);
  and (_29486_, _29485_, _29483_);
  or (_29487_, _29486_, _12763_);
  or (_29488_, _29487_, _29482_);
  and (_29489_, _29488_, _29276_);
  or (_29490_, _29489_, _11061_);
  or (_29491_, _12117_, _11060_);
  and (_29493_, _29491_, _11090_);
  and (_29494_, _29493_, _29490_);
  and (_29495_, _29273_, _11089_);
  or (_29496_, _29495_, _06588_);
  or (_29497_, _29496_, _29494_);
  nand (_29498_, _08207_, _06588_);
  and (_29499_, _29498_, _29497_);
  or (_29500_, _29499_, _05966_);
  nand (_29501_, _15518_, _05966_);
  and (_29502_, _29501_, _06596_);
  and (_29504_, _29502_, _29500_);
  or (_29505_, _29300_, _12959_);
  or (_29506_, _12258_, _12958_);
  and (_29507_, _29506_, _06460_);
  and (_29508_, _29507_, _29505_);
  or (_29509_, _29508_, _12779_);
  or (_29510_, _29509_, _29504_);
  and (_29511_, _29510_, _29275_);
  or (_29512_, _29511_, _12094_);
  or (_29513_, _12117_, _11204_);
  and (_29515_, _29513_, _12968_);
  and (_29516_, _29515_, _29512_);
  and (_29517_, _29273_, _11243_);
  or (_29518_, _29517_, _06305_);
  or (_29519_, _29518_, _29516_);
  nand (_29520_, _08207_, _06305_);
  and (_29521_, _29520_, _29519_);
  or (_29522_, _29521_, _05971_);
  nand (_29523_, _15518_, _05971_);
  and (_29524_, _29523_, _12978_);
  and (_29526_, _29524_, _29522_);
  or (_29527_, _12258_, _12959_);
  or (_29528_, _29300_, _12958_);
  and (_29529_, _29528_, _29527_);
  and (_29530_, _29529_, _06487_);
  or (_29531_, _29530_, _12988_);
  or (_29532_, _29531_, _29526_);
  or (_29533_, _29273_, _12987_);
  and (_29534_, _29533_, _07037_);
  and (_29535_, _29534_, _29532_);
  nand (_29537_, _12117_, _06606_);
  nand (_29538_, _29537_, _12994_);
  or (_29539_, _29538_, _29535_);
  or (_29540_, _29273_, _12994_);
  and (_29541_, _29540_, _09463_);
  and (_29542_, _29541_, _29539_);
  nor (_29543_, _06650_, _09463_);
  or (_29544_, _29543_, _05969_);
  or (_29545_, _29544_, _29542_);
  nand (_29546_, _15518_, _05969_);
  and (_29548_, _29546_, _06807_);
  and (_29549_, _29548_, _29545_);
  and (_29550_, _29529_, _06234_);
  or (_29551_, _29550_, _13012_);
  or (_29552_, _29551_, _29549_);
  or (_29553_, _29273_, _13011_);
  and (_29554_, _29553_, _06196_);
  and (_29555_, _29554_, _29552_);
  nand (_29556_, _12117_, _06195_);
  nand (_29557_, _29556_, _13019_);
  or (_29559_, _29557_, _29555_);
  or (_29560_, _29273_, _13019_);
  and (_29561_, _29560_, _13023_);
  and (_29562_, _29561_, _29559_);
  nor (_29563_, _06650_, _13023_);
  or (_29564_, _29563_, _05963_);
  or (_29565_, _29564_, _29562_);
  nand (_29566_, _15518_, _05963_);
  and (_29567_, _29566_, _13031_);
  and (_29568_, _29567_, _29565_);
  or (_29570_, _29568_, _29274_);
  or (_29571_, _29570_, _01379_);
  or (_29572_, _01375_, \uc8051golden_1.PC [13]);
  and (_29573_, _29572_, _42545_);
  and (_42991_, _29573_, _29571_);
  nor (_29574_, _29270_, \uc8051golden_1.PC [14]);
  nor (_29575_, _29574_, _12104_);
  nor (_29576_, _29575_, _12968_);
  nor (_29577_, _12752_, _15722_);
  nor (_29578_, _12731_, _15722_);
  nor (_29580_, _12700_, _15722_);
  nor (_29581_, _12676_, _15722_);
  and (_29582_, _15722_, _06406_);
  and (_29583_, _12362_, _12256_);
  nor (_29584_, _29583_, _12363_);
  or (_29585_, _29584_, _12466_);
  or (_29586_, _12464_, _12251_);
  and (_29587_, _29586_, _06401_);
  and (_29588_, _29587_, _29585_);
  and (_29589_, _12476_, _12111_);
  and (_29591_, _12207_, _12115_);
  nor (_29592_, _29591_, _12208_);
  and (_29593_, _29592_, _12474_);
  nor (_29594_, _29593_, _29589_);
  nand (_29595_, _29594_, _08643_);
  not (_29596_, _29575_);
  and (_29597_, _29596_, _12481_);
  nor (_29598_, _12481_, _12111_);
  nor (_29599_, _29598_, _29597_);
  nor (_29600_, _29599_, _25019_);
  nor (_29602_, _29596_, _12493_);
  not (_29603_, _29602_);
  and (_29604_, _15722_, _07199_);
  nor (_29605_, _29604_, _06854_);
  not (_29606_, _29605_);
  and (_29607_, _07333_, \uc8051golden_1.PC [14]);
  nor (_29608_, _29607_, _07199_);
  nor (_29609_, _29608_, _29606_);
  nor (_29610_, _29609_, _06790_);
  and (_29611_, _29610_, _29603_);
  nor (_29613_, _29611_, _29600_);
  nor (_29614_, _29613_, _08643_);
  not (_29615_, _29614_);
  and (_29616_, _29615_, _12497_);
  and (_29617_, _29616_, _29595_);
  or (_29618_, _29617_, _29588_);
  and (_29619_, _29618_, _12458_);
  nor (_29620_, _29596_, _12503_);
  or (_29621_, _29620_, _12502_);
  or (_29622_, _29621_, _29619_);
  nor (_29624_, _12455_, _12111_);
  nor (_29625_, _29624_, _12510_);
  nand (_29626_, _29625_, _29622_);
  and (_29627_, _29575_, _12510_);
  nor (_29628_, _29627_, _06406_);
  and (_29629_, _29628_, _29626_);
  or (_29630_, _29629_, _29582_);
  nand (_29631_, _29630_, _12517_);
  nor (_29632_, _29575_, _12517_);
  nor (_29633_, _29632_, _12524_);
  nand (_29635_, _29633_, _29631_);
  nor (_29636_, _12523_, _15722_);
  nor (_29637_, _29636_, _12450_);
  and (_29638_, _29637_, _29635_);
  and (_29639_, _12444_, _12251_);
  not (_29640_, _29584_);
  nor (_29641_, _29640_, _12444_);
  or (_29642_, _29641_, _29639_);
  nor (_29643_, _29642_, _12449_);
  or (_29644_, _29643_, _29638_);
  nand (_29646_, _29644_, _12411_);
  or (_29647_, _12407_, _12252_);
  nand (_29648_, _29584_, _12407_);
  and (_29649_, _29648_, _06457_);
  nand (_29650_, _29649_, _29647_);
  and (_29651_, _29650_, _06842_);
  and (_29652_, _29651_, _29646_);
  and (_29653_, _12546_, _12251_);
  nor (_29654_, _29640_, _12546_);
  nor (_29655_, _29654_, _29653_);
  nor (_29657_, _29655_, _06842_);
  or (_29658_, _29657_, _29652_);
  nand (_29659_, _29658_, _12534_);
  and (_29660_, _12251_, _12249_);
  and (_29661_, _29584_, _26421_);
  or (_29662_, _29661_, _29660_);
  and (_29663_, _29662_, _06482_);
  nor (_29664_, _29663_, _12237_);
  and (_29665_, _29664_, _29659_);
  nor (_29666_, _29575_, _12238_);
  or (_29668_, _29666_, _29665_);
  and (_29669_, _29668_, _12570_);
  nor (_29670_, _12570_, _12111_);
  or (_29671_, _29670_, _29669_);
  nand (_29672_, _29671_, _12576_);
  nor (_29673_, _29575_, _12576_);
  nor (_29674_, _29673_, _12583_);
  nand (_29675_, _29674_, _29672_);
  nor (_29676_, _12582_, _15722_);
  nor (_29677_, _29676_, _12594_);
  nand (_29679_, _29677_, _29675_);
  nor (_29680_, _29575_, _12588_);
  nor (_29681_, _29680_, _12593_);
  nand (_29682_, _29681_, _29679_);
  nor (_29683_, _15722_, _12592_);
  nor (_29684_, _29683_, _06022_);
  nand (_29685_, _29684_, _29682_);
  nor (_29686_, _29575_, _06023_);
  nor (_29687_, _29686_, _12603_);
  nand (_29688_, _29687_, _29685_);
  nor (_29690_, _12602_, _15722_);
  nor (_29691_, _29690_, _06472_);
  nand (_29692_, _29691_, _29688_);
  and (_29693_, _12252_, _06472_);
  nor (_29694_, _29693_, _13788_);
  nand (_29695_, _29694_, _29692_);
  nor (_29696_, _15722_, _06294_);
  nor (_29697_, _29696_, _06015_);
  nand (_29698_, _29697_, _29695_);
  and (_29699_, _12252_, _06015_);
  nor (_29700_, _29699_, _12620_);
  nand (_29701_, _29700_, _29698_);
  and (_29702_, _29575_, _12620_);
  nor (_29703_, _29702_, _12619_);
  nand (_29704_, _29703_, _29701_);
  nor (_29705_, _12618_, _12111_);
  nor (_29706_, _29705_, _12624_);
  and (_29707_, _29706_, _29704_);
  and (_29708_, _29592_, _12624_);
  nor (_29709_, _29708_, _29707_);
  or (_29712_, _29709_, _09013_);
  or (_29713_, _15722_, _09012_);
  and (_29714_, _29713_, _06276_);
  nand (_29715_, _29714_, _29712_);
  and (_29716_, _12252_, _06275_);
  nor (_29717_, _29716_, _10933_);
  nand (_29718_, _29717_, _29715_);
  and (_29719_, _12111_, _10933_);
  nor (_29720_, _29719_, _12639_);
  nand (_29721_, _29720_, _29718_);
  nor (_29723_, _12669_, \uc8051golden_1.DPH [6]);
  nor (_29724_, _29723_, _12670_);
  nor (_29725_, _29724_, _12640_);
  nor (_29726_, _29725_, _12677_);
  and (_29727_, _29726_, _29721_);
  or (_29728_, _29727_, _29581_);
  nand (_29729_, _29728_, _12681_);
  and (_29730_, _12111_, _11297_);
  and (_29731_, _29592_, _12687_);
  or (_29732_, _29731_, _29730_);
  and (_29734_, _29732_, _12680_);
  nor (_29735_, _29734_, _12685_);
  nand (_29736_, _29735_, _29729_);
  nor (_29737_, _29575_, _12233_);
  nor (_29738_, _29737_, _12228_);
  nand (_29739_, _29738_, _29736_);
  nor (_29740_, _15722_, _12227_);
  nor (_29741_, _29740_, _06474_);
  nand (_29742_, _29741_, _29739_);
  and (_29743_, _12252_, _06474_);
  nor (_29745_, _29743_, _12701_);
  and (_29746_, _29745_, _29742_);
  or (_29747_, _29746_, _29580_);
  nand (_29748_, _29747_, _12705_);
  and (_29749_, _12111_, _12687_);
  and (_29750_, _29592_, _11297_);
  or (_29751_, _29750_, _29749_);
  and (_29752_, _29751_, _12704_);
  nor (_29753_, _29752_, _12723_);
  nand (_29754_, _29753_, _29748_);
  nor (_29756_, _29575_, _12719_);
  nor (_29757_, _29756_, _12722_);
  nand (_29758_, _29757_, _29754_);
  nor (_29759_, _15722_, _12721_);
  nor (_29760_, _29759_, _06478_);
  nand (_29761_, _29760_, _29758_);
  and (_29762_, _12252_, _06478_);
  nor (_29763_, _29762_, _12732_);
  and (_29764_, _29763_, _29761_);
  or (_29765_, _29764_, _29578_);
  nand (_29767_, _29765_, _12736_);
  and (_29768_, _12111_, \uc8051golden_1.PSW [7]);
  and (_29769_, _29592_, _10524_);
  or (_29770_, _29769_, _29768_);
  and (_29771_, _29770_, _12735_);
  nor (_29772_, _29771_, _12224_);
  nand (_29773_, _29772_, _29767_);
  and (_29774_, _29596_, _12224_);
  nor (_29775_, _29774_, _11019_);
  nand (_29776_, _29775_, _29773_);
  nor (_29778_, _15722_, _11018_);
  nor (_29779_, _29778_, _06479_);
  nand (_29780_, _29779_, _29776_);
  and (_29781_, _12252_, _06479_);
  nor (_29782_, _29781_, _12753_);
  and (_29783_, _29782_, _29780_);
  or (_29784_, _29783_, _29577_);
  nand (_29785_, _29784_, _12756_);
  and (_29786_, _12111_, _10524_);
  and (_29787_, _29592_, \uc8051golden_1.PSW [7]);
  or (_29789_, _29787_, _29786_);
  and (_29790_, _29789_, _12217_);
  nor (_29791_, _29790_, _12763_);
  nand (_29792_, _29791_, _29785_);
  nor (_29793_, _29575_, _12761_);
  nor (_29794_, _29793_, _11061_);
  nand (_29795_, _29794_, _29792_);
  nor (_29796_, _15722_, _11060_);
  nor (_29797_, _29796_, _11089_);
  nand (_29798_, _29797_, _29795_);
  nor (_29800_, _29575_, _11090_);
  nor (_29801_, _29800_, _06588_);
  and (_29802_, _29801_, _29798_);
  nor (_29803_, _08118_, _13881_);
  or (_29804_, _29803_, _05966_);
  or (_29805_, _29804_, _29802_);
  and (_29806_, _15722_, _05966_);
  nor (_29807_, _29806_, _06460_);
  nand (_29808_, _29807_, _29805_);
  and (_29809_, _29640_, _12958_);
  nor (_29811_, _12251_, _12958_);
  or (_29812_, _29811_, _06596_);
  or (_29813_, _29812_, _29809_);
  and (_29814_, _29813_, _12108_);
  nand (_29815_, _29814_, _29808_);
  nor (_29816_, _29575_, _12108_);
  nor (_29817_, _29816_, _12094_);
  nand (_29818_, _29817_, _29815_);
  nor (_29819_, _15722_, _11204_);
  nor (_29820_, _29819_, _11243_);
  and (_29822_, _29820_, _29818_);
  or (_29823_, _29822_, _29576_);
  nand (_29824_, _29823_, _06306_);
  and (_29825_, _08118_, _06305_);
  nor (_29826_, _29825_, _05971_);
  and (_29827_, _29826_, _29824_);
  and (_29828_, _12111_, _05971_);
  or (_29829_, _29828_, _06487_);
  nor (_29830_, _29829_, _29827_);
  and (_29831_, _12252_, _12958_);
  nor (_29833_, _29584_, _12958_);
  nor (_29834_, _29833_, _29831_);
  nor (_29835_, _29834_, _12978_);
  or (_29836_, _29835_, _29830_);
  and (_29837_, _29836_, _12987_);
  nor (_29838_, _29575_, _12987_);
  or (_29839_, _29838_, _29837_);
  nand (_29840_, _29839_, _07037_);
  nand (_29841_, _15722_, _06606_);
  and (_29842_, _29841_, _12994_);
  nand (_29844_, _29842_, _29840_);
  and (_29845_, _29575_, _12995_);
  nor (_29846_, _29845_, _06465_);
  nand (_29847_, _29846_, _29844_);
  and (_29848_, _06465_, _06340_);
  nor (_29849_, _29848_, _05969_);
  nand (_29850_, _29849_, _29847_);
  and (_29851_, _12111_, _05969_);
  nor (_29852_, _29851_, _06234_);
  nand (_29853_, _29852_, _29850_);
  nor (_29855_, _29834_, _06807_);
  nor (_29856_, _29855_, _13012_);
  nand (_29857_, _29856_, _29853_);
  and (_29858_, _29575_, _13012_);
  nor (_29859_, _29858_, _06195_);
  nand (_29860_, _29859_, _29857_);
  and (_29861_, _15722_, _06195_);
  nor (_29862_, _29861_, _13020_);
  nand (_29863_, _29862_, _29860_);
  and (_29864_, _29575_, _13020_);
  nor (_29866_, _29864_, _06475_);
  and (_29867_, _29866_, _29863_);
  and (_29868_, _06475_, _06340_);
  or (_29869_, _29868_, _05963_);
  nor (_29870_, _29869_, _29867_);
  and (_29871_, _12111_, _05963_);
  or (_29872_, _29871_, _13030_);
  nor (_29873_, _29872_, _29870_);
  nor (_29874_, _29575_, _13031_);
  nor (_29875_, _29874_, _29873_);
  or (_29877_, _29875_, _01379_);
  or (_29878_, _01375_, \uc8051golden_1.PC [14]);
  and (_29879_, _29878_, _42545_);
  and (_42992_, _29879_, _29877_);
  nand (_29880_, _11225_, _07931_);
  and (_29881_, _13040_, \uc8051golden_1.P2 [0]);
  nor (_29882_, _29881_, _07276_);
  nand (_29883_, _29882_, _29880_);
  and (_29884_, _07931_, _07473_);
  or (_29885_, _29884_, _29881_);
  or (_29887_, _29885_, _06293_);
  nor (_29888_, _08521_, _13040_);
  or (_29889_, _29888_, _29881_);
  or (_29890_, _29889_, _07210_);
  and (_29891_, _07931_, \uc8051golden_1.ACC [0]);
  or (_29892_, _29891_, _29881_);
  and (_29893_, _29892_, _07199_);
  and (_29894_, _07200_, \uc8051golden_1.P2 [0]);
  or (_29895_, _29894_, _06401_);
  or (_29896_, _29895_, _29893_);
  and (_29898_, _29896_, _06396_);
  and (_29899_, _29898_, _29890_);
  and (_29900_, _13048_, \uc8051golden_1.P2 [0]);
  and (_29901_, _14339_, _08608_);
  or (_29902_, _29901_, _29900_);
  and (_29903_, _29902_, _06395_);
  or (_29904_, _29903_, _29899_);
  and (_29905_, _29904_, _07221_);
  and (_29906_, _29885_, _06399_);
  or (_29907_, _29906_, _06406_);
  or (_29909_, _29907_, _29905_);
  or (_29910_, _29892_, _06414_);
  and (_29911_, _29910_, _06844_);
  and (_29912_, _29911_, _29909_);
  and (_29913_, _29881_, _06393_);
  or (_29914_, _29913_, _06387_);
  or (_29915_, _29914_, _29912_);
  or (_29916_, _29889_, _07245_);
  and (_29917_, _29916_, _06446_);
  and (_29918_, _29917_, _29915_);
  and (_29920_, _14371_, _08608_);
  or (_29921_, _29920_, _29900_);
  and (_29922_, _29921_, _06300_);
  or (_29923_, _29922_, _10059_);
  or (_29924_, _29923_, _29918_);
  and (_29925_, _29924_, _29887_);
  or (_29926_, _29925_, _06281_);
  and (_29927_, _07931_, _09446_);
  or (_29928_, _29881_, _06282_);
  or (_29929_, _29928_, _29927_);
  and (_29931_, _29929_, _29926_);
  or (_29932_, _29931_, _06015_);
  and (_29933_, _14426_, _07931_);
  or (_29934_, _29881_, _06279_);
  or (_29935_, _29934_, _29933_);
  and (_29936_, _29935_, _06276_);
  and (_29937_, _29936_, _29932_);
  and (_29938_, _07931_, _08817_);
  or (_29939_, _29938_, _29881_);
  and (_29940_, _29939_, _06275_);
  or (_29942_, _29940_, _06474_);
  or (_29943_, _29942_, _29937_);
  and (_29944_, _14324_, _07931_);
  or (_29945_, _29944_, _29881_);
  or (_29946_, _29945_, _07282_);
  and (_29947_, _29946_, _07284_);
  and (_29948_, _29947_, _29943_);
  nor (_29949_, _12538_, _13040_);
  or (_29950_, _29949_, _29881_);
  and (_29951_, _29880_, _06582_);
  and (_29953_, _29951_, _29950_);
  or (_29954_, _29953_, _29948_);
  and (_29955_, _29954_, _07279_);
  nand (_29956_, _29939_, _06478_);
  nor (_29957_, _29956_, _29888_);
  or (_29958_, _29957_, _06569_);
  or (_29959_, _29958_, _29955_);
  and (_29960_, _29959_, _29883_);
  or (_29961_, _29960_, _06479_);
  and (_29962_, _14320_, _07931_);
  or (_29964_, _29881_, _09043_);
  or (_29965_, _29964_, _29962_);
  and (_29966_, _29965_, _09048_);
  and (_29967_, _29966_, _29961_);
  and (_29968_, _29950_, _06572_);
  or (_29969_, _29968_, _06606_);
  or (_29970_, _29969_, _29967_);
  or (_29971_, _29889_, _07037_);
  and (_29972_, _29971_, _29970_);
  or (_29973_, _29972_, _06234_);
  or (_29975_, _29881_, _06807_);
  and (_29976_, _29975_, _29973_);
  or (_29977_, _29976_, _06195_);
  or (_29978_, _29889_, _06196_);
  and (_29979_, _29978_, _01375_);
  and (_29980_, _29979_, _29977_);
  nor (_29981_, \uc8051golden_1.P2 [0], rst);
  nor (_29982_, _29981_, _01382_);
  or (_42993_, _29982_, _29980_);
  and (_29983_, _13040_, \uc8051golden_1.P2 [1]);
  nor (_29985_, _11223_, _13040_);
  or (_29986_, _29985_, _29983_);
  or (_29987_, _29986_, _09048_);
  nand (_29988_, _07931_, _07090_);
  or (_29989_, _07931_, \uc8051golden_1.P2 [1]);
  and (_29990_, _29989_, _06275_);
  and (_29991_, _29990_, _29988_);
  nor (_29992_, _13040_, _07196_);
  or (_29993_, _29992_, _29983_);
  or (_29994_, _29993_, _07221_);
  and (_29996_, _14532_, _07931_);
  not (_29997_, _29996_);
  and (_29998_, _29997_, _29989_);
  or (_29999_, _29998_, _07210_);
  and (_30000_, _07931_, \uc8051golden_1.ACC [1]);
  or (_30001_, _30000_, _29983_);
  and (_30002_, _30001_, _07199_);
  and (_30003_, _07200_, \uc8051golden_1.P2 [1]);
  or (_30004_, _30003_, _06401_);
  or (_30005_, _30004_, _30002_);
  and (_30007_, _30005_, _06396_);
  and (_30008_, _30007_, _29999_);
  and (_30009_, _13048_, \uc8051golden_1.P2 [1]);
  and (_30010_, _14514_, _08608_);
  or (_30011_, _30010_, _30009_);
  and (_30012_, _30011_, _06395_);
  or (_30013_, _30012_, _06399_);
  or (_30014_, _30013_, _30008_);
  and (_30015_, _30014_, _29994_);
  or (_30016_, _30015_, _06406_);
  or (_30018_, _30001_, _06414_);
  and (_30019_, _30018_, _06844_);
  and (_30020_, _30019_, _30016_);
  and (_30021_, _14517_, _08608_);
  or (_30022_, _30021_, _30009_);
  and (_30023_, _30022_, _06393_);
  or (_30024_, _30023_, _06387_);
  or (_30025_, _30024_, _30020_);
  and (_30026_, _30010_, _14513_);
  or (_30027_, _30009_, _07245_);
  or (_30029_, _30027_, _30026_);
  and (_30030_, _30029_, _06446_);
  and (_30031_, _30030_, _30025_);
  or (_30032_, _30009_, _14560_);
  and (_30033_, _30032_, _06300_);
  and (_30034_, _30033_, _30011_);
  or (_30035_, _30034_, _10059_);
  or (_30036_, _30035_, _30031_);
  or (_30037_, _29993_, _06293_);
  and (_30038_, _30037_, _30036_);
  or (_30040_, _30038_, _06281_);
  and (_30041_, _07931_, _09445_);
  or (_30042_, _29983_, _06282_);
  or (_30043_, _30042_, _30041_);
  and (_30044_, _30043_, _06279_);
  and (_30045_, _30044_, _30040_);
  and (_30046_, _14615_, _07931_);
  or (_30047_, _30046_, _29983_);
  and (_30048_, _30047_, _06015_);
  or (_30049_, _30048_, _30045_);
  and (_30051_, _30049_, _06276_);
  or (_30052_, _30051_, _29991_);
  and (_30053_, _30052_, _07282_);
  or (_30054_, _14507_, _13040_);
  and (_30055_, _29989_, _06474_);
  and (_30056_, _30055_, _30054_);
  or (_30057_, _30056_, _06582_);
  or (_30058_, _30057_, _30053_);
  nand (_30059_, _11222_, _07931_);
  and (_30060_, _30059_, _29986_);
  or (_30062_, _30060_, _07284_);
  and (_30063_, _30062_, _07279_);
  and (_30064_, _30063_, _30058_);
  or (_30065_, _14505_, _13040_);
  and (_30066_, _29989_, _06478_);
  and (_30067_, _30066_, _30065_);
  or (_30068_, _30067_, _06569_);
  or (_30069_, _30068_, _30064_);
  nor (_30070_, _29983_, _07276_);
  nand (_30071_, _30070_, _30059_);
  and (_30073_, _30071_, _09043_);
  and (_30074_, _30073_, _30069_);
  or (_30075_, _29988_, _08477_);
  and (_30076_, _29989_, _06479_);
  and (_30077_, _30076_, _30075_);
  or (_30078_, _30077_, _06572_);
  or (_30079_, _30078_, _30074_);
  and (_30080_, _30079_, _29987_);
  or (_30081_, _30080_, _06606_);
  or (_30082_, _29998_, _07037_);
  and (_30084_, _30082_, _06807_);
  and (_30085_, _30084_, _30081_);
  and (_30086_, _30022_, _06234_);
  or (_30087_, _30086_, _06195_);
  or (_30088_, _30087_, _30085_);
  or (_30089_, _29983_, _06196_);
  or (_30090_, _30089_, _29996_);
  and (_30091_, _30090_, _01375_);
  and (_30092_, _30091_, _30088_);
  nor (_30093_, \uc8051golden_1.P2 [1], rst);
  nor (_30095_, _30093_, _01382_);
  or (_42994_, _30095_, _30092_);
  and (_30096_, _13040_, \uc8051golden_1.P2 [2]);
  nor (_30097_, _13040_, _07623_);
  or (_30098_, _30097_, _30096_);
  or (_30099_, _30098_, _06293_);
  or (_30100_, _30098_, _07221_);
  and (_30101_, _14754_, _07931_);
  or (_30102_, _30101_, _30096_);
  or (_30103_, _30102_, _07210_);
  and (_30105_, _07931_, \uc8051golden_1.ACC [2]);
  or (_30106_, _30105_, _30096_);
  and (_30107_, _30106_, _07199_);
  and (_30108_, _07200_, \uc8051golden_1.P2 [2]);
  or (_30109_, _30108_, _06401_);
  or (_30110_, _30109_, _30107_);
  and (_30111_, _30110_, _06396_);
  and (_30112_, _30111_, _30103_);
  and (_30113_, _13048_, \uc8051golden_1.P2 [2]);
  and (_30114_, _14751_, _08608_);
  or (_30116_, _30114_, _30113_);
  and (_30117_, _30116_, _06395_);
  or (_30118_, _30117_, _06399_);
  or (_30119_, _30118_, _30112_);
  and (_30120_, _30119_, _30100_);
  or (_30121_, _30120_, _06406_);
  or (_30122_, _30106_, _06414_);
  and (_30123_, _30122_, _06844_);
  and (_30124_, _30123_, _30121_);
  and (_30125_, _14749_, _08608_);
  or (_30127_, _30125_, _30113_);
  and (_30128_, _30127_, _06393_);
  or (_30129_, _30128_, _06387_);
  or (_30130_, _30129_, _30124_);
  and (_30131_, _30114_, _14778_);
  or (_30132_, _30113_, _07245_);
  or (_30133_, _30132_, _30131_);
  and (_30134_, _30133_, _06446_);
  and (_30135_, _30134_, _30130_);
  and (_30136_, _14793_, _08608_);
  or (_30138_, _30136_, _30113_);
  and (_30139_, _30138_, _06300_);
  or (_30140_, _30139_, _10059_);
  or (_30141_, _30140_, _30135_);
  and (_30142_, _30141_, _30099_);
  or (_30143_, _30142_, _06281_);
  and (_30144_, _07931_, _09444_);
  or (_30145_, _30096_, _06282_);
  or (_30146_, _30145_, _30144_);
  and (_30147_, _30146_, _06279_);
  and (_30149_, _30147_, _30143_);
  and (_30150_, _14848_, _07931_);
  or (_30151_, _30150_, _30096_);
  and (_30152_, _30151_, _06015_);
  or (_30153_, _30152_, _06275_);
  or (_30154_, _30153_, _30149_);
  and (_30155_, _07931_, _08994_);
  or (_30156_, _30155_, _30096_);
  or (_30157_, _30156_, _06276_);
  and (_30158_, _30157_, _30154_);
  or (_30160_, _30158_, _06474_);
  and (_30161_, _14744_, _07931_);
  or (_30162_, _30161_, _30096_);
  or (_30163_, _30162_, _07282_);
  and (_30164_, _30163_, _07284_);
  and (_30165_, _30164_, _30160_);
  and (_30166_, _11221_, _07931_);
  or (_30167_, _30166_, _30096_);
  and (_30168_, _30167_, _06582_);
  or (_30169_, _30168_, _30165_);
  and (_30171_, _30169_, _07279_);
  or (_30172_, _30096_, _08433_);
  and (_30173_, _30156_, _06478_);
  and (_30174_, _30173_, _30172_);
  or (_30175_, _30174_, _30171_);
  and (_30176_, _30175_, _07276_);
  and (_30177_, _30106_, _06569_);
  and (_30178_, _30177_, _30172_);
  or (_30179_, _30178_, _06479_);
  or (_30180_, _30179_, _30176_);
  and (_30182_, _14741_, _07931_);
  or (_30183_, _30096_, _09043_);
  or (_30184_, _30183_, _30182_);
  and (_30185_, _30184_, _09048_);
  and (_30186_, _30185_, _30180_);
  nor (_30187_, _11220_, _13040_);
  or (_30188_, _30187_, _30096_);
  and (_30189_, _30188_, _06572_);
  or (_30190_, _30189_, _06606_);
  or (_30191_, _30190_, _30186_);
  or (_30193_, _30102_, _07037_);
  and (_30194_, _30193_, _06807_);
  and (_30195_, _30194_, _30191_);
  and (_30196_, _30127_, _06234_);
  or (_30197_, _30196_, _06195_);
  or (_30198_, _30197_, _30195_);
  and (_30199_, _14917_, _07931_);
  or (_30200_, _30096_, _06196_);
  or (_30201_, _30200_, _30199_);
  and (_30202_, _30201_, _01375_);
  and (_30204_, _30202_, _30198_);
  nor (_30205_, \uc8051golden_1.P2 [2], rst);
  nor (_30206_, _30205_, _01382_);
  or (_42995_, _30206_, _30204_);
  and (_30207_, _13040_, \uc8051golden_1.P2 [3]);
  nor (_30208_, _13040_, _07775_);
  or (_30209_, _30208_, _30207_);
  or (_30210_, _30209_, _06293_);
  and (_30211_, _14947_, _07931_);
  or (_30212_, _30211_, _30207_);
  or (_30214_, _30212_, _07210_);
  and (_30215_, _07931_, \uc8051golden_1.ACC [3]);
  or (_30216_, _30215_, _30207_);
  and (_30217_, _30216_, _07199_);
  and (_30218_, _07200_, \uc8051golden_1.P2 [3]);
  or (_30219_, _30218_, _06401_);
  or (_30220_, _30219_, _30217_);
  and (_30221_, _30220_, _06396_);
  and (_30222_, _30221_, _30214_);
  and (_30223_, _13048_, \uc8051golden_1.P2 [3]);
  and (_30225_, _14951_, _08608_);
  or (_30226_, _30225_, _30223_);
  and (_30227_, _30226_, _06395_);
  or (_30228_, _30227_, _06399_);
  or (_30229_, _30228_, _30222_);
  or (_30230_, _30209_, _07221_);
  and (_30231_, _30230_, _30229_);
  or (_30232_, _30231_, _06406_);
  or (_30233_, _30216_, _06414_);
  and (_30234_, _30233_, _06844_);
  and (_30236_, _30234_, _30232_);
  and (_30237_, _14961_, _08608_);
  or (_30238_, _30237_, _30223_);
  and (_30239_, _30238_, _06393_);
  or (_30240_, _30239_, _06387_);
  or (_30241_, _30240_, _30236_);
  or (_30242_, _30223_, _14968_);
  and (_30243_, _30242_, _30226_);
  or (_30244_, _30243_, _07245_);
  and (_30245_, _30244_, _06446_);
  and (_30247_, _30245_, _30241_);
  and (_30248_, _14985_, _08608_);
  or (_30249_, _30248_, _30223_);
  and (_30250_, _30249_, _06300_);
  or (_30251_, _30250_, _10059_);
  or (_30252_, _30251_, _30247_);
  and (_30253_, _30252_, _30210_);
  or (_30254_, _30253_, _06281_);
  and (_30255_, _07931_, _09443_);
  or (_30256_, _30207_, _06282_);
  or (_30258_, _30256_, _30255_);
  and (_30259_, _30258_, _06279_);
  and (_30260_, _30259_, _30254_);
  and (_30261_, _15039_, _07931_);
  or (_30262_, _30261_, _30207_);
  and (_30263_, _30262_, _06015_);
  or (_30264_, _30263_, _06275_);
  or (_30265_, _30264_, _30260_);
  and (_30266_, _07931_, _08815_);
  or (_30267_, _30266_, _30207_);
  or (_30269_, _30267_, _06276_);
  and (_30270_, _30269_, _30265_);
  or (_30271_, _30270_, _06474_);
  and (_30272_, _14934_, _07931_);
  or (_30273_, _30272_, _30207_);
  or (_30274_, _30273_, _07282_);
  and (_30275_, _30274_, _07284_);
  and (_30276_, _30275_, _30271_);
  and (_30277_, _12535_, _07931_);
  or (_30278_, _30277_, _30207_);
  and (_30280_, _30278_, _06582_);
  or (_30281_, _30280_, _30276_);
  and (_30282_, _30281_, _07279_);
  or (_30283_, _30207_, _08389_);
  and (_30284_, _30267_, _06478_);
  and (_30285_, _30284_, _30283_);
  or (_30286_, _30285_, _30282_);
  and (_30287_, _30286_, _07276_);
  and (_30288_, _30216_, _06569_);
  and (_30289_, _30288_, _30283_);
  or (_30291_, _30289_, _06479_);
  or (_30292_, _30291_, _30287_);
  and (_30293_, _14931_, _07931_);
  or (_30294_, _30207_, _09043_);
  or (_30295_, _30294_, _30293_);
  and (_30296_, _30295_, _09048_);
  and (_30297_, _30296_, _30292_);
  nor (_30298_, _11218_, _13040_);
  or (_30299_, _30298_, _30207_);
  and (_30300_, _30299_, _06572_);
  or (_30302_, _30300_, _06606_);
  or (_30303_, _30302_, _30297_);
  or (_30304_, _30212_, _07037_);
  and (_30305_, _30304_, _06807_);
  and (_30306_, _30305_, _30303_);
  and (_30307_, _30238_, _06234_);
  or (_30308_, _30307_, _06195_);
  or (_30309_, _30308_, _30306_);
  and (_30310_, _15113_, _07931_);
  or (_30311_, _30207_, _06196_);
  or (_30313_, _30311_, _30310_);
  and (_30314_, _30313_, _01375_);
  and (_30315_, _30314_, _30309_);
  nor (_30316_, \uc8051golden_1.P2 [3], rst);
  nor (_30317_, _30316_, _01382_);
  or (_42996_, _30317_, _30315_);
  and (_30318_, _13040_, \uc8051golden_1.P2 [4]);
  nor (_30319_, _13040_, _08301_);
  or (_30320_, _30319_, _30318_);
  or (_30321_, _30320_, _06293_);
  and (_30322_, _15130_, _07931_);
  or (_30323_, _30322_, _30318_);
  or (_30324_, _30323_, _07210_);
  and (_30325_, _07931_, \uc8051golden_1.ACC [4]);
  or (_30326_, _30325_, _30318_);
  and (_30327_, _30326_, _07199_);
  and (_30328_, _07200_, \uc8051golden_1.P2 [4]);
  or (_30329_, _30328_, _06401_);
  or (_30330_, _30329_, _30327_);
  and (_30331_, _30330_, _06396_);
  and (_30334_, _30331_, _30324_);
  and (_30335_, _13048_, \uc8051golden_1.P2 [4]);
  and (_30336_, _15139_, _08608_);
  or (_30337_, _30336_, _30335_);
  and (_30338_, _30337_, _06395_);
  or (_30339_, _30338_, _06399_);
  or (_30340_, _30339_, _30334_);
  or (_30341_, _30320_, _07221_);
  and (_30342_, _30341_, _30340_);
  or (_30343_, _30342_, _06406_);
  or (_30345_, _30326_, _06414_);
  and (_30346_, _30345_, _06844_);
  and (_30347_, _30346_, _30343_);
  and (_30348_, _15168_, _08608_);
  or (_30349_, _30348_, _30335_);
  and (_30350_, _30349_, _06393_);
  or (_30351_, _30350_, _06387_);
  or (_30352_, _30351_, _30347_);
  or (_30353_, _30335_, _15138_);
  and (_30354_, _30353_, _30337_);
  or (_30356_, _30354_, _07245_);
  and (_30357_, _30356_, _06446_);
  and (_30358_, _30357_, _30352_);
  and (_30359_, _15189_, _08608_);
  or (_30360_, _30359_, _30335_);
  and (_30361_, _30360_, _06300_);
  or (_30362_, _30361_, _10059_);
  or (_30363_, _30362_, _30358_);
  and (_30364_, _30363_, _30321_);
  or (_30365_, _30364_, _06281_);
  and (_30367_, _07931_, _09442_);
  or (_30368_, _30318_, _06282_);
  or (_30369_, _30368_, _30367_);
  and (_30370_, _30369_, _06279_);
  and (_30371_, _30370_, _30365_);
  and (_30372_, _15243_, _07931_);
  or (_30373_, _30372_, _30318_);
  and (_30374_, _30373_, _06015_);
  or (_30375_, _30374_, _06275_);
  or (_30376_, _30375_, _30371_);
  and (_30378_, _08883_, _07931_);
  or (_30379_, _30378_, _30318_);
  or (_30380_, _30379_, _06276_);
  and (_30381_, _30380_, _30376_);
  or (_30382_, _30381_, _06474_);
  and (_30383_, _15135_, _07931_);
  or (_30384_, _30383_, _30318_);
  or (_30385_, _30384_, _07282_);
  and (_30386_, _30385_, _07284_);
  and (_30387_, _30386_, _30382_);
  and (_30389_, _11216_, _07931_);
  or (_30390_, _30389_, _30318_);
  and (_30391_, _30390_, _06582_);
  or (_30392_, _30391_, _30387_);
  and (_30393_, _30392_, _07279_);
  or (_30394_, _30318_, _08345_);
  and (_30395_, _30379_, _06478_);
  and (_30396_, _30395_, _30394_);
  or (_30397_, _30396_, _30393_);
  and (_30398_, _30397_, _07276_);
  and (_30400_, _30326_, _06569_);
  and (_30401_, _30400_, _30394_);
  or (_30402_, _30401_, _06479_);
  or (_30403_, _30402_, _30398_);
  and (_30404_, _15134_, _07931_);
  or (_30405_, _30318_, _09043_);
  or (_30406_, _30405_, _30404_);
  and (_30407_, _30406_, _09048_);
  and (_30408_, _30407_, _30403_);
  nor (_30409_, _11215_, _13040_);
  or (_30411_, _30409_, _30318_);
  and (_30412_, _30411_, _06572_);
  or (_30413_, _30412_, _06606_);
  or (_30414_, _30413_, _30408_);
  or (_30415_, _30323_, _07037_);
  and (_30416_, _30415_, _06807_);
  and (_30417_, _30416_, _30414_);
  and (_30418_, _30349_, _06234_);
  or (_30419_, _30418_, _06195_);
  or (_30420_, _30419_, _30417_);
  and (_30422_, _15315_, _07931_);
  or (_30423_, _30318_, _06196_);
  or (_30424_, _30423_, _30422_);
  and (_30425_, _30424_, _01375_);
  and (_30426_, _30425_, _30420_);
  nor (_30427_, \uc8051golden_1.P2 [4], rst);
  nor (_30428_, _30427_, _01382_);
  or (_42997_, _30428_, _30426_);
  and (_30429_, _13040_, \uc8051golden_1.P2 [5]);
  nor (_30430_, _13040_, _08207_);
  or (_30432_, _30430_, _30429_);
  or (_30433_, _30432_, _06293_);
  and (_30434_, _15348_, _07931_);
  or (_30435_, _30434_, _30429_);
  or (_30436_, _30435_, _07210_);
  and (_30437_, _07931_, \uc8051golden_1.ACC [5]);
  or (_30438_, _30437_, _30429_);
  and (_30439_, _30438_, _07199_);
  and (_30440_, _07200_, \uc8051golden_1.P2 [5]);
  or (_30441_, _30440_, _06401_);
  or (_30443_, _30441_, _30439_);
  and (_30444_, _30443_, _06396_);
  and (_30445_, _30444_, _30436_);
  and (_30446_, _13048_, \uc8051golden_1.P2 [5]);
  and (_30447_, _15341_, _08608_);
  or (_30448_, _30447_, _30446_);
  and (_30449_, _30448_, _06395_);
  or (_30450_, _30449_, _06399_);
  or (_30451_, _30450_, _30445_);
  or (_30452_, _30432_, _07221_);
  and (_30454_, _30452_, _30451_);
  or (_30455_, _30454_, _06406_);
  or (_30456_, _30438_, _06414_);
  and (_30457_, _30456_, _06844_);
  and (_30458_, _30457_, _30455_);
  and (_30459_, _15345_, _08608_);
  or (_30460_, _30459_, _30446_);
  and (_30461_, _30460_, _06393_);
  or (_30462_, _30461_, _06387_);
  or (_30463_, _30462_, _30458_);
  or (_30465_, _30446_, _15378_);
  and (_30466_, _30465_, _30448_);
  or (_30467_, _30466_, _07245_);
  and (_30468_, _30467_, _06446_);
  and (_30469_, _30468_, _30463_);
  or (_30470_, _30446_, _15342_);
  and (_30471_, _30470_, _06300_);
  and (_30472_, _30471_, _30448_);
  or (_30473_, _30472_, _10059_);
  or (_30474_, _30473_, _30469_);
  and (_30476_, _30474_, _30433_);
  or (_30477_, _30476_, _06281_);
  and (_30478_, _07931_, _09441_);
  or (_30479_, _30429_, _06282_);
  or (_30480_, _30479_, _30478_);
  and (_30481_, _30480_, _06279_);
  and (_30482_, _30481_, _30477_);
  and (_30483_, _15446_, _07931_);
  or (_30484_, _30483_, _30429_);
  and (_30485_, _30484_, _06015_);
  or (_30487_, _30485_, _06275_);
  or (_30488_, _30487_, _30482_);
  and (_30489_, _08958_, _07931_);
  or (_30490_, _30489_, _30429_);
  or (_30491_, _30490_, _06276_);
  and (_30492_, _30491_, _30488_);
  or (_30493_, _30492_, _06474_);
  and (_30494_, _15338_, _07931_);
  or (_30495_, _30494_, _30429_);
  or (_30496_, _30495_, _07282_);
  and (_30498_, _30496_, _07284_);
  and (_30499_, _30498_, _30493_);
  and (_30500_, _12542_, _07931_);
  or (_30501_, _30500_, _30429_);
  and (_30502_, _30501_, _06582_);
  or (_30503_, _30502_, _30499_);
  and (_30504_, _30503_, _07279_);
  or (_30505_, _30429_, _08256_);
  and (_30506_, _30490_, _06478_);
  and (_30507_, _30506_, _30505_);
  or (_30509_, _30507_, _30504_);
  and (_30510_, _30509_, _07276_);
  and (_30511_, _30438_, _06569_);
  and (_30512_, _30511_, _30505_);
  or (_30513_, _30512_, _06479_);
  or (_30514_, _30513_, _30510_);
  and (_30515_, _15335_, _07931_);
  or (_30516_, _30429_, _09043_);
  or (_30517_, _30516_, _30515_);
  and (_30518_, _30517_, _09048_);
  and (_30520_, _30518_, _30514_);
  nor (_30521_, _11212_, _13040_);
  or (_30522_, _30521_, _30429_);
  and (_30523_, _30522_, _06572_);
  or (_30524_, _30523_, _06606_);
  or (_30525_, _30524_, _30520_);
  or (_30526_, _30435_, _07037_);
  and (_30527_, _30526_, _06807_);
  and (_30528_, _30527_, _30525_);
  and (_30529_, _30460_, _06234_);
  or (_30531_, _30529_, _06195_);
  or (_30532_, _30531_, _30528_);
  and (_30533_, _15509_, _07931_);
  or (_30534_, _30429_, _06196_);
  or (_30535_, _30534_, _30533_);
  and (_30536_, _30535_, _01375_);
  and (_30537_, _30536_, _30532_);
  nor (_30538_, \uc8051golden_1.P2 [5], rst);
  nor (_30539_, _30538_, _01382_);
  or (_42998_, _30539_, _30537_);
  and (_30541_, _13040_, \uc8051golden_1.P2 [6]);
  nor (_30542_, _13040_, _08118_);
  or (_30543_, _30542_, _30541_);
  or (_30544_, _30543_, _06293_);
  and (_30545_, _15550_, _07931_);
  or (_30546_, _30545_, _30541_);
  or (_30547_, _30546_, _07210_);
  and (_30548_, _07931_, \uc8051golden_1.ACC [6]);
  or (_30549_, _30548_, _30541_);
  and (_30550_, _30549_, _07199_);
  and (_30552_, _07200_, \uc8051golden_1.P2 [6]);
  or (_30553_, _30552_, _06401_);
  or (_30554_, _30553_, _30550_);
  and (_30555_, _30554_, _06396_);
  and (_30556_, _30555_, _30547_);
  and (_30557_, _13048_, \uc8051golden_1.P2 [6]);
  and (_30558_, _15535_, _08608_);
  or (_30559_, _30558_, _30557_);
  and (_30560_, _30559_, _06395_);
  or (_30561_, _30560_, _06399_);
  or (_30563_, _30561_, _30556_);
  or (_30564_, _30543_, _07221_);
  and (_30565_, _30564_, _30563_);
  or (_30566_, _30565_, _06406_);
  or (_30567_, _30549_, _06414_);
  and (_30568_, _30567_, _06844_);
  and (_30569_, _30568_, _30566_);
  and (_30570_, _15561_, _08608_);
  or (_30571_, _30570_, _30557_);
  and (_30572_, _30571_, _06393_);
  or (_30574_, _30572_, _06387_);
  or (_30575_, _30574_, _30569_);
  or (_30576_, _30557_, _15568_);
  and (_30577_, _30576_, _30559_);
  or (_30578_, _30577_, _07245_);
  and (_30579_, _30578_, _06446_);
  and (_30580_, _30579_, _30575_);
  and (_30581_, _15585_, _08608_);
  or (_30582_, _30581_, _30557_);
  and (_30583_, _30582_, _06300_);
  or (_30585_, _30583_, _10059_);
  or (_30586_, _30585_, _30580_);
  and (_30587_, _30586_, _30544_);
  or (_30588_, _30587_, _06281_);
  and (_30589_, _07931_, _09440_);
  or (_30590_, _30541_, _06282_);
  or (_30591_, _30590_, _30589_);
  and (_30592_, _30591_, _06279_);
  and (_30593_, _30592_, _30588_);
  and (_30594_, _15639_, _07931_);
  or (_30596_, _30594_, _30541_);
  and (_30597_, _30596_, _06015_);
  or (_30598_, _30597_, _06275_);
  or (_30599_, _30598_, _30593_);
  and (_30600_, _15646_, _07931_);
  or (_30601_, _30600_, _30541_);
  or (_30602_, _30601_, _06276_);
  and (_30603_, _30602_, _30599_);
  or (_30604_, _30603_, _06474_);
  and (_30605_, _15531_, _07931_);
  or (_30607_, _30605_, _30541_);
  or (_30608_, _30607_, _07282_);
  and (_30609_, _30608_, _07284_);
  and (_30610_, _30609_, _30604_);
  and (_30611_, _11210_, _07931_);
  or (_30612_, _30611_, _30541_);
  and (_30613_, _30612_, _06582_);
  or (_30614_, _30613_, _30610_);
  and (_30615_, _30614_, _07279_);
  or (_30616_, _30541_, _08162_);
  and (_30618_, _30601_, _06478_);
  and (_30619_, _30618_, _30616_);
  or (_30620_, _30619_, _30615_);
  and (_30621_, _30620_, _07276_);
  and (_30622_, _30549_, _06569_);
  and (_30623_, _30622_, _30616_);
  or (_30624_, _30623_, _06479_);
  or (_30625_, _30624_, _30621_);
  and (_30626_, _15528_, _07931_);
  or (_30627_, _30541_, _09043_);
  or (_30629_, _30627_, _30626_);
  and (_30630_, _30629_, _09048_);
  and (_30631_, _30630_, _30625_);
  nor (_30632_, _11209_, _13040_);
  or (_30633_, _30632_, _30541_);
  and (_30634_, _30633_, _06572_);
  or (_30635_, _30634_, _06606_);
  or (_30636_, _30635_, _30631_);
  or (_30637_, _30546_, _07037_);
  and (_30638_, _30637_, _06807_);
  and (_30640_, _30638_, _30636_);
  and (_30641_, _30571_, _06234_);
  or (_30642_, _30641_, _06195_);
  or (_30643_, _30642_, _30640_);
  and (_30644_, _15713_, _07931_);
  or (_30645_, _30541_, _06196_);
  or (_30646_, _30645_, _30644_);
  and (_30647_, _30646_, _01375_);
  and (_30648_, _30647_, _30643_);
  nor (_30649_, \uc8051golden_1.P2 [6], rst);
  nor (_30651_, _30649_, _01382_);
  or (_42999_, _30651_, _30648_);
  and (_30652_, _07945_, \uc8051golden_1.ACC [0]);
  and (_30653_, _30652_, _08521_);
  and (_30654_, _13143_, \uc8051golden_1.P3 [0]);
  or (_30655_, _30654_, _07276_);
  or (_30656_, _30655_, _30653_);
  and (_30657_, _07945_, _07473_);
  or (_30658_, _30657_, _30654_);
  or (_30659_, _30658_, _06293_);
  nor (_30661_, _08521_, _13143_);
  or (_30662_, _30661_, _30654_);
  or (_30663_, _30662_, _07210_);
  or (_30664_, _30652_, _30654_);
  and (_30665_, _30664_, _07199_);
  and (_30666_, _07200_, \uc8051golden_1.P3 [0]);
  or (_30667_, _30666_, _06401_);
  or (_30668_, _30667_, _30665_);
  and (_30669_, _30668_, _06396_);
  and (_30670_, _30669_, _30663_);
  and (_30672_, _13151_, \uc8051golden_1.P3 [0]);
  and (_30673_, _14339_, _08598_);
  or (_30674_, _30673_, _30672_);
  and (_30675_, _30674_, _06395_);
  or (_30676_, _30675_, _30670_);
  and (_30677_, _30676_, _07221_);
  and (_30678_, _30658_, _06399_);
  or (_30679_, _30678_, _06406_);
  or (_30680_, _30679_, _30677_);
  or (_30681_, _30664_, _06414_);
  and (_30683_, _30681_, _06844_);
  and (_30684_, _30683_, _30680_);
  and (_30685_, _30654_, _06393_);
  or (_30686_, _30685_, _06387_);
  or (_30687_, _30686_, _30684_);
  or (_30688_, _30662_, _07245_);
  and (_30689_, _30688_, _06446_);
  and (_30690_, _30689_, _30687_);
  and (_30691_, _14371_, _08598_);
  or (_30692_, _30691_, _30672_);
  and (_30694_, _30692_, _06300_);
  or (_30695_, _30694_, _10059_);
  or (_30696_, _30695_, _30690_);
  and (_30697_, _30696_, _30659_);
  or (_30698_, _30697_, _06281_);
  and (_30699_, _07945_, _09446_);
  or (_30700_, _30654_, _06282_);
  or (_30701_, _30700_, _30699_);
  and (_30702_, _30701_, _30698_);
  or (_30703_, _30702_, _06015_);
  and (_30705_, _14426_, _07945_);
  or (_30706_, _30654_, _06279_);
  or (_30707_, _30706_, _30705_);
  and (_30708_, _30707_, _06276_);
  and (_30709_, _30708_, _30703_);
  and (_30710_, _07945_, _08817_);
  or (_30711_, _30710_, _30654_);
  and (_30712_, _30711_, _06275_);
  or (_30713_, _30712_, _06474_);
  or (_30714_, _30713_, _30709_);
  and (_30716_, _14324_, _07945_);
  or (_30717_, _30716_, _30654_);
  or (_30718_, _30717_, _07282_);
  and (_30719_, _30718_, _07284_);
  and (_30720_, _30719_, _30714_);
  nor (_30721_, _12538_, _13143_);
  or (_30722_, _30721_, _30654_);
  nor (_30723_, _30653_, _07284_);
  and (_30724_, _30723_, _30722_);
  or (_30725_, _30724_, _30720_);
  and (_30727_, _30725_, _07279_);
  nand (_30728_, _30711_, _06478_);
  nor (_30729_, _30728_, _30661_);
  or (_30730_, _30729_, _06569_);
  or (_30731_, _30730_, _30727_);
  and (_30732_, _30731_, _30656_);
  or (_30733_, _30732_, _06479_);
  and (_30734_, _14320_, _07945_);
  or (_30735_, _30734_, _30654_);
  or (_30736_, _30735_, _09043_);
  and (_30738_, _30736_, _09048_);
  and (_30739_, _30738_, _30733_);
  and (_30740_, _30722_, _06572_);
  or (_30741_, _30740_, _06606_);
  or (_30742_, _30741_, _30739_);
  or (_30743_, _30662_, _07037_);
  and (_30744_, _30743_, _30742_);
  or (_30745_, _30744_, _06234_);
  or (_30746_, _30654_, _06807_);
  and (_30747_, _30746_, _30745_);
  or (_30749_, _30747_, _06195_);
  or (_30750_, _30662_, _06196_);
  and (_30751_, _30750_, _01375_);
  and (_30752_, _30751_, _30749_);
  nor (_30753_, \uc8051golden_1.P3 [0], rst);
  nor (_30754_, _30753_, _01382_);
  or (_43001_, _30754_, _30752_);
  and (_30755_, _13143_, \uc8051golden_1.P3 [1]);
  nor (_30756_, _11223_, _13143_);
  or (_30757_, _30756_, _30755_);
  or (_30759_, _30757_, _09048_);
  nand (_30760_, _07945_, _07090_);
  or (_30761_, _07945_, \uc8051golden_1.P3 [1]);
  and (_30762_, _30761_, _06275_);
  and (_30763_, _30762_, _30760_);
  nor (_30764_, _13143_, _07196_);
  or (_30765_, _30764_, _30755_);
  or (_30766_, _30765_, _07221_);
  and (_30767_, _14532_, _07945_);
  not (_30768_, _30767_);
  and (_30770_, _30768_, _30761_);
  or (_30771_, _30770_, _07210_);
  and (_30772_, _07945_, \uc8051golden_1.ACC [1]);
  or (_30773_, _30772_, _30755_);
  and (_30774_, _30773_, _07199_);
  and (_30775_, _07200_, \uc8051golden_1.P3 [1]);
  or (_30776_, _30775_, _06401_);
  or (_30777_, _30776_, _30774_);
  and (_30778_, _30777_, _06396_);
  and (_30779_, _30778_, _30771_);
  and (_30781_, _13151_, \uc8051golden_1.P3 [1]);
  and (_30782_, _14514_, _08598_);
  or (_30783_, _30782_, _30781_);
  and (_30784_, _30783_, _06395_);
  or (_30785_, _30784_, _06399_);
  or (_30786_, _30785_, _30779_);
  and (_30787_, _30786_, _30766_);
  or (_30788_, _30787_, _06406_);
  or (_30789_, _30773_, _06414_);
  and (_30790_, _30789_, _06844_);
  and (_30792_, _30790_, _30788_);
  and (_30793_, _14517_, _08598_);
  or (_30794_, _30793_, _30781_);
  and (_30795_, _30794_, _06393_);
  or (_30796_, _30795_, _06387_);
  or (_30797_, _30796_, _30792_);
  and (_30798_, _30782_, _14513_);
  or (_30799_, _30781_, _07245_);
  or (_30800_, _30799_, _30798_);
  and (_30801_, _30800_, _06446_);
  and (_30803_, _30801_, _30797_);
  or (_30804_, _30781_, _14560_);
  and (_30805_, _30804_, _06300_);
  and (_30806_, _30805_, _30783_);
  or (_30807_, _30806_, _10059_);
  or (_30808_, _30807_, _30803_);
  or (_30809_, _30765_, _06293_);
  and (_30810_, _30809_, _30808_);
  or (_30811_, _30810_, _06281_);
  and (_30812_, _07945_, _09445_);
  or (_30814_, _30755_, _06282_);
  or (_30815_, _30814_, _30812_);
  and (_30816_, _30815_, _06279_);
  and (_30817_, _30816_, _30811_);
  and (_30818_, _14615_, _07945_);
  or (_30819_, _30818_, _30755_);
  and (_30820_, _30819_, _06015_);
  or (_30821_, _30820_, _30817_);
  and (_30822_, _30821_, _06276_);
  or (_30823_, _30822_, _30763_);
  and (_30825_, _30823_, _07282_);
  or (_30826_, _14507_, _13143_);
  and (_30827_, _30761_, _06474_);
  and (_30828_, _30827_, _30826_);
  or (_30829_, _30828_, _06582_);
  or (_30830_, _30829_, _30825_);
  and (_30831_, _11224_, _07945_);
  or (_30832_, _30831_, _30755_);
  or (_30833_, _30832_, _07284_);
  and (_30834_, _30833_, _07279_);
  and (_30836_, _30834_, _30830_);
  or (_30837_, _14505_, _13143_);
  and (_30838_, _30761_, _06478_);
  and (_30839_, _30838_, _30837_);
  or (_30840_, _30839_, _06569_);
  or (_30841_, _30840_, _30836_);
  and (_30842_, _30772_, _08477_);
  or (_30843_, _30755_, _07276_);
  or (_30844_, _30843_, _30842_);
  and (_30845_, _30844_, _09043_);
  and (_30847_, _30845_, _30841_);
  or (_30848_, _30760_, _08477_);
  and (_30849_, _30761_, _06479_);
  and (_30850_, _30849_, _30848_);
  or (_30851_, _30850_, _06572_);
  or (_30852_, _30851_, _30847_);
  and (_30853_, _30852_, _30759_);
  or (_30854_, _30853_, _06606_);
  or (_30855_, _30770_, _07037_);
  and (_30856_, _30855_, _06807_);
  and (_30858_, _30856_, _30854_);
  and (_30859_, _30794_, _06234_);
  or (_30860_, _30859_, _06195_);
  or (_30861_, _30860_, _30858_);
  or (_30862_, _30755_, _06196_);
  or (_30863_, _30862_, _30767_);
  and (_30864_, _30863_, _01375_);
  and (_30865_, _30864_, _30861_);
  nor (_30866_, \uc8051golden_1.P3 [1], rst);
  nor (_30867_, _30866_, _01382_);
  or (_43002_, _30867_, _30865_);
  and (_30869_, _13143_, \uc8051golden_1.P3 [2]);
  nor (_30870_, _13143_, _07623_);
  or (_30871_, _30870_, _30869_);
  or (_30872_, _30871_, _06293_);
  or (_30873_, _30871_, _07221_);
  and (_30874_, _14754_, _07945_);
  or (_30875_, _30874_, _30869_);
  or (_30876_, _30875_, _07210_);
  and (_30877_, _07945_, \uc8051golden_1.ACC [2]);
  or (_30879_, _30877_, _30869_);
  and (_30880_, _30879_, _07199_);
  and (_30881_, _07200_, \uc8051golden_1.P3 [2]);
  or (_30882_, _30881_, _06401_);
  or (_30883_, _30882_, _30880_);
  and (_30884_, _30883_, _06396_);
  and (_30885_, _30884_, _30876_);
  and (_30886_, _13151_, \uc8051golden_1.P3 [2]);
  and (_30887_, _14751_, _08598_);
  or (_30888_, _30887_, _30886_);
  and (_30890_, _30888_, _06395_);
  or (_30891_, _30890_, _06399_);
  or (_30892_, _30891_, _30885_);
  and (_30893_, _30892_, _30873_);
  or (_30894_, _30893_, _06406_);
  or (_30895_, _30879_, _06414_);
  and (_30896_, _30895_, _06844_);
  and (_30897_, _30896_, _30894_);
  and (_30898_, _14749_, _08598_);
  or (_30899_, _30898_, _30886_);
  and (_30901_, _30899_, _06393_);
  or (_30902_, _30901_, _06387_);
  or (_30903_, _30902_, _30897_);
  and (_30904_, _30887_, _14778_);
  or (_30905_, _30886_, _07245_);
  or (_30906_, _30905_, _30904_);
  and (_30907_, _30906_, _06446_);
  and (_30908_, _30907_, _30903_);
  and (_30909_, _14793_, _08598_);
  or (_30910_, _30909_, _30886_);
  and (_30912_, _30910_, _06300_);
  or (_30913_, _30912_, _10059_);
  or (_30914_, _30913_, _30908_);
  and (_30915_, _30914_, _30872_);
  or (_30916_, _30915_, _06281_);
  and (_30917_, _07945_, _09444_);
  or (_30918_, _30869_, _06282_);
  or (_30919_, _30918_, _30917_);
  and (_30920_, _30919_, _06279_);
  and (_30921_, _30920_, _30916_);
  and (_30923_, _14848_, _07945_);
  or (_30924_, _30923_, _30869_);
  and (_30925_, _30924_, _06015_);
  or (_30926_, _30925_, _06275_);
  or (_30927_, _30926_, _30921_);
  and (_30928_, _07945_, _08994_);
  or (_30929_, _30928_, _30869_);
  or (_30930_, _30929_, _06276_);
  and (_30931_, _30930_, _30927_);
  or (_30932_, _30931_, _06474_);
  and (_30934_, _14744_, _07945_);
  or (_30935_, _30934_, _30869_);
  or (_30936_, _30935_, _07282_);
  and (_30937_, _30936_, _07284_);
  and (_30938_, _30937_, _30932_);
  and (_30939_, _11221_, _07945_);
  or (_30940_, _30939_, _30869_);
  and (_30941_, _30940_, _06582_);
  or (_30942_, _30941_, _30938_);
  and (_30943_, _30942_, _07279_);
  or (_30945_, _30869_, _08433_);
  and (_30946_, _30929_, _06478_);
  and (_30947_, _30946_, _30945_);
  or (_30948_, _30947_, _30943_);
  and (_30949_, _30948_, _07276_);
  and (_30950_, _30879_, _06569_);
  and (_30951_, _30950_, _30945_);
  or (_30952_, _30951_, _06479_);
  or (_30953_, _30952_, _30949_);
  and (_30954_, _14741_, _07945_);
  or (_30956_, _30869_, _09043_);
  or (_30957_, _30956_, _30954_);
  and (_30958_, _30957_, _09048_);
  and (_30959_, _30958_, _30953_);
  nor (_30960_, _11220_, _13143_);
  or (_30961_, _30960_, _30869_);
  and (_30962_, _30961_, _06572_);
  or (_30963_, _30962_, _06606_);
  or (_30964_, _30963_, _30959_);
  or (_30965_, _30875_, _07037_);
  and (_30967_, _30965_, _06807_);
  and (_30968_, _30967_, _30964_);
  and (_30969_, _30899_, _06234_);
  or (_30970_, _30969_, _06195_);
  or (_30971_, _30970_, _30968_);
  and (_30972_, _14917_, _07945_);
  or (_30973_, _30869_, _06196_);
  or (_30974_, _30973_, _30972_);
  and (_30975_, _30974_, _01375_);
  and (_30976_, _30975_, _30971_);
  nor (_30978_, \uc8051golden_1.P3 [2], rst);
  nor (_30979_, _30978_, _01382_);
  or (_43003_, _30979_, _30976_);
  nor (_30980_, \uc8051golden_1.P3 [3], rst);
  nor (_30981_, _30980_, _01382_);
  and (_30982_, _13143_, \uc8051golden_1.P3 [3]);
  nor (_30983_, _13143_, _07775_);
  or (_30984_, _30983_, _30982_);
  or (_30985_, _30984_, _06293_);
  and (_30986_, _14947_, _07945_);
  or (_30988_, _30986_, _30982_);
  or (_30989_, _30988_, _07210_);
  and (_30990_, _07945_, \uc8051golden_1.ACC [3]);
  or (_30991_, _30990_, _30982_);
  and (_30992_, _30991_, _07199_);
  and (_30993_, _07200_, \uc8051golden_1.P3 [3]);
  or (_30994_, _30993_, _06401_);
  or (_30995_, _30994_, _30992_);
  and (_30996_, _30995_, _06396_);
  and (_30997_, _30996_, _30989_);
  and (_30999_, _13151_, \uc8051golden_1.P3 [3]);
  and (_31000_, _14951_, _08598_);
  or (_31001_, _31000_, _30999_);
  and (_31002_, _31001_, _06395_);
  or (_31003_, _31002_, _06399_);
  or (_31004_, _31003_, _30997_);
  or (_31005_, _30984_, _07221_);
  and (_31006_, _31005_, _31004_);
  or (_31007_, _31006_, _06406_);
  or (_31008_, _30991_, _06414_);
  and (_31010_, _31008_, _06844_);
  and (_31011_, _31010_, _31007_);
  and (_31012_, _14961_, _08598_);
  or (_31013_, _31012_, _30999_);
  and (_31014_, _31013_, _06393_);
  or (_31015_, _31014_, _06387_);
  or (_31016_, _31015_, _31011_);
  or (_31017_, _30999_, _14968_);
  and (_31018_, _31017_, _31001_);
  or (_31019_, _31018_, _07245_);
  and (_31021_, _31019_, _06446_);
  and (_31022_, _31021_, _31016_);
  and (_31023_, _14985_, _08598_);
  or (_31024_, _31023_, _30999_);
  and (_31025_, _31024_, _06300_);
  or (_31026_, _31025_, _10059_);
  or (_31027_, _31026_, _31022_);
  and (_31028_, _31027_, _30985_);
  or (_31029_, _31028_, _06281_);
  and (_31030_, _07945_, _09443_);
  or (_31032_, _30982_, _06282_);
  or (_31033_, _31032_, _31030_);
  and (_31034_, _31033_, _06279_);
  and (_31035_, _31034_, _31029_);
  and (_31036_, _15039_, _07945_);
  or (_31037_, _31036_, _30982_);
  and (_31038_, _31037_, _06015_);
  or (_31039_, _31038_, _06275_);
  or (_31040_, _31039_, _31035_);
  and (_31041_, _07945_, _08815_);
  or (_31044_, _31041_, _30982_);
  or (_31045_, _31044_, _06276_);
  and (_31046_, _31045_, _31040_);
  or (_31047_, _31046_, _06474_);
  and (_31048_, _14934_, _07945_);
  or (_31049_, _31048_, _30982_);
  or (_31050_, _31049_, _07282_);
  and (_31051_, _31050_, _07284_);
  and (_31052_, _31051_, _31047_);
  and (_31053_, _12535_, _07945_);
  or (_31055_, _31053_, _30982_);
  and (_31056_, _31055_, _06582_);
  or (_31057_, _31056_, _31052_);
  and (_31058_, _31057_, _07279_);
  or (_31059_, _30982_, _08389_);
  and (_31060_, _31044_, _06478_);
  and (_31061_, _31060_, _31059_);
  or (_31062_, _31061_, _31058_);
  and (_31063_, _31062_, _07276_);
  and (_31064_, _30991_, _06569_);
  and (_31067_, _31064_, _31059_);
  or (_31068_, _31067_, _06479_);
  or (_31069_, _31068_, _31063_);
  and (_31070_, _14931_, _07945_);
  or (_31071_, _30982_, _09043_);
  or (_31072_, _31071_, _31070_);
  and (_31073_, _31072_, _09048_);
  and (_31074_, _31073_, _31069_);
  nor (_31075_, _11218_, _13143_);
  or (_31076_, _31075_, _30982_);
  and (_31078_, _31076_, _06572_);
  or (_31079_, _31078_, _06606_);
  or (_31080_, _31079_, _31074_);
  or (_31081_, _30988_, _07037_);
  and (_31082_, _31081_, _06807_);
  and (_31083_, _31082_, _31080_);
  and (_31084_, _31013_, _06234_);
  or (_31085_, _31084_, _06195_);
  or (_31086_, _31085_, _31083_);
  and (_31087_, _15113_, _07945_);
  or (_31090_, _30982_, _06196_);
  or (_31091_, _31090_, _31087_);
  and (_31092_, _31091_, _01375_);
  and (_31093_, _31092_, _31086_);
  or (_43004_, _31093_, _30981_);
  and (_31094_, _13143_, \uc8051golden_1.P3 [4]);
  nor (_31095_, _13143_, _08301_);
  or (_31096_, _31095_, _31094_);
  or (_31097_, _31096_, _06293_);
  and (_31098_, _15130_, _07945_);
  or (_31100_, _31098_, _31094_);
  or (_31101_, _31100_, _07210_);
  and (_31102_, _07945_, \uc8051golden_1.ACC [4]);
  or (_31103_, _31102_, _31094_);
  and (_31104_, _31103_, _07199_);
  and (_31105_, _07200_, \uc8051golden_1.P3 [4]);
  or (_31106_, _31105_, _06401_);
  or (_31107_, _31106_, _31104_);
  and (_31108_, _31107_, _06396_);
  and (_31109_, _31108_, _31101_);
  and (_31112_, _13151_, \uc8051golden_1.P3 [4]);
  and (_31113_, _15139_, _08598_);
  or (_31114_, _31113_, _31112_);
  and (_31115_, _31114_, _06395_);
  or (_31116_, _31115_, _06399_);
  or (_31117_, _31116_, _31109_);
  or (_31118_, _31096_, _07221_);
  and (_31119_, _31118_, _31117_);
  or (_31120_, _31119_, _06406_);
  or (_31121_, _31103_, _06414_);
  and (_31123_, _31121_, _06844_);
  and (_31124_, _31123_, _31120_);
  and (_31125_, _15168_, _08598_);
  or (_31126_, _31125_, _31112_);
  and (_31127_, _31126_, _06393_);
  or (_31128_, _31127_, _06387_);
  or (_31129_, _31128_, _31124_);
  or (_31130_, _31112_, _15138_);
  and (_31131_, _31130_, _31114_);
  or (_31132_, _31131_, _07245_);
  and (_31134_, _31132_, _06446_);
  and (_31135_, _31134_, _31129_);
  and (_31136_, _15189_, _08598_);
  or (_31137_, _31136_, _31112_);
  and (_31138_, _31137_, _06300_);
  or (_31139_, _31138_, _10059_);
  or (_31140_, _31139_, _31135_);
  and (_31141_, _31140_, _31097_);
  or (_31142_, _31141_, _06281_);
  and (_31143_, _07945_, _09442_);
  or (_31145_, _31094_, _06282_);
  or (_31146_, _31145_, _31143_);
  and (_31147_, _31146_, _06279_);
  and (_31148_, _31147_, _31142_);
  and (_31149_, _15243_, _07945_);
  or (_31150_, _31149_, _31094_);
  and (_31151_, _31150_, _06015_);
  or (_31152_, _31151_, _06275_);
  or (_31153_, _31152_, _31148_);
  and (_31154_, _08883_, _07945_);
  or (_31155_, _31154_, _31094_);
  or (_31156_, _31155_, _06276_);
  and (_31157_, _31156_, _31153_);
  or (_31158_, _31157_, _06474_);
  and (_31159_, _15135_, _07945_);
  or (_31160_, _31159_, _31094_);
  or (_31161_, _31160_, _07282_);
  and (_31162_, _31161_, _07284_);
  and (_31163_, _31162_, _31158_);
  and (_31164_, _11216_, _07945_);
  or (_31167_, _31164_, _31094_);
  and (_31168_, _31167_, _06582_);
  or (_31169_, _31168_, _31163_);
  and (_31170_, _31169_, _07279_);
  or (_31171_, _31094_, _08345_);
  and (_31172_, _31155_, _06478_);
  and (_31173_, _31172_, _31171_);
  or (_31174_, _31173_, _31170_);
  and (_31175_, _31174_, _07276_);
  and (_31176_, _31103_, _06569_);
  and (_31177_, _31176_, _31171_);
  or (_31178_, _31177_, _06479_);
  or (_31179_, _31178_, _31175_);
  and (_31180_, _15134_, _07945_);
  or (_31181_, _31094_, _09043_);
  or (_31182_, _31181_, _31180_);
  and (_31183_, _31182_, _09048_);
  and (_31184_, _31183_, _31179_);
  nor (_31185_, _11215_, _13143_);
  or (_31186_, _31185_, _31094_);
  and (_31189_, _31186_, _06572_);
  or (_31190_, _31189_, _06606_);
  or (_31191_, _31190_, _31184_);
  or (_31192_, _31100_, _07037_);
  and (_31193_, _31192_, _06807_);
  and (_31194_, _31193_, _31191_);
  and (_31195_, _31126_, _06234_);
  or (_31196_, _31195_, _06195_);
  or (_31197_, _31196_, _31194_);
  and (_31198_, _15315_, _07945_);
  or (_31199_, _31094_, _06196_);
  or (_31200_, _31199_, _31198_);
  and (_31201_, _31200_, _01375_);
  and (_31202_, _31201_, _31197_);
  nor (_31203_, \uc8051golden_1.P3 [4], rst);
  nor (_31204_, _31203_, _01382_);
  or (_43005_, _31204_, _31202_);
  and (_31205_, _13143_, \uc8051golden_1.P3 [5]);
  nor (_31206_, _13143_, _08207_);
  or (_31207_, _31206_, _31205_);
  or (_31210_, _31207_, _06293_);
  and (_31211_, _15348_, _07945_);
  or (_31212_, _31211_, _31205_);
  or (_31213_, _31212_, _07210_);
  and (_31214_, _07945_, \uc8051golden_1.ACC [5]);
  or (_31215_, _31214_, _31205_);
  and (_31216_, _31215_, _07199_);
  and (_31217_, _07200_, \uc8051golden_1.P3 [5]);
  or (_31218_, _31217_, _06401_);
  or (_31219_, _31218_, _31216_);
  and (_31220_, _31219_, _06396_);
  and (_31221_, _31220_, _31213_);
  and (_31222_, _13151_, \uc8051golden_1.P3 [5]);
  and (_31223_, _15341_, _08598_);
  or (_31224_, _31223_, _31222_);
  and (_31225_, _31224_, _06395_);
  or (_31226_, _31225_, _06399_);
  or (_31227_, _31226_, _31221_);
  or (_31228_, _31207_, _07221_);
  and (_31229_, _31228_, _31227_);
  or (_31232_, _31229_, _06406_);
  or (_31233_, _31215_, _06414_);
  and (_31234_, _31233_, _06844_);
  and (_31235_, _31234_, _31232_);
  and (_31236_, _15345_, _08598_);
  or (_31237_, _31236_, _31222_);
  and (_31238_, _31237_, _06393_);
  or (_31239_, _31238_, _06387_);
  or (_31240_, _31239_, _31235_);
  or (_31241_, _31222_, _15378_);
  and (_31242_, _31241_, _31224_);
  or (_31243_, _31242_, _07245_);
  and (_31244_, _31243_, _06446_);
  and (_31245_, _31244_, _31240_);
  or (_31246_, _31222_, _15342_);
  and (_31247_, _31246_, _06300_);
  and (_31248_, _31247_, _31224_);
  or (_31249_, _31248_, _10059_);
  or (_31250_, _31249_, _31245_);
  and (_31251_, _31250_, _31210_);
  or (_31254_, _31251_, _06281_);
  and (_31255_, _07945_, _09441_);
  or (_31256_, _31205_, _06282_);
  or (_31257_, _31256_, _31255_);
  and (_31258_, _31257_, _06279_);
  and (_31259_, _31258_, _31254_);
  and (_31260_, _15446_, _07945_);
  or (_31261_, _31260_, _31205_);
  and (_31262_, _31261_, _06015_);
  or (_31263_, _31262_, _06275_);
  or (_31264_, _31263_, _31259_);
  and (_31265_, _08958_, _07945_);
  or (_31266_, _31265_, _31205_);
  or (_31267_, _31266_, _06276_);
  and (_31268_, _31267_, _31264_);
  or (_31269_, _31268_, _06474_);
  and (_31270_, _15338_, _07945_);
  or (_31271_, _31270_, _31205_);
  or (_31272_, _31271_, _07282_);
  and (_31273_, _31272_, _07284_);
  and (_31276_, _31273_, _31269_);
  and (_31277_, _12542_, _07945_);
  or (_31278_, _31277_, _31205_);
  and (_31279_, _31278_, _06582_);
  or (_31280_, _31279_, _31276_);
  and (_31281_, _31280_, _07279_);
  or (_31282_, _31205_, _08256_);
  and (_31283_, _31266_, _06478_);
  and (_31284_, _31283_, _31282_);
  or (_31285_, _31284_, _31281_);
  and (_31286_, _31285_, _07276_);
  and (_31287_, _31215_, _06569_);
  and (_31288_, _31287_, _31282_);
  or (_31289_, _31288_, _06479_);
  or (_31290_, _31289_, _31286_);
  and (_31291_, _15335_, _07945_);
  or (_31292_, _31205_, _09043_);
  or (_31293_, _31292_, _31291_);
  and (_31294_, _31293_, _09048_);
  and (_31295_, _31294_, _31290_);
  nor (_31298_, _11212_, _13143_);
  or (_31299_, _31298_, _31205_);
  and (_31300_, _31299_, _06572_);
  or (_31301_, _31300_, _06606_);
  or (_31302_, _31301_, _31295_);
  or (_31303_, _31212_, _07037_);
  and (_31304_, _31303_, _06807_);
  and (_31305_, _31304_, _31302_);
  and (_31306_, _31237_, _06234_);
  or (_31307_, _31306_, _06195_);
  or (_31308_, _31307_, _31305_);
  and (_31309_, _15509_, _07945_);
  or (_31310_, _31205_, _06196_);
  or (_31311_, _31310_, _31309_);
  and (_31312_, _31311_, _01375_);
  and (_31313_, _31312_, _31308_);
  nor (_31314_, \uc8051golden_1.P3 [5], rst);
  nor (_31315_, _31314_, _01382_);
  or (_43006_, _31315_, _31313_);
  and (_31316_, _13143_, \uc8051golden_1.P3 [6]);
  nor (_31319_, _13143_, _08118_);
  or (_31320_, _31319_, _31316_);
  or (_31321_, _31320_, _06293_);
  and (_31322_, _15550_, _07945_);
  or (_31323_, _31322_, _31316_);
  or (_31324_, _31323_, _07210_);
  and (_31325_, _07945_, \uc8051golden_1.ACC [6]);
  or (_31326_, _31325_, _31316_);
  and (_31327_, _31326_, _07199_);
  and (_31328_, _07200_, \uc8051golden_1.P3 [6]);
  or (_31329_, _31328_, _06401_);
  or (_31330_, _31329_, _31327_);
  and (_31331_, _31330_, _06396_);
  and (_31332_, _31331_, _31324_);
  and (_31333_, _13151_, \uc8051golden_1.P3 [6]);
  and (_31334_, _15535_, _08598_);
  or (_31335_, _31334_, _31333_);
  and (_31336_, _31335_, _06395_);
  or (_31337_, _31336_, _06399_);
  or (_31338_, _31337_, _31332_);
  or (_31341_, _31320_, _07221_);
  and (_31342_, _31341_, _31338_);
  or (_31343_, _31342_, _06406_);
  or (_31344_, _31326_, _06414_);
  and (_31345_, _31344_, _06844_);
  and (_31346_, _31345_, _31343_);
  and (_31347_, _15561_, _08598_);
  or (_31348_, _31347_, _31333_);
  and (_31349_, _31348_, _06393_);
  or (_31350_, _31349_, _06387_);
  or (_31351_, _31350_, _31346_);
  or (_31352_, _31333_, _15568_);
  and (_31353_, _31352_, _31335_);
  or (_31354_, _31353_, _07245_);
  and (_31355_, _31354_, _06446_);
  and (_31356_, _31355_, _31351_);
  and (_31357_, _15585_, _08598_);
  or (_31358_, _31357_, _31333_);
  and (_31359_, _31358_, _06300_);
  or (_31360_, _31359_, _10059_);
  or (_31363_, _31360_, _31356_);
  and (_31364_, _31363_, _31321_);
  or (_31365_, _31364_, _06281_);
  and (_31366_, _07945_, _09440_);
  or (_31367_, _31316_, _06282_);
  or (_31368_, _31367_, _31366_);
  and (_31369_, _31368_, _06279_);
  and (_31370_, _31369_, _31365_);
  and (_31371_, _15639_, _07945_);
  or (_31372_, _31371_, _31316_);
  and (_31373_, _31372_, _06015_);
  or (_31374_, _31373_, _06275_);
  or (_31375_, _31374_, _31370_);
  and (_31376_, _15646_, _07945_);
  or (_31377_, _31376_, _31316_);
  or (_31378_, _31377_, _06276_);
  and (_31379_, _31378_, _31375_);
  or (_31380_, _31379_, _06474_);
  and (_31381_, _15531_, _07945_);
  or (_31382_, _31381_, _31316_);
  or (_31385_, _31382_, _07282_);
  and (_31386_, _31385_, _07284_);
  and (_31387_, _31386_, _31380_);
  and (_31388_, _11210_, _07945_);
  or (_31389_, _31388_, _31316_);
  and (_31390_, _31389_, _06582_);
  or (_31391_, _31390_, _31387_);
  and (_31392_, _31391_, _07279_);
  or (_31393_, _31316_, _08162_);
  and (_31394_, _31377_, _06478_);
  and (_31395_, _31394_, _31393_);
  or (_31396_, _31395_, _31392_);
  and (_31397_, _31396_, _07276_);
  and (_31398_, _31326_, _06569_);
  and (_31399_, _31398_, _31393_);
  or (_31400_, _31399_, _06479_);
  or (_31401_, _31400_, _31397_);
  and (_31402_, _15528_, _07945_);
  or (_31403_, _31316_, _09043_);
  or (_31404_, _31403_, _31402_);
  and (_31407_, _31404_, _09048_);
  and (_31408_, _31407_, _31401_);
  nor (_31409_, _11209_, _13143_);
  or (_31410_, _31409_, _31316_);
  and (_31411_, _31410_, _06572_);
  or (_31412_, _31411_, _06606_);
  or (_31413_, _31412_, _31408_);
  or (_31414_, _31323_, _07037_);
  and (_31415_, _31414_, _06807_);
  and (_31416_, _31415_, _31413_);
  and (_31417_, _31348_, _06234_);
  or (_31418_, _31417_, _06195_);
  or (_31419_, _31418_, _31416_);
  and (_31420_, _15713_, _07945_);
  or (_31421_, _31316_, _06196_);
  or (_31422_, _31421_, _31420_);
  and (_31423_, _31422_, _01375_);
  and (_31424_, _31423_, _31419_);
  nor (_31425_, \uc8051golden_1.P3 [6], rst);
  nor (_31426_, _31425_, _01382_);
  or (_43007_, _31426_, _31424_);
  nand (_31429_, _11225_, _08019_);
  not (_31430_, \uc8051golden_1.P0 [0]);
  nor (_31431_, _08019_, _31430_);
  nor (_31432_, _31431_, _07276_);
  nand (_31433_, _31432_, _31429_);
  and (_31434_, _08019_, _07473_);
  or (_31435_, _31434_, _31431_);
  or (_31436_, _31435_, _06293_);
  nor (_31437_, _08521_, _13246_);
  or (_31438_, _31437_, _31431_);
  or (_31439_, _31438_, _07210_);
  and (_31440_, _08019_, \uc8051golden_1.ACC [0]);
  or (_31441_, _31440_, _31431_);
  and (_31442_, _31441_, _07199_);
  nor (_31443_, _07199_, _31430_);
  or (_31444_, _31443_, _06401_);
  or (_31445_, _31444_, _31442_);
  and (_31446_, _31445_, _06396_);
  and (_31447_, _31446_, _31439_);
  nor (_31450_, _07959_, _31430_);
  and (_31451_, _14339_, _07959_);
  or (_31452_, _31451_, _31450_);
  and (_31453_, _31452_, _06395_);
  or (_31454_, _31453_, _31447_);
  and (_31455_, _31454_, _07221_);
  and (_31456_, _31435_, _06399_);
  or (_31457_, _31456_, _06406_);
  or (_31458_, _31457_, _31455_);
  or (_31459_, _31441_, _06414_);
  and (_31460_, _31459_, _06844_);
  and (_31461_, _31460_, _31458_);
  and (_31462_, _31431_, _06393_);
  or (_31463_, _31462_, _06387_);
  or (_31464_, _31463_, _31461_);
  or (_31465_, _31438_, _07245_);
  and (_31466_, _31465_, _06446_);
  and (_31467_, _31466_, _31464_);
  and (_31468_, _14371_, _07959_);
  or (_31469_, _31468_, _31450_);
  and (_31472_, _31469_, _06300_);
  or (_31473_, _31472_, _10059_);
  or (_31474_, _31473_, _31467_);
  and (_31475_, _31474_, _31436_);
  or (_31476_, _31475_, _06281_);
  and (_31477_, _08019_, _09446_);
  or (_31478_, _31431_, _06282_);
  or (_31479_, _31478_, _31477_);
  and (_31480_, _31479_, _31476_);
  or (_31481_, _31480_, _06015_);
  and (_31482_, _14426_, _08019_);
  or (_31483_, _31431_, _06279_);
  or (_31484_, _31483_, _31482_);
  and (_31485_, _31484_, _06276_);
  and (_31486_, _31485_, _31481_);
  and (_31487_, _08019_, _08817_);
  or (_31488_, _31487_, _31431_);
  and (_31489_, _31488_, _06275_);
  or (_31490_, _31489_, _06474_);
  or (_31491_, _31490_, _31486_);
  and (_31494_, _14324_, _08019_);
  or (_31495_, _31494_, _31431_);
  or (_31496_, _31495_, _07282_);
  and (_31497_, _31496_, _07284_);
  and (_31498_, _31497_, _31491_);
  nor (_31499_, _12538_, _13246_);
  or (_31500_, _31499_, _31431_);
  and (_31501_, _31429_, _06582_);
  and (_31502_, _31501_, _31500_);
  or (_31503_, _31502_, _31498_);
  and (_31504_, _31503_, _07279_);
  nand (_31505_, _31488_, _06478_);
  nor (_31506_, _31505_, _31437_);
  or (_31507_, _31506_, _06569_);
  or (_31508_, _31507_, _31504_);
  and (_31509_, _31508_, _31433_);
  or (_31510_, _31509_, _06479_);
  and (_31511_, _14320_, _08019_);
  or (_31512_, _31511_, _31431_);
  or (_31513_, _31512_, _09043_);
  and (_31516_, _31513_, _09048_);
  and (_31517_, _31516_, _31510_);
  and (_31518_, _31500_, _06572_);
  or (_31519_, _31518_, _06606_);
  or (_31520_, _31519_, _31517_);
  or (_31521_, _31438_, _07037_);
  and (_31522_, _31521_, _31520_);
  or (_31523_, _31522_, _06234_);
  or (_31524_, _31431_, _06807_);
  and (_31525_, _31524_, _31523_);
  or (_31526_, _31525_, _06195_);
  or (_31527_, _31438_, _06196_);
  and (_31528_, _31527_, _01375_);
  and (_31529_, _31528_, _31526_);
  nor (_31530_, \uc8051golden_1.P0 [0], rst);
  nor (_31531_, _31530_, _01382_);
  or (_43009_, _31531_, _31529_);
  not (_31532_, \uc8051golden_1.P0 [1]);
  nor (_31533_, _08019_, _31532_);
  nor (_31534_, _11223_, _13246_);
  or (_31537_, _31534_, _31533_);
  or (_31538_, _31537_, _09048_);
  nor (_31539_, _13246_, _07196_);
  or (_31540_, _31539_, _31533_);
  or (_31541_, _31540_, _07221_);
  or (_31542_, _08019_, \uc8051golden_1.P0 [1]);
  and (_31543_, _14532_, _08019_);
  not (_31544_, _31543_);
  and (_31545_, _31544_, _31542_);
  or (_31546_, _31545_, _07210_);
  and (_31547_, _08019_, \uc8051golden_1.ACC [1]);
  or (_31548_, _31547_, _31533_);
  and (_31549_, _31548_, _07199_);
  nor (_31550_, _07199_, _31532_);
  or (_31551_, _31550_, _06401_);
  or (_31552_, _31551_, _31549_);
  and (_31553_, _31552_, _06396_);
  and (_31554_, _31553_, _31546_);
  nor (_31555_, _07959_, _31532_);
  and (_31556_, _14514_, _07959_);
  or (_31559_, _31556_, _31555_);
  and (_31560_, _31559_, _06395_);
  or (_31561_, _31560_, _06399_);
  or (_31562_, _31561_, _31554_);
  and (_31563_, _31562_, _31541_);
  or (_31564_, _31563_, _06406_);
  or (_31565_, _31548_, _06414_);
  and (_31566_, _31565_, _06844_);
  and (_31567_, _31566_, _31564_);
  and (_31568_, _14517_, _07959_);
  or (_31569_, _31568_, _31555_);
  and (_31570_, _31569_, _06393_);
  or (_31571_, _31570_, _06387_);
  or (_31572_, _31571_, _31567_);
  and (_31573_, _31556_, _14513_);
  or (_31574_, _31555_, _07245_);
  or (_31575_, _31574_, _31573_);
  and (_31576_, _31575_, _06446_);
  and (_31577_, _31576_, _31572_);
  or (_31578_, _31555_, _14560_);
  and (_31581_, _31578_, _06300_);
  and (_31582_, _31581_, _31559_);
  or (_31583_, _31582_, _10059_);
  or (_31584_, _31583_, _31577_);
  or (_31585_, _31540_, _06293_);
  and (_31586_, _31585_, _31584_);
  or (_31587_, _31586_, _06281_);
  and (_31588_, _08019_, _09445_);
  or (_31589_, _31533_, _06282_);
  or (_31590_, _31589_, _31588_);
  and (_31591_, _31590_, _06279_);
  and (_31592_, _31591_, _31587_);
  and (_31593_, _14615_, _08019_);
  or (_31594_, _31593_, _31533_);
  and (_31595_, _31594_, _06015_);
  or (_31596_, _31595_, _31592_);
  and (_31597_, _31596_, _06276_);
  nand (_31598_, _08019_, _07090_);
  and (_31599_, _31542_, _06275_);
  and (_31600_, _31599_, _31598_);
  or (_31603_, _31600_, _31597_);
  and (_31604_, _31603_, _07282_);
  or (_31605_, _14507_, _13246_);
  and (_31606_, _31542_, _06474_);
  and (_31607_, _31606_, _31605_);
  or (_31608_, _31607_, _06582_);
  or (_31609_, _31608_, _31604_);
  nand (_31610_, _11222_, _08019_);
  and (_31611_, _31610_, _31537_);
  or (_31612_, _31611_, _07284_);
  and (_31613_, _31612_, _07279_);
  and (_31614_, _31613_, _31609_);
  or (_31615_, _14505_, _13246_);
  and (_31616_, _31542_, _06478_);
  and (_31617_, _31616_, _31615_);
  or (_31618_, _31617_, _06569_);
  or (_31619_, _31618_, _31614_);
  nor (_31620_, _31533_, _07276_);
  nand (_31621_, _31620_, _31610_);
  and (_31622_, _31621_, _09043_);
  and (_31625_, _31622_, _31619_);
  or (_31626_, _31598_, _08477_);
  and (_31627_, _31542_, _06479_);
  and (_31628_, _31627_, _31626_);
  or (_31629_, _31628_, _06572_);
  or (_31630_, _31629_, _31625_);
  and (_31631_, _31630_, _31538_);
  or (_31632_, _31631_, _06606_);
  or (_31633_, _31545_, _07037_);
  and (_31634_, _31633_, _06807_);
  and (_31635_, _31634_, _31632_);
  and (_31636_, _31569_, _06234_);
  or (_31637_, _31636_, _06195_);
  or (_31638_, _31637_, _31635_);
  or (_31639_, _31533_, _06196_);
  or (_31640_, _31639_, _31543_);
  and (_31641_, _31640_, _01375_);
  and (_31642_, _31641_, _31638_);
  nor (_31643_, \uc8051golden_1.P0 [1], rst);
  nor (_31644_, _31643_, _01382_);
  or (_43010_, _31644_, _31642_);
  and (_31647_, _13246_, \uc8051golden_1.P0 [2]);
  nor (_31648_, _13246_, _07623_);
  or (_31649_, _31648_, _31647_);
  or (_31650_, _31649_, _06293_);
  or (_31651_, _31649_, _07221_);
  and (_31652_, _14754_, _08019_);
  or (_31653_, _31652_, _31647_);
  or (_31654_, _31653_, _07210_);
  and (_31655_, _08019_, \uc8051golden_1.ACC [2]);
  or (_31656_, _31655_, _31647_);
  and (_31657_, _31656_, _07199_);
  and (_31658_, _07200_, \uc8051golden_1.P0 [2]);
  or (_31659_, _31658_, _06401_);
  or (_31660_, _31659_, _31657_);
  and (_31661_, _31660_, _06396_);
  and (_31662_, _31661_, _31654_);
  and (_31663_, _13254_, \uc8051golden_1.P0 [2]);
  and (_31664_, _14751_, _07959_);
  or (_31665_, _31664_, _31663_);
  and (_31668_, _31665_, _06395_);
  or (_31669_, _31668_, _06399_);
  or (_31670_, _31669_, _31662_);
  and (_31671_, _31670_, _31651_);
  or (_31672_, _31671_, _06406_);
  or (_31673_, _31656_, _06414_);
  and (_31674_, _31673_, _06844_);
  and (_31675_, _31674_, _31672_);
  and (_31676_, _14749_, _07959_);
  or (_31677_, _31676_, _31663_);
  and (_31678_, _31677_, _06393_);
  or (_31679_, _31678_, _06387_);
  or (_31680_, _31679_, _31675_);
  and (_31681_, _31664_, _14778_);
  or (_31682_, _31663_, _07245_);
  or (_31683_, _31682_, _31681_);
  and (_31684_, _31683_, _06446_);
  and (_31685_, _31684_, _31680_);
  and (_31686_, _14793_, _07959_);
  or (_31687_, _31686_, _31663_);
  and (_31690_, _31687_, _06300_);
  or (_31691_, _31690_, _10059_);
  or (_31692_, _31691_, _31685_);
  and (_31693_, _31692_, _31650_);
  or (_31694_, _31693_, _06281_);
  and (_31695_, _08019_, _09444_);
  or (_31696_, _31647_, _06282_);
  or (_31697_, _31696_, _31695_);
  and (_31698_, _31697_, _06279_);
  and (_31699_, _31698_, _31694_);
  and (_31700_, _14848_, _08019_);
  or (_31701_, _31700_, _31647_);
  and (_31702_, _31701_, _06015_);
  or (_31703_, _31702_, _06275_);
  or (_31704_, _31703_, _31699_);
  and (_31705_, _08019_, _08994_);
  or (_31706_, _31705_, _31647_);
  or (_31707_, _31706_, _06276_);
  and (_31708_, _31707_, _31704_);
  or (_31709_, _31708_, _06474_);
  and (_31712_, _14744_, _08019_);
  or (_31713_, _31712_, _31647_);
  or (_31714_, _31713_, _07282_);
  and (_31715_, _31714_, _07284_);
  and (_31716_, _31715_, _31709_);
  and (_31717_, _11221_, _08019_);
  or (_31718_, _31717_, _31647_);
  and (_31719_, _31718_, _06582_);
  or (_31720_, _31719_, _31716_);
  and (_31721_, _31720_, _07279_);
  or (_31722_, _31647_, _08433_);
  and (_31723_, _31706_, _06478_);
  and (_31724_, _31723_, _31722_);
  or (_31725_, _31724_, _31721_);
  and (_31726_, _31725_, _07276_);
  and (_31727_, _31656_, _06569_);
  and (_31728_, _31727_, _31722_);
  or (_31729_, _31728_, _06479_);
  or (_31730_, _31729_, _31726_);
  and (_31731_, _14741_, _08019_);
  or (_31734_, _31647_, _09043_);
  or (_31735_, _31734_, _31731_);
  and (_31736_, _31735_, _09048_);
  and (_31737_, _31736_, _31730_);
  nor (_31738_, _11220_, _13246_);
  or (_31739_, _31738_, _31647_);
  and (_31740_, _31739_, _06572_);
  or (_31741_, _31740_, _06606_);
  or (_31742_, _31741_, _31737_);
  or (_31743_, _31653_, _07037_);
  and (_31744_, _31743_, _06807_);
  and (_31745_, _31744_, _31742_);
  and (_31746_, _31677_, _06234_);
  or (_31747_, _31746_, _06195_);
  or (_31748_, _31747_, _31745_);
  and (_31749_, _14917_, _08019_);
  or (_31750_, _31647_, _06196_);
  or (_31751_, _31750_, _31749_);
  and (_31752_, _31751_, _01375_);
  and (_31753_, _31752_, _31748_);
  nor (_31756_, \uc8051golden_1.P0 [2], rst);
  nor (_31757_, _31756_, _01382_);
  or (_43011_, _31757_, _31753_);
  and (_31758_, _13246_, \uc8051golden_1.P0 [3]);
  nor (_31759_, _13246_, _07775_);
  or (_31760_, _31759_, _31758_);
  or (_31761_, _31760_, _06293_);
  and (_31762_, _14947_, _08019_);
  or (_31763_, _31762_, _31758_);
  or (_31764_, _31763_, _07210_);
  and (_31766_, _08019_, \uc8051golden_1.ACC [3]);
  or (_31767_, _31766_, _31758_);
  and (_31768_, _31767_, _07199_);
  and (_31769_, _07200_, \uc8051golden_1.P0 [3]);
  or (_31770_, _31769_, _06401_);
  or (_31771_, _31770_, _31768_);
  and (_31772_, _31771_, _06396_);
  and (_31773_, _31772_, _31764_);
  and (_31774_, _13254_, \uc8051golden_1.P0 [3]);
  and (_31775_, _14951_, _07959_);
  or (_31777_, _31775_, _31774_);
  and (_31778_, _31777_, _06395_);
  or (_31779_, _31778_, _06399_);
  or (_31780_, _31779_, _31773_);
  or (_31781_, _31760_, _07221_);
  and (_31782_, _31781_, _31780_);
  or (_31783_, _31782_, _06406_);
  or (_31784_, _31767_, _06414_);
  and (_31785_, _31784_, _06844_);
  and (_31786_, _31785_, _31783_);
  and (_31788_, _14961_, _07959_);
  or (_31789_, _31788_, _31774_);
  and (_31790_, _31789_, _06393_);
  or (_31791_, _31790_, _06387_);
  or (_31792_, _31791_, _31786_);
  or (_31793_, _31774_, _14968_);
  and (_31794_, _31793_, _31777_);
  or (_31795_, _31794_, _07245_);
  and (_31796_, _31795_, _06446_);
  and (_31797_, _31796_, _31792_);
  and (_31799_, _14985_, _07959_);
  or (_31800_, _31799_, _31774_);
  and (_31801_, _31800_, _06300_);
  or (_31802_, _31801_, _10059_);
  or (_31803_, _31802_, _31797_);
  and (_31804_, _31803_, _31761_);
  or (_31805_, _31804_, _06281_);
  and (_31806_, _08019_, _09443_);
  or (_31807_, _31758_, _06282_);
  or (_31808_, _31807_, _31806_);
  and (_31810_, _31808_, _06279_);
  and (_31811_, _31810_, _31805_);
  and (_31812_, _15039_, _08019_);
  or (_31813_, _31812_, _31758_);
  and (_31814_, _31813_, _06015_);
  or (_31815_, _31814_, _06275_);
  or (_31816_, _31815_, _31811_);
  and (_31817_, _08019_, _08815_);
  or (_31818_, _31817_, _31758_);
  or (_31819_, _31818_, _06276_);
  and (_31821_, _31819_, _31816_);
  or (_31822_, _31821_, _06474_);
  and (_31823_, _14934_, _08019_);
  or (_31824_, _31823_, _31758_);
  or (_31825_, _31824_, _07282_);
  and (_31826_, _31825_, _07284_);
  and (_31827_, _31826_, _31822_);
  and (_31828_, _12535_, _08019_);
  or (_31829_, _31828_, _31758_);
  and (_31830_, _31829_, _06582_);
  or (_31832_, _31830_, _31827_);
  and (_31833_, _31832_, _07279_);
  or (_31834_, _31758_, _08389_);
  and (_31835_, _31818_, _06478_);
  and (_31836_, _31835_, _31834_);
  or (_31837_, _31836_, _31833_);
  and (_31838_, _31837_, _07276_);
  and (_31839_, _31767_, _06569_);
  and (_31840_, _31839_, _31834_);
  or (_31841_, _31840_, _06479_);
  or (_31843_, _31841_, _31838_);
  and (_31844_, _14931_, _08019_);
  or (_31845_, _31758_, _09043_);
  or (_31846_, _31845_, _31844_);
  and (_31847_, _31846_, _09048_);
  and (_31848_, _31847_, _31843_);
  nor (_31849_, _11218_, _13246_);
  or (_31850_, _31849_, _31758_);
  and (_31851_, _31850_, _06572_);
  or (_31852_, _31851_, _06606_);
  or (_31853_, _31852_, _31848_);
  or (_31854_, _31763_, _07037_);
  and (_31855_, _31854_, _06807_);
  and (_31856_, _31855_, _31853_);
  and (_31857_, _31789_, _06234_);
  or (_31858_, _31857_, _06195_);
  or (_31859_, _31858_, _31856_);
  and (_31860_, _15113_, _08019_);
  or (_31861_, _31758_, _06196_);
  or (_31862_, _31861_, _31860_);
  and (_31864_, _31862_, _01375_);
  and (_31865_, _31864_, _31859_);
  nor (_31866_, \uc8051golden_1.P0 [3], rst);
  nor (_31867_, _31866_, _01382_);
  or (_43012_, _31867_, _31865_);
  nor (_31868_, \uc8051golden_1.P0 [4], rst);
  nor (_31869_, _31868_, _01382_);
  and (_31870_, _13246_, \uc8051golden_1.P0 [4]);
  nor (_31871_, _13246_, _08301_);
  or (_31872_, _31871_, _31870_);
  or (_31874_, _31872_, _06293_);
  and (_31875_, _15130_, _08019_);
  or (_31876_, _31875_, _31870_);
  or (_31877_, _31876_, _07210_);
  and (_31878_, _08019_, \uc8051golden_1.ACC [4]);
  or (_31879_, _31878_, _31870_);
  and (_31880_, _31879_, _07199_);
  and (_31881_, _07200_, \uc8051golden_1.P0 [4]);
  or (_31882_, _31881_, _06401_);
  or (_31883_, _31882_, _31880_);
  and (_31885_, _31883_, _06396_);
  and (_31886_, _31885_, _31877_);
  and (_31887_, _13254_, \uc8051golden_1.P0 [4]);
  and (_31888_, _15139_, _07959_);
  or (_31889_, _31888_, _31887_);
  and (_31890_, _31889_, _06395_);
  or (_31891_, _31890_, _06399_);
  or (_31892_, _31891_, _31886_);
  or (_31893_, _31872_, _07221_);
  and (_31894_, _31893_, _31892_);
  or (_31896_, _31894_, _06406_);
  or (_31897_, _31879_, _06414_);
  and (_31898_, _31897_, _06844_);
  and (_31899_, _31898_, _31896_);
  and (_31900_, _15168_, _07959_);
  or (_31901_, _31900_, _31887_);
  and (_31902_, _31901_, _06393_);
  or (_31903_, _31902_, _06387_);
  or (_31904_, _31903_, _31899_);
  or (_31905_, _31887_, _15138_);
  and (_31907_, _31905_, _31889_);
  or (_31908_, _31907_, _07245_);
  and (_31909_, _31908_, _06446_);
  and (_31910_, _31909_, _31904_);
  and (_31911_, _15189_, _07959_);
  or (_31912_, _31911_, _31887_);
  and (_31913_, _31912_, _06300_);
  or (_31914_, _31913_, _10059_);
  or (_31915_, _31914_, _31910_);
  and (_31916_, _31915_, _31874_);
  or (_31918_, _31916_, _06281_);
  and (_31919_, _08019_, _09442_);
  or (_31920_, _31870_, _06282_);
  or (_31921_, _31920_, _31919_);
  and (_31922_, _31921_, _06279_);
  and (_31923_, _31922_, _31918_);
  and (_31924_, _15243_, _08019_);
  or (_31925_, _31924_, _31870_);
  and (_31926_, _31925_, _06015_);
  or (_31927_, _31926_, _06275_);
  or (_31929_, _31927_, _31923_);
  and (_31930_, _08883_, _08019_);
  or (_31931_, _31930_, _31870_);
  or (_31932_, _31931_, _06276_);
  and (_31933_, _31932_, _31929_);
  or (_31934_, _31933_, _06474_);
  and (_31935_, _15135_, _08019_);
  or (_31936_, _31935_, _31870_);
  or (_31937_, _31936_, _07282_);
  and (_31938_, _31937_, _07284_);
  and (_31940_, _31938_, _31934_);
  and (_31941_, _11216_, _08019_);
  or (_31942_, _31941_, _31870_);
  and (_31943_, _31942_, _06582_);
  or (_31944_, _31943_, _31940_);
  and (_31945_, _31944_, _07279_);
  or (_31946_, _31870_, _08345_);
  and (_31947_, _31931_, _06478_);
  and (_31948_, _31947_, _31946_);
  or (_31949_, _31948_, _31945_);
  and (_31951_, _31949_, _07276_);
  and (_31952_, _31879_, _06569_);
  and (_31953_, _31952_, _31946_);
  or (_31954_, _31953_, _06479_);
  or (_31955_, _31954_, _31951_);
  and (_31956_, _15134_, _08019_);
  or (_31957_, _31870_, _09043_);
  or (_31958_, _31957_, _31956_);
  and (_31959_, _31958_, _09048_);
  and (_31960_, _31959_, _31955_);
  nor (_31962_, _11215_, _13246_);
  or (_31963_, _31962_, _31870_);
  and (_31964_, _31963_, _06572_);
  or (_31965_, _31964_, _06606_);
  or (_31966_, _31965_, _31960_);
  or (_31967_, _31876_, _07037_);
  and (_31968_, _31967_, _06807_);
  and (_31969_, _31968_, _31966_);
  and (_31970_, _31901_, _06234_);
  or (_31971_, _31970_, _06195_);
  or (_31973_, _31971_, _31969_);
  and (_31974_, _15315_, _08019_);
  or (_31975_, _31870_, _06196_);
  or (_31976_, _31975_, _31974_);
  and (_31977_, _31976_, _01375_);
  and (_31978_, _31977_, _31973_);
  or (_43013_, _31978_, _31869_);
  and (_31979_, _13246_, \uc8051golden_1.P0 [5]);
  nor (_31980_, _13246_, _08207_);
  or (_31981_, _31980_, _31979_);
  or (_31983_, _31981_, _06293_);
  and (_31984_, _15348_, _08019_);
  or (_31985_, _31984_, _31979_);
  or (_31986_, _31985_, _07210_);
  and (_31987_, _08019_, \uc8051golden_1.ACC [5]);
  or (_31988_, _31987_, _31979_);
  and (_31989_, _31988_, _07199_);
  and (_31990_, _07200_, \uc8051golden_1.P0 [5]);
  or (_31991_, _31990_, _06401_);
  or (_31992_, _31991_, _31989_);
  and (_31994_, _31992_, _06396_);
  and (_31995_, _31994_, _31986_);
  and (_31996_, _13254_, \uc8051golden_1.P0 [5]);
  and (_31997_, _15341_, _07959_);
  or (_31998_, _31997_, _31996_);
  and (_31999_, _31998_, _06395_);
  or (_32000_, _31999_, _06399_);
  or (_32001_, _32000_, _31995_);
  or (_32002_, _31981_, _07221_);
  and (_32003_, _32002_, _32001_);
  or (_32005_, _32003_, _06406_);
  or (_32006_, _31988_, _06414_);
  and (_32007_, _32006_, _06844_);
  and (_32008_, _32007_, _32005_);
  and (_32009_, _15345_, _07959_);
  or (_32010_, _32009_, _31996_);
  and (_32011_, _32010_, _06393_);
  or (_32012_, _32011_, _06387_);
  or (_32013_, _32012_, _32008_);
  or (_32014_, _31996_, _15378_);
  and (_32016_, _32014_, _31998_);
  or (_32017_, _32016_, _07245_);
  and (_32018_, _32017_, _06446_);
  and (_32019_, _32018_, _32013_);
  or (_32020_, _31996_, _15342_);
  and (_32021_, _32020_, _06300_);
  and (_32022_, _32021_, _31998_);
  or (_32023_, _32022_, _10059_);
  or (_32024_, _32023_, _32019_);
  and (_32025_, _32024_, _31983_);
  or (_32027_, _32025_, _06281_);
  and (_32028_, _08019_, _09441_);
  or (_32029_, _31979_, _06282_);
  or (_32030_, _32029_, _32028_);
  and (_32031_, _32030_, _06279_);
  and (_32032_, _32031_, _32027_);
  and (_32033_, _15446_, _08019_);
  or (_32034_, _32033_, _31979_);
  and (_32035_, _32034_, _06015_);
  or (_32036_, _32035_, _06275_);
  or (_32038_, _32036_, _32032_);
  and (_32039_, _08958_, _08019_);
  or (_32040_, _32039_, _31979_);
  or (_32041_, _32040_, _06276_);
  and (_32042_, _32041_, _32038_);
  or (_32043_, _32042_, _06474_);
  and (_32044_, _15338_, _08019_);
  or (_32045_, _32044_, _31979_);
  or (_32046_, _32045_, _07282_);
  and (_32047_, _32046_, _07284_);
  and (_32049_, _32047_, _32043_);
  and (_32050_, _12542_, _08019_);
  or (_32051_, _32050_, _31979_);
  and (_32052_, _32051_, _06582_);
  or (_32053_, _32052_, _32049_);
  and (_32054_, _32053_, _07279_);
  or (_32055_, _31979_, _08256_);
  and (_32056_, _32040_, _06478_);
  and (_32057_, _32056_, _32055_);
  or (_32058_, _32057_, _32054_);
  and (_32060_, _32058_, _07276_);
  and (_32061_, _31988_, _06569_);
  and (_32062_, _32061_, _32055_);
  or (_32063_, _32062_, _06479_);
  or (_32064_, _32063_, _32060_);
  and (_32065_, _15335_, _08019_);
  or (_32066_, _31979_, _09043_);
  or (_32067_, _32066_, _32065_);
  and (_32068_, _32067_, _09048_);
  and (_32069_, _32068_, _32064_);
  nor (_32071_, _11212_, _13246_);
  or (_32072_, _32071_, _31979_);
  and (_32073_, _32072_, _06572_);
  or (_32074_, _32073_, _06606_);
  or (_32075_, _32074_, _32069_);
  or (_32076_, _31985_, _07037_);
  and (_32077_, _32076_, _06807_);
  and (_32078_, _32077_, _32075_);
  and (_32079_, _32010_, _06234_);
  or (_32080_, _32079_, _06195_);
  or (_32082_, _32080_, _32078_);
  and (_32083_, _15509_, _08019_);
  or (_32084_, _31979_, _06196_);
  or (_32085_, _32084_, _32083_);
  and (_32086_, _32085_, _01375_);
  and (_32087_, _32086_, _32082_);
  nor (_32088_, \uc8051golden_1.P0 [5], rst);
  nor (_32089_, _32088_, _01382_);
  or (_43014_, _32089_, _32087_);
  and (_32092_, _13246_, \uc8051golden_1.P0 [6]);
  nor (_32095_, _13246_, _08118_);
  or (_32097_, _32095_, _32092_);
  or (_32099_, _32097_, _06293_);
  and (_32101_, _15550_, _08019_);
  or (_32103_, _32101_, _32092_);
  or (_32105_, _32103_, _07210_);
  and (_32107_, _08019_, \uc8051golden_1.ACC [6]);
  or (_32109_, _32107_, _32092_);
  and (_32110_, _32109_, _07199_);
  and (_32111_, _07200_, \uc8051golden_1.P0 [6]);
  or (_32113_, _32111_, _06401_);
  or (_32114_, _32113_, _32110_);
  and (_32115_, _32114_, _06396_);
  and (_32116_, _32115_, _32105_);
  and (_32117_, _13254_, \uc8051golden_1.P0 [6]);
  and (_32118_, _15535_, _07959_);
  or (_32119_, _32118_, _32117_);
  and (_32120_, _32119_, _06395_);
  or (_32121_, _32120_, _06399_);
  or (_32122_, _32121_, _32116_);
  or (_32124_, _32097_, _07221_);
  and (_32125_, _32124_, _32122_);
  or (_32126_, _32125_, _06406_);
  or (_32127_, _32109_, _06414_);
  and (_32128_, _32127_, _06844_);
  and (_32129_, _32128_, _32126_);
  and (_32130_, _15561_, _07959_);
  or (_32131_, _32130_, _32117_);
  and (_32132_, _32131_, _06393_);
  or (_32133_, _32132_, _06387_);
  or (_32135_, _32133_, _32129_);
  or (_32136_, _32117_, _15568_);
  and (_32137_, _32136_, _32119_);
  or (_32138_, _32137_, _07245_);
  and (_32139_, _32138_, _06446_);
  and (_32140_, _32139_, _32135_);
  and (_32141_, _15585_, _07959_);
  or (_32142_, _32141_, _32117_);
  and (_32143_, _32142_, _06300_);
  or (_32144_, _32143_, _10059_);
  or (_32146_, _32144_, _32140_);
  and (_32147_, _32146_, _32099_);
  or (_32148_, _32147_, _06281_);
  and (_32149_, _08019_, _09440_);
  or (_32150_, _32092_, _06282_);
  or (_32151_, _32150_, _32149_);
  and (_32152_, _32151_, _06279_);
  and (_32153_, _32152_, _32148_);
  and (_32154_, _15639_, _08019_);
  or (_32155_, _32154_, _32092_);
  and (_32157_, _32155_, _06015_);
  or (_32158_, _32157_, _06275_);
  or (_32159_, _32158_, _32153_);
  and (_32160_, _15646_, _08019_);
  or (_32161_, _32160_, _32092_);
  or (_32162_, _32161_, _06276_);
  and (_32163_, _32162_, _32159_);
  or (_32164_, _32163_, _06474_);
  and (_32165_, _15531_, _08019_);
  or (_32166_, _32165_, _32092_);
  or (_32168_, _32166_, _07282_);
  and (_32169_, _32168_, _07284_);
  and (_32170_, _32169_, _32164_);
  and (_32171_, _11210_, _08019_);
  or (_32172_, _32171_, _32092_);
  and (_32173_, _32172_, _06582_);
  or (_32174_, _32173_, _32170_);
  and (_32175_, _32174_, _07279_);
  or (_32176_, _32092_, _08162_);
  and (_32177_, _32161_, _06478_);
  and (_32179_, _32177_, _32176_);
  or (_32180_, _32179_, _32175_);
  and (_32181_, _32180_, _07276_);
  and (_32182_, _32109_, _06569_);
  and (_32183_, _32182_, _32176_);
  or (_32184_, _32183_, _06479_);
  or (_32185_, _32184_, _32181_);
  and (_32186_, _15528_, _08019_);
  or (_32187_, _32092_, _09043_);
  or (_32188_, _32187_, _32186_);
  and (_32190_, _32188_, _09048_);
  and (_32191_, _32190_, _32185_);
  nor (_32192_, _11209_, _13246_);
  or (_32193_, _32192_, _32092_);
  and (_32194_, _32193_, _06572_);
  or (_32195_, _32194_, _06606_);
  or (_32196_, _32195_, _32191_);
  or (_32197_, _32103_, _07037_);
  and (_32198_, _32197_, _06807_);
  and (_32199_, _32198_, _32196_);
  and (_32201_, _32131_, _06234_);
  or (_32202_, _32201_, _06195_);
  or (_32203_, _32202_, _32199_);
  and (_32204_, _15713_, _08019_);
  or (_32205_, _32092_, _06196_);
  or (_32206_, _32205_, _32204_);
  and (_32207_, _32206_, _01375_);
  and (_32208_, _32207_, _32203_);
  nor (_32209_, \uc8051golden_1.P0 [6], rst);
  nor (_32210_, _32209_, _01382_);
  or (_43015_, _32210_, _32208_);
  nor (_32212_, \uc8051golden_1.P1 [0], rst);
  nor (_32213_, _32212_, _01382_);
  nand (_32214_, _11225_, _07970_);
  and (_32215_, _13351_, \uc8051golden_1.P1 [0]);
  nor (_32216_, _32215_, _07276_);
  nand (_32217_, _32216_, _32214_);
  and (_32218_, _07970_, _07473_);
  or (_32219_, _32218_, _32215_);
  or (_32220_, _32219_, _06293_);
  nor (_32222_, _08521_, _13351_);
  or (_32223_, _32222_, _32215_);
  or (_32224_, _32223_, _07210_);
  and (_32225_, _07970_, \uc8051golden_1.ACC [0]);
  or (_32226_, _32225_, _32215_);
  and (_32227_, _32226_, _07199_);
  and (_32228_, _07200_, \uc8051golden_1.P1 [0]);
  or (_32229_, _32228_, _06401_);
  or (_32230_, _32229_, _32227_);
  and (_32231_, _32230_, _06396_);
  and (_32233_, _32231_, _32224_);
  and (_32234_, _13359_, \uc8051golden_1.P1 [0]);
  and (_32235_, _14339_, _08626_);
  or (_32236_, _32235_, _32234_);
  and (_32237_, _32236_, _06395_);
  or (_32238_, _32237_, _32233_);
  and (_32239_, _32238_, _07221_);
  and (_32240_, _32219_, _06399_);
  or (_32241_, _32240_, _06406_);
  or (_32242_, _32241_, _32239_);
  or (_32244_, _32226_, _06414_);
  and (_32245_, _32244_, _06844_);
  and (_32246_, _32245_, _32242_);
  and (_32247_, _32215_, _06393_);
  or (_32248_, _32247_, _06387_);
  or (_32249_, _32248_, _32246_);
  or (_32250_, _32223_, _07245_);
  and (_32251_, _32250_, _06446_);
  and (_32252_, _32251_, _32249_);
  and (_32253_, _14371_, _08626_);
  or (_32255_, _32253_, _32234_);
  and (_32256_, _32255_, _06300_);
  or (_32257_, _32256_, _10059_);
  or (_32258_, _32257_, _32252_);
  and (_32259_, _32258_, _32220_);
  or (_32260_, _32259_, _06281_);
  and (_32261_, _07970_, _09446_);
  or (_32262_, _32215_, _06282_);
  or (_32263_, _32262_, _32261_);
  and (_32264_, _32263_, _32260_);
  or (_32266_, _32264_, _06015_);
  and (_32267_, _14426_, _07970_);
  or (_32268_, _32215_, _06279_);
  or (_32269_, _32268_, _32267_);
  and (_32270_, _32269_, _06276_);
  and (_32271_, _32270_, _32266_);
  and (_32272_, _07970_, _08817_);
  or (_32273_, _32272_, _32215_);
  and (_32274_, _32273_, _06275_);
  or (_32275_, _32274_, _06474_);
  or (_32277_, _32275_, _32271_);
  and (_32278_, _14324_, _07970_);
  or (_32279_, _32278_, _32215_);
  or (_32280_, _32279_, _07282_);
  and (_32281_, _32280_, _07284_);
  and (_32282_, _32281_, _32277_);
  nor (_32283_, _12538_, _13351_);
  or (_32284_, _32283_, _32215_);
  and (_32285_, _32214_, _06582_);
  and (_32286_, _32285_, _32284_);
  or (_32288_, _32286_, _32282_);
  and (_32289_, _32288_, _07279_);
  nand (_32290_, _32273_, _06478_);
  nor (_32291_, _32290_, _32222_);
  or (_32292_, _32291_, _06569_);
  or (_32293_, _32292_, _32289_);
  and (_32294_, _32293_, _32217_);
  or (_32295_, _32294_, _06479_);
  and (_32296_, _14320_, _07970_);
  or (_32297_, _32215_, _09043_);
  or (_32299_, _32297_, _32296_);
  and (_32300_, _32299_, _09048_);
  and (_32301_, _32300_, _32295_);
  and (_32302_, _32284_, _06572_);
  or (_32303_, _32302_, _06606_);
  or (_32304_, _32303_, _32301_);
  or (_32305_, _32223_, _07037_);
  and (_32306_, _32305_, _32304_);
  or (_32307_, _32306_, _06234_);
  or (_32308_, _32215_, _06807_);
  and (_32310_, _32308_, _32307_);
  or (_32311_, _32310_, _06195_);
  or (_32312_, _32223_, _06196_);
  and (_32313_, _32312_, _01375_);
  and (_32314_, _32313_, _32311_);
  or (_43017_, _32314_, _32213_);
  and (_32315_, _13351_, \uc8051golden_1.P1 [1]);
  nor (_32316_, _11223_, _13351_);
  or (_32317_, _32316_, _32315_);
  or (_32318_, _32317_, _09048_);
  nand (_32320_, _07970_, _07090_);
  or (_32321_, _07970_, \uc8051golden_1.P1 [1]);
  and (_32322_, _32321_, _06275_);
  and (_32323_, _32322_, _32320_);
  nor (_32324_, _13351_, _07196_);
  or (_32325_, _32324_, _32315_);
  or (_32326_, _32325_, _07221_);
  and (_32327_, _14532_, _07970_);
  not (_32328_, _32327_);
  and (_32329_, _32328_, _32321_);
  or (_32331_, _32329_, _07210_);
  and (_32332_, _07970_, \uc8051golden_1.ACC [1]);
  or (_32333_, _32332_, _32315_);
  and (_32334_, _32333_, _07199_);
  and (_32335_, _07200_, \uc8051golden_1.P1 [1]);
  or (_32336_, _32335_, _06401_);
  or (_32337_, _32336_, _32334_);
  and (_32338_, _32337_, _06396_);
  and (_32339_, _32338_, _32331_);
  and (_32340_, _13359_, \uc8051golden_1.P1 [1]);
  and (_32342_, _14514_, _08626_);
  or (_32343_, _32342_, _32340_);
  and (_32344_, _32343_, _06395_);
  or (_32345_, _32344_, _06399_);
  or (_32346_, _32345_, _32339_);
  and (_32347_, _32346_, _32326_);
  or (_32348_, _32347_, _06406_);
  or (_32349_, _32333_, _06414_);
  and (_32350_, _32349_, _06844_);
  and (_32351_, _32350_, _32348_);
  and (_32353_, _14517_, _08626_);
  or (_32354_, _32353_, _32340_);
  and (_32355_, _32354_, _06393_);
  or (_32356_, _32355_, _06387_);
  or (_32357_, _32356_, _32351_);
  and (_32358_, _32342_, _14513_);
  or (_32359_, _32340_, _07245_);
  or (_32360_, _32359_, _32358_);
  and (_32361_, _32360_, _06446_);
  and (_32362_, _32361_, _32357_);
  or (_32364_, _32340_, _14560_);
  and (_32365_, _32364_, _06300_);
  and (_32366_, _32365_, _32343_);
  or (_32367_, _32366_, _10059_);
  or (_32368_, _32367_, _32362_);
  or (_32369_, _32325_, _06293_);
  and (_32370_, _32369_, _32368_);
  or (_32371_, _32370_, _06281_);
  and (_32372_, _07970_, _09445_);
  or (_32373_, _32315_, _06282_);
  or (_32375_, _32373_, _32372_);
  and (_32376_, _32375_, _06279_);
  and (_32377_, _32376_, _32371_);
  and (_32378_, _14615_, _07970_);
  or (_32379_, _32378_, _32315_);
  and (_32380_, _32379_, _06015_);
  or (_32381_, _32380_, _32377_);
  and (_32382_, _32381_, _06276_);
  or (_32383_, _32382_, _32323_);
  and (_32384_, _32383_, _07282_);
  or (_32386_, _14507_, _13351_);
  and (_32387_, _32321_, _06474_);
  and (_32388_, _32387_, _32386_);
  or (_32389_, _32388_, _06582_);
  or (_32390_, _32389_, _32384_);
  and (_32391_, _11224_, _07970_);
  or (_32392_, _32391_, _32315_);
  or (_32393_, _32392_, _07284_);
  and (_32394_, _32393_, _07279_);
  and (_32395_, _32394_, _32390_);
  or (_32397_, _14505_, _13351_);
  and (_32398_, _32321_, _06478_);
  and (_32399_, _32398_, _32397_);
  or (_32400_, _32399_, _06569_);
  or (_32401_, _32400_, _32395_);
  and (_32402_, _32332_, _08477_);
  or (_32403_, _32315_, _07276_);
  or (_32404_, _32403_, _32402_);
  and (_32405_, _32404_, _09043_);
  and (_32406_, _32405_, _32401_);
  or (_32408_, _32320_, _08477_);
  and (_32409_, _32321_, _06479_);
  and (_32410_, _32409_, _32408_);
  or (_32411_, _32410_, _06572_);
  or (_32412_, _32411_, _32406_);
  and (_32413_, _32412_, _32318_);
  or (_32414_, _32413_, _06606_);
  or (_32415_, _32329_, _07037_);
  and (_32416_, _32415_, _06807_);
  and (_32417_, _32416_, _32414_);
  and (_32418_, _32354_, _06234_);
  or (_32419_, _32418_, _06195_);
  or (_32420_, _32419_, _32417_);
  or (_32421_, _32315_, _06196_);
  or (_32422_, _32421_, _32327_);
  and (_32423_, _32422_, _01375_);
  and (_32424_, _32423_, _32420_);
  nor (_32425_, \uc8051golden_1.P1 [1], rst);
  nor (_32426_, _32425_, _01382_);
  or (_43018_, _32426_, _32424_);
  and (_32428_, _13351_, \uc8051golden_1.P1 [2]);
  nor (_32429_, _13351_, _07623_);
  or (_32430_, _32429_, _32428_);
  or (_32431_, _32430_, _06293_);
  and (_32432_, _32430_, _06399_);
  and (_32433_, _13359_, \uc8051golden_1.P1 [2]);
  and (_32434_, _14751_, _08626_);
  or (_32435_, _32434_, _32433_);
  or (_32436_, _32435_, _06396_);
  and (_32437_, _14754_, _07970_);
  or (_32439_, _32437_, _32428_);
  and (_32440_, _32439_, _06401_);
  and (_32441_, _07200_, \uc8051golden_1.P1 [2]);
  and (_32442_, _07970_, \uc8051golden_1.ACC [2]);
  or (_32443_, _32442_, _32428_);
  and (_32444_, _32443_, _07199_);
  or (_32445_, _32444_, _32441_);
  and (_32446_, _32445_, _07210_);
  or (_32447_, _32446_, _06395_);
  or (_32448_, _32447_, _32440_);
  and (_32450_, _32448_, _32436_);
  and (_32451_, _32450_, _07221_);
  or (_32452_, _32451_, _32432_);
  or (_32453_, _32452_, _06406_);
  or (_32454_, _32443_, _06414_);
  and (_32455_, _32454_, _06844_);
  and (_32456_, _32455_, _32453_);
  and (_32457_, _14749_, _08626_);
  or (_32458_, _32457_, _32433_);
  and (_32459_, _32458_, _06393_);
  or (_32461_, _32459_, _06387_);
  or (_32462_, _32461_, _32456_);
  or (_32463_, _32433_, _14778_);
  and (_32464_, _32463_, _32435_);
  or (_32465_, _32464_, _07245_);
  and (_32466_, _32465_, _06446_);
  and (_32467_, _32466_, _32462_);
  and (_32468_, _14793_, _08626_);
  or (_32469_, _32468_, _32433_);
  and (_32470_, _32469_, _06300_);
  or (_32472_, _32470_, _10059_);
  or (_32473_, _32472_, _32467_);
  and (_32474_, _32473_, _32431_);
  or (_32475_, _32474_, _06281_);
  and (_32476_, _07970_, _09444_);
  or (_32477_, _32428_, _06282_);
  or (_32478_, _32477_, _32476_);
  and (_32479_, _32478_, _06279_);
  and (_32480_, _32479_, _32475_);
  and (_32481_, _14848_, _07970_);
  or (_32483_, _32481_, _32428_);
  and (_32484_, _32483_, _06015_);
  or (_32485_, _32484_, _06275_);
  or (_32486_, _32485_, _32480_);
  and (_32487_, _07970_, _08994_);
  or (_32488_, _32487_, _32428_);
  or (_32489_, _32488_, _06276_);
  and (_32490_, _32489_, _32486_);
  or (_32491_, _32490_, _06474_);
  and (_32492_, _14744_, _07970_);
  or (_32494_, _32492_, _32428_);
  or (_32495_, _32494_, _07282_);
  and (_32496_, _32495_, _07284_);
  and (_32497_, _32496_, _32491_);
  and (_32498_, _11221_, _07970_);
  or (_32499_, _32498_, _32428_);
  and (_32500_, _32499_, _06582_);
  or (_32501_, _32500_, _32497_);
  and (_32502_, _32501_, _07279_);
  or (_32503_, _32428_, _08433_);
  and (_32505_, _32488_, _06478_);
  and (_32506_, _32505_, _32503_);
  or (_32507_, _32506_, _32502_);
  and (_32508_, _32507_, _07276_);
  and (_32509_, _32443_, _06569_);
  and (_32510_, _32509_, _32503_);
  or (_32511_, _32510_, _06479_);
  or (_32512_, _32511_, _32508_);
  and (_32513_, _14741_, _07970_);
  or (_32514_, _32428_, _09043_);
  or (_32516_, _32514_, _32513_);
  and (_32517_, _32516_, _09048_);
  and (_32518_, _32517_, _32512_);
  nor (_32519_, _11220_, _13351_);
  or (_32520_, _32519_, _32428_);
  and (_32521_, _32520_, _06572_);
  or (_32522_, _32521_, _06606_);
  or (_32523_, _32522_, _32518_);
  or (_32524_, _32439_, _07037_);
  and (_32525_, _32524_, _06807_);
  and (_32527_, _32525_, _32523_);
  and (_32528_, _32458_, _06234_);
  or (_32529_, _32528_, _06195_);
  or (_32530_, _32529_, _32527_);
  and (_32531_, _14917_, _07970_);
  or (_32532_, _32428_, _06196_);
  or (_32533_, _32532_, _32531_);
  and (_32534_, _32533_, _01375_);
  and (_32535_, _32534_, _32530_);
  nor (_32536_, \uc8051golden_1.P1 [2], rst);
  nor (_32538_, _32536_, _01382_);
  or (_43019_, _32538_, _32535_);
  and (_32539_, _13351_, \uc8051golden_1.P1 [3]);
  nor (_32540_, _13351_, _07775_);
  or (_32541_, _32540_, _32539_);
  or (_32542_, _32541_, _06293_);
  and (_32543_, _14947_, _07970_);
  or (_32544_, _32543_, _32539_);
  or (_32545_, _32544_, _07210_);
  and (_32546_, _07970_, \uc8051golden_1.ACC [3]);
  or (_32548_, _32546_, _32539_);
  and (_32549_, _32548_, _07199_);
  and (_32550_, _07200_, \uc8051golden_1.P1 [3]);
  or (_32551_, _32550_, _06401_);
  or (_32552_, _32551_, _32549_);
  and (_32553_, _32552_, _06396_);
  and (_32554_, _32553_, _32545_);
  and (_32555_, _13359_, \uc8051golden_1.P1 [3]);
  and (_32556_, _14951_, _08626_);
  or (_32557_, _32556_, _32555_);
  and (_32559_, _32557_, _06395_);
  or (_32560_, _32559_, _06399_);
  or (_32561_, _32560_, _32554_);
  or (_32562_, _32541_, _07221_);
  and (_32563_, _32562_, _32561_);
  or (_32564_, _32563_, _06406_);
  or (_32565_, _32548_, _06414_);
  and (_32566_, _32565_, _06844_);
  and (_32567_, _32566_, _32564_);
  and (_32568_, _14961_, _08626_);
  or (_32570_, _32568_, _32555_);
  and (_32571_, _32570_, _06393_);
  or (_32572_, _32571_, _06387_);
  or (_32573_, _32572_, _32567_);
  or (_32574_, _32555_, _14968_);
  and (_32575_, _32574_, _32557_);
  or (_32576_, _32575_, _07245_);
  and (_32577_, _32576_, _06446_);
  and (_32578_, _32577_, _32573_);
  and (_32579_, _14985_, _08626_);
  or (_32581_, _32579_, _32555_);
  and (_32582_, _32581_, _06300_);
  or (_32583_, _32582_, _10059_);
  or (_32584_, _32583_, _32578_);
  and (_32585_, _32584_, _32542_);
  or (_32586_, _32585_, _06281_);
  and (_32587_, _07970_, _09443_);
  or (_32588_, _32539_, _06282_);
  or (_32589_, _32588_, _32587_);
  and (_32590_, _32589_, _06279_);
  and (_32592_, _32590_, _32586_);
  and (_32593_, _15039_, _07970_);
  or (_32594_, _32593_, _32539_);
  and (_32595_, _32594_, _06015_);
  or (_32596_, _32595_, _06275_);
  or (_32597_, _32596_, _32592_);
  and (_32598_, _07970_, _08815_);
  or (_32599_, _32598_, _32539_);
  or (_32600_, _32599_, _06276_);
  and (_32601_, _32600_, _32597_);
  or (_32603_, _32601_, _06474_);
  and (_32604_, _14934_, _07970_);
  or (_32605_, _32604_, _32539_);
  or (_32606_, _32605_, _07282_);
  and (_32607_, _32606_, _07284_);
  and (_32608_, _32607_, _32603_);
  and (_32609_, _12535_, _07970_);
  or (_32610_, _32609_, _32539_);
  and (_32611_, _32610_, _06582_);
  or (_32612_, _32611_, _32608_);
  and (_32614_, _32612_, _07279_);
  or (_32615_, _32539_, _08389_);
  and (_32616_, _32599_, _06478_);
  and (_32617_, _32616_, _32615_);
  or (_32618_, _32617_, _32614_);
  and (_32619_, _32618_, _07276_);
  and (_32620_, _32548_, _06569_);
  and (_32621_, _32620_, _32615_);
  or (_32622_, _32621_, _06479_);
  or (_32623_, _32622_, _32619_);
  and (_32625_, _14931_, _07970_);
  or (_32626_, _32539_, _09043_);
  or (_32627_, _32626_, _32625_);
  and (_32628_, _32627_, _09048_);
  and (_32629_, _32628_, _32623_);
  nor (_32630_, _11218_, _13351_);
  or (_32631_, _32630_, _32539_);
  and (_32632_, _32631_, _06572_);
  or (_32633_, _32632_, _06606_);
  or (_32634_, _32633_, _32629_);
  or (_32636_, _32544_, _07037_);
  and (_32637_, _32636_, _06807_);
  and (_32638_, _32637_, _32634_);
  and (_32639_, _32570_, _06234_);
  or (_32640_, _32639_, _06195_);
  or (_32641_, _32640_, _32638_);
  and (_32642_, _15113_, _07970_);
  or (_32643_, _32539_, _06196_);
  or (_32644_, _32643_, _32642_);
  and (_32645_, _32644_, _01375_);
  and (_32647_, _32645_, _32641_);
  nor (_32648_, \uc8051golden_1.P1 [3], rst);
  nor (_32649_, _32648_, _01382_);
  or (_43020_, _32649_, _32647_);
  nor (_32650_, \uc8051golden_1.P1 [4], rst);
  nor (_32651_, _32650_, _01382_);
  and (_32652_, _13351_, \uc8051golden_1.P1 [4]);
  nor (_32653_, _13351_, _08301_);
  or (_32654_, _32653_, _32652_);
  or (_32655_, _32654_, _06293_);
  and (_32657_, _15130_, _07970_);
  or (_32658_, _32657_, _32652_);
  or (_32659_, _32658_, _07210_);
  and (_32660_, _07970_, \uc8051golden_1.ACC [4]);
  or (_32661_, _32660_, _32652_);
  and (_32662_, _32661_, _07199_);
  and (_32663_, _07200_, \uc8051golden_1.P1 [4]);
  or (_32664_, _32663_, _06401_);
  or (_32665_, _32664_, _32662_);
  and (_32666_, _32665_, _06396_);
  and (_32668_, _32666_, _32659_);
  and (_32669_, _13359_, \uc8051golden_1.P1 [4]);
  and (_32670_, _15139_, _08626_);
  or (_32671_, _32670_, _32669_);
  and (_32672_, _32671_, _06395_);
  or (_32673_, _32672_, _06399_);
  or (_32674_, _32673_, _32668_);
  or (_32675_, _32654_, _07221_);
  and (_32676_, _32675_, _32674_);
  or (_32677_, _32676_, _06406_);
  or (_32679_, _32661_, _06414_);
  and (_32680_, _32679_, _06844_);
  and (_32681_, _32680_, _32677_);
  and (_32682_, _15168_, _08626_);
  or (_32683_, _32682_, _32669_);
  and (_32684_, _32683_, _06393_);
  or (_32685_, _32684_, _06387_);
  or (_32686_, _32685_, _32681_);
  or (_32687_, _32669_, _15138_);
  and (_32688_, _32687_, _32671_);
  or (_32690_, _32688_, _07245_);
  and (_32691_, _32690_, _06446_);
  and (_32692_, _32691_, _32686_);
  and (_32693_, _15189_, _08626_);
  or (_32694_, _32693_, _32669_);
  and (_32695_, _32694_, _06300_);
  or (_32696_, _32695_, _10059_);
  or (_32697_, _32696_, _32692_);
  and (_32698_, _32697_, _32655_);
  or (_32699_, _32698_, _06281_);
  and (_32701_, _07970_, _09442_);
  or (_32702_, _32652_, _06282_);
  or (_32703_, _32702_, _32701_);
  and (_32704_, _32703_, _06279_);
  and (_32705_, _32704_, _32699_);
  and (_32706_, _15243_, _07970_);
  or (_32707_, _32706_, _32652_);
  and (_32708_, _32707_, _06015_);
  or (_32709_, _32708_, _06275_);
  or (_32710_, _32709_, _32705_);
  and (_32712_, _08883_, _07970_);
  or (_32713_, _32712_, _32652_);
  or (_32714_, _32713_, _06276_);
  and (_32715_, _32714_, _32710_);
  or (_32716_, _32715_, _06474_);
  and (_32717_, _15135_, _07970_);
  or (_32718_, _32717_, _32652_);
  or (_32719_, _32718_, _07282_);
  and (_32720_, _32719_, _07284_);
  and (_32721_, _32720_, _32716_);
  and (_32723_, _11216_, _07970_);
  or (_32724_, _32723_, _32652_);
  and (_32725_, _32724_, _06582_);
  or (_32726_, _32725_, _32721_);
  and (_32727_, _32726_, _07279_);
  or (_32728_, _32652_, _08345_);
  and (_32729_, _32713_, _06478_);
  and (_32730_, _32729_, _32728_);
  or (_32731_, _32730_, _32727_);
  and (_32732_, _32731_, _07276_);
  and (_32734_, _32661_, _06569_);
  and (_32735_, _32734_, _32728_);
  or (_32736_, _32735_, _06479_);
  or (_32737_, _32736_, _32732_);
  and (_32738_, _15134_, _07970_);
  or (_32739_, _32652_, _09043_);
  or (_32740_, _32739_, _32738_);
  and (_32741_, _32740_, _09048_);
  and (_32742_, _32741_, _32737_);
  nor (_32743_, _11215_, _13351_);
  or (_32745_, _32743_, _32652_);
  and (_32746_, _32745_, _06572_);
  or (_32747_, _32746_, _06606_);
  or (_32748_, _32747_, _32742_);
  or (_32749_, _32658_, _07037_);
  and (_32750_, _32749_, _06807_);
  and (_32751_, _32750_, _32748_);
  and (_32752_, _32683_, _06234_);
  or (_32753_, _32752_, _06195_);
  or (_32754_, _32753_, _32751_);
  and (_32756_, _15315_, _07970_);
  or (_32757_, _32652_, _06196_);
  or (_32758_, _32757_, _32756_);
  and (_32759_, _32758_, _01375_);
  and (_32760_, _32759_, _32754_);
  or (_43021_, _32760_, _32651_);
  and (_32761_, _13351_, \uc8051golden_1.P1 [5]);
  nor (_32762_, _13351_, _08207_);
  or (_32763_, _32762_, _32761_);
  or (_32764_, _32763_, _06293_);
  and (_32766_, _15348_, _07970_);
  or (_32767_, _32766_, _32761_);
  or (_32768_, _32767_, _07210_);
  and (_32769_, _07970_, \uc8051golden_1.ACC [5]);
  or (_32770_, _32769_, _32761_);
  and (_32771_, _32770_, _07199_);
  and (_32772_, _07200_, \uc8051golden_1.P1 [5]);
  or (_32773_, _32772_, _06401_);
  or (_32774_, _32773_, _32771_);
  and (_32775_, _32774_, _06396_);
  and (_32777_, _32775_, _32768_);
  and (_32778_, _13359_, \uc8051golden_1.P1 [5]);
  and (_32779_, _15341_, _08626_);
  or (_32780_, _32779_, _32778_);
  and (_32781_, _32780_, _06395_);
  or (_32782_, _32781_, _06399_);
  or (_32783_, _32782_, _32777_);
  or (_32784_, _32763_, _07221_);
  and (_32785_, _32784_, _32783_);
  or (_32786_, _32785_, _06406_);
  or (_32788_, _32770_, _06414_);
  and (_32789_, _32788_, _06844_);
  and (_32790_, _32789_, _32786_);
  and (_32791_, _15345_, _08626_);
  or (_32792_, _32791_, _32778_);
  and (_32793_, _32792_, _06393_);
  or (_32794_, _32793_, _06387_);
  or (_32795_, _32794_, _32790_);
  or (_32796_, _32778_, _15378_);
  and (_32797_, _32796_, _32780_);
  or (_32799_, _32797_, _07245_);
  and (_32800_, _32799_, _06446_);
  and (_32801_, _32800_, _32795_);
  or (_32802_, _32778_, _15342_);
  and (_32803_, _32802_, _06300_);
  and (_32804_, _32803_, _32780_);
  or (_32805_, _32804_, _10059_);
  or (_32806_, _32805_, _32801_);
  and (_32807_, _32806_, _32764_);
  or (_32808_, _32807_, _06281_);
  and (_32810_, _07970_, _09441_);
  or (_32811_, _32761_, _06282_);
  or (_32812_, _32811_, _32810_);
  and (_32813_, _32812_, _06279_);
  and (_32814_, _32813_, _32808_);
  and (_32815_, _15446_, _07970_);
  or (_32816_, _32815_, _32761_);
  and (_32817_, _32816_, _06015_);
  or (_32818_, _32817_, _06275_);
  or (_32819_, _32818_, _32814_);
  and (_32821_, _08958_, _07970_);
  or (_32822_, _32821_, _32761_);
  or (_32823_, _32822_, _06276_);
  and (_32824_, _32823_, _32819_);
  or (_32825_, _32824_, _06474_);
  and (_32826_, _15338_, _07970_);
  or (_32827_, _32826_, _32761_);
  or (_32828_, _32827_, _07282_);
  and (_32829_, _32828_, _07284_);
  and (_32830_, _32829_, _32825_);
  and (_32832_, _12542_, _07970_);
  or (_32833_, _32832_, _32761_);
  and (_32834_, _32833_, _06582_);
  or (_32835_, _32834_, _32830_);
  and (_32836_, _32835_, _07279_);
  or (_32837_, _32761_, _08256_);
  and (_32838_, _32822_, _06478_);
  and (_32839_, _32838_, _32837_);
  or (_32840_, _32839_, _32836_);
  and (_32841_, _32840_, _07276_);
  and (_32843_, _32770_, _06569_);
  and (_32844_, _32843_, _32837_);
  or (_32845_, _32844_, _06479_);
  or (_32846_, _32845_, _32841_);
  and (_32847_, _15335_, _07970_);
  or (_32848_, _32761_, _09043_);
  or (_32849_, _32848_, _32847_);
  and (_32850_, _32849_, _09048_);
  and (_32851_, _32850_, _32846_);
  nor (_32852_, _11212_, _13351_);
  or (_32854_, _32852_, _32761_);
  and (_32855_, _32854_, _06572_);
  or (_32856_, _32855_, _06606_);
  or (_32857_, _32856_, _32851_);
  or (_32858_, _32767_, _07037_);
  and (_32859_, _32858_, _06807_);
  and (_32860_, _32859_, _32857_);
  and (_32861_, _32792_, _06234_);
  or (_32862_, _32861_, _06195_);
  or (_32863_, _32862_, _32860_);
  and (_32865_, _15509_, _07970_);
  or (_32866_, _32761_, _06196_);
  or (_32867_, _32866_, _32865_);
  and (_32868_, _32867_, _01375_);
  and (_32869_, _32868_, _32863_);
  nor (_32870_, \uc8051golden_1.P1 [5], rst);
  nor (_32871_, _32870_, _01382_);
  or (_43022_, _32871_, _32869_);
  and (_32872_, _13351_, \uc8051golden_1.P1 [6]);
  nor (_32873_, _13351_, _08118_);
  or (_32875_, _32873_, _32872_);
  or (_32876_, _32875_, _06293_);
  and (_32877_, _15550_, _07970_);
  or (_32878_, _32877_, _32872_);
  or (_32879_, _32878_, _07210_);
  and (_32880_, _07970_, \uc8051golden_1.ACC [6]);
  or (_32881_, _32880_, _32872_);
  and (_32882_, _32881_, _07199_);
  and (_32883_, _07200_, \uc8051golden_1.P1 [6]);
  or (_32884_, _32883_, _06401_);
  or (_32886_, _32884_, _32882_);
  and (_32887_, _32886_, _06396_);
  and (_32888_, _32887_, _32879_);
  and (_32889_, _13359_, \uc8051golden_1.P1 [6]);
  and (_32890_, _15535_, _08626_);
  or (_32891_, _32890_, _32889_);
  and (_32892_, _32891_, _06395_);
  or (_32893_, _32892_, _06399_);
  or (_32894_, _32893_, _32888_);
  or (_32895_, _32875_, _07221_);
  and (_32897_, _32895_, _32894_);
  or (_32898_, _32897_, _06406_);
  or (_32899_, _32881_, _06414_);
  and (_32900_, _32899_, _06844_);
  and (_32901_, _32900_, _32898_);
  and (_32902_, _15561_, _08626_);
  or (_32903_, _32902_, _32889_);
  and (_32904_, _32903_, _06393_);
  or (_32905_, _32904_, _06387_);
  or (_32906_, _32905_, _32901_);
  or (_32908_, _32889_, _15568_);
  and (_32909_, _32908_, _32891_);
  or (_32910_, _32909_, _07245_);
  and (_32911_, _32910_, _06446_);
  and (_32912_, _32911_, _32906_);
  and (_32913_, _15585_, _08626_);
  or (_32914_, _32913_, _32889_);
  and (_32915_, _32914_, _06300_);
  or (_32916_, _32915_, _10059_);
  or (_32917_, _32916_, _32912_);
  and (_32919_, _32917_, _32876_);
  or (_32920_, _32919_, _06281_);
  and (_32921_, _07970_, _09440_);
  or (_32922_, _32872_, _06282_);
  or (_32923_, _32922_, _32921_);
  and (_32924_, _32923_, _06279_);
  and (_32925_, _32924_, _32920_);
  and (_32926_, _15639_, _07970_);
  or (_32927_, _32926_, _32872_);
  and (_32928_, _32927_, _06015_);
  or (_32930_, _32928_, _06275_);
  or (_32931_, _32930_, _32925_);
  and (_32932_, _15646_, _07970_);
  or (_32933_, _32932_, _32872_);
  or (_32934_, _32933_, _06276_);
  and (_32935_, _32934_, _32931_);
  or (_32936_, _32935_, _06474_);
  and (_32937_, _15531_, _07970_);
  or (_32938_, _32937_, _32872_);
  or (_32939_, _32938_, _07282_);
  and (_32941_, _32939_, _07284_);
  and (_32942_, _32941_, _32936_);
  and (_32943_, _11210_, _07970_);
  or (_32944_, _32943_, _32872_);
  and (_32945_, _32944_, _06582_);
  or (_32946_, _32945_, _32942_);
  and (_32947_, _32946_, _07279_);
  or (_32948_, _32872_, _08162_);
  and (_32949_, _32933_, _06478_);
  and (_32950_, _32949_, _32948_);
  or (_32952_, _32950_, _32947_);
  and (_32953_, _32952_, _07276_);
  and (_32954_, _32881_, _06569_);
  and (_32955_, _32954_, _32948_);
  or (_32956_, _32955_, _06479_);
  or (_32957_, _32956_, _32953_);
  and (_32958_, _15528_, _07970_);
  or (_32959_, _32872_, _09043_);
  or (_32960_, _32959_, _32958_);
  and (_32961_, _32960_, _09048_);
  and (_32963_, _32961_, _32957_);
  nor (_32964_, _11209_, _13351_);
  or (_32965_, _32964_, _32872_);
  and (_32966_, _32965_, _06572_);
  or (_32967_, _32966_, _06606_);
  or (_32968_, _32967_, _32963_);
  or (_32969_, _32878_, _07037_);
  and (_32970_, _32969_, _06807_);
  and (_32971_, _32970_, _32968_);
  and (_32972_, _32903_, _06234_);
  or (_32974_, _32972_, _06195_);
  or (_32975_, _32974_, _32971_);
  and (_32976_, _15713_, _07970_);
  or (_32977_, _32872_, _06196_);
  or (_32978_, _32977_, _32976_);
  and (_32979_, _32978_, _01375_);
  and (_32980_, _32979_, _32975_);
  nor (_32981_, \uc8051golden_1.P1 [6], rst);
  nor (_32982_, _32981_, _01382_);
  or (_43023_, _32982_, _32980_);
  not (_32984_, \uc8051golden_1.IP [0]);
  nor (_32985_, _01375_, _32984_);
  nand (_32986_, _11225_, _07999_);
  nor (_32987_, _07999_, _32984_);
  nor (_32988_, _32987_, _07276_);
  nand (_32989_, _32988_, _32986_);
  nor (_32990_, _08521_, _13453_);
  or (_32991_, _32990_, _32987_);
  and (_32992_, _32991_, _06401_);
  nor (_32993_, _07199_, _32984_);
  and (_32995_, _07999_, \uc8051golden_1.ACC [0]);
  or (_32996_, _32995_, _32987_);
  and (_32997_, _32996_, _07199_);
  or (_32998_, _32997_, _32993_);
  and (_32999_, _32998_, _07210_);
  or (_33000_, _32999_, _06395_);
  or (_33001_, _33000_, _32992_);
  and (_33002_, _14339_, _08614_);
  nor (_33003_, _08614_, _32984_);
  or (_33004_, _33003_, _06396_);
  or (_33006_, _33004_, _33002_);
  and (_33007_, _33006_, _07221_);
  and (_33008_, _33007_, _33001_);
  and (_33009_, _07999_, _07473_);
  or (_33010_, _33009_, _32987_);
  and (_33011_, _33010_, _06399_);
  or (_33012_, _33011_, _06406_);
  or (_33013_, _33012_, _33008_);
  or (_33014_, _32996_, _06414_);
  and (_33015_, _33014_, _06844_);
  and (_33017_, _33015_, _33013_);
  and (_33018_, _32987_, _06393_);
  or (_33019_, _33018_, _06387_);
  or (_33020_, _33019_, _33017_);
  or (_33021_, _32991_, _07245_);
  and (_33022_, _33021_, _06446_);
  and (_33023_, _33022_, _33020_);
  and (_33024_, _14371_, _08614_);
  or (_33025_, _33024_, _33003_);
  and (_33026_, _33025_, _06300_);
  or (_33028_, _33026_, _10059_);
  or (_33029_, _33028_, _33023_);
  or (_33030_, _33010_, _06293_);
  and (_33031_, _33030_, _33029_);
  or (_33032_, _33031_, _06281_);
  and (_33033_, _07999_, _09446_);
  or (_33034_, _32987_, _06282_);
  or (_33035_, _33034_, _33033_);
  and (_33036_, _33035_, _06279_);
  and (_33037_, _33036_, _33032_);
  and (_33039_, _14426_, _07999_);
  or (_33040_, _33039_, _32987_);
  and (_33041_, _33040_, _06015_);
  or (_33042_, _33041_, _06275_);
  or (_33043_, _33042_, _33037_);
  and (_33044_, _07999_, _08817_);
  or (_33045_, _33044_, _32987_);
  or (_33046_, _33045_, _06276_);
  and (_33047_, _33046_, _33043_);
  or (_33048_, _33047_, _06474_);
  and (_33050_, _14324_, _07999_);
  or (_33051_, _33050_, _32987_);
  or (_33052_, _33051_, _07282_);
  and (_33053_, _33052_, _07284_);
  and (_33054_, _33053_, _33048_);
  nor (_33055_, _12538_, _13453_);
  or (_33056_, _33055_, _32987_);
  and (_33057_, _32986_, _06582_);
  and (_33058_, _33057_, _33056_);
  or (_33059_, _33058_, _33054_);
  and (_33061_, _33059_, _07279_);
  nand (_33062_, _33045_, _06478_);
  nor (_33063_, _33062_, _32990_);
  or (_33064_, _33063_, _06569_);
  or (_33065_, _33064_, _33061_);
  and (_33066_, _33065_, _32989_);
  or (_33067_, _33066_, _06479_);
  and (_33068_, _14320_, _07999_);
  or (_33069_, _33068_, _32987_);
  or (_33070_, _33069_, _09043_);
  and (_33072_, _33070_, _09048_);
  and (_33073_, _33072_, _33067_);
  and (_33074_, _33056_, _06572_);
  or (_33075_, _33074_, _06606_);
  or (_33076_, _33075_, _33073_);
  or (_33077_, _32991_, _07037_);
  and (_33078_, _33077_, _33076_);
  or (_33079_, _33078_, _06234_);
  or (_33080_, _32987_, _06807_);
  and (_33081_, _33080_, _33079_);
  or (_33083_, _33081_, _06195_);
  or (_33084_, _32991_, _06196_);
  and (_33085_, _33084_, _01375_);
  and (_33086_, _33085_, _33083_);
  or (_33087_, _33086_, _32985_);
  and (_43025_, _33087_, _42545_);
  not (_33088_, \uc8051golden_1.IP [1]);
  nor (_33089_, _01375_, _33088_);
  nor (_33090_, _07999_, _33088_);
  nor (_33091_, _11223_, _13453_);
  or (_33093_, _33091_, _33090_);
  or (_33094_, _33093_, _09048_);
  nand (_33095_, _07999_, _07090_);
  or (_33096_, _07999_, \uc8051golden_1.IP [1]);
  and (_33097_, _33096_, _06275_);
  and (_33098_, _33097_, _33095_);
  nor (_33099_, _13453_, _07196_);
  or (_33100_, _33099_, _33090_);
  or (_33101_, _33100_, _07221_);
  and (_33102_, _14532_, _07999_);
  not (_33103_, _33102_);
  and (_33104_, _33103_, _33096_);
  or (_33105_, _33104_, _07210_);
  and (_33106_, _07999_, \uc8051golden_1.ACC [1]);
  or (_33107_, _33106_, _33090_);
  and (_33108_, _33107_, _07199_);
  nor (_33109_, _07199_, _33088_);
  or (_33110_, _33109_, _06401_);
  or (_33111_, _33110_, _33108_);
  and (_33112_, _33111_, _06396_);
  and (_33114_, _33112_, _33105_);
  nor (_33115_, _08614_, _33088_);
  and (_33116_, _14514_, _08614_);
  or (_33117_, _33116_, _33115_);
  and (_33118_, _33117_, _06395_);
  or (_33119_, _33118_, _06399_);
  or (_33120_, _33119_, _33114_);
  and (_33121_, _33120_, _33101_);
  or (_33122_, _33121_, _06406_);
  or (_33123_, _33107_, _06414_);
  and (_33125_, _33123_, _06844_);
  and (_33126_, _33125_, _33122_);
  and (_33127_, _14517_, _08614_);
  or (_33128_, _33127_, _33115_);
  and (_33129_, _33128_, _06393_);
  or (_33130_, _33129_, _06387_);
  or (_33131_, _33130_, _33126_);
  and (_33132_, _33116_, _14513_);
  or (_33133_, _33115_, _07245_);
  or (_33134_, _33133_, _33132_);
  and (_33136_, _33134_, _06446_);
  and (_33137_, _33136_, _33131_);
  or (_33138_, _33115_, _14560_);
  and (_33139_, _33138_, _06300_);
  and (_33140_, _33139_, _33117_);
  or (_33141_, _33140_, _10059_);
  or (_33142_, _33141_, _33137_);
  or (_33143_, _33100_, _06293_);
  and (_33144_, _33143_, _33142_);
  or (_33145_, _33144_, _06281_);
  and (_33147_, _07999_, _09445_);
  or (_33148_, _33090_, _06282_);
  or (_33149_, _33148_, _33147_);
  and (_33150_, _33149_, _06279_);
  and (_33151_, _33150_, _33145_);
  and (_33152_, _14615_, _07999_);
  or (_33153_, _33152_, _33090_);
  and (_33154_, _33153_, _06015_);
  or (_33155_, _33154_, _33151_);
  and (_33156_, _33155_, _06276_);
  or (_33158_, _33156_, _33098_);
  and (_33159_, _33158_, _07282_);
  or (_33160_, _14507_, _13453_);
  and (_33161_, _33096_, _06474_);
  and (_33162_, _33161_, _33160_);
  or (_33163_, _33162_, _06582_);
  or (_33164_, _33163_, _33159_);
  nand (_33165_, _11222_, _07999_);
  and (_33166_, _33165_, _33093_);
  or (_33167_, _33166_, _07284_);
  and (_33169_, _33167_, _07279_);
  and (_33170_, _33169_, _33164_);
  or (_33171_, _14505_, _13453_);
  and (_33172_, _33096_, _06478_);
  and (_33173_, _33172_, _33171_);
  or (_33174_, _33173_, _06569_);
  or (_33175_, _33174_, _33170_);
  nor (_33176_, _33090_, _07276_);
  nand (_33177_, _33176_, _33165_);
  and (_33178_, _33177_, _09043_);
  and (_33180_, _33178_, _33175_);
  or (_33181_, _33095_, _08477_);
  and (_33182_, _33096_, _06479_);
  and (_33183_, _33182_, _33181_);
  or (_33184_, _33183_, _06572_);
  or (_33185_, _33184_, _33180_);
  and (_33186_, _33185_, _33094_);
  or (_33187_, _33186_, _06606_);
  or (_33188_, _33104_, _07037_);
  and (_33189_, _33188_, _06807_);
  and (_33191_, _33189_, _33187_);
  and (_33192_, _33128_, _06234_);
  or (_33193_, _33192_, _06195_);
  or (_33194_, _33193_, _33191_);
  or (_33195_, _33090_, _06196_);
  or (_33196_, _33195_, _33102_);
  and (_33197_, _33196_, _01375_);
  and (_33198_, _33197_, _33194_);
  or (_33199_, _33198_, _33089_);
  and (_43026_, _33199_, _42545_);
  and (_33201_, _01379_, \uc8051golden_1.IP [2]);
  and (_33202_, _13453_, \uc8051golden_1.IP [2]);
  nor (_33203_, _13453_, _07623_);
  or (_33204_, _33203_, _33202_);
  or (_33205_, _33204_, _06293_);
  or (_33206_, _33204_, _07221_);
  and (_33207_, _14754_, _07999_);
  or (_33208_, _33207_, _33202_);
  or (_33209_, _33208_, _07210_);
  and (_33210_, _07999_, \uc8051golden_1.ACC [2]);
  or (_33212_, _33210_, _33202_);
  and (_33213_, _33212_, _07199_);
  and (_33214_, _07200_, \uc8051golden_1.IP [2]);
  or (_33215_, _33214_, _06401_);
  or (_33216_, _33215_, _33213_);
  and (_33217_, _33216_, _06396_);
  and (_33218_, _33217_, _33209_);
  and (_33219_, _13461_, \uc8051golden_1.IP [2]);
  and (_33220_, _14751_, _08614_);
  or (_33221_, _33220_, _33219_);
  and (_33223_, _33221_, _06395_);
  or (_33224_, _33223_, _06399_);
  or (_33225_, _33224_, _33218_);
  and (_33226_, _33225_, _33206_);
  or (_33227_, _33226_, _06406_);
  or (_33228_, _33212_, _06414_);
  and (_33229_, _33228_, _06844_);
  and (_33230_, _33229_, _33227_);
  and (_33231_, _14749_, _08614_);
  or (_33232_, _33231_, _33219_);
  and (_33234_, _33232_, _06393_);
  or (_33235_, _33234_, _06387_);
  or (_33236_, _33235_, _33230_);
  and (_33237_, _33220_, _14778_);
  or (_33238_, _33219_, _07245_);
  or (_33239_, _33238_, _33237_);
  and (_33240_, _33239_, _06446_);
  and (_33241_, _33240_, _33236_);
  and (_33242_, _14793_, _08614_);
  or (_33243_, _33242_, _33219_);
  and (_33245_, _33243_, _06300_);
  or (_33246_, _33245_, _10059_);
  or (_33247_, _33246_, _33241_);
  and (_33248_, _33247_, _33205_);
  or (_33249_, _33248_, _06281_);
  and (_33250_, _07999_, _09444_);
  or (_33251_, _33202_, _06282_);
  or (_33252_, _33251_, _33250_);
  and (_33253_, _33252_, _06279_);
  and (_33254_, _33253_, _33249_);
  and (_33256_, _14848_, _07999_);
  or (_33257_, _33256_, _33202_);
  and (_33258_, _33257_, _06015_);
  or (_33259_, _33258_, _06275_);
  or (_33260_, _33259_, _33254_);
  and (_33261_, _07999_, _08994_);
  or (_33262_, _33261_, _33202_);
  or (_33263_, _33262_, _06276_);
  and (_33264_, _33263_, _33260_);
  or (_33265_, _33264_, _06474_);
  and (_33267_, _14744_, _07999_);
  or (_33268_, _33267_, _33202_);
  or (_33269_, _33268_, _07282_);
  and (_33270_, _33269_, _07284_);
  and (_33271_, _33270_, _33265_);
  and (_33272_, _11221_, _07999_);
  or (_33273_, _33272_, _33202_);
  and (_33274_, _33273_, _06582_);
  or (_33275_, _33274_, _33271_);
  and (_33276_, _33275_, _07279_);
  or (_33278_, _33202_, _08433_);
  and (_33279_, _33262_, _06478_);
  and (_33280_, _33279_, _33278_);
  or (_33281_, _33280_, _33276_);
  and (_33282_, _33281_, _07276_);
  and (_33283_, _33212_, _06569_);
  and (_33284_, _33283_, _33278_);
  or (_33285_, _33284_, _06479_);
  or (_33286_, _33285_, _33282_);
  and (_33287_, _14741_, _07999_);
  or (_33289_, _33202_, _09043_);
  or (_33290_, _33289_, _33287_);
  and (_33291_, _33290_, _09048_);
  and (_33292_, _33291_, _33286_);
  nor (_33293_, _11220_, _13453_);
  or (_33294_, _33293_, _33202_);
  and (_33295_, _33294_, _06572_);
  or (_33296_, _33295_, _06606_);
  or (_33297_, _33296_, _33292_);
  or (_33298_, _33208_, _07037_);
  and (_33300_, _33298_, _06807_);
  and (_33301_, _33300_, _33297_);
  and (_33302_, _33232_, _06234_);
  or (_33303_, _33302_, _06195_);
  or (_33304_, _33303_, _33301_);
  and (_33305_, _14917_, _07999_);
  or (_33306_, _33202_, _06196_);
  or (_33307_, _33306_, _33305_);
  and (_33308_, _33307_, _01375_);
  and (_33309_, _33308_, _33304_);
  or (_33311_, _33309_, _33201_);
  and (_43027_, _33311_, _42545_);
  and (_33312_, _01379_, \uc8051golden_1.IP [3]);
  and (_33313_, _13453_, \uc8051golden_1.IP [3]);
  nor (_33314_, _13453_, _07775_);
  or (_33315_, _33314_, _33313_);
  or (_33316_, _33315_, _06293_);
  and (_33317_, _14947_, _07999_);
  or (_33318_, _33317_, _33313_);
  or (_33319_, _33318_, _07210_);
  and (_33321_, _07999_, \uc8051golden_1.ACC [3]);
  or (_33322_, _33321_, _33313_);
  and (_33323_, _33322_, _07199_);
  and (_33324_, _07200_, \uc8051golden_1.IP [3]);
  or (_33325_, _33324_, _06401_);
  or (_33326_, _33325_, _33323_);
  and (_33327_, _33326_, _06396_);
  and (_33328_, _33327_, _33319_);
  and (_33329_, _13461_, \uc8051golden_1.IP [3]);
  and (_33330_, _14951_, _08614_);
  or (_33332_, _33330_, _33329_);
  and (_33333_, _33332_, _06395_);
  or (_33334_, _33333_, _06399_);
  or (_33335_, _33334_, _33328_);
  or (_33336_, _33315_, _07221_);
  and (_33337_, _33336_, _33335_);
  or (_33338_, _33337_, _06406_);
  or (_33339_, _33322_, _06414_);
  and (_33340_, _33339_, _06844_);
  and (_33341_, _33340_, _33338_);
  and (_33343_, _14961_, _08614_);
  or (_33344_, _33343_, _33329_);
  and (_33345_, _33344_, _06393_);
  or (_33346_, _33345_, _06387_);
  or (_33347_, _33346_, _33341_);
  or (_33348_, _33329_, _14968_);
  and (_33349_, _33348_, _33332_);
  or (_33350_, _33349_, _07245_);
  and (_33351_, _33350_, _06446_);
  and (_33352_, _33351_, _33347_);
  and (_33354_, _14985_, _08614_);
  or (_33355_, _33354_, _33329_);
  and (_33356_, _33355_, _06300_);
  or (_33357_, _33356_, _10059_);
  or (_33358_, _33357_, _33352_);
  and (_33359_, _33358_, _33316_);
  or (_33360_, _33359_, _06281_);
  and (_33361_, _07999_, _09443_);
  or (_33362_, _33313_, _06282_);
  or (_33363_, _33362_, _33361_);
  and (_33365_, _33363_, _06279_);
  and (_33366_, _33365_, _33360_);
  and (_33367_, _15039_, _07999_);
  or (_33368_, _33367_, _33313_);
  and (_33369_, _33368_, _06015_);
  or (_33370_, _33369_, _06275_);
  or (_33371_, _33370_, _33366_);
  and (_33372_, _07999_, _08815_);
  or (_33373_, _33372_, _33313_);
  or (_33374_, _33373_, _06276_);
  and (_33376_, _33374_, _33371_);
  or (_33377_, _33376_, _06474_);
  and (_33378_, _14934_, _07999_);
  or (_33379_, _33378_, _33313_);
  or (_33380_, _33379_, _07282_);
  and (_33381_, _33380_, _07284_);
  and (_33382_, _33381_, _33377_);
  and (_33383_, _12535_, _07999_);
  or (_33384_, _33383_, _33313_);
  and (_33385_, _33384_, _06582_);
  or (_33387_, _33385_, _33382_);
  and (_33388_, _33387_, _07279_);
  or (_33389_, _33313_, _08389_);
  and (_33390_, _33373_, _06478_);
  and (_33391_, _33390_, _33389_);
  or (_33392_, _33391_, _33388_);
  and (_33393_, _33392_, _07276_);
  and (_33394_, _33322_, _06569_);
  and (_33395_, _33394_, _33389_);
  or (_33396_, _33395_, _06479_);
  or (_33398_, _33396_, _33393_);
  and (_33399_, _14931_, _07999_);
  or (_33400_, _33313_, _09043_);
  or (_33401_, _33400_, _33399_);
  and (_33402_, _33401_, _09048_);
  and (_33403_, _33402_, _33398_);
  nor (_33404_, _11218_, _13453_);
  or (_33405_, _33404_, _33313_);
  and (_33406_, _33405_, _06572_);
  or (_33407_, _33406_, _06606_);
  or (_33409_, _33407_, _33403_);
  or (_33410_, _33318_, _07037_);
  and (_33411_, _33410_, _06807_);
  and (_33412_, _33411_, _33409_);
  and (_33413_, _33344_, _06234_);
  or (_33414_, _33413_, _06195_);
  or (_33415_, _33414_, _33412_);
  and (_33416_, _15113_, _07999_);
  or (_33417_, _33313_, _06196_);
  or (_33418_, _33417_, _33416_);
  and (_33420_, _33418_, _01375_);
  and (_33421_, _33420_, _33415_);
  or (_33422_, _33421_, _33312_);
  and (_43028_, _33422_, _42545_);
  and (_33423_, _01379_, \uc8051golden_1.IP [4]);
  and (_33424_, _13453_, \uc8051golden_1.IP [4]);
  nor (_33425_, _13453_, _08301_);
  or (_33426_, _33425_, _33424_);
  or (_33427_, _33426_, _06293_);
  and (_33428_, _15130_, _07999_);
  or (_33430_, _33428_, _33424_);
  or (_33431_, _33430_, _07210_);
  and (_33432_, _07999_, \uc8051golden_1.ACC [4]);
  or (_33433_, _33432_, _33424_);
  and (_33434_, _33433_, _07199_);
  and (_33435_, _07200_, \uc8051golden_1.IP [4]);
  or (_33436_, _33435_, _06401_);
  or (_33437_, _33436_, _33434_);
  and (_33438_, _33437_, _06396_);
  and (_33439_, _33438_, _33431_);
  and (_33441_, _13461_, \uc8051golden_1.IP [4]);
  and (_33442_, _15139_, _08614_);
  or (_33443_, _33442_, _33441_);
  and (_33444_, _33443_, _06395_);
  or (_33445_, _33444_, _06399_);
  or (_33446_, _33445_, _33439_);
  or (_33447_, _33426_, _07221_);
  and (_33448_, _33447_, _33446_);
  or (_33449_, _33448_, _06406_);
  or (_33450_, _33433_, _06414_);
  and (_33452_, _33450_, _06844_);
  and (_33453_, _33452_, _33449_);
  and (_33454_, _15168_, _08614_);
  or (_33455_, _33454_, _33441_);
  and (_33456_, _33455_, _06393_);
  or (_33457_, _33456_, _06387_);
  or (_33458_, _33457_, _33453_);
  or (_33459_, _33441_, _15138_);
  and (_33460_, _33459_, _33443_);
  or (_33461_, _33460_, _07245_);
  and (_33463_, _33461_, _06446_);
  and (_33464_, _33463_, _33458_);
  and (_33465_, _15189_, _08614_);
  or (_33466_, _33465_, _33441_);
  and (_33467_, _33466_, _06300_);
  or (_33468_, _33467_, _10059_);
  or (_33469_, _33468_, _33464_);
  and (_33470_, _33469_, _33427_);
  or (_33471_, _33470_, _06281_);
  and (_33472_, _07999_, _09442_);
  or (_33474_, _33424_, _06282_);
  or (_33475_, _33474_, _33472_);
  and (_33476_, _33475_, _06279_);
  and (_33477_, _33476_, _33471_);
  and (_33478_, _15243_, _07999_);
  or (_33479_, _33478_, _33424_);
  and (_33480_, _33479_, _06015_);
  or (_33481_, _33480_, _06275_);
  or (_33482_, _33481_, _33477_);
  and (_33483_, _08883_, _07999_);
  or (_33485_, _33483_, _33424_);
  or (_33486_, _33485_, _06276_);
  and (_33487_, _33486_, _33482_);
  or (_33488_, _33487_, _06474_);
  and (_33489_, _15135_, _07999_);
  or (_33490_, _33489_, _33424_);
  or (_33491_, _33490_, _07282_);
  and (_33492_, _33491_, _07284_);
  and (_33493_, _33492_, _33488_);
  and (_33494_, _11216_, _07999_);
  or (_33496_, _33494_, _33424_);
  and (_33497_, _33496_, _06582_);
  or (_33498_, _33497_, _33493_);
  and (_33499_, _33498_, _07279_);
  or (_33500_, _33424_, _08345_);
  and (_33501_, _33485_, _06478_);
  and (_33502_, _33501_, _33500_);
  or (_33503_, _33502_, _33499_);
  and (_33504_, _33503_, _07276_);
  and (_33505_, _33433_, _06569_);
  and (_33507_, _33505_, _33500_);
  or (_33508_, _33507_, _06479_);
  or (_33509_, _33508_, _33504_);
  and (_33510_, _15134_, _07999_);
  or (_33511_, _33424_, _09043_);
  or (_33512_, _33511_, _33510_);
  and (_33513_, _33512_, _09048_);
  and (_33514_, _33513_, _33509_);
  nor (_33515_, _11215_, _13453_);
  or (_33516_, _33515_, _33424_);
  and (_33518_, _33516_, _06572_);
  or (_33519_, _33518_, _06606_);
  or (_33520_, _33519_, _33514_);
  or (_33521_, _33430_, _07037_);
  and (_33522_, _33521_, _06807_);
  and (_33523_, _33522_, _33520_);
  and (_33524_, _33455_, _06234_);
  or (_33525_, _33524_, _06195_);
  or (_33526_, _33525_, _33523_);
  and (_33527_, _15315_, _07999_);
  or (_33529_, _33424_, _06196_);
  or (_33530_, _33529_, _33527_);
  and (_33531_, _33530_, _01375_);
  and (_33532_, _33531_, _33526_);
  or (_33533_, _33532_, _33423_);
  and (_43029_, _33533_, _42545_);
  and (_33534_, _01379_, \uc8051golden_1.IP [5]);
  and (_33535_, _13453_, \uc8051golden_1.IP [5]);
  nor (_33536_, _13453_, _08207_);
  or (_33537_, _33536_, _33535_);
  or (_33539_, _33537_, _06293_);
  and (_33540_, _15348_, _07999_);
  or (_33541_, _33540_, _33535_);
  or (_33542_, _33541_, _07210_);
  and (_33543_, _07999_, \uc8051golden_1.ACC [5]);
  or (_33544_, _33543_, _33535_);
  and (_33545_, _33544_, _07199_);
  and (_33546_, _07200_, \uc8051golden_1.IP [5]);
  or (_33547_, _33546_, _06401_);
  or (_33548_, _33547_, _33545_);
  and (_33550_, _33548_, _06396_);
  and (_33551_, _33550_, _33542_);
  and (_33552_, _13461_, \uc8051golden_1.IP [5]);
  and (_33553_, _15341_, _08614_);
  or (_33554_, _33553_, _33552_);
  and (_33555_, _33554_, _06395_);
  or (_33556_, _33555_, _06399_);
  or (_33557_, _33556_, _33551_);
  or (_33558_, _33537_, _07221_);
  and (_33559_, _33558_, _33557_);
  or (_33561_, _33559_, _06406_);
  or (_33562_, _33544_, _06414_);
  and (_33563_, _33562_, _06844_);
  and (_33564_, _33563_, _33561_);
  and (_33565_, _15345_, _08614_);
  or (_33566_, _33565_, _33552_);
  and (_33567_, _33566_, _06393_);
  or (_33568_, _33567_, _06387_);
  or (_33569_, _33568_, _33564_);
  or (_33570_, _33552_, _15378_);
  and (_33572_, _33570_, _33554_);
  or (_33573_, _33572_, _07245_);
  and (_33574_, _33573_, _06446_);
  and (_33575_, _33574_, _33569_);
  or (_33576_, _33552_, _15342_);
  and (_33577_, _33576_, _06300_);
  and (_33578_, _33577_, _33554_);
  or (_33579_, _33578_, _10059_);
  or (_33580_, _33579_, _33575_);
  and (_33581_, _33580_, _33539_);
  or (_33583_, _33581_, _06281_);
  and (_33584_, _07999_, _09441_);
  or (_33585_, _33535_, _06282_);
  or (_33586_, _33585_, _33584_);
  and (_33587_, _33586_, _06279_);
  and (_33588_, _33587_, _33583_);
  and (_33589_, _15446_, _07999_);
  or (_33590_, _33589_, _33535_);
  and (_33591_, _33590_, _06015_);
  or (_33592_, _33591_, _06275_);
  or (_33594_, _33592_, _33588_);
  and (_33595_, _08958_, _07999_);
  or (_33596_, _33595_, _33535_);
  or (_33597_, _33596_, _06276_);
  and (_33598_, _33597_, _33594_);
  or (_33599_, _33598_, _06474_);
  and (_33600_, _15338_, _07999_);
  or (_33601_, _33600_, _33535_);
  or (_33602_, _33601_, _07282_);
  and (_33603_, _33602_, _07284_);
  and (_33605_, _33603_, _33599_);
  and (_33606_, _12542_, _07999_);
  or (_33607_, _33606_, _33535_);
  and (_33608_, _33607_, _06582_);
  or (_33609_, _33608_, _33605_);
  and (_33610_, _33609_, _07279_);
  or (_33611_, _33535_, _08256_);
  and (_33612_, _33596_, _06478_);
  and (_33613_, _33612_, _33611_);
  or (_33614_, _33613_, _33610_);
  and (_33616_, _33614_, _07276_);
  and (_33617_, _33544_, _06569_);
  and (_33618_, _33617_, _33611_);
  or (_33619_, _33618_, _06479_);
  or (_33620_, _33619_, _33616_);
  and (_33621_, _15335_, _07999_);
  or (_33622_, _33535_, _09043_);
  or (_33623_, _33622_, _33621_);
  and (_33624_, _33623_, _09048_);
  and (_33625_, _33624_, _33620_);
  nor (_33627_, _11212_, _13453_);
  or (_33628_, _33627_, _33535_);
  and (_33629_, _33628_, _06572_);
  or (_33630_, _33629_, _06606_);
  or (_33631_, _33630_, _33625_);
  or (_33632_, _33541_, _07037_);
  and (_33633_, _33632_, _06807_);
  and (_33634_, _33633_, _33631_);
  and (_33635_, _33566_, _06234_);
  or (_33636_, _33635_, _06195_);
  or (_33638_, _33636_, _33634_);
  and (_33639_, _15509_, _07999_);
  or (_33640_, _33535_, _06196_);
  or (_33641_, _33640_, _33639_);
  and (_33642_, _33641_, _01375_);
  and (_33643_, _33642_, _33638_);
  or (_33644_, _33643_, _33534_);
  and (_43030_, _33644_, _42545_);
  and (_33645_, _01379_, \uc8051golden_1.IP [6]);
  and (_33646_, _13453_, \uc8051golden_1.IP [6]);
  nor (_33648_, _13453_, _08118_);
  or (_33649_, _33648_, _33646_);
  or (_33650_, _33649_, _06293_);
  and (_33651_, _15550_, _07999_);
  or (_33652_, _33651_, _33646_);
  or (_33653_, _33652_, _07210_);
  and (_33654_, _07999_, \uc8051golden_1.ACC [6]);
  or (_33655_, _33654_, _33646_);
  and (_33656_, _33655_, _07199_);
  and (_33657_, _07200_, \uc8051golden_1.IP [6]);
  or (_33659_, _33657_, _06401_);
  or (_33660_, _33659_, _33656_);
  and (_33661_, _33660_, _06396_);
  and (_33662_, _33661_, _33653_);
  and (_33663_, _13461_, \uc8051golden_1.IP [6]);
  and (_33664_, _15535_, _08614_);
  or (_33665_, _33664_, _33663_);
  and (_33666_, _33665_, _06395_);
  or (_33667_, _33666_, _06399_);
  or (_33668_, _33667_, _33662_);
  or (_33670_, _33649_, _07221_);
  and (_33671_, _33670_, _33668_);
  or (_33672_, _33671_, _06406_);
  or (_33673_, _33655_, _06414_);
  and (_33674_, _33673_, _06844_);
  and (_33675_, _33674_, _33672_);
  and (_33676_, _15561_, _08614_);
  or (_33677_, _33676_, _33663_);
  and (_33678_, _33677_, _06393_);
  or (_33679_, _33678_, _06387_);
  or (_33681_, _33679_, _33675_);
  or (_33682_, _33663_, _15568_);
  and (_33683_, _33682_, _33665_);
  or (_33684_, _33683_, _07245_);
  and (_33685_, _33684_, _06446_);
  and (_33686_, _33685_, _33681_);
  and (_33687_, _15585_, _08614_);
  or (_33688_, _33687_, _33663_);
  and (_33689_, _33688_, _06300_);
  or (_33690_, _33689_, _10059_);
  or (_33692_, _33690_, _33686_);
  and (_33693_, _33692_, _33650_);
  or (_33694_, _33693_, _06281_);
  and (_33695_, _07999_, _09440_);
  or (_33696_, _33646_, _06282_);
  or (_33697_, _33696_, _33695_);
  and (_33698_, _33697_, _06279_);
  and (_33699_, _33698_, _33694_);
  and (_33700_, _15639_, _07999_);
  or (_33701_, _33700_, _33646_);
  and (_33703_, _33701_, _06015_);
  or (_33704_, _33703_, _06275_);
  or (_33705_, _33704_, _33699_);
  and (_33706_, _15646_, _07999_);
  or (_33707_, _33706_, _33646_);
  or (_33708_, _33707_, _06276_);
  and (_33709_, _33708_, _33705_);
  or (_33710_, _33709_, _06474_);
  and (_33711_, _15531_, _07999_);
  or (_33712_, _33711_, _33646_);
  or (_33714_, _33712_, _07282_);
  and (_33715_, _33714_, _07284_);
  and (_33716_, _33715_, _33710_);
  and (_33717_, _11210_, _07999_);
  or (_33718_, _33717_, _33646_);
  and (_33719_, _33718_, _06582_);
  or (_33720_, _33719_, _33716_);
  and (_33721_, _33720_, _07279_);
  or (_33722_, _33646_, _08162_);
  and (_33723_, _33707_, _06478_);
  and (_33725_, _33723_, _33722_);
  or (_33726_, _33725_, _33721_);
  and (_33727_, _33726_, _07276_);
  and (_33728_, _33655_, _06569_);
  and (_33729_, _33728_, _33722_);
  or (_33730_, _33729_, _06479_);
  or (_33731_, _33730_, _33727_);
  and (_33732_, _15528_, _07999_);
  or (_33733_, _33646_, _09043_);
  or (_33734_, _33733_, _33732_);
  and (_33736_, _33734_, _09048_);
  and (_33737_, _33736_, _33731_);
  nor (_33738_, _11209_, _13453_);
  or (_33739_, _33738_, _33646_);
  and (_33740_, _33739_, _06572_);
  or (_33741_, _33740_, _06606_);
  or (_33742_, _33741_, _33737_);
  or (_33743_, _33652_, _07037_);
  and (_33744_, _33743_, _06807_);
  and (_33745_, _33744_, _33742_);
  and (_33747_, _33677_, _06234_);
  or (_33748_, _33747_, _06195_);
  or (_33749_, _33748_, _33745_);
  and (_33750_, _15713_, _07999_);
  or (_33751_, _33646_, _06196_);
  or (_33752_, _33751_, _33750_);
  and (_33753_, _33752_, _01375_);
  and (_33754_, _33753_, _33749_);
  or (_33755_, _33754_, _33645_);
  and (_43031_, _33755_, _42545_);
  not (_33757_, \uc8051golden_1.IE [0]);
  nor (_33758_, _01375_, _33757_);
  nand (_33759_, _11225_, _07948_);
  nor (_33760_, _07948_, _33757_);
  nor (_33761_, _33760_, _07276_);
  nand (_33762_, _33761_, _33759_);
  and (_33763_, _07948_, _07473_);
  or (_33764_, _33763_, _33760_);
  or (_33765_, _33764_, _06293_);
  nor (_33766_, _08521_, _13556_);
  or (_33768_, _33766_, _33760_);
  or (_33769_, _33768_, _07210_);
  and (_33770_, _07948_, \uc8051golden_1.ACC [0]);
  or (_33771_, _33770_, _33760_);
  and (_33772_, _33771_, _07199_);
  nor (_33773_, _07199_, _33757_);
  or (_33774_, _33773_, _06401_);
  or (_33775_, _33774_, _33772_);
  and (_33776_, _33775_, _06396_);
  and (_33777_, _33776_, _33769_);
  nor (_33779_, _08603_, _33757_);
  and (_33780_, _14339_, _08603_);
  or (_33781_, _33780_, _33779_);
  and (_33782_, _33781_, _06395_);
  or (_33783_, _33782_, _33777_);
  and (_33784_, _33783_, _07221_);
  and (_33785_, _33764_, _06399_);
  or (_33786_, _33785_, _06406_);
  or (_33787_, _33786_, _33784_);
  or (_33788_, _33771_, _06414_);
  and (_33790_, _33788_, _06844_);
  and (_33791_, _33790_, _33787_);
  and (_33792_, _33760_, _06393_);
  or (_33793_, _33792_, _06387_);
  or (_33794_, _33793_, _33791_);
  or (_33795_, _33768_, _07245_);
  and (_33796_, _33795_, _06446_);
  and (_33797_, _33796_, _33794_);
  and (_33798_, _14371_, _08603_);
  or (_33799_, _33798_, _33779_);
  and (_33801_, _33799_, _06300_);
  or (_33802_, _33801_, _10059_);
  or (_33803_, _33802_, _33797_);
  and (_33804_, _33803_, _33765_);
  or (_33805_, _33804_, _06281_);
  and (_33806_, _07948_, _09446_);
  or (_33807_, _33760_, _06282_);
  or (_33808_, _33807_, _33806_);
  and (_33809_, _33808_, _33805_);
  or (_33810_, _33809_, _06015_);
  and (_33812_, _14426_, _07948_);
  or (_33813_, _33760_, _06279_);
  or (_33814_, _33813_, _33812_);
  and (_33815_, _33814_, _06276_);
  and (_33816_, _33815_, _33810_);
  and (_33817_, _07948_, _08817_);
  or (_33818_, _33817_, _33760_);
  and (_33819_, _33818_, _06275_);
  or (_33820_, _33819_, _06474_);
  or (_33821_, _33820_, _33816_);
  and (_33823_, _14324_, _07948_);
  or (_33824_, _33823_, _33760_);
  or (_33825_, _33824_, _07282_);
  and (_33826_, _33825_, _07284_);
  and (_33827_, _33826_, _33821_);
  nor (_33828_, _12538_, _13556_);
  or (_33829_, _33828_, _33760_);
  and (_33830_, _33759_, _06582_);
  and (_33831_, _33830_, _33829_);
  or (_33832_, _33831_, _33827_);
  and (_33833_, _33832_, _07279_);
  nand (_33834_, _33818_, _06478_);
  nor (_33835_, _33834_, _33766_);
  or (_33836_, _33835_, _06569_);
  or (_33837_, _33836_, _33833_);
  and (_33838_, _33837_, _33762_);
  or (_33839_, _33838_, _06479_);
  and (_33840_, _14320_, _07948_);
  or (_33841_, _33760_, _09043_);
  or (_33842_, _33841_, _33840_);
  and (_33844_, _33842_, _09048_);
  and (_33845_, _33844_, _33839_);
  and (_33846_, _33829_, _06572_);
  or (_33847_, _33846_, _06606_);
  or (_33848_, _33847_, _33845_);
  or (_33849_, _33768_, _07037_);
  and (_33850_, _33849_, _33848_);
  or (_33851_, _33850_, _06234_);
  or (_33852_, _33760_, _06807_);
  and (_33853_, _33852_, _33851_);
  or (_33855_, _33853_, _06195_);
  or (_33856_, _33768_, _06196_);
  and (_33857_, _33856_, _01375_);
  and (_33858_, _33857_, _33855_);
  or (_33859_, _33858_, _33758_);
  and (_43032_, _33859_, _42545_);
  not (_33860_, \uc8051golden_1.IE [1]);
  nor (_33861_, _01375_, _33860_);
  nor (_33862_, _07948_, _33860_);
  nor (_33863_, _11223_, _13556_);
  or (_33865_, _33863_, _33862_);
  or (_33866_, _33865_, _09048_);
  nand (_33867_, _07948_, _07090_);
  or (_33868_, _07948_, \uc8051golden_1.IE [1]);
  and (_33869_, _33868_, _06275_);
  and (_33870_, _33869_, _33867_);
  nor (_33871_, _13556_, _07196_);
  or (_33872_, _33871_, _33862_);
  and (_33873_, _33872_, _06399_);
  nor (_33874_, _08603_, _33860_);
  and (_33876_, _14514_, _08603_);
  or (_33877_, _33876_, _33874_);
  or (_33878_, _33877_, _06396_);
  and (_33879_, _14532_, _07948_);
  not (_33880_, _33879_);
  and (_33881_, _33880_, _33868_);
  and (_33882_, _33881_, _06401_);
  nor (_33883_, _07199_, _33860_);
  and (_33884_, _07948_, \uc8051golden_1.ACC [1]);
  or (_33885_, _33884_, _33862_);
  and (_33887_, _33885_, _07199_);
  or (_33888_, _33887_, _33883_);
  and (_33889_, _33888_, _07210_);
  or (_33890_, _33889_, _06395_);
  or (_33891_, _33890_, _33882_);
  and (_33892_, _33891_, _33878_);
  and (_33893_, _33892_, _07221_);
  or (_33894_, _33893_, _33873_);
  or (_33895_, _33894_, _06406_);
  or (_33896_, _33885_, _06414_);
  and (_33898_, _33896_, _06844_);
  and (_33899_, _33898_, _33895_);
  and (_33900_, _14517_, _08603_);
  or (_33901_, _33900_, _33874_);
  and (_33902_, _33901_, _06393_);
  or (_33903_, _33902_, _06387_);
  or (_33904_, _33903_, _33899_);
  or (_33905_, _33874_, _14513_);
  and (_33906_, _33905_, _33877_);
  or (_33907_, _33906_, _07245_);
  and (_33909_, _33907_, _06446_);
  and (_33910_, _33909_, _33904_);
  or (_33911_, _33874_, _14560_);
  and (_33912_, _33911_, _06300_);
  and (_33913_, _33912_, _33877_);
  or (_33914_, _33913_, _10059_);
  or (_33915_, _33914_, _33910_);
  or (_33916_, _33872_, _06293_);
  and (_33917_, _33916_, _33915_);
  or (_33918_, _33917_, _06281_);
  and (_33920_, _07948_, _09445_);
  or (_33921_, _33862_, _06282_);
  or (_33922_, _33921_, _33920_);
  and (_33923_, _33922_, _06279_);
  and (_33924_, _33923_, _33918_);
  and (_33925_, _14615_, _07948_);
  or (_33926_, _33925_, _33862_);
  and (_33927_, _33926_, _06015_);
  or (_33928_, _33927_, _33924_);
  and (_33929_, _33928_, _06276_);
  or (_33931_, _33929_, _33870_);
  and (_33932_, _33931_, _07282_);
  or (_33933_, _14507_, _13556_);
  and (_33934_, _33868_, _06474_);
  and (_33935_, _33934_, _33933_);
  or (_33936_, _33935_, _06582_);
  or (_33937_, _33936_, _33932_);
  nand (_33938_, _11222_, _07948_);
  and (_33939_, _33938_, _33865_);
  or (_33940_, _33939_, _07284_);
  and (_33942_, _33940_, _07279_);
  and (_33943_, _33942_, _33937_);
  or (_33944_, _14505_, _13556_);
  and (_33945_, _33868_, _06478_);
  and (_33946_, _33945_, _33944_);
  or (_33947_, _33946_, _06569_);
  or (_33948_, _33947_, _33943_);
  nor (_33949_, _33862_, _07276_);
  nand (_33950_, _33949_, _33938_);
  and (_33951_, _33950_, _09043_);
  and (_33953_, _33951_, _33948_);
  or (_33954_, _33867_, _08477_);
  and (_33955_, _33868_, _06479_);
  and (_33956_, _33955_, _33954_);
  or (_33957_, _33956_, _06572_);
  or (_33958_, _33957_, _33953_);
  and (_33959_, _33958_, _33866_);
  or (_33960_, _33959_, _06606_);
  or (_33961_, _33881_, _07037_);
  and (_33962_, _33961_, _06807_);
  and (_33964_, _33962_, _33960_);
  and (_33965_, _33901_, _06234_);
  or (_33966_, _33965_, _06195_);
  or (_33967_, _33966_, _33964_);
  or (_33968_, _33862_, _06196_);
  or (_33969_, _33968_, _33879_);
  and (_33970_, _33969_, _01375_);
  and (_33971_, _33970_, _33967_);
  or (_33972_, _33971_, _33861_);
  and (_43034_, _33972_, _42545_);
  and (_33974_, _01379_, \uc8051golden_1.IE [2]);
  and (_33975_, _13556_, \uc8051golden_1.IE [2]);
  nor (_33976_, _13556_, _07623_);
  or (_33977_, _33976_, _33975_);
  or (_33978_, _33977_, _06293_);
  or (_33979_, _33977_, _07221_);
  and (_33980_, _14754_, _07948_);
  or (_33981_, _33980_, _33975_);
  or (_33982_, _33981_, _07210_);
  and (_33983_, _07948_, \uc8051golden_1.ACC [2]);
  or (_33985_, _33983_, _33975_);
  and (_33986_, _33985_, _07199_);
  and (_33987_, _07200_, \uc8051golden_1.IE [2]);
  or (_33988_, _33987_, _06401_);
  or (_33989_, _33988_, _33986_);
  and (_33990_, _33989_, _06396_);
  and (_33991_, _33990_, _33982_);
  and (_33992_, _13564_, \uc8051golden_1.IE [2]);
  and (_33993_, _14751_, _08603_);
  or (_33994_, _33993_, _33992_);
  and (_33996_, _33994_, _06395_);
  or (_33997_, _33996_, _06399_);
  or (_33998_, _33997_, _33991_);
  and (_33999_, _33998_, _33979_);
  or (_34000_, _33999_, _06406_);
  or (_34001_, _33985_, _06414_);
  and (_34002_, _34001_, _06844_);
  and (_34003_, _34002_, _34000_);
  and (_34004_, _14749_, _08603_);
  or (_34005_, _34004_, _33992_);
  and (_34007_, _34005_, _06393_);
  or (_34008_, _34007_, _06387_);
  or (_34009_, _34008_, _34003_);
  and (_34010_, _33993_, _14778_);
  or (_34011_, _33992_, _07245_);
  or (_34012_, _34011_, _34010_);
  and (_34013_, _34012_, _06446_);
  and (_34014_, _34013_, _34009_);
  and (_34015_, _14793_, _08603_);
  or (_34016_, _34015_, _33992_);
  and (_34018_, _34016_, _06300_);
  or (_34019_, _34018_, _10059_);
  or (_34020_, _34019_, _34014_);
  and (_34021_, _34020_, _33978_);
  or (_34022_, _34021_, _06281_);
  and (_34023_, _07948_, _09444_);
  or (_34024_, _33975_, _06282_);
  or (_34025_, _34024_, _34023_);
  and (_34026_, _34025_, _06279_);
  and (_34027_, _34026_, _34022_);
  and (_34029_, _14848_, _07948_);
  or (_34030_, _34029_, _33975_);
  and (_34031_, _34030_, _06015_);
  or (_34032_, _34031_, _06275_);
  or (_34033_, _34032_, _34027_);
  and (_34034_, _07948_, _08994_);
  or (_34035_, _34034_, _33975_);
  or (_34036_, _34035_, _06276_);
  and (_34037_, _34036_, _34033_);
  or (_34038_, _34037_, _06474_);
  and (_34040_, _14744_, _07948_);
  or (_34041_, _34040_, _33975_);
  or (_34042_, _34041_, _07282_);
  and (_34043_, _34042_, _07284_);
  and (_34044_, _34043_, _34038_);
  and (_34045_, _11221_, _07948_);
  or (_34046_, _34045_, _33975_);
  and (_34047_, _34046_, _06582_);
  or (_34048_, _34047_, _34044_);
  and (_34049_, _34048_, _07279_);
  or (_34051_, _33975_, _08433_);
  and (_34052_, _34035_, _06478_);
  and (_34053_, _34052_, _34051_);
  or (_34054_, _34053_, _34049_);
  and (_34055_, _34054_, _07276_);
  and (_34056_, _33985_, _06569_);
  and (_34057_, _34056_, _34051_);
  or (_34058_, _34057_, _06479_);
  or (_34059_, _34058_, _34055_);
  and (_34060_, _14741_, _07948_);
  or (_34062_, _33975_, _09043_);
  or (_34063_, _34062_, _34060_);
  and (_34064_, _34063_, _09048_);
  and (_34065_, _34064_, _34059_);
  nor (_34066_, _11220_, _13556_);
  or (_34067_, _34066_, _33975_);
  and (_34068_, _34067_, _06572_);
  or (_34069_, _34068_, _06606_);
  or (_34070_, _34069_, _34065_);
  or (_34071_, _33981_, _07037_);
  and (_34073_, _34071_, _06807_);
  and (_34074_, _34073_, _34070_);
  and (_34075_, _34005_, _06234_);
  or (_34076_, _34075_, _06195_);
  or (_34077_, _34076_, _34074_);
  and (_34078_, _14917_, _07948_);
  or (_34079_, _33975_, _06196_);
  or (_34080_, _34079_, _34078_);
  and (_34081_, _34080_, _01375_);
  and (_34082_, _34081_, _34077_);
  or (_34084_, _34082_, _33974_);
  and (_43035_, _34084_, _42545_);
  and (_34085_, _01379_, \uc8051golden_1.IE [3]);
  and (_34086_, _13556_, \uc8051golden_1.IE [3]);
  nor (_34087_, _13556_, _07775_);
  or (_34088_, _34087_, _34086_);
  or (_34089_, _34088_, _06293_);
  and (_34090_, _14947_, _07948_);
  or (_34091_, _34090_, _34086_);
  or (_34092_, _34091_, _07210_);
  and (_34094_, _07948_, \uc8051golden_1.ACC [3]);
  or (_34095_, _34094_, _34086_);
  and (_34096_, _34095_, _07199_);
  and (_34097_, _07200_, \uc8051golden_1.IE [3]);
  or (_34098_, _34097_, _06401_);
  or (_34099_, _34098_, _34096_);
  and (_34100_, _34099_, _06396_);
  and (_34101_, _34100_, _34092_);
  and (_34102_, _13564_, \uc8051golden_1.IE [3]);
  and (_34103_, _14951_, _08603_);
  or (_34105_, _34103_, _34102_);
  and (_34106_, _34105_, _06395_);
  or (_34107_, _34106_, _06399_);
  or (_34108_, _34107_, _34101_);
  or (_34109_, _34088_, _07221_);
  and (_34110_, _34109_, _34108_);
  or (_34111_, _34110_, _06406_);
  or (_34112_, _34095_, _06414_);
  and (_34113_, _34112_, _06844_);
  and (_34114_, _34113_, _34111_);
  and (_34116_, _14961_, _08603_);
  or (_34117_, _34116_, _34102_);
  and (_34118_, _34117_, _06393_);
  or (_34119_, _34118_, _06387_);
  or (_34120_, _34119_, _34114_);
  or (_34121_, _34102_, _14968_);
  and (_34122_, _34121_, _34105_);
  or (_34123_, _34122_, _07245_);
  and (_34124_, _34123_, _06446_);
  and (_34125_, _34124_, _34120_);
  and (_34127_, _14985_, _08603_);
  or (_34128_, _34127_, _34102_);
  and (_34129_, _34128_, _06300_);
  or (_34130_, _34129_, _10059_);
  or (_34131_, _34130_, _34125_);
  and (_34132_, _34131_, _34089_);
  or (_34133_, _34132_, _06281_);
  and (_34134_, _07948_, _09443_);
  or (_34135_, _34086_, _06282_);
  or (_34136_, _34135_, _34134_);
  and (_34138_, _34136_, _06279_);
  and (_34139_, _34138_, _34133_);
  and (_34140_, _15039_, _07948_);
  or (_34141_, _34140_, _34086_);
  and (_34142_, _34141_, _06015_);
  or (_34143_, _34142_, _06275_);
  or (_34144_, _34143_, _34139_);
  and (_34145_, _07948_, _08815_);
  or (_34146_, _34145_, _34086_);
  or (_34147_, _34146_, _06276_);
  and (_34149_, _34147_, _34144_);
  or (_34150_, _34149_, _06474_);
  and (_34151_, _14934_, _07948_);
  or (_34152_, _34151_, _34086_);
  or (_34153_, _34152_, _07282_);
  and (_34154_, _34153_, _07284_);
  and (_34155_, _34154_, _34150_);
  and (_34156_, _12535_, _07948_);
  or (_34157_, _34156_, _34086_);
  and (_34158_, _34157_, _06582_);
  or (_34160_, _34158_, _34155_);
  and (_34161_, _34160_, _07279_);
  or (_34162_, _34086_, _08389_);
  and (_34163_, _34146_, _06478_);
  and (_34164_, _34163_, _34162_);
  or (_34165_, _34164_, _34161_);
  and (_34166_, _34165_, _07276_);
  and (_34167_, _34095_, _06569_);
  and (_34168_, _34167_, _34162_);
  or (_34169_, _34168_, _06479_);
  or (_34171_, _34169_, _34166_);
  and (_34172_, _14931_, _07948_);
  or (_34173_, _34086_, _09043_);
  or (_34174_, _34173_, _34172_);
  and (_34175_, _34174_, _09048_);
  and (_34176_, _34175_, _34171_);
  nor (_34177_, _11218_, _13556_);
  or (_34178_, _34177_, _34086_);
  and (_34179_, _34178_, _06572_);
  or (_34180_, _34179_, _06606_);
  or (_34182_, _34180_, _34176_);
  or (_34183_, _34091_, _07037_);
  and (_34184_, _34183_, _06807_);
  and (_34185_, _34184_, _34182_);
  and (_34186_, _34117_, _06234_);
  or (_34187_, _34186_, _06195_);
  or (_34188_, _34187_, _34185_);
  and (_34189_, _15113_, _07948_);
  or (_34190_, _34086_, _06196_);
  or (_34191_, _34190_, _34189_);
  and (_34193_, _34191_, _01375_);
  and (_34194_, _34193_, _34188_);
  or (_34195_, _34194_, _34085_);
  and (_43036_, _34195_, _42545_);
  and (_34196_, _01379_, \uc8051golden_1.IE [4]);
  and (_34197_, _13556_, \uc8051golden_1.IE [4]);
  nor (_34198_, _13556_, _08301_);
  or (_34199_, _34198_, _34197_);
  or (_34200_, _34199_, _06293_);
  and (_34201_, _15130_, _07948_);
  or (_34203_, _34201_, _34197_);
  or (_34204_, _34203_, _07210_);
  and (_34205_, _07948_, \uc8051golden_1.ACC [4]);
  or (_34206_, _34205_, _34197_);
  and (_34207_, _34206_, _07199_);
  and (_34208_, _07200_, \uc8051golden_1.IE [4]);
  or (_34209_, _34208_, _06401_);
  or (_34210_, _34209_, _34207_);
  and (_34211_, _34210_, _06396_);
  and (_34212_, _34211_, _34204_);
  and (_34214_, _13564_, \uc8051golden_1.IE [4]);
  and (_34215_, _15139_, _08603_);
  or (_34216_, _34215_, _34214_);
  and (_34217_, _34216_, _06395_);
  or (_34218_, _34217_, _06399_);
  or (_34219_, _34218_, _34212_);
  or (_34220_, _34199_, _07221_);
  and (_34221_, _34220_, _34219_);
  or (_34222_, _34221_, _06406_);
  or (_34223_, _34206_, _06414_);
  and (_34225_, _34223_, _06844_);
  and (_34226_, _34225_, _34222_);
  and (_34227_, _15168_, _08603_);
  or (_34228_, _34227_, _34214_);
  and (_34229_, _34228_, _06393_);
  or (_34230_, _34229_, _06387_);
  or (_34231_, _34230_, _34226_);
  or (_34232_, _34214_, _15138_);
  and (_34233_, _34232_, _34216_);
  or (_34234_, _34233_, _07245_);
  and (_34236_, _34234_, _06446_);
  and (_34237_, _34236_, _34231_);
  and (_34238_, _15189_, _08603_);
  or (_34239_, _34238_, _34214_);
  and (_34240_, _34239_, _06300_);
  or (_34241_, _34240_, _10059_);
  or (_34242_, _34241_, _34237_);
  and (_34243_, _34242_, _34200_);
  or (_34244_, _34243_, _06281_);
  and (_34245_, _07948_, _09442_);
  or (_34247_, _34197_, _06282_);
  or (_34248_, _34247_, _34245_);
  and (_34249_, _34248_, _06279_);
  and (_34250_, _34249_, _34244_);
  and (_34251_, _15243_, _07948_);
  or (_34252_, _34251_, _34197_);
  and (_34253_, _34252_, _06015_);
  or (_34254_, _34253_, _06275_);
  or (_34255_, _34254_, _34250_);
  and (_34256_, _08883_, _07948_);
  or (_34258_, _34256_, _34197_);
  or (_34259_, _34258_, _06276_);
  and (_34260_, _34259_, _34255_);
  or (_34261_, _34260_, _06474_);
  and (_34262_, _15135_, _07948_);
  or (_34263_, _34262_, _34197_);
  or (_34264_, _34263_, _07282_);
  and (_34265_, _34264_, _07284_);
  and (_34266_, _34265_, _34261_);
  and (_34267_, _11216_, _07948_);
  or (_34269_, _34267_, _34197_);
  and (_34270_, _34269_, _06582_);
  or (_34271_, _34270_, _34266_);
  and (_34272_, _34271_, _07279_);
  or (_34273_, _34197_, _08345_);
  and (_34274_, _34258_, _06478_);
  and (_34275_, _34274_, _34273_);
  or (_34276_, _34275_, _34272_);
  and (_34277_, _34276_, _07276_);
  and (_34278_, _34206_, _06569_);
  and (_34280_, _34278_, _34273_);
  or (_34281_, _34280_, _06479_);
  or (_34282_, _34281_, _34277_);
  and (_34283_, _15134_, _07948_);
  or (_34284_, _34197_, _09043_);
  or (_34285_, _34284_, _34283_);
  and (_34286_, _34285_, _09048_);
  and (_34287_, _34286_, _34282_);
  nor (_34288_, _11215_, _13556_);
  or (_34289_, _34288_, _34197_);
  and (_34291_, _34289_, _06572_);
  or (_34292_, _34291_, _06606_);
  or (_34293_, _34292_, _34287_);
  or (_34294_, _34203_, _07037_);
  and (_34295_, _34294_, _06807_);
  and (_34296_, _34295_, _34293_);
  and (_34297_, _34228_, _06234_);
  or (_34298_, _34297_, _06195_);
  or (_34299_, _34298_, _34296_);
  and (_34300_, _15315_, _07948_);
  or (_34302_, _34197_, _06196_);
  or (_34303_, _34302_, _34300_);
  and (_34304_, _34303_, _01375_);
  and (_34305_, _34304_, _34299_);
  or (_34306_, _34305_, _34196_);
  and (_43037_, _34306_, _42545_);
  and (_34307_, _01379_, \uc8051golden_1.IE [5]);
  and (_34308_, _13556_, \uc8051golden_1.IE [5]);
  nor (_34309_, _13556_, _08207_);
  or (_34310_, _34309_, _34308_);
  or (_34312_, _34310_, _06293_);
  and (_34313_, _15348_, _07948_);
  or (_34314_, _34313_, _34308_);
  or (_34315_, _34314_, _07210_);
  and (_34316_, _07948_, \uc8051golden_1.ACC [5]);
  or (_34317_, _34316_, _34308_);
  and (_34318_, _34317_, _07199_);
  and (_34319_, _07200_, \uc8051golden_1.IE [5]);
  or (_34320_, _34319_, _06401_);
  or (_34321_, _34320_, _34318_);
  and (_34323_, _34321_, _06396_);
  and (_34324_, _34323_, _34315_);
  and (_34325_, _13564_, \uc8051golden_1.IE [5]);
  and (_34326_, _15341_, _08603_);
  or (_34327_, _34326_, _34325_);
  and (_34328_, _34327_, _06395_);
  or (_34329_, _34328_, _06399_);
  or (_34330_, _34329_, _34324_);
  or (_34331_, _34310_, _07221_);
  and (_34332_, _34331_, _34330_);
  or (_34334_, _34332_, _06406_);
  or (_34335_, _34317_, _06414_);
  and (_34336_, _34335_, _06844_);
  and (_34337_, _34336_, _34334_);
  and (_34338_, _15345_, _08603_);
  or (_34339_, _34338_, _34325_);
  and (_34340_, _34339_, _06393_);
  or (_34341_, _34340_, _06387_);
  or (_34342_, _34341_, _34337_);
  or (_34343_, _34325_, _15378_);
  and (_34345_, _34343_, _34327_);
  or (_34346_, _34345_, _07245_);
  and (_34347_, _34346_, _06446_);
  and (_34348_, _34347_, _34342_);
  or (_34349_, _34325_, _15342_);
  and (_34350_, _34349_, _06300_);
  and (_34351_, _34350_, _34327_);
  or (_34352_, _34351_, _10059_);
  or (_34353_, _34352_, _34348_);
  and (_34354_, _34353_, _34312_);
  or (_34356_, _34354_, _06281_);
  and (_34357_, _07948_, _09441_);
  or (_34358_, _34308_, _06282_);
  or (_34359_, _34358_, _34357_);
  and (_34360_, _34359_, _06279_);
  and (_34361_, _34360_, _34356_);
  and (_34362_, _15446_, _07948_);
  or (_34363_, _34362_, _34308_);
  and (_34364_, _34363_, _06015_);
  or (_34365_, _34364_, _06275_);
  or (_34367_, _34365_, _34361_);
  and (_34368_, _08958_, _07948_);
  or (_34369_, _34368_, _34308_);
  or (_34370_, _34369_, _06276_);
  and (_34371_, _34370_, _34367_);
  or (_34372_, _34371_, _06474_);
  and (_34373_, _15338_, _07948_);
  or (_34374_, _34373_, _34308_);
  or (_34375_, _34374_, _07282_);
  and (_34376_, _34375_, _07284_);
  and (_34378_, _34376_, _34372_);
  and (_34379_, _12542_, _07948_);
  or (_34380_, _34379_, _34308_);
  and (_34381_, _34380_, _06582_);
  or (_34382_, _34381_, _34378_);
  and (_34383_, _34382_, _07279_);
  or (_34384_, _34308_, _08256_);
  and (_34385_, _34369_, _06478_);
  and (_34386_, _34385_, _34384_);
  or (_34387_, _34386_, _34383_);
  and (_34389_, _34387_, _07276_);
  and (_34390_, _34317_, _06569_);
  and (_34391_, _34390_, _34384_);
  or (_34392_, _34391_, _06479_);
  or (_34393_, _34392_, _34389_);
  and (_34394_, _15335_, _07948_);
  or (_34395_, _34308_, _09043_);
  or (_34396_, _34395_, _34394_);
  and (_34397_, _34396_, _09048_);
  and (_34398_, _34397_, _34393_);
  nor (_34400_, _11212_, _13556_);
  or (_34401_, _34400_, _34308_);
  and (_34402_, _34401_, _06572_);
  or (_34403_, _34402_, _06606_);
  or (_34404_, _34403_, _34398_);
  or (_34405_, _34314_, _07037_);
  and (_34406_, _34405_, _06807_);
  and (_34407_, _34406_, _34404_);
  and (_34408_, _34339_, _06234_);
  or (_34409_, _34408_, _06195_);
  or (_34411_, _34409_, _34407_);
  and (_34412_, _15509_, _07948_);
  or (_34413_, _34308_, _06196_);
  or (_34414_, _34413_, _34412_);
  and (_34415_, _34414_, _01375_);
  and (_34416_, _34415_, _34411_);
  or (_34417_, _34416_, _34307_);
  and (_43038_, _34417_, _42545_);
  and (_34418_, _01379_, \uc8051golden_1.IE [6]);
  and (_34419_, _13556_, \uc8051golden_1.IE [6]);
  nor (_34421_, _13556_, _08118_);
  or (_34422_, _34421_, _34419_);
  or (_34423_, _34422_, _06293_);
  and (_34424_, _15550_, _07948_);
  or (_34425_, _34424_, _34419_);
  or (_34426_, _34425_, _07210_);
  and (_34427_, _07948_, \uc8051golden_1.ACC [6]);
  or (_34428_, _34427_, _34419_);
  and (_34429_, _34428_, _07199_);
  and (_34430_, _07200_, \uc8051golden_1.IE [6]);
  or (_34432_, _34430_, _06401_);
  or (_34433_, _34432_, _34429_);
  and (_34434_, _34433_, _06396_);
  and (_34435_, _34434_, _34426_);
  and (_34436_, _13564_, \uc8051golden_1.IE [6]);
  and (_34437_, _15535_, _08603_);
  or (_34438_, _34437_, _34436_);
  and (_34439_, _34438_, _06395_);
  or (_34440_, _34439_, _06399_);
  or (_34441_, _34440_, _34435_);
  or (_34443_, _34422_, _07221_);
  and (_34444_, _34443_, _34441_);
  or (_34445_, _34444_, _06406_);
  or (_34446_, _34428_, _06414_);
  and (_34447_, _34446_, _06844_);
  and (_34448_, _34447_, _34445_);
  and (_34449_, _15561_, _08603_);
  or (_34450_, _34449_, _34436_);
  and (_34451_, _34450_, _06393_);
  or (_34452_, _34451_, _06387_);
  or (_34454_, _34452_, _34448_);
  or (_34455_, _34436_, _15568_);
  and (_34456_, _34455_, _34438_);
  or (_34457_, _34456_, _07245_);
  and (_34458_, _34457_, _06446_);
  and (_34459_, _34458_, _34454_);
  and (_34460_, _15585_, _08603_);
  or (_34461_, _34460_, _34436_);
  and (_34462_, _34461_, _06300_);
  or (_34463_, _34462_, _10059_);
  or (_34465_, _34463_, _34459_);
  and (_34466_, _34465_, _34423_);
  or (_34467_, _34466_, _06281_);
  and (_34468_, _07948_, _09440_);
  or (_34469_, _34419_, _06282_);
  or (_34470_, _34469_, _34468_);
  and (_34471_, _34470_, _06279_);
  and (_34472_, _34471_, _34467_);
  and (_34473_, _15639_, _07948_);
  or (_34474_, _34473_, _34419_);
  and (_34476_, _34474_, _06015_);
  or (_34477_, _34476_, _06275_);
  or (_34478_, _34477_, _34472_);
  and (_34479_, _15646_, _07948_);
  or (_34480_, _34479_, _34419_);
  or (_34481_, _34480_, _06276_);
  and (_34482_, _34481_, _34478_);
  or (_34483_, _34482_, _06474_);
  and (_34484_, _15531_, _07948_);
  or (_34485_, _34484_, _34419_);
  or (_34487_, _34485_, _07282_);
  and (_34488_, _34487_, _07284_);
  and (_34489_, _34488_, _34483_);
  and (_34490_, _11210_, _07948_);
  or (_34491_, _34490_, _34419_);
  and (_34492_, _34491_, _06582_);
  or (_34493_, _34492_, _34489_);
  and (_34494_, _34493_, _07279_);
  or (_34495_, _34419_, _08162_);
  and (_34496_, _34480_, _06478_);
  and (_34498_, _34496_, _34495_);
  or (_34499_, _34498_, _34494_);
  and (_34500_, _34499_, _07276_);
  and (_34501_, _34428_, _06569_);
  and (_34502_, _34501_, _34495_);
  or (_34503_, _34502_, _06479_);
  or (_34504_, _34503_, _34500_);
  and (_34505_, _15528_, _07948_);
  or (_34506_, _34419_, _09043_);
  or (_34507_, _34506_, _34505_);
  and (_34509_, _34507_, _09048_);
  and (_34510_, _34509_, _34504_);
  nor (_34511_, _11209_, _13556_);
  or (_34512_, _34511_, _34419_);
  and (_34513_, _34512_, _06572_);
  or (_34514_, _34513_, _06606_);
  or (_34515_, _34514_, _34510_);
  or (_34516_, _34425_, _07037_);
  and (_34517_, _34516_, _06807_);
  and (_34518_, _34517_, _34515_);
  and (_34520_, _34450_, _06234_);
  or (_34521_, _34520_, _06195_);
  or (_34522_, _34521_, _34518_);
  and (_34523_, _15713_, _07948_);
  or (_34524_, _34419_, _06196_);
  or (_34525_, _34524_, _34523_);
  and (_34526_, _34525_, _01375_);
  and (_34527_, _34526_, _34522_);
  or (_34528_, _34527_, _34418_);
  and (_43039_, _34528_, _42545_);
  not (_34530_, \uc8051golden_1.SCON [0]);
  nor (_34531_, _01375_, _34530_);
  nand (_34532_, _11225_, _07972_);
  nor (_34533_, _07972_, _34530_);
  nor (_34534_, _34533_, _07276_);
  nand (_34535_, _34534_, _34532_);
  and (_34536_, _07972_, _07473_);
  or (_34537_, _34536_, _34533_);
  or (_34538_, _34537_, _06293_);
  nor (_34539_, _08521_, _13664_);
  or (_34541_, _34539_, _34533_);
  or (_34542_, _34541_, _07210_);
  and (_34543_, _07972_, \uc8051golden_1.ACC [0]);
  or (_34544_, _34543_, _34533_);
  and (_34545_, _34544_, _07199_);
  nor (_34546_, _07199_, _34530_);
  or (_34547_, _34546_, _06401_);
  or (_34548_, _34547_, _34545_);
  and (_34549_, _34548_, _06396_);
  and (_34550_, _34549_, _34542_);
  nor (_34551_, _08606_, _34530_);
  and (_34552_, _14339_, _08606_);
  or (_34553_, _34552_, _34551_);
  and (_34554_, _34553_, _06395_);
  or (_34555_, _34554_, _34550_);
  and (_34556_, _34555_, _07221_);
  and (_34557_, _34537_, _06399_);
  or (_34558_, _34557_, _06406_);
  or (_34559_, _34558_, _34556_);
  or (_34560_, _34544_, _06414_);
  and (_34562_, _34560_, _06844_);
  and (_34563_, _34562_, _34559_);
  and (_34564_, _34533_, _06393_);
  or (_34565_, _34564_, _06387_);
  or (_34566_, _34565_, _34563_);
  or (_34567_, _34541_, _07245_);
  and (_34568_, _34567_, _06446_);
  and (_34569_, _34568_, _34566_);
  and (_34570_, _14371_, _08606_);
  or (_34571_, _34570_, _34551_);
  and (_34573_, _34571_, _06300_);
  or (_34574_, _34573_, _10059_);
  or (_34575_, _34574_, _34569_);
  and (_34576_, _34575_, _34538_);
  or (_34577_, _34576_, _06281_);
  and (_34578_, _07972_, _09446_);
  or (_34579_, _34533_, _06282_);
  or (_34580_, _34579_, _34578_);
  and (_34581_, _34580_, _34577_);
  or (_34582_, _34581_, _06015_);
  and (_34584_, _14426_, _07972_);
  or (_34585_, _34533_, _06279_);
  or (_34586_, _34585_, _34584_);
  and (_34587_, _34586_, _06276_);
  and (_34588_, _34587_, _34582_);
  and (_34589_, _07972_, _08817_);
  or (_34590_, _34589_, _34533_);
  and (_34591_, _34590_, _06275_);
  or (_34592_, _34591_, _06474_);
  or (_34593_, _34592_, _34588_);
  and (_34595_, _14324_, _07972_);
  or (_34596_, _34595_, _34533_);
  or (_34597_, _34596_, _07282_);
  and (_34598_, _34597_, _07284_);
  and (_34599_, _34598_, _34593_);
  nor (_34600_, _12538_, _13664_);
  or (_34601_, _34600_, _34533_);
  and (_34602_, _34532_, _06582_);
  and (_34603_, _34602_, _34601_);
  or (_34604_, _34603_, _34599_);
  and (_34606_, _34604_, _07279_);
  nand (_34607_, _34590_, _06478_);
  nor (_34608_, _34607_, _34539_);
  or (_34609_, _34608_, _06569_);
  or (_34610_, _34609_, _34606_);
  and (_34611_, _34610_, _34535_);
  or (_34612_, _34611_, _06479_);
  and (_34613_, _14320_, _07972_);
  or (_34614_, _34613_, _34533_);
  or (_34615_, _34614_, _09043_);
  and (_34617_, _34615_, _09048_);
  and (_34618_, _34617_, _34612_);
  and (_34619_, _34601_, _06572_);
  or (_34620_, _34619_, _06606_);
  or (_34621_, _34620_, _34618_);
  or (_34622_, _34541_, _07037_);
  and (_34623_, _34622_, _34621_);
  or (_34624_, _34623_, _06234_);
  or (_34625_, _34533_, _06807_);
  and (_34626_, _34625_, _34624_);
  or (_34628_, _34626_, _06195_);
  or (_34629_, _34541_, _06196_);
  and (_34630_, _34629_, _01375_);
  and (_34631_, _34630_, _34628_);
  or (_34632_, _34631_, _34531_);
  and (_43041_, _34632_, _42545_);
  not (_34633_, \uc8051golden_1.SCON [1]);
  nor (_34634_, _01375_, _34633_);
  nor (_34635_, _07972_, _34633_);
  nor (_34636_, _11223_, _13664_);
  or (_34638_, _34636_, _34635_);
  or (_34639_, _34638_, _09048_);
  nand (_34640_, _07972_, _07090_);
  or (_34641_, _07972_, \uc8051golden_1.SCON [1]);
  and (_34642_, _34641_, _06275_);
  and (_34643_, _34642_, _34640_);
  nor (_34644_, _13664_, _07196_);
  or (_34645_, _34644_, _34635_);
  or (_34646_, _34645_, _07221_);
  and (_34647_, _14532_, _07972_);
  not (_34649_, _34647_);
  and (_34650_, _34649_, _34641_);
  or (_34651_, _34650_, _07210_);
  and (_34652_, _07972_, \uc8051golden_1.ACC [1]);
  or (_34653_, _34652_, _34635_);
  and (_34654_, _34653_, _07199_);
  nor (_34655_, _07199_, _34633_);
  or (_34656_, _34655_, _06401_);
  or (_34657_, _34656_, _34654_);
  and (_34658_, _34657_, _06396_);
  and (_34660_, _34658_, _34651_);
  nor (_34661_, _08606_, _34633_);
  and (_34662_, _14514_, _08606_);
  or (_34663_, _34662_, _34661_);
  and (_34664_, _34663_, _06395_);
  or (_34665_, _34664_, _06399_);
  or (_34666_, _34665_, _34660_);
  and (_34667_, _34666_, _34646_);
  or (_34668_, _34667_, _06406_);
  or (_34669_, _34653_, _06414_);
  and (_34671_, _34669_, _06844_);
  and (_34672_, _34671_, _34668_);
  and (_34673_, _14517_, _08606_);
  or (_34674_, _34673_, _34661_);
  and (_34675_, _34674_, _06393_);
  or (_34676_, _34675_, _06387_);
  or (_34677_, _34676_, _34672_);
  and (_34678_, _34662_, _14513_);
  or (_34679_, _34661_, _07245_);
  or (_34680_, _34679_, _34678_);
  and (_34682_, _34680_, _06446_);
  and (_34683_, _34682_, _34677_);
  or (_34684_, _34661_, _14560_);
  and (_34685_, _34684_, _06300_);
  and (_34686_, _34685_, _34663_);
  or (_34687_, _34686_, _10059_);
  or (_34688_, _34687_, _34683_);
  or (_34689_, _34645_, _06293_);
  and (_34690_, _34689_, _34688_);
  or (_34691_, _34690_, _06281_);
  and (_34693_, _07972_, _09445_);
  or (_34694_, _34635_, _06282_);
  or (_34695_, _34694_, _34693_);
  and (_34696_, _34695_, _06279_);
  and (_34697_, _34696_, _34691_);
  and (_34698_, _14615_, _07972_);
  or (_34699_, _34698_, _34635_);
  and (_34700_, _34699_, _06015_);
  or (_34701_, _34700_, _34697_);
  and (_34702_, _34701_, _06276_);
  or (_34704_, _34702_, _34643_);
  and (_34705_, _34704_, _07282_);
  or (_34706_, _14507_, _13664_);
  and (_34707_, _34641_, _06474_);
  and (_34708_, _34707_, _34706_);
  or (_34709_, _34708_, _06582_);
  or (_34710_, _34709_, _34705_);
  nand (_34711_, _11222_, _07972_);
  and (_34712_, _34711_, _34638_);
  or (_34713_, _34712_, _07284_);
  and (_34715_, _34713_, _07279_);
  and (_34716_, _34715_, _34710_);
  or (_34717_, _14505_, _13664_);
  and (_34718_, _34641_, _06478_);
  and (_34719_, _34718_, _34717_);
  or (_34720_, _34719_, _06569_);
  or (_34721_, _34720_, _34716_);
  nor (_34722_, _34635_, _07276_);
  nand (_34723_, _34722_, _34711_);
  and (_34724_, _34723_, _09043_);
  and (_34726_, _34724_, _34721_);
  or (_34727_, _34640_, _08477_);
  and (_34728_, _34641_, _06479_);
  and (_34729_, _34728_, _34727_);
  or (_34730_, _34729_, _06572_);
  or (_34731_, _34730_, _34726_);
  and (_34732_, _34731_, _34639_);
  or (_34733_, _34732_, _06606_);
  or (_34734_, _34650_, _07037_);
  and (_34735_, _34734_, _06807_);
  and (_34737_, _34735_, _34733_);
  and (_34738_, _34674_, _06234_);
  or (_34739_, _34738_, _06195_);
  or (_34740_, _34739_, _34737_);
  or (_34741_, _34635_, _06196_);
  or (_34742_, _34741_, _34647_);
  and (_34743_, _34742_, _01375_);
  and (_34744_, _34743_, _34740_);
  or (_34745_, _34744_, _34634_);
  and (_43042_, _34745_, _42545_);
  and (_34747_, _01379_, \uc8051golden_1.SCON [2]);
  and (_34748_, _13664_, \uc8051golden_1.SCON [2]);
  nor (_34749_, _13664_, _07623_);
  or (_34750_, _34749_, _34748_);
  or (_34751_, _34750_, _06293_);
  or (_34752_, _34750_, _07221_);
  and (_34753_, _14754_, _07972_);
  or (_34754_, _34753_, _34748_);
  or (_34755_, _34754_, _07210_);
  and (_34756_, _07972_, \uc8051golden_1.ACC [2]);
  or (_34758_, _34756_, _34748_);
  and (_34759_, _34758_, _07199_);
  and (_34760_, _07200_, \uc8051golden_1.SCON [2]);
  or (_34761_, _34760_, _06401_);
  or (_34762_, _34761_, _34759_);
  and (_34763_, _34762_, _06396_);
  and (_34764_, _34763_, _34755_);
  and (_34765_, _13673_, \uc8051golden_1.SCON [2]);
  and (_34766_, _14751_, _08606_);
  or (_34767_, _34766_, _34765_);
  and (_34769_, _34767_, _06395_);
  or (_34770_, _34769_, _06399_);
  or (_34771_, _34770_, _34764_);
  and (_34772_, _34771_, _34752_);
  or (_34773_, _34772_, _06406_);
  or (_34774_, _34758_, _06414_);
  and (_34775_, _34774_, _06844_);
  and (_34776_, _34775_, _34773_);
  and (_34777_, _14749_, _08606_);
  or (_34778_, _34777_, _34765_);
  and (_34780_, _34778_, _06393_);
  or (_34781_, _34780_, _06387_);
  or (_34782_, _34781_, _34776_);
  and (_34783_, _34766_, _14778_);
  or (_34784_, _34765_, _07245_);
  or (_34785_, _34784_, _34783_);
  and (_34786_, _34785_, _06446_);
  and (_34787_, _34786_, _34782_);
  and (_34788_, _14793_, _08606_);
  or (_34789_, _34788_, _34765_);
  and (_34791_, _34789_, _06300_);
  or (_34792_, _34791_, _10059_);
  or (_34793_, _34792_, _34787_);
  and (_34794_, _34793_, _34751_);
  or (_34795_, _34794_, _06281_);
  and (_34796_, _07972_, _09444_);
  or (_34797_, _34748_, _06282_);
  or (_34798_, _34797_, _34796_);
  and (_34799_, _34798_, _06279_);
  and (_34800_, _34799_, _34795_);
  and (_34802_, _14848_, _07972_);
  or (_34803_, _34802_, _34748_);
  and (_34804_, _34803_, _06015_);
  or (_34805_, _34804_, _06275_);
  or (_34806_, _34805_, _34800_);
  and (_34807_, _07972_, _08994_);
  or (_34808_, _34807_, _34748_);
  or (_34809_, _34808_, _06276_);
  and (_34810_, _34809_, _34806_);
  or (_34811_, _34810_, _06474_);
  and (_34813_, _14744_, _07972_);
  or (_34814_, _34813_, _34748_);
  or (_34815_, _34814_, _07282_);
  and (_34816_, _34815_, _07284_);
  and (_34817_, _34816_, _34811_);
  and (_34818_, _11221_, _07972_);
  or (_34819_, _34818_, _34748_);
  and (_34820_, _34819_, _06582_);
  or (_34821_, _34820_, _34817_);
  and (_34822_, _34821_, _07279_);
  or (_34824_, _34748_, _08433_);
  and (_34825_, _34808_, _06478_);
  and (_34826_, _34825_, _34824_);
  or (_34827_, _34826_, _34822_);
  and (_34828_, _34827_, _07276_);
  and (_34829_, _34758_, _06569_);
  and (_34830_, _34829_, _34824_);
  or (_34831_, _34830_, _06479_);
  or (_34832_, _34831_, _34828_);
  and (_34833_, _14741_, _07972_);
  or (_34835_, _34748_, _09043_);
  or (_34836_, _34835_, _34833_);
  and (_34837_, _34836_, _09048_);
  and (_34838_, _34837_, _34832_);
  nor (_34839_, _11220_, _13664_);
  or (_34840_, _34839_, _34748_);
  and (_34841_, _34840_, _06572_);
  or (_34842_, _34841_, _06606_);
  or (_34843_, _34842_, _34838_);
  or (_34844_, _34754_, _07037_);
  and (_34846_, _34844_, _06807_);
  and (_34847_, _34846_, _34843_);
  and (_34848_, _34778_, _06234_);
  or (_34849_, _34848_, _06195_);
  or (_34850_, _34849_, _34847_);
  and (_34851_, _14917_, _07972_);
  or (_34852_, _34748_, _06196_);
  or (_34853_, _34852_, _34851_);
  and (_34854_, _34853_, _01375_);
  and (_34855_, _34854_, _34850_);
  or (_34857_, _34855_, _34747_);
  and (_43043_, _34857_, _42545_);
  and (_34858_, _01379_, \uc8051golden_1.SCON [3]);
  and (_34859_, _13664_, \uc8051golden_1.SCON [3]);
  nor (_34860_, _13664_, _07775_);
  or (_34861_, _34860_, _34859_);
  or (_34862_, _34861_, _06293_);
  and (_34863_, _14947_, _07972_);
  or (_34864_, _34863_, _34859_);
  or (_34865_, _34864_, _07210_);
  and (_34867_, _07972_, \uc8051golden_1.ACC [3]);
  or (_34868_, _34867_, _34859_);
  and (_34869_, _34868_, _07199_);
  and (_34870_, _07200_, \uc8051golden_1.SCON [3]);
  or (_34871_, _34870_, _06401_);
  or (_34872_, _34871_, _34869_);
  and (_34873_, _34872_, _06396_);
  and (_34874_, _34873_, _34865_);
  and (_34875_, _13673_, \uc8051golden_1.SCON [3]);
  and (_34876_, _14951_, _08606_);
  or (_34878_, _34876_, _34875_);
  and (_34879_, _34878_, _06395_);
  or (_34880_, _34879_, _06399_);
  or (_34881_, _34880_, _34874_);
  or (_34882_, _34861_, _07221_);
  and (_34883_, _34882_, _34881_);
  or (_34884_, _34883_, _06406_);
  or (_34885_, _34868_, _06414_);
  and (_34886_, _34885_, _06844_);
  and (_34887_, _34886_, _34884_);
  and (_34889_, _14961_, _08606_);
  or (_34890_, _34889_, _34875_);
  and (_34891_, _34890_, _06393_);
  or (_34892_, _34891_, _06387_);
  or (_34893_, _34892_, _34887_);
  or (_34894_, _34875_, _14968_);
  and (_34895_, _34894_, _34878_);
  or (_34896_, _34895_, _07245_);
  and (_34897_, _34896_, _06446_);
  and (_34898_, _34897_, _34893_);
  and (_34900_, _14985_, _08606_);
  or (_34901_, _34900_, _34875_);
  and (_34902_, _34901_, _06300_);
  or (_34903_, _34902_, _10059_);
  or (_34904_, _34903_, _34898_);
  and (_34905_, _34904_, _34862_);
  or (_34906_, _34905_, _06281_);
  and (_34907_, _07972_, _09443_);
  or (_34908_, _34859_, _06282_);
  or (_34909_, _34908_, _34907_);
  and (_34911_, _34909_, _06279_);
  and (_34912_, _34911_, _34906_);
  and (_34913_, _15039_, _07972_);
  or (_34914_, _34913_, _34859_);
  and (_34915_, _34914_, _06015_);
  or (_34916_, _34915_, _06275_);
  or (_34917_, _34916_, _34912_);
  and (_34918_, _07972_, _08815_);
  or (_34919_, _34918_, _34859_);
  or (_34920_, _34919_, _06276_);
  and (_34922_, _34920_, _34917_);
  or (_34923_, _34922_, _06474_);
  and (_34924_, _14934_, _07972_);
  or (_34925_, _34924_, _34859_);
  or (_34926_, _34925_, _07282_);
  and (_34927_, _34926_, _07284_);
  and (_34928_, _34927_, _34923_);
  and (_34929_, _12535_, _07972_);
  or (_34930_, _34929_, _34859_);
  and (_34931_, _34930_, _06582_);
  or (_34933_, _34931_, _34928_);
  and (_34934_, _34933_, _07279_);
  or (_34935_, _34859_, _08389_);
  and (_34936_, _34919_, _06478_);
  and (_34937_, _34936_, _34935_);
  or (_34938_, _34937_, _34934_);
  and (_34939_, _34938_, _07276_);
  and (_34940_, _34868_, _06569_);
  and (_34941_, _34940_, _34935_);
  or (_34942_, _34941_, _06479_);
  or (_34944_, _34942_, _34939_);
  and (_34945_, _14931_, _07972_);
  or (_34946_, _34859_, _09043_);
  or (_34947_, _34946_, _34945_);
  and (_34948_, _34947_, _09048_);
  and (_34949_, _34948_, _34944_);
  nor (_34950_, _11218_, _13664_);
  or (_34951_, _34950_, _34859_);
  and (_34952_, _34951_, _06572_);
  or (_34953_, _34952_, _06606_);
  or (_34955_, _34953_, _34949_);
  or (_34956_, _34864_, _07037_);
  and (_34957_, _34956_, _06807_);
  and (_34958_, _34957_, _34955_);
  and (_34959_, _34890_, _06234_);
  or (_34960_, _34959_, _06195_);
  or (_34961_, _34960_, _34958_);
  and (_34962_, _15113_, _07972_);
  or (_34963_, _34859_, _06196_);
  or (_34964_, _34963_, _34962_);
  and (_34966_, _34964_, _01375_);
  and (_34967_, _34966_, _34961_);
  or (_34968_, _34967_, _34858_);
  and (_43044_, _34968_, _42545_);
  and (_34969_, _01379_, \uc8051golden_1.SCON [4]);
  and (_34970_, _13664_, \uc8051golden_1.SCON [4]);
  nor (_34971_, _13664_, _08301_);
  or (_34972_, _34971_, _34970_);
  or (_34973_, _34972_, _06293_);
  and (_34974_, _15130_, _07972_);
  or (_34976_, _34974_, _34970_);
  or (_34977_, _34976_, _07210_);
  and (_34978_, _07972_, \uc8051golden_1.ACC [4]);
  or (_34979_, _34978_, _34970_);
  and (_34980_, _34979_, _07199_);
  and (_34981_, _07200_, \uc8051golden_1.SCON [4]);
  or (_34982_, _34981_, _06401_);
  or (_34983_, _34982_, _34980_);
  and (_34984_, _34983_, _06396_);
  and (_34985_, _34984_, _34977_);
  and (_34987_, _13673_, \uc8051golden_1.SCON [4]);
  and (_34988_, _15139_, _08606_);
  or (_34989_, _34988_, _34987_);
  and (_34990_, _34989_, _06395_);
  or (_34991_, _34990_, _06399_);
  or (_34992_, _34991_, _34985_);
  or (_34993_, _34972_, _07221_);
  and (_34994_, _34993_, _34992_);
  or (_34995_, _34994_, _06406_);
  or (_34996_, _34979_, _06414_);
  and (_34998_, _34996_, _06844_);
  and (_34999_, _34998_, _34995_);
  and (_35000_, _15168_, _08606_);
  or (_35001_, _35000_, _34987_);
  and (_35002_, _35001_, _06393_);
  or (_35003_, _35002_, _06387_);
  or (_35004_, _35003_, _34999_);
  or (_35005_, _34987_, _15138_);
  and (_35006_, _35005_, _34989_);
  or (_35007_, _35006_, _07245_);
  and (_35009_, _35007_, _06446_);
  and (_35010_, _35009_, _35004_);
  and (_35011_, _15189_, _08606_);
  or (_35012_, _35011_, _34987_);
  and (_35013_, _35012_, _06300_);
  or (_35014_, _35013_, _10059_);
  or (_35015_, _35014_, _35010_);
  and (_35016_, _35015_, _34973_);
  or (_35017_, _35016_, _06281_);
  and (_35018_, _07972_, _09442_);
  or (_35020_, _34970_, _06282_);
  or (_35021_, _35020_, _35018_);
  and (_35022_, _35021_, _06279_);
  and (_35023_, _35022_, _35017_);
  and (_35024_, _15243_, _07972_);
  or (_35025_, _35024_, _34970_);
  and (_35026_, _35025_, _06015_);
  or (_35027_, _35026_, _06275_);
  or (_35028_, _35027_, _35023_);
  and (_35029_, _08883_, _07972_);
  or (_35031_, _35029_, _34970_);
  or (_35032_, _35031_, _06276_);
  and (_35033_, _35032_, _35028_);
  or (_35034_, _35033_, _06474_);
  and (_35035_, _15135_, _07972_);
  or (_35036_, _35035_, _34970_);
  or (_35037_, _35036_, _07282_);
  and (_35038_, _35037_, _07284_);
  and (_35039_, _35038_, _35034_);
  and (_35040_, _11216_, _07972_);
  or (_35042_, _35040_, _34970_);
  and (_35043_, _35042_, _06582_);
  or (_35044_, _35043_, _35039_);
  and (_35045_, _35044_, _07279_);
  or (_35046_, _34970_, _08345_);
  and (_35047_, _35031_, _06478_);
  and (_35048_, _35047_, _35046_);
  or (_35049_, _35048_, _35045_);
  and (_35050_, _35049_, _07276_);
  and (_35051_, _34979_, _06569_);
  and (_35053_, _35051_, _35046_);
  or (_35054_, _35053_, _06479_);
  or (_35055_, _35054_, _35050_);
  and (_35056_, _15134_, _07972_);
  or (_35057_, _34970_, _09043_);
  or (_35058_, _35057_, _35056_);
  and (_35059_, _35058_, _09048_);
  and (_35060_, _35059_, _35055_);
  nor (_35061_, _11215_, _13664_);
  or (_35062_, _35061_, _34970_);
  and (_35064_, _35062_, _06572_);
  or (_35065_, _35064_, _06606_);
  or (_35066_, _35065_, _35060_);
  or (_35067_, _34976_, _07037_);
  and (_35068_, _35067_, _06807_);
  and (_35069_, _35068_, _35066_);
  and (_35070_, _35001_, _06234_);
  or (_35071_, _35070_, _06195_);
  or (_35072_, _35071_, _35069_);
  and (_35073_, _15315_, _07972_);
  or (_35075_, _34970_, _06196_);
  or (_35076_, _35075_, _35073_);
  and (_35077_, _35076_, _01375_);
  and (_35078_, _35077_, _35072_);
  or (_35079_, _35078_, _34969_);
  and (_43045_, _35079_, _42545_);
  and (_35080_, _01379_, \uc8051golden_1.SCON [5]);
  and (_35081_, _13664_, \uc8051golden_1.SCON [5]);
  nor (_35082_, _13664_, _08207_);
  or (_35083_, _35082_, _35081_);
  or (_35085_, _35083_, _06293_);
  and (_35086_, _15348_, _07972_);
  or (_35087_, _35086_, _35081_);
  or (_35088_, _35087_, _07210_);
  and (_35089_, _07972_, \uc8051golden_1.ACC [5]);
  or (_35090_, _35089_, _35081_);
  and (_35091_, _35090_, _07199_);
  and (_35092_, _07200_, \uc8051golden_1.SCON [5]);
  or (_35093_, _35092_, _06401_);
  or (_35094_, _35093_, _35091_);
  and (_35096_, _35094_, _06396_);
  and (_35097_, _35096_, _35088_);
  and (_35098_, _13673_, \uc8051golden_1.SCON [5]);
  and (_35099_, _15341_, _08606_);
  or (_35100_, _35099_, _35098_);
  and (_35101_, _35100_, _06395_);
  or (_35102_, _35101_, _06399_);
  or (_35103_, _35102_, _35097_);
  or (_35104_, _35083_, _07221_);
  and (_35105_, _35104_, _35103_);
  or (_35107_, _35105_, _06406_);
  or (_35108_, _35090_, _06414_);
  and (_35109_, _35108_, _06844_);
  and (_35110_, _35109_, _35107_);
  and (_35111_, _15345_, _08606_);
  or (_35112_, _35111_, _35098_);
  and (_35113_, _35112_, _06393_);
  or (_35114_, _35113_, _06387_);
  or (_35115_, _35114_, _35110_);
  or (_35116_, _35098_, _15378_);
  and (_35118_, _35116_, _35100_);
  or (_35119_, _35118_, _07245_);
  and (_35120_, _35119_, _06446_);
  and (_35121_, _35120_, _35115_);
  or (_35122_, _35098_, _15342_);
  and (_35123_, _35122_, _06300_);
  and (_35124_, _35123_, _35100_);
  or (_35125_, _35124_, _10059_);
  or (_35126_, _35125_, _35121_);
  and (_35127_, _35126_, _35085_);
  or (_35129_, _35127_, _06281_);
  and (_35130_, _07972_, _09441_);
  or (_35131_, _35081_, _06282_);
  or (_35132_, _35131_, _35130_);
  and (_35133_, _35132_, _06279_);
  and (_35134_, _35133_, _35129_);
  and (_35135_, _15446_, _07972_);
  or (_35136_, _35135_, _35081_);
  and (_35137_, _35136_, _06015_);
  or (_35138_, _35137_, _06275_);
  or (_35140_, _35138_, _35134_);
  and (_35141_, _08958_, _07972_);
  or (_35142_, _35141_, _35081_);
  or (_35143_, _35142_, _06276_);
  and (_35144_, _35143_, _35140_);
  or (_35145_, _35144_, _06474_);
  and (_35146_, _15338_, _07972_);
  or (_35147_, _35146_, _35081_);
  or (_35148_, _35147_, _07282_);
  and (_35149_, _35148_, _07284_);
  and (_35151_, _35149_, _35145_);
  and (_35152_, _12542_, _07972_);
  or (_35153_, _35152_, _35081_);
  and (_35154_, _35153_, _06582_);
  or (_35155_, _35154_, _35151_);
  and (_35156_, _35155_, _07279_);
  or (_35157_, _35081_, _08256_);
  and (_35158_, _35142_, _06478_);
  and (_35159_, _35158_, _35157_);
  or (_35160_, _35159_, _35156_);
  and (_35162_, _35160_, _07276_);
  and (_35163_, _35090_, _06569_);
  and (_35164_, _35163_, _35157_);
  or (_35165_, _35164_, _06479_);
  or (_35166_, _35165_, _35162_);
  and (_35167_, _15335_, _07972_);
  or (_35168_, _35081_, _09043_);
  or (_35169_, _35168_, _35167_);
  and (_35170_, _35169_, _09048_);
  and (_35171_, _35170_, _35166_);
  nor (_35173_, _11212_, _13664_);
  or (_35174_, _35173_, _35081_);
  and (_35175_, _35174_, _06572_);
  or (_35176_, _35175_, _06606_);
  or (_35177_, _35176_, _35171_);
  or (_35178_, _35087_, _07037_);
  and (_35179_, _35178_, _06807_);
  and (_35180_, _35179_, _35177_);
  and (_35181_, _35112_, _06234_);
  or (_35182_, _35181_, _06195_);
  or (_35184_, _35182_, _35180_);
  and (_35185_, _15509_, _07972_);
  or (_35186_, _35081_, _06196_);
  or (_35187_, _35186_, _35185_);
  and (_35188_, _35187_, _01375_);
  and (_35189_, _35188_, _35184_);
  or (_35190_, _35189_, _35080_);
  and (_43046_, _35190_, _42545_);
  and (_35191_, _01379_, \uc8051golden_1.SCON [6]);
  and (_35192_, _13664_, \uc8051golden_1.SCON [6]);
  nor (_35194_, _13664_, _08118_);
  or (_35195_, _35194_, _35192_);
  or (_35196_, _35195_, _06293_);
  and (_35197_, _15550_, _07972_);
  or (_35198_, _35197_, _35192_);
  or (_35199_, _35198_, _07210_);
  and (_35200_, _07972_, \uc8051golden_1.ACC [6]);
  or (_35201_, _35200_, _35192_);
  and (_35202_, _35201_, _07199_);
  and (_35203_, _07200_, \uc8051golden_1.SCON [6]);
  or (_35205_, _35203_, _06401_);
  or (_35206_, _35205_, _35202_);
  and (_35207_, _35206_, _06396_);
  and (_35208_, _35207_, _35199_);
  and (_35209_, _13673_, \uc8051golden_1.SCON [6]);
  and (_35210_, _15535_, _08606_);
  or (_35211_, _35210_, _35209_);
  and (_35212_, _35211_, _06395_);
  or (_35213_, _35212_, _06399_);
  or (_35214_, _35213_, _35208_);
  or (_35216_, _35195_, _07221_);
  and (_35217_, _35216_, _35214_);
  or (_35218_, _35217_, _06406_);
  or (_35219_, _35201_, _06414_);
  and (_35220_, _35219_, _06844_);
  and (_35221_, _35220_, _35218_);
  and (_35222_, _15561_, _08606_);
  or (_35223_, _35222_, _35209_);
  and (_35224_, _35223_, _06393_);
  or (_35225_, _35224_, _06387_);
  or (_35227_, _35225_, _35221_);
  or (_35228_, _35209_, _15568_);
  and (_35229_, _35228_, _35211_);
  or (_35230_, _35229_, _07245_);
  and (_35231_, _35230_, _06446_);
  and (_35232_, _35231_, _35227_);
  and (_35233_, _15585_, _08606_);
  or (_35234_, _35233_, _35209_);
  and (_35235_, _35234_, _06300_);
  or (_35236_, _35235_, _10059_);
  or (_35238_, _35236_, _35232_);
  and (_35239_, _35238_, _35196_);
  or (_35240_, _35239_, _06281_);
  and (_35241_, _07972_, _09440_);
  or (_35242_, _35192_, _06282_);
  or (_35243_, _35242_, _35241_);
  and (_35244_, _35243_, _06279_);
  and (_35245_, _35244_, _35240_);
  and (_35246_, _15639_, _07972_);
  or (_35247_, _35246_, _35192_);
  and (_35249_, _35247_, _06015_);
  or (_35250_, _35249_, _06275_);
  or (_35251_, _35250_, _35245_);
  and (_35252_, _15646_, _07972_);
  or (_35253_, _35252_, _35192_);
  or (_35254_, _35253_, _06276_);
  and (_35255_, _35254_, _35251_);
  or (_35256_, _35255_, _06474_);
  and (_35257_, _15531_, _07972_);
  or (_35258_, _35257_, _35192_);
  or (_35260_, _35258_, _07282_);
  and (_35261_, _35260_, _07284_);
  and (_35262_, _35261_, _35256_);
  and (_35263_, _11210_, _07972_);
  or (_35264_, _35263_, _35192_);
  and (_35265_, _35264_, _06582_);
  or (_35266_, _35265_, _35262_);
  and (_35267_, _35266_, _07279_);
  or (_35268_, _35192_, _08162_);
  and (_35269_, _35253_, _06478_);
  and (_35271_, _35269_, _35268_);
  or (_35272_, _35271_, _35267_);
  and (_35273_, _35272_, _07276_);
  and (_35274_, _35201_, _06569_);
  and (_35275_, _35274_, _35268_);
  or (_35276_, _35275_, _06479_);
  or (_35277_, _35276_, _35273_);
  and (_35278_, _15528_, _07972_);
  or (_35279_, _35192_, _09043_);
  or (_35280_, _35279_, _35278_);
  and (_35282_, _35280_, _09048_);
  and (_35283_, _35282_, _35277_);
  nor (_35284_, _11209_, _13664_);
  or (_35285_, _35284_, _35192_);
  and (_35286_, _35285_, _06572_);
  or (_35287_, _35286_, _06606_);
  or (_35288_, _35287_, _35283_);
  or (_35289_, _35198_, _07037_);
  and (_35290_, _35289_, _06807_);
  and (_35291_, _35290_, _35288_);
  and (_35293_, _35223_, _06234_);
  or (_35294_, _35293_, _06195_);
  or (_35295_, _35294_, _35291_);
  and (_35296_, _15713_, _07972_);
  or (_35297_, _35192_, _06196_);
  or (_35298_, _35297_, _35296_);
  and (_35299_, _35298_, _01375_);
  and (_35300_, _35299_, _35295_);
  or (_35301_, _35300_, _35191_);
  and (_43047_, _35301_, _42545_);
  nor (_35303_, _01375_, _06270_);
  nor (_35304_, _07956_, _06270_);
  and (_35305_, _07956_, \uc8051golden_1.ACC [0]);
  and (_35306_, _35305_, _08521_);
  or (_35307_, _35306_, _35304_);
  or (_35308_, _35307_, _07276_);
  nor (_35309_, _08521_, _13789_);
  or (_35310_, _35309_, _35304_);
  or (_35311_, _35310_, _07210_);
  or (_35312_, _35305_, _35304_);
  and (_35314_, _35312_, _07199_);
  nor (_35315_, _07199_, _06270_);
  or (_35316_, _35315_, _06401_);
  or (_35317_, _35316_, _35314_);
  and (_35318_, _35317_, _07221_);
  nand (_35319_, _35318_, _35311_);
  nand (_35320_, _35319_, _06871_);
  or (_35321_, _35312_, _06414_);
  and (_35322_, _35321_, _07785_);
  and (_35323_, _35322_, _35320_);
  nand (_35325_, _07510_, _06293_);
  or (_35326_, _35325_, _35323_);
  and (_35327_, _08236_, _07473_);
  or (_35328_, _35304_, _06293_);
  or (_35329_, _35328_, _35327_);
  and (_35330_, _35329_, _35326_);
  or (_35331_, _35330_, _06281_);
  or (_35332_, _35304_, _06282_);
  and (_35333_, _07956_, _09446_);
  or (_35334_, _35333_, _35332_);
  and (_35336_, _35334_, _35331_);
  or (_35337_, _35336_, _06015_);
  and (_35338_, _14426_, _08236_);
  or (_35339_, _35304_, _06279_);
  or (_35340_, _35339_, _35338_);
  and (_35341_, _35340_, _06276_);
  and (_35342_, _35341_, _35337_);
  and (_35343_, _07956_, _08817_);
  or (_35344_, _35343_, _35304_);
  and (_35345_, _35344_, _06275_);
  or (_35347_, _35345_, _06474_);
  or (_35348_, _35347_, _35342_);
  and (_35349_, _14324_, _07956_);
  or (_35350_, _35349_, _35304_);
  or (_35351_, _35350_, _07282_);
  and (_35352_, _35351_, _07284_);
  and (_35353_, _35352_, _35348_);
  nor (_35354_, _12538_, _13789_);
  or (_35355_, _35354_, _35304_);
  nor (_35356_, _35306_, _07284_);
  and (_35358_, _35356_, _35355_);
  or (_35359_, _35358_, _35353_);
  and (_35360_, _35359_, _07279_);
  nand (_35361_, _35344_, _06478_);
  nor (_35362_, _35361_, _35309_);
  or (_35363_, _35362_, _06569_);
  or (_35364_, _35363_, _35360_);
  and (_35365_, _35364_, _35308_);
  or (_35366_, _35365_, _06479_);
  and (_35367_, _14320_, _07956_);
  or (_35368_, _35367_, _35304_);
  or (_35369_, _35368_, _09043_);
  and (_35370_, _35369_, _09048_);
  and (_35371_, _35370_, _35366_);
  and (_35372_, _35355_, _06572_);
  or (_35373_, _35372_, _19434_);
  or (_35374_, _35373_, _35371_);
  or (_35375_, _35310_, _06700_);
  and (_35376_, _35375_, _01375_);
  and (_35377_, _35376_, _35374_);
  or (_35379_, _35377_, _35303_);
  and (_43048_, _35379_, _42545_);
  nand (_35380_, _08236_, _07090_);
  or (_35381_, _35380_, _08477_);
  or (_35382_, _07956_, \uc8051golden_1.SP [1]);
  and (_35383_, _35382_, _06479_);
  and (_35384_, _35383_, _35381_);
  and (_35385_, _11222_, _08236_);
  nor (_35386_, _07956_, _06268_);
  or (_35387_, _35386_, _07276_);
  or (_35389_, _35387_, _35385_);
  and (_35390_, _14532_, _08236_);
  not (_35391_, _35390_);
  and (_35392_, _35391_, _35382_);
  or (_35393_, _35392_, _07210_);
  nand (_35394_, _06790_, \uc8051golden_1.SP [1]);
  and (_35395_, _07956_, \uc8051golden_1.ACC [1]);
  or (_35396_, _35395_, _35386_);
  and (_35397_, _35396_, _07199_);
  nor (_35398_, _07199_, _06268_);
  or (_35400_, _35398_, _06790_);
  or (_35401_, _35400_, _35397_);
  and (_35402_, _35401_, _35394_);
  or (_35403_, _35402_, _06401_);
  and (_35404_, _35403_, _05997_);
  and (_35405_, _35404_, _35393_);
  nor (_35406_, _05997_, \uc8051golden_1.SP [1]);
  or (_35407_, _35406_, _06399_);
  or (_35408_, _35407_, _35405_);
  nand (_35409_, _06399_, _06273_);
  and (_35411_, _35409_, _35408_);
  or (_35412_, _35411_, _06406_);
  or (_35413_, _35396_, _06414_);
  and (_35414_, _35413_, _07785_);
  and (_35415_, _35414_, _35412_);
  not (_35416_, _07350_);
  or (_35417_, _35416_, _07243_);
  or (_35418_, _35417_, _35415_);
  or (_35419_, _07350_, _06268_);
  and (_35420_, _35419_, _06293_);
  and (_35422_, _35420_, _35418_);
  nand (_35423_, _08236_, _07196_);
  and (_35424_, _35382_, _10059_);
  and (_35425_, _35424_, _35423_);
  or (_35426_, _35425_, _06281_);
  or (_35427_, _35426_, _35422_);
  or (_35428_, _35386_, _06282_);
  and (_35429_, _07956_, _09445_);
  or (_35430_, _35429_, _35428_);
  and (_35431_, _35430_, _06279_);
  and (_35433_, _35431_, _35427_);
  and (_35434_, _35382_, _06015_);
  or (_35435_, _14615_, _13789_);
  and (_35436_, _35435_, _35434_);
  or (_35437_, _35436_, _35433_);
  and (_35438_, _35437_, _06276_);
  and (_35439_, _35382_, _06275_);
  and (_35440_, _35439_, _35380_);
  or (_35441_, _35440_, _05943_);
  or (_35442_, _35441_, _35438_);
  nand (_35444_, _05943_, \uc8051golden_1.SP [1]);
  and (_35445_, _35444_, _07282_);
  and (_35446_, _35445_, _35442_);
  or (_35447_, _14507_, _13789_);
  and (_35448_, _35382_, _06474_);
  and (_35449_, _35448_, _35447_);
  or (_35450_, _35449_, _06582_);
  or (_35451_, _35450_, _35446_);
  and (_35452_, _11224_, _07956_);
  or (_35453_, _35452_, _35386_);
  or (_35455_, _35453_, _07284_);
  and (_35456_, _35455_, _07279_);
  and (_35457_, _35456_, _35451_);
  or (_35458_, _14505_, _13789_);
  and (_35459_, _35382_, _06478_);
  and (_35460_, _35459_, _35458_);
  or (_35461_, _35460_, _06569_);
  or (_35462_, _35461_, _35457_);
  and (_35463_, _35462_, _35389_);
  or (_35464_, _35463_, _05956_);
  nand (_35466_, _05956_, \uc8051golden_1.SP [1]);
  and (_35467_, _35466_, _09043_);
  and (_35468_, _35467_, _35464_);
  or (_35469_, _35468_, _35384_);
  and (_35470_, _35469_, _09048_);
  nor (_35471_, _11223_, _13789_);
  or (_35472_, _35471_, _35386_);
  and (_35473_, _35472_, _06572_);
  or (_35474_, _35473_, _06588_);
  or (_35475_, _35474_, _35470_);
  nand (_35477_, _35475_, _07121_);
  nor (_35478_, _06305_, _05966_);
  nand (_35479_, _35478_, _35477_);
  or (_35480_, _35478_, _06268_);
  and (_35481_, _35480_, _07037_);
  and (_35482_, _35481_, _35479_);
  and (_35483_, _35392_, _06606_);
  or (_35484_, _35483_, _07887_);
  or (_35485_, _35484_, _35482_);
  or (_35486_, _07312_, _06268_);
  and (_35488_, _35486_, _06196_);
  and (_35489_, _35488_, _35485_);
  or (_35490_, _35390_, _35386_);
  and (_35491_, _35490_, _06195_);
  or (_35492_, _35491_, _01379_);
  or (_35493_, _35492_, _35489_);
  or (_35494_, _01375_, \uc8051golden_1.SP [1]);
  and (_35495_, _35494_, _42545_);
  and (_43049_, _35495_, _35493_);
  nor (_35496_, _01375_, _06738_);
  nand (_35498_, _14714_, _05943_);
  nor (_35499_, _13789_, _07623_);
  nor (_35500_, _07956_, _06738_);
  or (_35501_, _35500_, _06293_);
  or (_35502_, _35501_, _35499_);
  or (_35503_, _07659_, _07349_);
  and (_35504_, _14754_, _08236_);
  or (_35505_, _35504_, _35500_);
  or (_35506_, _35505_, _07210_);
  and (_35507_, _07956_, \uc8051golden_1.ACC [2]);
  or (_35509_, _35507_, _35500_);
  or (_35510_, _35509_, _07200_);
  or (_35511_, _07199_, \uc8051golden_1.SP [2]);
  and (_35512_, _35511_, _07366_);
  and (_35513_, _35512_, _35510_);
  and (_35514_, _07912_, _06790_);
  or (_35515_, _35514_, _06401_);
  or (_35516_, _35515_, _35513_);
  and (_35517_, _35516_, _05997_);
  and (_35518_, _35517_, _35506_);
  nor (_35520_, _14714_, _05997_);
  or (_35521_, _35520_, _06399_);
  or (_35522_, _35521_, _35518_);
  nand (_35523_, _08677_, _06399_);
  and (_35524_, _35523_, _35522_);
  or (_35525_, _35524_, _06406_);
  or (_35526_, _35509_, _06414_);
  and (_35527_, _35526_, _07785_);
  and (_35528_, _35527_, _35525_);
  or (_35529_, _35528_, _35503_);
  nor (_35531_, _07912_, _05994_);
  nor (_35532_, _35531_, _06017_);
  and (_35533_, _35532_, _35529_);
  nand (_35534_, _07912_, _06017_);
  nand (_35535_, _35534_, _06293_);
  or (_35536_, _35535_, _35533_);
  and (_35537_, _35536_, _35502_);
  or (_35538_, _35537_, _06281_);
  or (_35539_, _35500_, _06282_);
  and (_35540_, _07956_, _09444_);
  or (_35542_, _35540_, _35539_);
  and (_35543_, _35542_, _06279_);
  and (_35544_, _35543_, _35538_);
  and (_35545_, _14848_, _07956_);
  or (_35546_, _35545_, _35500_);
  and (_35547_, _35546_, _06015_);
  or (_35548_, _35547_, _06275_);
  or (_35549_, _35548_, _35544_);
  and (_35550_, _07956_, _08994_);
  or (_35551_, _35550_, _35500_);
  or (_35553_, _35551_, _06276_);
  and (_35554_, _35553_, _35549_);
  or (_35555_, _35554_, _05943_);
  and (_35556_, _35555_, _35498_);
  or (_35557_, _35556_, _06474_);
  and (_35558_, _14744_, _07956_);
  or (_35559_, _35558_, _35500_);
  or (_35560_, _35559_, _07282_);
  and (_35561_, _35560_, _07284_);
  and (_35562_, _35561_, _35557_);
  and (_35564_, _11221_, _07956_);
  or (_35565_, _35564_, _35500_);
  and (_35566_, _35565_, _06582_);
  or (_35567_, _35566_, _35562_);
  and (_35568_, _35567_, _07279_);
  or (_35569_, _35500_, _08433_);
  and (_35570_, _35551_, _06478_);
  and (_35571_, _35570_, _35569_);
  or (_35572_, _35571_, _35568_);
  and (_35573_, _35572_, _12731_);
  and (_35575_, _35509_, _06569_);
  and (_35576_, _35575_, _35569_);
  and (_35577_, _07912_, _05956_);
  or (_35578_, _35577_, _06479_);
  or (_35579_, _35578_, _35576_);
  or (_35580_, _35579_, _35573_);
  and (_35581_, _14741_, _07956_);
  or (_35582_, _35581_, _35500_);
  or (_35583_, _35582_, _09043_);
  and (_35584_, _35583_, _35580_);
  or (_35586_, _35584_, _06572_);
  nor (_35587_, _11220_, _13789_);
  or (_35588_, _35587_, _35500_);
  or (_35589_, _35588_, _09048_);
  and (_35590_, _35589_, _13881_);
  and (_35591_, _35590_, _35586_);
  and (_35592_, _14714_, _06588_);
  or (_35593_, _35592_, _05966_);
  or (_35594_, _35593_, _35591_);
  nand (_35595_, _14714_, _05966_);
  and (_35597_, _35595_, _06306_);
  and (_35598_, _35597_, _35594_);
  and (_35599_, _14714_, _06305_);
  or (_35600_, _35599_, _06606_);
  or (_35601_, _35600_, _35598_);
  or (_35602_, _35505_, _07037_);
  and (_35603_, _35602_, _07312_);
  and (_35604_, _35603_, _35601_);
  nor (_35605_, _14714_, _07312_);
  or (_35606_, _35605_, _06195_);
  or (_35608_, _35606_, _35604_);
  and (_35609_, _14917_, _08236_);
  or (_35610_, _35500_, _06196_);
  or (_35611_, _35610_, _35609_);
  and (_35612_, _35611_, _01375_);
  and (_35613_, _35612_, _35608_);
  or (_35614_, _35613_, _35496_);
  and (_43050_, _35614_, _42545_);
  nor (_35615_, _01375_, _06398_);
  or (_35616_, _07915_, _07312_);
  nand (_35618_, _14718_, _05966_);
  nand (_35619_, _14718_, _05943_);
  nor (_35620_, _13789_, _07775_);
  nor (_35621_, _07956_, _06398_);
  or (_35622_, _35621_, _06281_);
  or (_35623_, _35622_, _35620_);
  and (_35624_, _35623_, _13788_);
  and (_35625_, _14947_, _08236_);
  or (_35626_, _35625_, _35621_);
  or (_35627_, _35626_, _07210_);
  and (_35629_, _07956_, \uc8051golden_1.ACC [3]);
  or (_35630_, _35629_, _35621_);
  or (_35631_, _35630_, _07200_);
  or (_35632_, _07199_, \uc8051golden_1.SP [3]);
  and (_35633_, _35632_, _07366_);
  and (_35634_, _35633_, _35631_);
  and (_35635_, _07915_, _06790_);
  or (_35636_, _35635_, _06401_);
  or (_35637_, _35636_, _35634_);
  and (_35638_, _35637_, _05997_);
  and (_35640_, _35638_, _35627_);
  nor (_35641_, _14718_, _05997_);
  or (_35642_, _35641_, _06399_);
  or (_35643_, _35642_, _35640_);
  nand (_35644_, _08666_, _06399_);
  and (_35645_, _35644_, _35643_);
  or (_35646_, _35645_, _06406_);
  or (_35647_, _35630_, _06414_);
  and (_35648_, _35647_, _07785_);
  and (_35649_, _35648_, _35646_);
  or (_35651_, _07827_, _35416_);
  or (_35652_, _35651_, _35649_);
  or (_35653_, _07915_, _07350_);
  and (_35654_, _35653_, _06293_);
  and (_35655_, _35654_, _35652_);
  or (_35656_, _35655_, _35624_);
  or (_35657_, _35621_, _06282_);
  and (_35658_, _07956_, _09443_);
  or (_35659_, _35658_, _35657_);
  and (_35660_, _35659_, _06279_);
  and (_35662_, _35660_, _35656_);
  and (_35663_, _15039_, _07956_);
  or (_35664_, _35663_, _35621_);
  and (_35665_, _35664_, _06015_);
  or (_35666_, _35665_, _06275_);
  or (_35667_, _35666_, _35662_);
  and (_35668_, _07956_, _08815_);
  or (_35669_, _35668_, _35621_);
  or (_35670_, _35669_, _06276_);
  and (_35671_, _35670_, _35667_);
  or (_35673_, _35671_, _05943_);
  and (_35674_, _35673_, _35619_);
  or (_35675_, _35674_, _06474_);
  and (_35676_, _14934_, _07956_);
  or (_35677_, _35676_, _35621_);
  or (_35678_, _35677_, _07282_);
  and (_35679_, _35678_, _07284_);
  and (_35680_, _35679_, _35675_);
  and (_35681_, _12535_, _07956_);
  or (_35682_, _35681_, _35621_);
  and (_35684_, _35682_, _06582_);
  or (_35685_, _35684_, _35680_);
  and (_35686_, _35685_, _07279_);
  or (_35687_, _35621_, _08389_);
  and (_35688_, _35669_, _06478_);
  and (_35689_, _35688_, _35687_);
  or (_35690_, _35689_, _35686_);
  and (_35691_, _35690_, _12731_);
  and (_35692_, _35630_, _06569_);
  and (_35693_, _35692_, _35687_);
  and (_35695_, _07915_, _05956_);
  or (_35696_, _35695_, _06479_);
  or (_35697_, _35696_, _35693_);
  or (_35698_, _35697_, _35691_);
  and (_35699_, _14931_, _08236_);
  or (_35700_, _35621_, _09043_);
  or (_35701_, _35700_, _35699_);
  and (_35702_, _35701_, _35698_);
  or (_35703_, _35702_, _06572_);
  nor (_35704_, _11218_, _13789_);
  or (_35706_, _35704_, _35621_);
  or (_35707_, _35706_, _09048_);
  and (_35708_, _35707_, _13881_);
  and (_35709_, _35708_, _35703_);
  nor (_35710_, _08663_, _06398_);
  or (_35711_, _35710_, _08664_);
  and (_35712_, _35711_, _06588_);
  or (_35713_, _35712_, _05966_);
  or (_35714_, _35713_, _35709_);
  and (_35715_, _35714_, _35618_);
  or (_35717_, _35715_, _06305_);
  or (_35718_, _35711_, _06306_);
  and (_35719_, _35718_, _07037_);
  and (_35720_, _35719_, _35717_);
  and (_35721_, _35626_, _06606_);
  or (_35722_, _35721_, _07887_);
  or (_35723_, _35722_, _35720_);
  and (_35724_, _35723_, _35616_);
  or (_35725_, _35724_, _06195_);
  and (_35726_, _15113_, _08236_);
  or (_35728_, _35621_, _06196_);
  or (_35729_, _35728_, _35726_);
  and (_35730_, _35729_, _01375_);
  and (_35731_, _35730_, _35725_);
  or (_35732_, _35731_, _35615_);
  and (_43052_, _35732_, _42545_);
  nor (_35733_, _01375_, _13813_);
  nor (_35734_, _07781_, \uc8051golden_1.SP [4]);
  nor (_35735_, _35734_, _13777_);
  or (_35736_, _35735_, _07312_);
  nor (_35738_, _13789_, _08301_);
  nor (_35739_, _07956_, _13813_);
  or (_35740_, _35739_, _06281_);
  or (_35741_, _35740_, _35738_);
  and (_35742_, _35741_, _13788_);
  and (_35743_, _15130_, _08236_);
  or (_35744_, _35743_, _35739_);
  or (_35745_, _35744_, _07210_);
  and (_35746_, _07956_, \uc8051golden_1.ACC [4]);
  or (_35747_, _35746_, _35739_);
  or (_35749_, _35747_, _07200_);
  or (_35750_, _07199_, \uc8051golden_1.SP [4]);
  and (_35751_, _35750_, _07366_);
  and (_35752_, _35751_, _35749_);
  and (_35753_, _35735_, _06790_);
  or (_35754_, _35753_, _06401_);
  or (_35755_, _35754_, _35752_);
  and (_35756_, _35755_, _05997_);
  and (_35757_, _35756_, _35745_);
  and (_35758_, _35735_, _07351_);
  or (_35760_, _35758_, _06399_);
  or (_35761_, _35760_, _35757_);
  and (_35762_, _13814_, _06270_);
  nor (_35763_, _08665_, _13813_);
  nor (_35764_, _35763_, _35762_);
  nand (_35765_, _35764_, _06399_);
  and (_35766_, _35765_, _35761_);
  or (_35767_, _35766_, _06406_);
  or (_35768_, _35747_, _06414_);
  and (_35769_, _35768_, _07785_);
  and (_35771_, _35769_, _35767_);
  and (_35772_, _07782_, \uc8051golden_1.SP [4]);
  nor (_35773_, _07782_, \uc8051golden_1.SP [4]);
  nor (_35774_, _35773_, _35772_);
  nand (_35775_, _35774_, _06419_);
  nand (_35776_, _35775_, _07350_);
  or (_35777_, _35776_, _35771_);
  or (_35778_, _35735_, _07350_);
  and (_35779_, _35778_, _06293_);
  and (_35780_, _35779_, _35777_);
  or (_35782_, _35780_, _35742_);
  or (_35783_, _35739_, _06282_);
  and (_35784_, _07956_, _09442_);
  or (_35785_, _35784_, _35783_);
  and (_35786_, _35785_, _06279_);
  and (_35787_, _35786_, _35782_);
  and (_35788_, _15243_, _07956_);
  or (_35789_, _35788_, _35739_);
  and (_35790_, _35789_, _06015_);
  or (_35791_, _35790_, _06275_);
  or (_35793_, _35791_, _35787_);
  and (_35794_, _08883_, _07956_);
  or (_35795_, _35794_, _35739_);
  or (_35796_, _35795_, _06276_);
  and (_35797_, _35796_, _35793_);
  or (_35798_, _35797_, _05943_);
  or (_35799_, _35735_, _13854_);
  and (_35800_, _35799_, _35798_);
  or (_35801_, _35800_, _06474_);
  and (_35802_, _15135_, _07956_);
  or (_35804_, _35802_, _35739_);
  or (_35805_, _35804_, _07282_);
  and (_35806_, _35805_, _07284_);
  and (_35807_, _35806_, _35801_);
  and (_35808_, _11216_, _07956_);
  or (_35809_, _35808_, _35739_);
  and (_35810_, _35809_, _06582_);
  or (_35811_, _35810_, _35807_);
  and (_35812_, _35811_, _07279_);
  or (_35813_, _35739_, _08345_);
  and (_35815_, _35795_, _06478_);
  and (_35816_, _35815_, _35813_);
  or (_35817_, _35816_, _35812_);
  and (_35818_, _35817_, _12731_);
  and (_35819_, _35747_, _06569_);
  and (_35820_, _35819_, _35813_);
  and (_35821_, _35735_, _05956_);
  or (_35822_, _35821_, _06479_);
  or (_35823_, _35822_, _35820_);
  or (_35824_, _35823_, _35818_);
  and (_35826_, _15134_, _07956_);
  or (_35827_, _35826_, _35739_);
  or (_35828_, _35827_, _09043_);
  and (_35829_, _35828_, _35824_);
  or (_35830_, _35829_, _06572_);
  nor (_35831_, _11215_, _13789_);
  or (_35832_, _35831_, _35739_);
  or (_35833_, _35832_, _09048_);
  and (_35834_, _35833_, _13881_);
  and (_35835_, _35834_, _35830_);
  nor (_35837_, _08664_, _13813_);
  or (_35838_, _35837_, _13814_);
  and (_35839_, _35838_, _06588_);
  or (_35840_, _35839_, _05966_);
  or (_35841_, _35840_, _35835_);
  or (_35842_, _35735_, _05967_);
  and (_35843_, _35842_, _35841_);
  or (_35844_, _35843_, _06305_);
  or (_35845_, _35838_, _06306_);
  and (_35846_, _35845_, _07037_);
  and (_35848_, _35846_, _35844_);
  and (_35849_, _35744_, _06606_);
  or (_35850_, _35849_, _07887_);
  or (_35851_, _35850_, _35848_);
  and (_35852_, _35851_, _35736_);
  or (_35853_, _35852_, _06195_);
  and (_35854_, _15315_, _08236_);
  or (_35855_, _35739_, _06196_);
  or (_35856_, _35855_, _35854_);
  and (_35857_, _35856_, _01375_);
  and (_35859_, _35857_, _35853_);
  or (_35860_, _35859_, _35733_);
  and (_43053_, _35860_, _42545_);
  nor (_35861_, _01375_, _13812_);
  nor (_35862_, _13777_, \uc8051golden_1.SP [5]);
  nor (_35863_, _35862_, _13778_);
  or (_35864_, _35863_, _07312_);
  nor (_35865_, _13789_, _08207_);
  nor (_35866_, _07956_, _13812_);
  or (_35867_, _35866_, _06281_);
  or (_35869_, _35867_, _35865_);
  and (_35870_, _35869_, _13788_);
  and (_35871_, _15348_, _08236_);
  or (_35872_, _35871_, _35866_);
  or (_35873_, _35872_, _07210_);
  and (_35874_, _07956_, \uc8051golden_1.ACC [5]);
  or (_35875_, _35874_, _35866_);
  or (_35876_, _35875_, _07200_);
  or (_35877_, _07199_, \uc8051golden_1.SP [5]);
  and (_35878_, _35877_, _07366_);
  and (_35880_, _35878_, _35876_);
  and (_35881_, _35863_, _06790_);
  or (_35882_, _35881_, _06401_);
  or (_35883_, _35882_, _35880_);
  and (_35884_, _35883_, _05997_);
  and (_35885_, _35884_, _35873_);
  and (_35886_, _35863_, _07351_);
  or (_35887_, _35886_, _06399_);
  or (_35888_, _35887_, _35885_);
  and (_35889_, _13815_, _06270_);
  nor (_35891_, _35762_, _13812_);
  nor (_35892_, _35891_, _35889_);
  nand (_35893_, _35892_, _06399_);
  and (_35894_, _35893_, _35888_);
  or (_35895_, _35894_, _06406_);
  or (_35896_, _35875_, _06414_);
  and (_35897_, _35896_, _07785_);
  and (_35898_, _35897_, _35895_);
  nor (_35899_, _35772_, \uc8051golden_1.SP [5]);
  nor (_35900_, _35899_, _13827_);
  nand (_35902_, _35900_, _06419_);
  nand (_35903_, _35902_, _07350_);
  or (_35904_, _35903_, _35898_);
  or (_35905_, _35863_, _07350_);
  and (_35906_, _35905_, _06293_);
  and (_35907_, _35906_, _35904_);
  or (_35908_, _35907_, _35870_);
  or (_35909_, _35866_, _06282_);
  and (_35910_, _07956_, _09441_);
  or (_35911_, _35910_, _35909_);
  and (_35913_, _35911_, _06279_);
  and (_35914_, _35913_, _35908_);
  and (_35915_, _15446_, _07956_);
  or (_35916_, _35915_, _35866_);
  and (_35917_, _35916_, _06015_);
  or (_35918_, _35917_, _06275_);
  or (_35919_, _35918_, _35914_);
  and (_35920_, _08958_, _07956_);
  or (_35921_, _35920_, _35866_);
  or (_35922_, _35921_, _06276_);
  and (_35924_, _35922_, _35919_);
  or (_35925_, _35924_, _05943_);
  or (_35926_, _35863_, _13854_);
  and (_35927_, _35926_, _35925_);
  or (_35928_, _35927_, _06474_);
  and (_35929_, _15338_, _07956_);
  or (_35930_, _35929_, _35866_);
  or (_35931_, _35930_, _07282_);
  and (_35932_, _35931_, _07284_);
  and (_35933_, _35932_, _35928_);
  and (_35935_, _12542_, _07956_);
  or (_35936_, _35935_, _35866_);
  and (_35937_, _35936_, _06582_);
  or (_35938_, _35937_, _35933_);
  and (_35939_, _35938_, _07279_);
  or (_35940_, _35866_, _08256_);
  and (_35941_, _35921_, _06478_);
  and (_35942_, _35941_, _35940_);
  or (_35943_, _35942_, _35939_);
  and (_35944_, _35943_, _12731_);
  and (_35946_, _35875_, _06569_);
  and (_35947_, _35946_, _35940_);
  and (_35948_, _35863_, _05956_);
  or (_35949_, _35948_, _06479_);
  or (_35950_, _35949_, _35947_);
  or (_35951_, _35950_, _35944_);
  and (_35952_, _15335_, _07956_);
  or (_35953_, _35952_, _35866_);
  or (_35954_, _35953_, _09043_);
  and (_35955_, _35954_, _35951_);
  or (_35957_, _35955_, _06572_);
  nor (_35958_, _11212_, _13789_);
  or (_35959_, _35958_, _35866_);
  or (_35960_, _35959_, _09048_);
  and (_35961_, _35960_, _13881_);
  and (_35962_, _35961_, _35957_);
  nor (_35963_, _13814_, _13812_);
  or (_35964_, _35963_, _13815_);
  and (_35965_, _35964_, _06588_);
  or (_35966_, _35965_, _05966_);
  or (_35968_, _35966_, _35962_);
  or (_35969_, _35863_, _05967_);
  and (_35970_, _35969_, _35968_);
  or (_35971_, _35970_, _06305_);
  or (_35972_, _35964_, _06306_);
  and (_35973_, _35972_, _07037_);
  and (_35974_, _35973_, _35971_);
  and (_35975_, _35872_, _06606_);
  or (_35976_, _35975_, _07887_);
  or (_35977_, _35976_, _35974_);
  and (_35979_, _35977_, _35864_);
  or (_35980_, _35979_, _06195_);
  and (_35981_, _15509_, _08236_);
  or (_35982_, _35866_, _06196_);
  or (_35983_, _35982_, _35981_);
  and (_35984_, _35983_, _01375_);
  and (_35985_, _35984_, _35980_);
  or (_35986_, _35985_, _35861_);
  and (_43054_, _35986_, _42545_);
  nor (_35987_, _01375_, _13811_);
  nor (_35989_, _13789_, _08118_);
  nor (_35990_, _07956_, _13811_);
  or (_35991_, _35990_, _06293_);
  or (_35992_, _35991_, _35989_);
  and (_35993_, _15550_, _08236_);
  or (_35994_, _35993_, _35990_);
  or (_35995_, _35994_, _07210_);
  and (_35996_, _07956_, \uc8051golden_1.ACC [6]);
  or (_35997_, _35996_, _35990_);
  or (_35998_, _35997_, _07200_);
  or (_36000_, _07199_, \uc8051golden_1.SP [6]);
  and (_36001_, _36000_, _07366_);
  and (_36002_, _36001_, _35998_);
  nor (_36003_, _13778_, \uc8051golden_1.SP [6]);
  nor (_36004_, _36003_, _13779_);
  and (_36005_, _36004_, _06790_);
  or (_36006_, _36005_, _06401_);
  or (_36007_, _36006_, _36002_);
  and (_36008_, _36007_, _05997_);
  and (_36009_, _36008_, _35995_);
  and (_36011_, _36004_, _07351_);
  or (_36012_, _36011_, _06399_);
  or (_36013_, _36012_, _36009_);
  nor (_36014_, _35889_, _13811_);
  nor (_36015_, _36014_, _13817_);
  nand (_36016_, _36015_, _06399_);
  and (_36017_, _36016_, _36013_);
  or (_36018_, _36017_, _06406_);
  or (_36019_, _35997_, _06414_);
  and (_36020_, _36019_, _07785_);
  and (_36022_, _36020_, _36018_);
  nor (_36023_, _13827_, \uc8051golden_1.SP [6]);
  nor (_36024_, _36023_, _13828_);
  and (_36025_, _36024_, _06419_);
  or (_36026_, _36025_, _36022_);
  and (_36027_, _36026_, _07350_);
  and (_36028_, _36004_, _35416_);
  or (_36029_, _36028_, _10059_);
  or (_36030_, _36029_, _36027_);
  and (_36031_, _36030_, _35992_);
  or (_36033_, _36031_, _06281_);
  or (_36034_, _35990_, _06282_);
  and (_36035_, _07956_, _09440_);
  or (_36036_, _36035_, _36034_);
  and (_36037_, _36036_, _06279_);
  and (_36038_, _36037_, _36033_);
  and (_36039_, _15639_, _07956_);
  or (_36040_, _36039_, _35990_);
  and (_36041_, _36040_, _06015_);
  or (_36042_, _36041_, _06275_);
  or (_36044_, _36042_, _36038_);
  and (_36045_, _15646_, _07956_);
  or (_36046_, _36045_, _35990_);
  or (_36047_, _36046_, _06276_);
  and (_36048_, _36047_, _36044_);
  or (_36049_, _36048_, _05943_);
  or (_36050_, _36004_, _13854_);
  and (_36051_, _36050_, _36049_);
  or (_36052_, _36051_, _06474_);
  and (_36053_, _15531_, _07956_);
  or (_36055_, _36053_, _35990_);
  or (_36056_, _36055_, _07282_);
  and (_36057_, _36056_, _07284_);
  and (_36058_, _36057_, _36052_);
  and (_36059_, _11210_, _07956_);
  or (_36060_, _36059_, _35990_);
  and (_36061_, _36060_, _06582_);
  or (_36062_, _36061_, _36058_);
  and (_36063_, _36062_, _07279_);
  or (_36064_, _35990_, _08162_);
  and (_36066_, _36046_, _06478_);
  and (_36067_, _36066_, _36064_);
  or (_36068_, _36067_, _36063_);
  and (_36069_, _36068_, _12731_);
  and (_36070_, _35997_, _06569_);
  and (_36071_, _36070_, _36064_);
  and (_36072_, _36004_, _05956_);
  or (_36073_, _36072_, _06479_);
  or (_36074_, _36073_, _36071_);
  or (_36075_, _36074_, _36069_);
  and (_36077_, _15528_, _07956_);
  or (_36078_, _36077_, _35990_);
  or (_36079_, _36078_, _09043_);
  and (_36080_, _36079_, _36075_);
  or (_36081_, _36080_, _06572_);
  nor (_36082_, _11209_, _13789_);
  or (_36083_, _36082_, _35990_);
  or (_36084_, _36083_, _09048_);
  and (_36085_, _36084_, _13881_);
  and (_36086_, _36085_, _36081_);
  nor (_36088_, _13815_, _13811_);
  or (_36089_, _36088_, _13816_);
  and (_36090_, _36089_, _06588_);
  or (_36091_, _36090_, _05966_);
  or (_36092_, _36091_, _36086_);
  or (_36093_, _36004_, _05967_);
  and (_36094_, _36093_, _06306_);
  and (_36095_, _36094_, _36092_);
  and (_36096_, _36089_, _06305_);
  or (_36097_, _36096_, _06606_);
  or (_36099_, _36097_, _36095_);
  or (_36100_, _35994_, _07037_);
  and (_36101_, _36100_, _07312_);
  and (_36102_, _36101_, _36099_);
  and (_36103_, _36004_, _07887_);
  or (_36104_, _36103_, _06195_);
  or (_36105_, _36104_, _36102_);
  and (_36106_, _15713_, _08236_);
  or (_36107_, _35990_, _06196_);
  or (_36108_, _36107_, _36106_);
  and (_36110_, _36108_, _01375_);
  and (_36111_, _36110_, _36105_);
  or (_36112_, _36111_, _35987_);
  and (_43055_, _36112_, _42545_);
  not (_36113_, \uc8051golden_1.SBUF [0]);
  nor (_36114_, _01375_, _36113_);
  nand (_36115_, _11225_, _07940_);
  nor (_36116_, _07940_, _36113_);
  nor (_36117_, _36116_, _07276_);
  nand (_36118_, _36117_, _36115_);
  and (_36120_, _07940_, _07473_);
  or (_36121_, _36120_, _36116_);
  or (_36122_, _36121_, _06293_);
  nor (_36123_, _08521_, _13910_);
  or (_36124_, _36123_, _36116_);
  or (_36125_, _36124_, _07210_);
  and (_36126_, _07940_, \uc8051golden_1.ACC [0]);
  or (_36127_, _36126_, _36116_);
  and (_36128_, _36127_, _07199_);
  nor (_36129_, _07199_, _36113_);
  or (_36130_, _36129_, _06401_);
  or (_36131_, _36130_, _36128_);
  and (_36132_, _36131_, _07221_);
  and (_36133_, _36132_, _36125_);
  and (_36134_, _36121_, _06399_);
  or (_36135_, _36134_, _36133_);
  and (_36136_, _36135_, _06414_);
  and (_36137_, _36127_, _06406_);
  or (_36138_, _36137_, _10059_);
  or (_36139_, _36138_, _36136_);
  and (_36141_, _36139_, _36122_);
  or (_36142_, _36141_, _06281_);
  and (_36143_, _07940_, _09446_);
  or (_36144_, _36116_, _06282_);
  or (_36145_, _36144_, _36143_);
  and (_36146_, _36145_, _36142_);
  or (_36147_, _36146_, _06015_);
  and (_36148_, _14426_, _07940_);
  or (_36149_, _36116_, _06279_);
  or (_36150_, _36149_, _36148_);
  and (_36152_, _36150_, _06276_);
  and (_36153_, _36152_, _36147_);
  and (_36154_, _07940_, _08817_);
  or (_36155_, _36154_, _36116_);
  and (_36156_, _36155_, _06275_);
  or (_36157_, _36156_, _06474_);
  or (_36158_, _36157_, _36153_);
  and (_36159_, _14324_, _07940_);
  or (_36160_, _36159_, _36116_);
  or (_36161_, _36160_, _07282_);
  and (_36163_, _36161_, _07284_);
  and (_36164_, _36163_, _36158_);
  nor (_36165_, _12538_, _13910_);
  or (_36166_, _36165_, _36116_);
  and (_36167_, _36115_, _06582_);
  and (_36168_, _36167_, _36166_);
  or (_36169_, _36168_, _36164_);
  and (_36170_, _36169_, _07279_);
  nand (_36171_, _36155_, _06478_);
  nor (_36172_, _36171_, _36123_);
  or (_36174_, _36172_, _06569_);
  or (_36175_, _36174_, _36170_);
  and (_36176_, _36175_, _36118_);
  or (_36177_, _36176_, _06479_);
  and (_36178_, _14320_, _07940_);
  or (_36179_, _36116_, _09043_);
  or (_36180_, _36179_, _36178_);
  and (_36181_, _36180_, _09048_);
  and (_36182_, _36181_, _36177_);
  and (_36183_, _36166_, _06572_);
  or (_36185_, _36183_, _19434_);
  or (_36186_, _36185_, _36182_);
  or (_36187_, _36124_, _06700_);
  and (_36188_, _36187_, _01375_);
  and (_36189_, _36188_, _36186_);
  or (_36190_, _36189_, _36114_);
  and (_43057_, _36190_, _42545_);
  not (_36191_, \uc8051golden_1.SBUF [1]);
  nor (_36192_, _01375_, _36191_);
  nand (_36193_, _07940_, _07090_);
  or (_36195_, _07940_, \uc8051golden_1.SBUF [1]);
  and (_36196_, _36195_, _06275_);
  and (_36197_, _36196_, _36193_);
  and (_36198_, _07940_, _09445_);
  nor (_36199_, _07940_, _36191_);
  or (_36200_, _36199_, _06282_);
  or (_36201_, _36200_, _36198_);
  nor (_36202_, _13910_, _07196_);
  or (_36203_, _36199_, _23891_);
  or (_36204_, _36203_, _36202_);
  and (_36206_, _07940_, \uc8051golden_1.ACC [1]);
  or (_36207_, _36206_, _36199_);
  and (_36208_, _36207_, _06406_);
  or (_36209_, _36208_, _10059_);
  and (_36210_, _14532_, _07940_);
  not (_36211_, _36210_);
  and (_36212_, _36211_, _36195_);
  and (_36213_, _36212_, _06401_);
  nor (_36214_, _07199_, _36191_);
  and (_36215_, _36207_, _07199_);
  or (_36217_, _36215_, _36214_);
  and (_36218_, _36217_, _07210_);
  or (_36219_, _36218_, _06399_);
  or (_36220_, _36219_, _36213_);
  and (_36221_, _36220_, _06414_);
  or (_36222_, _36221_, _36209_);
  and (_36223_, _36222_, _36204_);
  or (_36224_, _36223_, _06281_);
  and (_36225_, _36224_, _06279_);
  and (_36226_, _36225_, _36201_);
  or (_36228_, _14615_, _13910_);
  and (_36229_, _36195_, _06015_);
  and (_36230_, _36229_, _36228_);
  or (_36231_, _36230_, _36226_);
  and (_36232_, _36231_, _06276_);
  or (_36233_, _36232_, _36197_);
  and (_36234_, _36233_, _07282_);
  or (_36235_, _14507_, _13910_);
  and (_36236_, _36195_, _06474_);
  and (_36237_, _36236_, _36235_);
  or (_36239_, _36237_, _06582_);
  or (_36240_, _36239_, _36234_);
  nor (_36241_, _11223_, _13910_);
  or (_36242_, _36241_, _36199_);
  nand (_36243_, _11222_, _07940_);
  and (_36244_, _36243_, _36242_);
  or (_36245_, _36244_, _07284_);
  and (_36246_, _36245_, _07279_);
  and (_36247_, _36246_, _36240_);
  or (_36248_, _14505_, _13910_);
  and (_36250_, _36195_, _06478_);
  and (_36251_, _36250_, _36248_);
  or (_36252_, _36251_, _06569_);
  or (_36253_, _36252_, _36247_);
  nor (_36254_, _36199_, _07276_);
  nand (_36255_, _36254_, _36243_);
  and (_36256_, _36255_, _09043_);
  and (_36257_, _36256_, _36253_);
  or (_36258_, _36193_, _08477_);
  and (_36259_, _36195_, _06479_);
  and (_36261_, _36259_, _36258_);
  or (_36262_, _36261_, _06572_);
  or (_36263_, _36262_, _36257_);
  or (_36264_, _36242_, _09048_);
  and (_36265_, _36264_, _07037_);
  and (_36266_, _36265_, _36263_);
  and (_36267_, _36212_, _06606_);
  or (_36268_, _36267_, _06195_);
  or (_36269_, _36268_, _36266_);
  or (_36270_, _36199_, _06196_);
  or (_36272_, _36270_, _36210_);
  and (_36273_, _36272_, _01375_);
  and (_36274_, _36273_, _36269_);
  or (_36275_, _36274_, _36192_);
  and (_43058_, _36275_, _42545_);
  and (_36276_, _01379_, \uc8051golden_1.SBUF [2]);
  and (_36277_, _13910_, \uc8051golden_1.SBUF [2]);
  and (_36278_, _07940_, _08994_);
  or (_36279_, _36278_, _36277_);
  or (_36280_, _36279_, _06276_);
  and (_36282_, _07940_, _09444_);
  or (_36283_, _36282_, _36277_);
  and (_36284_, _36283_, _06281_);
  and (_36285_, _14754_, _07940_);
  or (_36286_, _36285_, _36277_);
  or (_36287_, _36286_, _07210_);
  and (_36288_, _07940_, \uc8051golden_1.ACC [2]);
  or (_36289_, _36288_, _36277_);
  and (_36290_, _36289_, _07199_);
  and (_36291_, _07200_, \uc8051golden_1.SBUF [2]);
  or (_36293_, _36291_, _06401_);
  or (_36294_, _36293_, _36290_);
  and (_36295_, _36294_, _07221_);
  and (_36296_, _36295_, _36287_);
  nor (_36297_, _13910_, _07623_);
  or (_36298_, _36297_, _36277_);
  and (_36299_, _36298_, _06399_);
  or (_36300_, _36299_, _36296_);
  and (_36301_, _36300_, _06414_);
  and (_36302_, _36289_, _06406_);
  or (_36304_, _36302_, _10059_);
  or (_36305_, _36304_, _36301_);
  and (_36306_, _36298_, _06282_);
  or (_36307_, _36306_, _06294_);
  and (_36308_, _36307_, _36305_);
  or (_36309_, _36308_, _06015_);
  or (_36310_, _36309_, _36284_);
  and (_36311_, _14848_, _07940_);
  or (_36312_, _36311_, _36277_);
  or (_36313_, _36312_, _06279_);
  and (_36315_, _36313_, _36310_);
  or (_36316_, _36315_, _06275_);
  and (_36317_, _36316_, _36280_);
  or (_36318_, _36317_, _06474_);
  and (_36319_, _14744_, _07940_);
  or (_36320_, _36277_, _07282_);
  or (_36321_, _36320_, _36319_);
  and (_36322_, _36321_, _07284_);
  and (_36323_, _36322_, _36318_);
  and (_36324_, _11221_, _07940_);
  or (_36326_, _36324_, _36277_);
  and (_36327_, _36326_, _06582_);
  or (_36328_, _36327_, _36323_);
  and (_36329_, _36328_, _07279_);
  or (_36330_, _36277_, _08433_);
  and (_36331_, _36279_, _06478_);
  and (_36332_, _36331_, _36330_);
  or (_36333_, _36332_, _36329_);
  and (_36334_, _36333_, _07276_);
  and (_36335_, _36289_, _06569_);
  and (_36337_, _36335_, _36330_);
  or (_36338_, _36337_, _06479_);
  or (_36339_, _36338_, _36334_);
  and (_36340_, _14741_, _07940_);
  or (_36341_, _36277_, _09043_);
  or (_36342_, _36341_, _36340_);
  and (_36343_, _36342_, _09048_);
  and (_36344_, _36343_, _36339_);
  nor (_36345_, _11220_, _13910_);
  or (_36346_, _36345_, _36277_);
  and (_36348_, _36346_, _06572_);
  or (_36349_, _36348_, _36344_);
  and (_36350_, _36349_, _07037_);
  and (_36351_, _36286_, _06606_);
  or (_36352_, _36351_, _06195_);
  or (_36353_, _36352_, _36350_);
  and (_36354_, _14917_, _07940_);
  or (_36355_, _36277_, _06196_);
  or (_36356_, _36355_, _36354_);
  and (_36357_, _36356_, _01375_);
  and (_36359_, _36357_, _36353_);
  or (_36360_, _36359_, _36276_);
  and (_43059_, _36360_, _42545_);
  and (_36361_, _13910_, \uc8051golden_1.SBUF [3]);
  and (_36362_, _14934_, _07940_);
  or (_36363_, _36362_, _36361_);
  and (_36364_, _36363_, _06474_);
  and (_36365_, _07940_, _09443_);
  or (_36366_, _36365_, _36361_);
  and (_36367_, _36366_, _06281_);
  and (_36369_, _14947_, _07940_);
  or (_36370_, _36369_, _36361_);
  or (_36371_, _36370_, _07210_);
  and (_36372_, _07940_, \uc8051golden_1.ACC [3]);
  or (_36373_, _36372_, _36361_);
  and (_36374_, _36373_, _07199_);
  and (_36375_, _07200_, \uc8051golden_1.SBUF [3]);
  or (_36376_, _36375_, _06401_);
  or (_36377_, _36376_, _36374_);
  and (_36378_, _36377_, _07221_);
  and (_36380_, _36378_, _36371_);
  nor (_36381_, _13910_, _07775_);
  or (_36382_, _36381_, _36361_);
  and (_36383_, _36382_, _06399_);
  or (_36384_, _36383_, _36380_);
  and (_36385_, _36384_, _06414_);
  and (_36386_, _36373_, _06406_);
  or (_36387_, _36386_, _10059_);
  or (_36388_, _36387_, _36385_);
  and (_36389_, _36382_, _06282_);
  or (_36391_, _36389_, _06294_);
  and (_36392_, _36391_, _36388_);
  or (_36393_, _36392_, _06015_);
  or (_36394_, _36393_, _36367_);
  and (_36395_, _15039_, _07940_);
  or (_36396_, _36395_, _36361_);
  or (_36397_, _36396_, _06279_);
  and (_36398_, _36397_, _36394_);
  or (_36399_, _36398_, _06275_);
  and (_36400_, _07940_, _08815_);
  or (_36402_, _36400_, _36361_);
  or (_36403_, _36402_, _06276_);
  and (_36404_, _36403_, _07282_);
  and (_36405_, _36404_, _36399_);
  or (_36406_, _36405_, _36364_);
  and (_36407_, _36406_, _07284_);
  and (_36408_, _12535_, _07940_);
  or (_36409_, _36408_, _36361_);
  and (_36410_, _36409_, _06582_);
  or (_36411_, _36410_, _36407_);
  and (_36413_, _36411_, _07279_);
  or (_36414_, _36361_, _08389_);
  and (_36415_, _36402_, _06478_);
  and (_36416_, _36415_, _36414_);
  or (_36417_, _36416_, _36413_);
  and (_36418_, _36417_, _07276_);
  and (_36419_, _36373_, _06569_);
  and (_36420_, _36419_, _36414_);
  or (_36421_, _36420_, _06479_);
  or (_36422_, _36421_, _36418_);
  and (_36424_, _14931_, _07940_);
  or (_36425_, _36361_, _09043_);
  or (_36426_, _36425_, _36424_);
  and (_36427_, _36426_, _09048_);
  and (_36428_, _36427_, _36422_);
  nor (_36429_, _11218_, _13910_);
  or (_36430_, _36429_, _36361_);
  and (_36431_, _36430_, _06572_);
  or (_36432_, _36431_, _06606_);
  or (_36433_, _36432_, _36428_);
  or (_36435_, _36370_, _07037_);
  and (_36436_, _36435_, _06196_);
  and (_36437_, _36436_, _36433_);
  and (_36438_, _15113_, _07940_);
  or (_36439_, _36438_, _36361_);
  and (_36440_, _36439_, _06195_);
  or (_36441_, _36440_, _01379_);
  or (_36442_, _36441_, _36437_);
  or (_36443_, _01375_, \uc8051golden_1.SBUF [3]);
  and (_36444_, _36443_, _42545_);
  and (_43060_, _36444_, _36442_);
  and (_36446_, _13910_, \uc8051golden_1.SBUF [4]);
  and (_36447_, _07940_, _09442_);
  or (_36448_, _36447_, _36446_);
  and (_36449_, _36448_, _06281_);
  and (_36450_, _15130_, _07940_);
  or (_36451_, _36450_, _36446_);
  or (_36452_, _36451_, _07210_);
  and (_36453_, _07940_, \uc8051golden_1.ACC [4]);
  or (_36454_, _36453_, _36446_);
  and (_36456_, _36454_, _07199_);
  and (_36457_, _07200_, \uc8051golden_1.SBUF [4]);
  or (_36458_, _36457_, _06401_);
  or (_36459_, _36458_, _36456_);
  and (_36460_, _36459_, _07221_);
  and (_36461_, _36460_, _36452_);
  nor (_36462_, _13910_, _08301_);
  or (_36463_, _36462_, _36446_);
  and (_36464_, _36463_, _06399_);
  or (_36465_, _36464_, _36461_);
  and (_36467_, _36465_, _06414_);
  and (_36468_, _36454_, _06406_);
  or (_36469_, _36468_, _10059_);
  or (_36470_, _36469_, _36467_);
  and (_36471_, _36463_, _06282_);
  or (_36472_, _36471_, _06294_);
  and (_36473_, _36472_, _36470_);
  or (_36474_, _36473_, _06015_);
  or (_36475_, _36474_, _36449_);
  and (_36476_, _15243_, _07940_);
  or (_36478_, _36446_, _06279_);
  or (_36479_, _36478_, _36476_);
  and (_36480_, _36479_, _06276_);
  and (_36481_, _36480_, _36475_);
  and (_36482_, _08883_, _07940_);
  or (_36483_, _36482_, _36446_);
  and (_36484_, _36483_, _06275_);
  or (_36485_, _36484_, _06474_);
  or (_36486_, _36485_, _36481_);
  and (_36487_, _15135_, _07940_);
  or (_36489_, _36446_, _07282_);
  or (_36490_, _36489_, _36487_);
  and (_36491_, _36490_, _07284_);
  and (_36492_, _36491_, _36486_);
  and (_36493_, _11216_, _07940_);
  or (_36494_, _36493_, _36446_);
  and (_36495_, _36494_, _06582_);
  or (_36496_, _36495_, _36492_);
  and (_36497_, _36496_, _07279_);
  or (_36498_, _36446_, _08345_);
  and (_36500_, _36483_, _06478_);
  and (_36501_, _36500_, _36498_);
  or (_36502_, _36501_, _36497_);
  and (_36503_, _36502_, _07276_);
  and (_36504_, _36454_, _06569_);
  and (_36505_, _36504_, _36498_);
  or (_36506_, _36505_, _06479_);
  or (_36507_, _36506_, _36503_);
  and (_36508_, _15134_, _07940_);
  or (_36509_, _36446_, _09043_);
  or (_36511_, _36509_, _36508_);
  and (_36512_, _36511_, _09048_);
  and (_36513_, _36512_, _36507_);
  nor (_36514_, _11215_, _13910_);
  or (_36515_, _36514_, _36446_);
  and (_36516_, _36515_, _06572_);
  or (_36517_, _36516_, _06606_);
  or (_36518_, _36517_, _36513_);
  or (_36519_, _36451_, _07037_);
  and (_36520_, _36519_, _06196_);
  and (_36522_, _36520_, _36518_);
  and (_36523_, _15315_, _07940_);
  or (_36524_, _36523_, _36446_);
  and (_36525_, _36524_, _06195_);
  or (_36526_, _36525_, _01379_);
  or (_36527_, _36526_, _36522_);
  or (_36528_, _01375_, \uc8051golden_1.SBUF [4]);
  and (_36529_, _36528_, _42545_);
  and (_43061_, _36529_, _36527_);
  and (_36530_, _13910_, \uc8051golden_1.SBUF [5]);
  nor (_36532_, _13910_, _08207_);
  or (_36533_, _36532_, _36530_);
  or (_36534_, _36533_, _06293_);
  and (_36535_, _15348_, _07940_);
  or (_36536_, _36535_, _36530_);
  or (_36537_, _36536_, _07210_);
  and (_36538_, _07940_, \uc8051golden_1.ACC [5]);
  or (_36539_, _36538_, _36530_);
  and (_36540_, _36539_, _07199_);
  and (_36541_, _07200_, \uc8051golden_1.SBUF [5]);
  or (_36543_, _36541_, _06401_);
  or (_36544_, _36543_, _36540_);
  and (_36545_, _36544_, _07221_);
  and (_36546_, _36545_, _36537_);
  and (_36547_, _36533_, _06399_);
  or (_36548_, _36547_, _36546_);
  and (_36549_, _36548_, _06414_);
  and (_36550_, _36539_, _06406_);
  or (_36551_, _36550_, _10059_);
  or (_36552_, _36551_, _36549_);
  and (_36554_, _36552_, _36534_);
  or (_36555_, _36554_, _06281_);
  and (_36556_, _07940_, _09441_);
  or (_36557_, _36530_, _06282_);
  or (_36558_, _36557_, _36556_);
  and (_36559_, _36558_, _06279_);
  and (_36560_, _36559_, _36555_);
  and (_36561_, _15446_, _07940_);
  or (_36562_, _36561_, _36530_);
  and (_36563_, _36562_, _06015_);
  or (_36565_, _36563_, _06275_);
  or (_36566_, _36565_, _36560_);
  and (_36567_, _08958_, _07940_);
  or (_36568_, _36567_, _36530_);
  or (_36569_, _36568_, _06276_);
  and (_36570_, _36569_, _36566_);
  or (_36571_, _36570_, _06474_);
  and (_36572_, _15338_, _07940_);
  or (_36573_, _36572_, _36530_);
  or (_36574_, _36573_, _07282_);
  and (_36576_, _36574_, _07284_);
  and (_36577_, _36576_, _36571_);
  and (_36578_, _12542_, _07940_);
  or (_36579_, _36578_, _36530_);
  and (_36580_, _36579_, _06582_);
  or (_36581_, _36580_, _36577_);
  and (_36582_, _36581_, _07279_);
  or (_36583_, _36530_, _08256_);
  and (_36584_, _36568_, _06478_);
  and (_36585_, _36584_, _36583_);
  or (_36587_, _36585_, _36582_);
  and (_36588_, _36587_, _07276_);
  and (_36589_, _36539_, _06569_);
  and (_36590_, _36589_, _36583_);
  or (_36591_, _36590_, _06479_);
  or (_36592_, _36591_, _36588_);
  and (_36593_, _15335_, _07940_);
  or (_36594_, _36530_, _09043_);
  or (_36595_, _36594_, _36593_);
  and (_36596_, _36595_, _09048_);
  and (_36598_, _36596_, _36592_);
  nor (_36599_, _11212_, _13910_);
  or (_36600_, _36599_, _36530_);
  and (_36601_, _36600_, _06572_);
  or (_36602_, _36601_, _06606_);
  or (_36603_, _36602_, _36598_);
  or (_36604_, _36536_, _07037_);
  and (_36605_, _36604_, _06196_);
  and (_36606_, _36605_, _36603_);
  and (_36607_, _15509_, _07940_);
  or (_36609_, _36607_, _36530_);
  and (_36610_, _36609_, _06195_);
  or (_36611_, _36610_, _01379_);
  or (_36612_, _36611_, _36606_);
  or (_36613_, _01375_, \uc8051golden_1.SBUF [5]);
  and (_36614_, _36613_, _42545_);
  and (_43062_, _36614_, _36612_);
  and (_36615_, _13910_, \uc8051golden_1.SBUF [6]);
  and (_36616_, _15531_, _07940_);
  or (_36617_, _36616_, _36615_);
  and (_36619_, _36617_, _06474_);
  and (_36620_, _15550_, _07940_);
  or (_36621_, _36620_, _36615_);
  or (_36622_, _36621_, _07210_);
  and (_36623_, _07940_, \uc8051golden_1.ACC [6]);
  or (_36624_, _36623_, _36615_);
  and (_36625_, _36624_, _07199_);
  and (_36626_, _07200_, \uc8051golden_1.SBUF [6]);
  or (_36627_, _36626_, _06401_);
  or (_36628_, _36627_, _36625_);
  and (_36630_, _36628_, _07221_);
  and (_36631_, _36630_, _36622_);
  nor (_36632_, _13910_, _08118_);
  or (_36633_, _36632_, _36615_);
  and (_36634_, _36633_, _06399_);
  or (_36635_, _36634_, _36631_);
  and (_36636_, _36635_, _06414_);
  and (_36637_, _36624_, _06406_);
  or (_36638_, _36637_, _10059_);
  or (_36639_, _36638_, _36636_);
  and (_36641_, _36633_, _06282_);
  or (_36642_, _36641_, _06294_);
  and (_36643_, _36642_, _36639_);
  and (_36644_, _07940_, _09440_);
  or (_36645_, _36644_, _36615_);
  and (_36646_, _36645_, _06281_);
  or (_36647_, _36646_, _06015_);
  or (_36648_, _36647_, _36643_);
  and (_36649_, _15639_, _07940_);
  or (_36650_, _36649_, _36615_);
  or (_36652_, _36650_, _06279_);
  and (_36653_, _36652_, _36648_);
  or (_36654_, _36653_, _06275_);
  and (_36655_, _15646_, _07940_);
  or (_36656_, _36655_, _36615_);
  or (_36657_, _36656_, _06276_);
  and (_36658_, _36657_, _07282_);
  and (_36659_, _36658_, _36654_);
  or (_36660_, _36659_, _36619_);
  and (_36661_, _36660_, _07284_);
  and (_36663_, _11210_, _07940_);
  or (_36664_, _36663_, _36615_);
  and (_36665_, _36664_, _06582_);
  or (_36666_, _36665_, _36661_);
  and (_36667_, _36666_, _07279_);
  or (_36668_, _36615_, _08162_);
  and (_36669_, _36656_, _06478_);
  and (_36670_, _36669_, _36668_);
  or (_36671_, _36670_, _36667_);
  and (_36672_, _36671_, _07276_);
  and (_36674_, _36624_, _06569_);
  and (_36675_, _36674_, _36668_);
  or (_36676_, _36675_, _06479_);
  or (_36677_, _36676_, _36672_);
  and (_36678_, _15528_, _07940_);
  or (_36679_, _36615_, _09043_);
  or (_36680_, _36679_, _36678_);
  and (_36681_, _36680_, _09048_);
  and (_36682_, _36681_, _36677_);
  nor (_36683_, _11209_, _13910_);
  or (_36685_, _36683_, _36615_);
  and (_36686_, _36685_, _06572_);
  or (_36687_, _36686_, _06606_);
  or (_36688_, _36687_, _36682_);
  or (_36689_, _36621_, _07037_);
  and (_36690_, _36689_, _06196_);
  and (_36691_, _36690_, _36688_);
  and (_36692_, _15713_, _07940_);
  or (_36693_, _36692_, _36615_);
  and (_36694_, _36693_, _06195_);
  or (_36696_, _36694_, _01379_);
  or (_36697_, _36696_, _36691_);
  or (_36698_, _01375_, \uc8051golden_1.SBUF [6]);
  and (_36699_, _36698_, _42545_);
  and (_43063_, _36699_, _36697_);
  not (_36700_, \uc8051golden_1.PSW [0]);
  nor (_36701_, _01375_, _36700_);
  nand (_36702_, _11225_, _07988_);
  nor (_36703_, _07988_, _36700_);
  nor (_36704_, _36703_, _07276_);
  nand (_36706_, _36704_, _36702_);
  and (_36707_, _07988_, _07473_);
  or (_36708_, _36707_, _36703_);
  or (_36709_, _36708_, _06293_);
  nor (_36710_, _08521_, _13994_);
  or (_36711_, _36710_, _36703_);
  or (_36712_, _36711_, _07210_);
  and (_36713_, _07988_, \uc8051golden_1.ACC [0]);
  or (_36714_, _36713_, _36703_);
  and (_36715_, _36714_, _07199_);
  nor (_36717_, _07199_, _36700_);
  or (_36718_, _36717_, _06401_);
  or (_36719_, _36718_, _36715_);
  and (_36720_, _36719_, _06396_);
  and (_36721_, _36720_, _36712_);
  nor (_36722_, _08612_, _36700_);
  and (_36723_, _14339_, _08612_);
  or (_36724_, _36723_, _36722_);
  and (_36725_, _36724_, _06395_);
  or (_36726_, _36725_, _36721_);
  and (_36728_, _36726_, _07221_);
  and (_36729_, _36708_, _06399_);
  or (_36730_, _36729_, _06406_);
  or (_36731_, _36730_, _36728_);
  or (_36732_, _36714_, _06414_);
  and (_36733_, _36732_, _06844_);
  and (_36734_, _36733_, _36731_);
  and (_36735_, _36703_, _06393_);
  or (_36736_, _36735_, _06387_);
  or (_36737_, _36736_, _36734_);
  or (_36739_, _36711_, _07245_);
  and (_36740_, _36739_, _06446_);
  and (_36741_, _36740_, _36737_);
  and (_36742_, _14371_, _08612_);
  or (_36743_, _36742_, _36722_);
  and (_36744_, _36743_, _06300_);
  or (_36745_, _36744_, _10059_);
  or (_36746_, _36745_, _36741_);
  and (_36747_, _36746_, _36709_);
  or (_36748_, _36747_, _06281_);
  and (_36750_, _07988_, _09446_);
  or (_36751_, _36703_, _06282_);
  or (_36752_, _36751_, _36750_);
  and (_36753_, _36752_, _36748_);
  or (_36754_, _36753_, _06015_);
  and (_36755_, _14426_, _07988_);
  or (_36756_, _36703_, _06279_);
  or (_36757_, _36756_, _36755_);
  and (_36758_, _36757_, _06276_);
  and (_36759_, _36758_, _36754_);
  and (_36761_, _07988_, _08817_);
  or (_36762_, _36761_, _36703_);
  and (_36763_, _36762_, _06275_);
  or (_36764_, _36763_, _06474_);
  or (_36765_, _36764_, _36759_);
  and (_36766_, _14324_, _07988_);
  or (_36767_, _36766_, _36703_);
  or (_36768_, _36767_, _07282_);
  and (_36769_, _36768_, _07284_);
  and (_36770_, _36769_, _36765_);
  nor (_36772_, _12538_, _13994_);
  or (_36773_, _36772_, _36703_);
  and (_36774_, _36702_, _06582_);
  and (_36775_, _36774_, _36773_);
  or (_36776_, _36775_, _36770_);
  and (_36777_, _36776_, _07279_);
  nand (_36778_, _36762_, _06478_);
  nor (_36779_, _36778_, _36710_);
  or (_36780_, _36779_, _06569_);
  or (_36781_, _36780_, _36777_);
  and (_36783_, _36781_, _36706_);
  or (_36784_, _36783_, _06479_);
  and (_36785_, _14320_, _07988_);
  or (_36786_, _36703_, _09043_);
  or (_36787_, _36786_, _36785_);
  and (_36788_, _36787_, _09048_);
  and (_36789_, _36788_, _36784_);
  and (_36790_, _36773_, _06572_);
  or (_36791_, _36790_, _06606_);
  or (_36792_, _36791_, _36789_);
  or (_36794_, _36711_, _07037_);
  and (_36795_, _36794_, _36792_);
  or (_36796_, _36795_, _06234_);
  or (_36797_, _36703_, _06807_);
  and (_36798_, _36797_, _36796_);
  or (_36799_, _36798_, _06195_);
  or (_36800_, _36711_, _06196_);
  and (_36801_, _36800_, _01375_);
  and (_36802_, _36801_, _36799_);
  or (_36803_, _36802_, _36701_);
  and (_43065_, _36803_, _42545_);
  not (_36805_, \uc8051golden_1.PSW [1]);
  nor (_36806_, _01375_, _36805_);
  nor (_36807_, _07988_, _36805_);
  nor (_36808_, _11223_, _13994_);
  or (_36809_, _36808_, _36807_);
  or (_36810_, _36809_, _09048_);
  nor (_36811_, _13994_, _07196_);
  or (_36812_, _36811_, _36807_);
  or (_36813_, _36812_, _06293_);
  or (_36815_, _36812_, _07221_);
  or (_36816_, _07988_, \uc8051golden_1.PSW [1]);
  and (_36817_, _14532_, _07988_);
  not (_36818_, _36817_);
  and (_36819_, _36818_, _36816_);
  or (_36820_, _36819_, _07210_);
  and (_36821_, _07988_, \uc8051golden_1.ACC [1]);
  or (_36822_, _36821_, _36807_);
  and (_36823_, _36822_, _07199_);
  nor (_36824_, _07199_, _36805_);
  or (_36826_, _36824_, _06401_);
  or (_36827_, _36826_, _36823_);
  and (_36828_, _36827_, _06396_);
  and (_36829_, _36828_, _36820_);
  nor (_36830_, _08612_, _36805_);
  and (_36831_, _14514_, _08612_);
  or (_36832_, _36831_, _36830_);
  and (_36833_, _36832_, _06395_);
  or (_36834_, _36833_, _06399_);
  or (_36835_, _36834_, _36829_);
  and (_36837_, _36835_, _36815_);
  or (_36838_, _36837_, _06406_);
  or (_36839_, _36822_, _06414_);
  and (_36840_, _36839_, _06844_);
  and (_36841_, _36840_, _36838_);
  and (_36842_, _14517_, _08612_);
  or (_36843_, _36842_, _36830_);
  and (_36844_, _36843_, _06393_);
  or (_36845_, _36844_, _06387_);
  or (_36846_, _36845_, _36841_);
  and (_36848_, _36831_, _14513_);
  or (_36849_, _36830_, _07245_);
  or (_36850_, _36849_, _36848_);
  and (_36851_, _36850_, _06446_);
  and (_36852_, _36851_, _36846_);
  or (_36853_, _36830_, _14560_);
  and (_36854_, _36853_, _06300_);
  and (_36855_, _36854_, _36832_);
  or (_36856_, _36855_, _10059_);
  or (_36857_, _36856_, _36852_);
  and (_36859_, _36857_, _36813_);
  or (_36860_, _36859_, _06281_);
  and (_36861_, _07988_, _09445_);
  or (_36862_, _36807_, _06282_);
  or (_36863_, _36862_, _36861_);
  and (_36864_, _36863_, _06279_);
  and (_36865_, _36864_, _36860_);
  or (_36866_, _14615_, _13994_);
  and (_36867_, _36816_, _06015_);
  and (_36868_, _36867_, _36866_);
  or (_36869_, _36868_, _36865_);
  and (_36870_, _36869_, _06276_);
  nand (_36871_, _07988_, _07090_);
  and (_36872_, _36816_, _06275_);
  and (_36873_, _36872_, _36871_);
  or (_36874_, _36873_, _36870_);
  and (_36875_, _36874_, _07282_);
  or (_36876_, _14507_, _13994_);
  and (_36877_, _36816_, _06474_);
  and (_36878_, _36877_, _36876_);
  or (_36880_, _36878_, _06582_);
  or (_36881_, _36880_, _36875_);
  nand (_36882_, _11222_, _07988_);
  and (_36883_, _36882_, _36809_);
  or (_36884_, _36883_, _07284_);
  and (_36885_, _36884_, _07279_);
  and (_36886_, _36885_, _36881_);
  or (_36887_, _14505_, _13994_);
  and (_36888_, _36816_, _06478_);
  and (_36889_, _36888_, _36887_);
  or (_36891_, _36889_, _06569_);
  or (_36892_, _36891_, _36886_);
  nor (_36893_, _36807_, _07276_);
  nand (_36894_, _36893_, _36882_);
  and (_36895_, _36894_, _09043_);
  and (_36896_, _36895_, _36892_);
  or (_36897_, _36871_, _08477_);
  and (_36898_, _36816_, _06479_);
  and (_36899_, _36898_, _36897_);
  or (_36900_, _36899_, _06572_);
  or (_36902_, _36900_, _36896_);
  and (_36903_, _36902_, _36810_);
  or (_36904_, _36903_, _06606_);
  or (_36905_, _36819_, _07037_);
  and (_36906_, _36905_, _06807_);
  and (_36907_, _36906_, _36904_);
  and (_36908_, _36843_, _06234_);
  or (_36909_, _36908_, _06195_);
  or (_36910_, _36909_, _36907_);
  or (_36911_, _36807_, _06196_);
  or (_36913_, _36911_, _36817_);
  and (_36914_, _36913_, _01375_);
  and (_36915_, _36914_, _36910_);
  or (_36916_, _36915_, _36806_);
  and (_43066_, _36916_, _42545_);
  and (_36917_, _01379_, \uc8051golden_1.PSW [2]);
  or (_36918_, _11157_, _10549_);
  nand (_36919_, _14269_, _11156_);
  and (_36920_, _36919_, _36918_);
  and (_36921_, _36920_, _11121_);
  and (_36923_, _13994_, \uc8051golden_1.PSW [2]);
  and (_36924_, _14744_, _07988_);
  or (_36925_, _36924_, _36923_);
  and (_36926_, _36925_, _06474_);
  nor (_36927_, _13994_, _07623_);
  or (_36928_, _36927_, _36923_);
  or (_36929_, _36928_, _06293_);
  and (_36930_, _36928_, _06399_);
  not (_36931_, _08612_);
  and (_36932_, _36931_, \uc8051golden_1.PSW [2]);
  and (_36934_, _14751_, _08612_);
  or (_36935_, _36934_, _36932_);
  or (_36936_, _36935_, _06396_);
  and (_36937_, _14754_, _07988_);
  or (_36938_, _36937_, _36923_);
  and (_36939_, _36938_, _06401_);
  and (_36940_, _07200_, \uc8051golden_1.PSW [2]);
  and (_36941_, _07988_, \uc8051golden_1.ACC [2]);
  or (_36942_, _36941_, _36923_);
  and (_36943_, _36942_, _07199_);
  or (_36945_, _36943_, _36940_);
  and (_36946_, _36945_, _07210_);
  or (_36947_, _36946_, _06395_);
  or (_36948_, _36947_, _36939_);
  and (_36949_, _36948_, _36936_);
  and (_36950_, _36949_, _07221_);
  or (_36951_, _36950_, _36930_);
  or (_36952_, _36951_, _06406_);
  or (_36953_, _36942_, _06414_);
  and (_36954_, _36953_, _06844_);
  and (_36956_, _36954_, _36952_);
  and (_36957_, _14749_, _08612_);
  or (_36958_, _36957_, _36932_);
  and (_36959_, _36958_, _06393_);
  or (_36960_, _36959_, _36956_);
  and (_36961_, _36960_, _07245_);
  or (_36962_, _36932_, _14778_);
  and (_36963_, _36935_, _06387_);
  and (_36964_, _36963_, _36962_);
  or (_36965_, _36964_, _36961_);
  and (_36967_, _36965_, _09544_);
  or (_36968_, _16568_, _16457_);
  or (_36969_, _36968_, _16680_);
  or (_36970_, _36969_, _16798_);
  or (_36971_, _36970_, _16916_);
  or (_36972_, _36971_, _17032_);
  or (_36973_, _36972_, _10055_);
  or (_36974_, _36973_, _17152_);
  and (_36975_, _36974_, _09538_);
  or (_36976_, _36975_, _14157_);
  or (_36978_, _36976_, _36967_);
  not (_36979_, _10809_);
  or (_36980_, _10743_, _08070_);
  nor (_36981_, _36980_, _08651_);
  and (_36982_, _36980_, _08651_);
  or (_36983_, _36982_, _36981_);
  and (_36984_, _36983_, _14166_);
  nor (_36985_, _36983_, _14166_);
  nor (_36986_, _36985_, _36984_);
  nor (_36987_, _36986_, _36979_);
  and (_36989_, _36986_, _36979_);
  or (_36990_, _36989_, _36987_);
  or (_36991_, _36990_, _10740_);
  and (_36992_, _36991_, _36978_);
  and (_36993_, _36992_, _12587_);
  nor (_36994_, _14275_, _14176_);
  nor (_36995_, _10474_, \uc8051golden_1.ACC [7]);
  or (_36996_, _36995_, _36994_);
  or (_36997_, _36996_, _14175_);
  nand (_36998_, _36996_, _14175_);
  and (_37000_, _36998_, _36997_);
  and (_37001_, _37000_, _10833_);
  nor (_37002_, _37000_, _10833_);
  or (_37003_, _37002_, _37001_);
  and (_37004_, _37003_, _12586_);
  or (_37005_, _37004_, _36993_);
  and (_37006_, _37005_, _06442_);
  nor (_37007_, _10581_, \uc8051golden_1.ACC [7]);
  nor (_37008_, _10580_, _14282_);
  nor (_37009_, _37008_, _37007_);
  nor (_37011_, _37009_, _10586_);
  nor (_37012_, _14012_, _10582_);
  or (_37013_, _37012_, _37011_);
  nand (_37014_, _37013_, _10635_);
  or (_37015_, _37013_, _10635_);
  and (_37016_, _37015_, _06437_);
  and (_37017_, _37016_, _37014_);
  or (_37018_, _37017_, _10572_);
  or (_37019_, _37018_, _37006_);
  nor (_37020_, _10844_, _14288_);
  nor (_37022_, _10846_, \uc8051golden_1.ACC [7]);
  nor (_37023_, _37022_, _37020_);
  not (_37024_, _37023_);
  or (_37025_, _37024_, _14189_);
  nand (_37026_, _37024_, _14189_);
  and (_37027_, _37026_, _37025_);
  and (_37028_, _37027_, _10904_);
  nor (_37029_, _37027_, _10904_);
  or (_37030_, _37029_, _37028_);
  or (_37031_, _37030_, _10573_);
  and (_37033_, _37031_, _06446_);
  and (_37034_, _37033_, _37019_);
  and (_37035_, _14793_, _08612_);
  or (_37036_, _37035_, _36932_);
  and (_37037_, _37036_, _06300_);
  or (_37038_, _37037_, _10059_);
  or (_37039_, _37038_, _37034_);
  and (_37040_, _37039_, _36929_);
  or (_37041_, _37040_, _06281_);
  and (_37042_, _07988_, _09444_);
  or (_37044_, _36923_, _06282_);
  or (_37045_, _37044_, _37042_);
  and (_37046_, _37045_, _06279_);
  and (_37047_, _37046_, _37041_);
  and (_37048_, _14848_, _07988_);
  or (_37049_, _37048_, _36923_);
  and (_37050_, _37049_, _06015_);
  or (_37051_, _37050_, _10072_);
  or (_37052_, _37051_, _37047_);
  nor (_37053_, \uc8051golden_1.B [1], \uc8051golden_1.B [0]);
  nand (_37055_, _37053_, _10100_);
  nand (_37056_, _37055_, _10072_);
  and (_37057_, _37056_, _37052_);
  or (_37058_, _37057_, _06275_);
  and (_37059_, _07988_, _08994_);
  or (_37060_, _37059_, _36923_);
  or (_37061_, _37060_, _06276_);
  and (_37062_, _37061_, _07282_);
  and (_37063_, _37062_, _37058_);
  or (_37064_, _37063_, _36926_);
  and (_37066_, _37064_, _07284_);
  and (_37067_, _11221_, _07988_);
  or (_37068_, _37067_, _36923_);
  and (_37069_, _37068_, _06582_);
  or (_37070_, _37069_, _37066_);
  and (_37071_, _37070_, _07279_);
  or (_37072_, _36923_, _08433_);
  and (_37073_, _37060_, _06478_);
  and (_37074_, _37073_, _37072_);
  or (_37075_, _37074_, _37071_);
  and (_37077_, _37075_, _07276_);
  and (_37078_, _36942_, _06569_);
  and (_37079_, _37078_, _37072_);
  or (_37080_, _37079_, _06479_);
  or (_37081_, _37080_, _37077_);
  and (_37082_, _14741_, _07988_);
  or (_37083_, _37082_, _36923_);
  or (_37084_, _37083_, _09043_);
  and (_37085_, _37084_, _09048_);
  and (_37086_, _37085_, _37081_);
  nor (_37088_, _11220_, _13994_);
  or (_37089_, _37088_, _36923_);
  and (_37090_, _37089_, _06572_);
  or (_37091_, _37090_, _11030_);
  or (_37092_, _37091_, _37086_);
  nor (_37093_, _36983_, _14241_);
  nor (_37094_, _37093_, _36981_);
  and (_37095_, _37094_, _11054_);
  and (_37096_, _36981_, _11051_);
  or (_37097_, _37096_, _11028_);
  or (_37099_, _37097_, _37095_);
  and (_37100_, _37099_, _37092_);
  or (_37101_, _37100_, _10471_);
  nor (_37102_, _36996_, _14247_);
  nor (_37103_, _37102_, _36994_);
  or (_37104_, _37103_, _10472_);
  and (_37105_, _37104_, _10544_);
  and (_37106_, _36994_, _06579_);
  and (_37107_, _37106_, _10539_);
  or (_37108_, _37107_, _37105_);
  and (_37110_, _37108_, _37101_);
  not (_37111_, _37009_);
  nor (_37112_, _37111_, _14253_);
  nor (_37113_, _37112_, _37008_);
  and (_37114_, _37113_, _11085_);
  and (_37115_, _37008_, _11082_);
  or (_37116_, _37115_, _37114_);
  and (_37117_, _37116_, _06578_);
  or (_37118_, _37117_, _11059_);
  or (_37119_, _37118_, _37110_);
  nor (_37121_, _37024_, _14259_);
  nor (_37122_, _37121_, _37020_);
  and (_37123_, _37122_, _11115_);
  and (_37124_, _37020_, _11112_);
  or (_37125_, _37124_, _37123_);
  or (_37126_, _37125_, _11091_);
  and (_37127_, _37126_, _11120_);
  and (_37128_, _37127_, _37119_);
  or (_37129_, _37128_, _36921_);
  and (_37130_, _37129_, _11165_);
  nand (_37132_, _11198_, _14275_);
  and (_37133_, _37132_, _14277_);
  or (_37134_, _37133_, _37130_);
  and (_37135_, _37134_, _11204_);
  or (_37136_, _11238_, _09033_);
  and (_37137_, _14284_, _37136_);
  nand (_37138_, _11274_, _14288_);
  and (_37139_, _37138_, _14291_);
  or (_37140_, _37139_, _06606_);
  or (_37141_, _37140_, _37137_);
  or (_37143_, _37141_, _37135_);
  or (_37144_, _36938_, _07037_);
  and (_37145_, _37144_, _06807_);
  and (_37146_, _37145_, _37143_);
  and (_37147_, _36958_, _06234_);
  or (_37148_, _37147_, _06195_);
  or (_37149_, _37148_, _37146_);
  and (_37150_, _14917_, _07988_);
  or (_37151_, _36923_, _06196_);
  or (_37152_, _37151_, _37150_);
  and (_37154_, _37152_, _01375_);
  and (_37155_, _37154_, _37149_);
  or (_37156_, _37155_, _36917_);
  and (_43067_, _37156_, _42545_);
  nor (_37157_, _01375_, _07789_);
  nor (_37158_, _07988_, _07789_);
  nor (_37159_, _13994_, _07775_);
  or (_37160_, _37159_, _37158_);
  or (_37161_, _37160_, _06293_);
  and (_37162_, _14947_, _07988_);
  or (_37164_, _37162_, _37158_);
  or (_37165_, _37164_, _07210_);
  and (_37166_, _07988_, \uc8051golden_1.ACC [3]);
  or (_37167_, _37166_, _37158_);
  and (_37168_, _37167_, _07199_);
  nor (_37169_, _07199_, _07789_);
  or (_37170_, _37169_, _06401_);
  or (_37171_, _37170_, _37168_);
  and (_37172_, _37171_, _06396_);
  and (_37173_, _37172_, _37165_);
  nor (_37175_, _08612_, _07789_);
  and (_37176_, _14951_, _08612_);
  or (_37177_, _37176_, _37175_);
  and (_37178_, _37177_, _06395_);
  or (_37179_, _37178_, _06399_);
  or (_37180_, _37179_, _37173_);
  or (_37181_, _37160_, _07221_);
  and (_37182_, _37181_, _37180_);
  or (_37183_, _37182_, _06406_);
  or (_37184_, _37167_, _06414_);
  and (_37186_, _37184_, _06844_);
  and (_37187_, _37186_, _37183_);
  and (_37188_, _14961_, _08612_);
  or (_37189_, _37188_, _37175_);
  and (_37190_, _37189_, _06393_);
  or (_37191_, _37190_, _06387_);
  or (_37192_, _37191_, _37187_);
  or (_37193_, _37175_, _14968_);
  and (_37194_, _37193_, _37177_);
  or (_37195_, _37194_, _07245_);
  and (_37197_, _37195_, _06446_);
  and (_37198_, _37197_, _37192_);
  and (_37199_, _14985_, _08612_);
  or (_37200_, _37199_, _37175_);
  and (_37201_, _37200_, _06300_);
  or (_37202_, _37201_, _10059_);
  or (_37203_, _37202_, _37198_);
  and (_37204_, _37203_, _37161_);
  or (_37205_, _37204_, _06281_);
  and (_37206_, _07988_, _09443_);
  or (_37208_, _37158_, _06282_);
  or (_37209_, _37208_, _37206_);
  and (_37210_, _37209_, _37205_);
  or (_37211_, _37210_, _06015_);
  and (_37212_, _15039_, _07988_);
  or (_37213_, _37158_, _06279_);
  or (_37214_, _37213_, _37212_);
  and (_37215_, _37214_, _06276_);
  and (_37216_, _37215_, _37211_);
  and (_37217_, _07988_, _08815_);
  or (_37219_, _37217_, _37158_);
  and (_37220_, _37219_, _06275_);
  or (_37221_, _37220_, _06474_);
  or (_37222_, _37221_, _37216_);
  and (_37223_, _14934_, _07988_);
  or (_37224_, _37223_, _37158_);
  or (_37225_, _37224_, _07282_);
  and (_37226_, _37225_, _07284_);
  and (_37227_, _37226_, _37222_);
  and (_37228_, _12535_, _07988_);
  or (_37230_, _37228_, _37158_);
  and (_37231_, _37230_, _06582_);
  or (_37232_, _37231_, _37227_);
  and (_37233_, _37232_, _07279_);
  or (_37234_, _37158_, _08389_);
  and (_37235_, _37219_, _06478_);
  and (_37236_, _37235_, _37234_);
  or (_37237_, _37236_, _37233_);
  and (_37238_, _37237_, _07276_);
  and (_37239_, _37167_, _06569_);
  and (_37241_, _37239_, _37234_);
  or (_37242_, _37241_, _06479_);
  or (_37243_, _37242_, _37238_);
  and (_37244_, _14931_, _07988_);
  or (_37245_, _37158_, _09043_);
  or (_37246_, _37245_, _37244_);
  and (_37247_, _37246_, _09048_);
  and (_37248_, _37247_, _37243_);
  nor (_37249_, _11218_, _13994_);
  or (_37250_, _37249_, _37158_);
  and (_37252_, _37250_, _06572_);
  or (_37253_, _37252_, _06606_);
  or (_37254_, _37253_, _37248_);
  or (_37255_, _37164_, _07037_);
  and (_37256_, _37255_, _06807_);
  and (_37257_, _37256_, _37254_);
  and (_37258_, _37189_, _06234_);
  or (_37259_, _37258_, _06195_);
  or (_37260_, _37259_, _37257_);
  and (_37261_, _15113_, _07988_);
  or (_37263_, _37158_, _06196_);
  or (_37264_, _37263_, _37261_);
  and (_37265_, _37264_, _01375_);
  and (_37266_, _37265_, _37260_);
  or (_37267_, _37266_, _37157_);
  and (_43068_, _37267_, _42545_);
  and (_37268_, _01379_, \uc8051golden_1.PSW [4]);
  and (_37269_, _36931_, \uc8051golden_1.PSW [4]);
  and (_37270_, _15168_, _08612_);
  or (_37271_, _37270_, _37269_);
  and (_37273_, _37271_, _06393_);
  and (_37274_, _13994_, \uc8051golden_1.PSW [4]);
  and (_37275_, _15130_, _07988_);
  or (_37276_, _37275_, _37274_);
  or (_37277_, _37276_, _07210_);
  and (_37278_, _07988_, \uc8051golden_1.ACC [4]);
  or (_37279_, _37278_, _37274_);
  and (_37280_, _37279_, _07199_);
  and (_37281_, _07200_, \uc8051golden_1.PSW [4]);
  or (_37282_, _37281_, _06401_);
  or (_37284_, _37282_, _37280_);
  and (_37285_, _37284_, _06396_);
  and (_37286_, _37285_, _37277_);
  and (_37287_, _15139_, _08612_);
  or (_37288_, _37287_, _37269_);
  and (_37289_, _37288_, _06395_);
  or (_37290_, _37289_, _06399_);
  or (_37291_, _37290_, _37286_);
  nor (_37292_, _13994_, _08301_);
  or (_37293_, _37292_, _37274_);
  or (_37295_, _37293_, _07221_);
  and (_37296_, _37295_, _37291_);
  or (_37297_, _37296_, _06406_);
  or (_37298_, _37279_, _06414_);
  and (_37299_, _37298_, _06844_);
  and (_37300_, _37299_, _37297_);
  or (_37301_, _37300_, _37273_);
  and (_37302_, _37301_, _07245_);
  or (_37303_, _37269_, _15138_);
  and (_37304_, _37303_, _06387_);
  and (_37306_, _37304_, _37288_);
  or (_37307_, _37306_, _37302_);
  and (_37308_, _37307_, _06446_);
  and (_37309_, _15189_, _08612_);
  or (_37310_, _37309_, _37269_);
  and (_37311_, _37310_, _06300_);
  or (_37312_, _37311_, _10059_);
  or (_37313_, _37312_, _37308_);
  or (_37314_, _37293_, _06293_);
  nand (_37315_, _37314_, _37313_);
  nor (_37317_, _37315_, _25765_);
  and (_37318_, _07988_, _09442_);
  or (_37319_, _37318_, _37274_);
  and (_37320_, _37319_, _25765_);
  or (_37321_, _37320_, _37317_);
  and (_37322_, _37321_, _25764_);
  and (_37323_, _37319_, _25763_);
  or (_37324_, _37323_, _06015_);
  or (_37325_, _37324_, _37322_);
  and (_37326_, _15243_, _07988_);
  or (_37328_, _37326_, _37274_);
  or (_37329_, _37328_, _06279_);
  and (_37330_, _37329_, _37325_);
  or (_37331_, _37330_, _06275_);
  and (_37332_, _08883_, _07988_);
  or (_37333_, _37332_, _37274_);
  or (_37334_, _37333_, _06276_);
  and (_37335_, _37334_, _07282_);
  and (_37336_, _37335_, _37331_);
  and (_37337_, _15135_, _07988_);
  or (_37339_, _37337_, _37274_);
  and (_37340_, _37339_, _06474_);
  or (_37341_, _37340_, _37336_);
  and (_37342_, _37341_, _07284_);
  and (_37343_, _11216_, _07988_);
  or (_37344_, _37343_, _37274_);
  and (_37345_, _37344_, _06582_);
  or (_37346_, _37345_, _37342_);
  and (_37347_, _37346_, _07279_);
  or (_37348_, _37274_, _08345_);
  and (_37350_, _37333_, _06478_);
  and (_37351_, _37350_, _37348_);
  or (_37352_, _37351_, _37347_);
  and (_37353_, _37352_, _07276_);
  and (_37354_, _37279_, _06569_);
  and (_37355_, _37354_, _37348_);
  or (_37356_, _37355_, _06479_);
  or (_37357_, _37356_, _37353_);
  and (_37358_, _15134_, _07988_);
  or (_37359_, _37274_, _09043_);
  or (_37361_, _37359_, _37358_);
  and (_37362_, _37361_, _09048_);
  and (_37363_, _37362_, _37357_);
  nor (_37364_, _11215_, _13994_);
  or (_37365_, _37364_, _37274_);
  and (_37366_, _37365_, _06572_);
  or (_37367_, _37366_, _06606_);
  or (_37368_, _37367_, _37363_);
  or (_37369_, _37276_, _07037_);
  and (_37370_, _37369_, _06807_);
  and (_37372_, _37370_, _37368_);
  and (_37373_, _37271_, _06234_);
  or (_37374_, _37373_, _06195_);
  or (_37375_, _37374_, _37372_);
  and (_37376_, _15315_, _07988_);
  or (_37377_, _37274_, _06196_);
  or (_37378_, _37377_, _37376_);
  and (_37379_, _37378_, _01375_);
  and (_37380_, _37379_, _37375_);
  or (_37381_, _37380_, _37268_);
  and (_43069_, _37381_, _42545_);
  and (_37383_, _01379_, \uc8051golden_1.PSW [5]);
  and (_37384_, _13994_, \uc8051golden_1.PSW [5]);
  and (_37385_, _15348_, _07988_);
  or (_37386_, _37385_, _37384_);
  or (_37387_, _37386_, _07210_);
  and (_37388_, _07988_, \uc8051golden_1.ACC [5]);
  or (_37389_, _37388_, _37384_);
  and (_37390_, _37389_, _07199_);
  and (_37391_, _07200_, \uc8051golden_1.PSW [5]);
  or (_37393_, _37391_, _06401_);
  or (_37394_, _37393_, _37390_);
  and (_37395_, _37394_, _06396_);
  and (_37396_, _37395_, _37387_);
  and (_37397_, _36931_, \uc8051golden_1.PSW [5]);
  and (_37398_, _15341_, _08612_);
  or (_37399_, _37398_, _37397_);
  and (_37400_, _37399_, _06395_);
  or (_37401_, _37400_, _06399_);
  or (_37402_, _37401_, _37396_);
  nor (_37404_, _13994_, _08207_);
  or (_37405_, _37404_, _37384_);
  or (_37406_, _37405_, _07221_);
  and (_37407_, _37406_, _37402_);
  or (_37408_, _37407_, _06406_);
  or (_37409_, _37389_, _06414_);
  and (_37410_, _37409_, _06844_);
  and (_37411_, _37410_, _37408_);
  and (_37412_, _15345_, _08612_);
  or (_37413_, _37412_, _37397_);
  and (_37415_, _37413_, _06393_);
  or (_37416_, _37415_, _06387_);
  or (_37417_, _37416_, _37411_);
  or (_37418_, _37397_, _15378_);
  and (_37419_, _37418_, _37399_);
  or (_37420_, _37419_, _07245_);
  and (_37421_, _37420_, _06446_);
  and (_37422_, _37421_, _37417_);
  or (_37423_, _37397_, _15342_);
  and (_37424_, _37423_, _06300_);
  and (_37426_, _37424_, _37399_);
  or (_37427_, _37426_, _10059_);
  or (_37428_, _37427_, _37422_);
  or (_37429_, _37405_, _06293_);
  and (_37430_, _37429_, _06282_);
  and (_37431_, _37430_, _37428_);
  and (_37432_, _07988_, _09441_);
  or (_37433_, _37432_, _37384_);
  and (_37434_, _37433_, _06281_);
  or (_37435_, _37434_, _06015_);
  or (_37437_, _37435_, _37431_);
  and (_37438_, _15446_, _07988_);
  or (_37439_, _37384_, _06279_);
  or (_37440_, _37439_, _37438_);
  and (_37441_, _37440_, _06276_);
  and (_37442_, _37441_, _37437_);
  and (_37443_, _08958_, _07988_);
  or (_37444_, _37443_, _37384_);
  and (_37445_, _37444_, _06275_);
  or (_37446_, _37445_, _06474_);
  or (_37448_, _37446_, _37442_);
  and (_37449_, _15338_, _07988_);
  or (_37450_, _37449_, _37384_);
  or (_37451_, _37450_, _07282_);
  and (_37452_, _37451_, _07284_);
  and (_37453_, _37452_, _37448_);
  and (_37454_, _12542_, _07988_);
  or (_37455_, _37454_, _37384_);
  and (_37456_, _37455_, _06582_);
  or (_37457_, _37456_, _37453_);
  and (_37459_, _37457_, _07279_);
  or (_37460_, _37384_, _08256_);
  and (_37461_, _37444_, _06478_);
  and (_37462_, _37461_, _37460_);
  or (_37463_, _37462_, _37459_);
  and (_37464_, _37463_, _07276_);
  and (_37465_, _37389_, _06569_);
  and (_37466_, _37465_, _37460_);
  or (_37467_, _37466_, _06479_);
  or (_37468_, _37467_, _37464_);
  and (_37470_, _15335_, _07988_);
  or (_37471_, _37384_, _09043_);
  or (_37472_, _37471_, _37470_);
  and (_37473_, _37472_, _09048_);
  and (_37474_, _37473_, _37468_);
  nor (_37475_, _11212_, _13994_);
  or (_37476_, _37475_, _37384_);
  and (_37477_, _37476_, _06572_);
  or (_37478_, _37477_, _06606_);
  or (_37479_, _37478_, _37474_);
  or (_37481_, _37386_, _07037_);
  and (_37482_, _37481_, _06807_);
  and (_37483_, _37482_, _37479_);
  and (_37484_, _37413_, _06234_);
  or (_37485_, _37484_, _06195_);
  or (_37486_, _37485_, _37483_);
  and (_37487_, _15509_, _07988_);
  or (_37488_, _37384_, _06196_);
  or (_37489_, _37488_, _37487_);
  and (_37490_, _37489_, _01375_);
  and (_37492_, _37490_, _37486_);
  or (_37493_, _37492_, _37383_);
  and (_43071_, _37493_, _42545_);
  nor (_37494_, _01375_, _18122_);
  or (_37495_, _11106_, _10842_);
  and (_37496_, _37495_, _11059_);
  and (_37497_, _06466_, _05965_);
  or (_37498_, _11045_, _10762_);
  nand (_37499_, _37498_, _37497_);
  nor (_37500_, _07988_, _18122_);
  nor (_37502_, _13994_, _08118_);
  or (_37503_, _37502_, _37500_);
  or (_37504_, _37503_, _06293_);
  or (_37505_, _10826_, _12587_);
  or (_37506_, _37505_, _10495_);
  nor (_37507_, _08612_, _18122_);
  and (_37508_, _15561_, _08612_);
  or (_37509_, _37508_, _37507_);
  and (_37510_, _37509_, _06393_);
  and (_37511_, _15550_, _07988_);
  or (_37513_, _37511_, _37500_);
  or (_37514_, _37513_, _07210_);
  and (_37515_, _07988_, \uc8051golden_1.ACC [6]);
  or (_37516_, _37515_, _37500_);
  and (_37517_, _37516_, _07199_);
  nor (_37518_, _07199_, _18122_);
  or (_37519_, _37518_, _06401_);
  or (_37520_, _37519_, _37517_);
  and (_37521_, _37520_, _06396_);
  and (_37522_, _37521_, _37514_);
  and (_37524_, _15535_, _08612_);
  or (_37525_, _37524_, _37507_);
  and (_37526_, _37525_, _06395_);
  or (_37527_, _37526_, _06399_);
  or (_37528_, _37527_, _37522_);
  or (_37529_, _37503_, _07221_);
  and (_37530_, _37529_, _37528_);
  or (_37531_, _37530_, _06406_);
  or (_37532_, _37516_, _06414_);
  and (_37533_, _37532_, _06844_);
  and (_37535_, _37533_, _37531_);
  or (_37536_, _37535_, _37510_);
  and (_37537_, _37536_, _07245_);
  or (_37538_, _37507_, _15568_);
  and (_37539_, _37538_, _06387_);
  and (_37540_, _37539_, _37525_);
  or (_37541_, _37540_, _14157_);
  or (_37542_, _37541_, _37537_);
  or (_37543_, _10762_, _10740_);
  or (_37544_, _37543_, _10796_);
  and (_37546_, _37544_, _37542_);
  or (_37547_, _37546_, _12586_);
  and (_37548_, _37547_, _06442_);
  and (_37549_, _37548_, _37506_);
  or (_37550_, _10577_, _10572_);
  or (_37551_, _37550_, _10628_);
  and (_37552_, _37551_, _12593_);
  or (_37553_, _37552_, _37549_);
  or (_37554_, _10842_, _10573_);
  or (_37555_, _37554_, _10894_);
  and (_37557_, _37555_, _06446_);
  and (_37558_, _37557_, _37553_);
  and (_37559_, _15585_, _08612_);
  or (_37560_, _37559_, _37507_);
  and (_37561_, _37560_, _06300_);
  or (_37562_, _37561_, _10059_);
  or (_37563_, _37562_, _37558_);
  and (_37564_, _37563_, _37504_);
  or (_37565_, _37564_, _06281_);
  and (_37566_, _07988_, _09440_);
  or (_37568_, _37500_, _06282_);
  or (_37569_, _37568_, _37566_);
  and (_37570_, _37569_, _06279_);
  and (_37571_, _37570_, _37565_);
  and (_37572_, _15639_, _07988_);
  or (_37573_, _37572_, _37500_);
  and (_37574_, _37573_, _06015_);
  or (_37575_, _37574_, _06275_);
  or (_37576_, _37575_, _37571_);
  and (_37577_, _15646_, _07988_);
  or (_37579_, _37577_, _37500_);
  or (_37580_, _37579_, _06276_);
  and (_37581_, _37580_, _37576_);
  or (_37582_, _37581_, _06474_);
  and (_37583_, _15531_, _07988_);
  or (_37584_, _37583_, _37500_);
  or (_37585_, _37584_, _07282_);
  and (_37586_, _37585_, _07284_);
  and (_37587_, _37586_, _37582_);
  and (_37588_, _11210_, _07988_);
  or (_37590_, _37588_, _37500_);
  and (_37591_, _37590_, _06582_);
  or (_37592_, _37591_, _37587_);
  and (_37593_, _37592_, _07279_);
  or (_37594_, _37500_, _08162_);
  and (_37595_, _37579_, _06478_);
  and (_37596_, _37595_, _37594_);
  or (_37597_, _37596_, _37593_);
  and (_37598_, _37597_, _07276_);
  and (_37599_, _37516_, _06569_);
  and (_37601_, _37599_, _37594_);
  or (_37602_, _37601_, _06479_);
  or (_37603_, _37602_, _37598_);
  and (_37604_, _15528_, _07988_);
  or (_37605_, _37604_, _37500_);
  or (_37606_, _37605_, _09043_);
  and (_37607_, _37606_, _37603_);
  or (_37608_, _37607_, _06572_);
  and (_37609_, _07378_, _05965_);
  nor (_37610_, _11209_, _13994_);
  or (_37612_, _37610_, _37500_);
  nor (_37613_, _37612_, _09048_);
  nor (_37614_, _37613_, _37609_);
  and (_37615_, _37614_, _37608_);
  and (_37616_, _37498_, _37609_);
  or (_37617_, _37616_, _06754_);
  or (_37618_, _37617_, _37615_);
  not (_37619_, _06754_);
  nor (_37620_, _37498_, _37619_);
  and (_37621_, _06289_, _05965_);
  nor (_37623_, _37621_, _37620_);
  and (_37624_, _37623_, _37618_);
  and (_37625_, _37621_, _37498_);
  nor (_37626_, _37625_, _37624_);
  or (_37627_, _37626_, _37497_);
  nand (_37628_, _37627_, _37499_);
  and (_37629_, _37628_, _06983_);
  and (_37630_, _37498_, _06982_);
  or (_37631_, _37630_, _37629_);
  and (_37632_, _37631_, _17464_);
  or (_37634_, _10533_, _10495_);
  and (_37635_, _37634_, _17463_);
  or (_37636_, _37635_, _37632_);
  and (_37637_, _37636_, _17687_);
  and (_37638_, _37634_, _06984_);
  or (_37639_, _37638_, _06578_);
  or (_37640_, _37639_, _37637_);
  or (_37641_, _10577_, _06579_);
  or (_37642_, _37641_, _11076_);
  and (_37643_, _37642_, _11091_);
  and (_37645_, _37643_, _37640_);
  or (_37646_, _37645_, _37496_);
  and (_37647_, _37646_, _11120_);
  and (_37648_, _11150_, _11121_);
  or (_37649_, _37648_, _11163_);
  or (_37650_, _37649_, _37647_);
  or (_37651_, _11192_, _11165_);
  and (_37652_, _37651_, _06308_);
  and (_37653_, _37652_, _37650_);
  or (_37654_, _11232_, _11203_);
  and (_37656_, _37654_, _12094_);
  or (_37657_, _37656_, _37653_);
  or (_37658_, _11268_, _14289_);
  and (_37659_, _37658_, _07037_);
  and (_37660_, _37659_, _37657_);
  and (_37661_, _37513_, _06606_);
  or (_37662_, _37661_, _37660_);
  and (_37663_, _37662_, _06807_);
  and (_37664_, _37509_, _06234_);
  or (_37665_, _37664_, _06195_);
  or (_37667_, _37665_, _37663_);
  and (_37668_, _15713_, _07988_);
  or (_37669_, _37500_, _06196_);
  or (_37670_, _37669_, _37668_);
  and (_37671_, _37670_, _01375_);
  and (_37672_, _37671_, _37667_);
  or (_37673_, _37672_, _37494_);
  and (_43072_, _37673_, _42545_);
  and (_37674_, _05962_, op0_cnst);
  or (_00000_, _37674_, rst);
  and (_37676_, _37674_, _01375_);
  and (_37677_, _25608_, _01987_);
  nor (_37678_, _25608_, _01987_);
  and (_37679_, _25962_, _01991_);
  nor (_37680_, _25962_, _01991_);
  or (_37681_, _37680_, _37679_);
  and (_37682_, _27696_, _02009_);
  nor (_37683_, _27696_, _02009_);
  or (_37684_, _37683_, _37682_);
  or (_37685_, _37684_, _37681_);
  nand (_37687_, _26651_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_37688_, _26651_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_37689_, _37688_, _37687_);
  and (_37690_, _27345_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_37691_, _27345_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_37692_, _28342_, _38214_);
  and (_37693_, _28342_, _38214_);
  or (_37694_, _37693_, _37692_);
  nand (_37695_, _28020_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_37696_, _28020_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_37698_, _37696_, _37695_);
  and (_37699_, _28954_, _38204_);
  nor (_37700_, _28954_, _38204_);
  or (_37701_, _37700_, _37699_);
  nor (_37702_, _29570_, _38230_);
  or (_37703_, _37702_, _37701_);
  nor (_37704_, _28654_, _38219_);
  nand (_37705_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_37706_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_37707_, _37706_, _37705_);
  or (_37709_, _29875_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_37710_, _29875_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_37711_, _37710_, _37709_);
  or (_37712_, _25232_, _01983_);
  nand (_37713_, _25232_, _01983_);
  and (_37714_, _37713_, _37712_);
  and (_37715_, _29266_, _38225_);
  nor (_37716_, _29266_, _38225_);
  or (_37717_, _37716_, _37715_);
  or (_37718_, _37717_, _37714_);
  or (_37720_, _37718_, _37711_);
  or (_37721_, _37720_, _37707_);
  or (_37722_, _37721_, _37704_);
  and (_37723_, _28654_, _38219_);
  and (_37724_, _29570_, _38230_);
  or (_37725_, _37724_, _37723_);
  or (_37726_, _37725_, _37722_);
  or (_37727_, _37726_, _37703_);
  or (_37728_, _37727_, _37698_);
  or (_37729_, _37728_, _37694_);
  or (_37731_, _37729_, _37691_);
  or (_37732_, _37731_, _37690_);
  and (_37733_, _26310_, _01995_);
  nor (_37734_, _26310_, _01995_);
  or (_37735_, _37734_, _37733_);
  nor (_37736_, _27002_, _02002_);
  and (_37737_, _27002_, _02002_);
  or (_37738_, _37737_, _37736_);
  or (_37739_, _37738_, _37735_);
  or (_37740_, _37739_, _37732_);
  or (_37742_, _37740_, _37689_);
  or (_37743_, _37742_, _37685_);
  or (_37744_, _37743_, _37678_);
  or (_37745_, _37744_, _37677_);
  and (property_invalid_pc, _37745_, _37676_);
  buf (_00543_, _42548_);
  buf (_03212_, _42545_);
  buf (_03257_, _42545_);
  buf (_03300_, _42545_);
  buf (_03347_, _42545_);
  buf (_03394_, _42545_);
  buf (_03444_, _42545_);
  buf (_03497_, _42545_);
  buf (_03550_, _42545_);
  buf (_03604_, _42545_);
  buf (_03657_, _42545_);
  buf (_03710_, _42545_);
  buf (_03763_, _42545_);
  buf (_03816_, _42545_);
  buf (_03870_, _42545_);
  buf (_03923_, _42545_);
  buf (_03974_, _42545_);
  buf (_38493_, _38389_);
  buf (_38495_, _38391_);
  buf (_38508_, _38389_);
  buf (_38509_, _38391_);
  buf (_38819_, _38409_);
  buf (_38820_, _38410_);
  buf (_38821_, _38412_);
  buf (_38822_, _38413_);
  buf (_38823_, _38414_);
  buf (_38824_, _38415_);
  buf (_38825_, _38416_);
  buf (_38826_, _38418_);
  buf (_38827_, _38419_);
  buf (_38828_, _38420_);
  buf (_38829_, _38421_);
  buf (_38830_, _38422_);
  buf (_38831_, _38424_);
  buf (_38832_, _38425_);
  buf (_38884_, _38409_);
  buf (_38885_, _38410_);
  buf (_38886_, _38412_);
  buf (_38887_, _38413_);
  buf (_38888_, _38414_);
  buf (_38889_, _38415_);
  buf (_38890_, _38416_);
  buf (_38891_, _38418_);
  buf (_38892_, _38419_);
  buf (_38894_, _38420_);
  buf (_38895_, _38421_);
  buf (_38896_, _38422_);
  buf (_38897_, _38424_);
  buf (_38898_, _38425_);
  buf (_39429_, _39204_);
  buf (_39586_, _39204_);
  dff (op0_cnst, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _03215_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _03218_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _03222_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _03225_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _03228_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _03232_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _03235_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _03209_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _03212_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _03260_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _03263_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _03267_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _03270_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _03274_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _03277_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _03280_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _03254_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _03257_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _03714_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _03718_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _03722_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _03726_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _03730_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _03734_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _03738_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _03707_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _03710_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _03767_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _03771_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _03775_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _03779_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _03783_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _03787_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _03791_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _03760_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _03763_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _03820_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _03824_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _03828_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _03832_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _03836_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _03840_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _03844_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _03813_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _03816_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _03874_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _03878_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _03882_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _03886_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _03890_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _03894_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _03898_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _03867_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _03870_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _03927_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _03931_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _03934_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _03938_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _03942_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _03946_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _03950_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _03920_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _03923_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _03978_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _03982_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _03986_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _03990_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _03994_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _03998_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _04002_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _03971_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _03974_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _03304_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _03307_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _03311_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _03314_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _03318_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _03321_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _03325_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _03297_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _03300_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _03350_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _03354_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _03357_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _03361_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _03364_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _03368_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _03373_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _03344_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _03347_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _03397_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _03400_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _03404_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _03407_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _03411_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _03415_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _03419_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _03391_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _03394_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _03448_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _03452_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _03456_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _03460_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _03464_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _03468_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _03472_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _03441_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _03444_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _03501_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _03505_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _03509_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _03513_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _03517_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _03521_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _03525_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _03494_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _03497_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _03554_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _03558_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _03562_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _03566_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _03570_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _03574_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _03578_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _03547_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _03550_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _03608_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _03612_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _03616_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _03620_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _03624_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _03628_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _03632_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _03600_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _03604_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _03661_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _03665_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _03669_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _03673_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _03677_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _03681_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _03685_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _03654_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _03657_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02915_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02928_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02952_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02975_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02998_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00950_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03010_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00925_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03021_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03034_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03045_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03058_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03070_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03081_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03091_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00968_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02351_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22121_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02542_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02736_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02964_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03166_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03371_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03603_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03848_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04074_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04170_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04270_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04369_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04468_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04563_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04662_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04760_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24280_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38401_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38403_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38404_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38405_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38406_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38407_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38408_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38388_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38409_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38410_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38412_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38413_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38414_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38415_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38416_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38389_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38418_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38419_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38420_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38421_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38422_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38424_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38425_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38391_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _32090_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _07747_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _32091_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _32094_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _07750_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _32096_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _32098_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _07753_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _32100_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _07756_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _32102_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _32104_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _32106_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _07759_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _32108_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _07762_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _07765_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _07824_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _07826_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _07729_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _07829_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _07832_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _07732_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _07835_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _07735_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _07838_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _07841_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _07844_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _07847_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _07850_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _07853_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _07856_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _07738_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _07741_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _07859_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _07744_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39204_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _39304_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _39305_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _39306_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _39307_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _39308_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _39309_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _39310_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39205_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _39311_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _39312_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _39313_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _39315_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _39316_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _39317_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _39318_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39206_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _39319_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _39320_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _39321_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _39322_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _39323_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _39324_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _39326_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39207_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _39327_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _39328_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _39329_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _39330_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _39331_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _39332_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _39333_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39209_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _39334_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _39335_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _39337_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _39338_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _39339_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _39340_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _39341_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _39210_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _39342_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _39343_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _39344_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _39345_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _39346_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _39348_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _39349_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _39211_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _39350_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _39351_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _39352_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _39353_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _39354_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _39355_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _39356_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _39212_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _39357_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _39358_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _39359_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _39360_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _39361_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _39362_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _39363_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _39213_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _38772_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _38773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _38774_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _38775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38491_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38565_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38567_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38568_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38569_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38571_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38572_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38573_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38574_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38575_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38576_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38577_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38578_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _38579_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _38580_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38450_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _38584_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _38585_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _38586_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _38587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _38588_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _38589_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _38590_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _38591_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _38592_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _38593_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _38594_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _38595_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _38596_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _38597_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _38598_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38451_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _38776_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _38777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _38778_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _38779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _38781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _38782_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _38783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _38784_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _38785_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _38786_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _38787_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _38788_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _38789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _38790_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _38792_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _38793_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _38794_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _38795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _38796_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _38797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _38798_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _38799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _38800_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _38801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _38803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _38804_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _38805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _38806_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _38807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _38808_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _38809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38516_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38489_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _38810_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _38812_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _38813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _38814_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _38815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _38816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _38818_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38492_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _38819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _38820_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _38821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _38822_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _38823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _38824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _38825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38493_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _38826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _38827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _38828_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _38829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _38830_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _38831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _38832_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38495_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38496_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38497_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _38833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _38834_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _38835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _38836_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _38837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _38839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _38840_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38498_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _38841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _38842_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _38843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _38844_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _38845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _38846_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _38847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _38848_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _38850_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _38851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _38852_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _38853_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _38854_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _38855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _38856_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38499_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _38857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _38858_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _38859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _38861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _38862_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _38863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _38864_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _38865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _38866_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _38867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _38868_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _38869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _38870_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _38872_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _38873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38501_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38502_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38504_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38503_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _38874_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _38875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _38876_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _38877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _38878_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _38879_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _38880_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38506_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _38881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _38883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38507_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _38884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _38885_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _38886_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _38887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _38888_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _38889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _38890_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38508_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _38891_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _38892_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _38894_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _38895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _38896_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _38897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _38898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38509_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _38510_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _38899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _38900_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _38901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _38902_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _38903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _38905_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _38906_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38511_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _38513_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38514_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _38907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _38908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _38909_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38515_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _38910_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _38911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _38912_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _38913_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _38914_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _38916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _38917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _38918_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _38919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _38920_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _38921_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _38922_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _38923_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _38924_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _38925_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _38927_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _38928_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _38929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _38930_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _38931_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _38932_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _38933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _38934_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _38935_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _38936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _38938_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _38939_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _38940_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _38941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _38942_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _38943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38517_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _38944_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _38945_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _38946_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _38947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _38949_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _38950_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _38951_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38518_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38519_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38521_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _38952_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _38953_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _38954_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _38955_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _38956_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _38957_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _38958_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _38960_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _38961_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _38962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _38963_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _38964_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _38965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _38966_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _38967_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38522_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38523_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38524_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38525_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _38968_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _38969_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _38971_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _38972_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _38973_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _38974_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _38975_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _38976_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _38977_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _38978_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _38979_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _38980_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _38982_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _38983_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _38984_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38526_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38527_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39584_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39604_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39605_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39606_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39607_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39608_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39609_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39610_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39585_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39586_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39611_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39613_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _02987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _02990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _02993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _02997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _02959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _02962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _02966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _02970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _02973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _02977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _02980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _02983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _02930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _02933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _02936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _02940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _02943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _02947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _02950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _02954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _02899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _02903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _02906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _02910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _02914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _02918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _02922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _02924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _02871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _02874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _02878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _02881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _02885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _02889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _02892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _02895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _02843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _02847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _02850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _02853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _02856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _02860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _02864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _02866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _02815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _02818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _02822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _02825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _02828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _02831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _02835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _02837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _02792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _02796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _02799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _02802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _02805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _02809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _02811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _03193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _03194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _03196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _03198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _03200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _03201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _03203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02573_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _39423_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _39505_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _39506_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _39507_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _39425_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39426_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39427_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39509_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39510_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39511_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39512_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39513_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39514_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39515_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39428_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39429_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19778_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19789_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19801_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19813_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17961_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08902_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08913_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08946_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08957_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13611_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13676_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12675_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13687_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _42549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _42548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _42545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42543_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _42541_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _42539_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _42537_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _42535_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42533_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42531_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _42493_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _42491_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _42489_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _42487_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _42484_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00171_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _42482_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00176_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00182_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00185_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _42479_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40232_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40238_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40240_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40251_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40253_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40255_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40257_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31054_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40259_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40263_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40265_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40267_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31077_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40272_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40274_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40276_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40278_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40280_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40284_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31099_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17359_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17370_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17381_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17392_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09507_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10669_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10713_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10724_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09528_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _40734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _40737_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41251_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41253_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _40740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41260_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41262_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41264_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41268_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41270_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _40743_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _40746_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _40749_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41273_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41277_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41283_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41285_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _40752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41287_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41288_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41292_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _40755_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _40758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41304_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41311_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _40761_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01625_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01628_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01631_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02117_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02120_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02124_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02125_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02127_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02129_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02171_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01207_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01208_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01210_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01213_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01215_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00567_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00543_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00546_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00551_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00554_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00556_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01227_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01229_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01231_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01233_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01235_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01241_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00564_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00572_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01246_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01248_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01252_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01260_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01262_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01264_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01268_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01270_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01272_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01274_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01276_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01278_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01280_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01283_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00588_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01285_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01287_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01291_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01295_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00591_);
  dff (\uc8051golden_1.IRAM[15] [0], _40544_);
  dff (\uc8051golden_1.IRAM[15] [1], _40545_);
  dff (\uc8051golden_1.IRAM[15] [2], _40547_);
  dff (\uc8051golden_1.IRAM[15] [3], _40548_);
  dff (\uc8051golden_1.IRAM[15] [4], _40549_);
  dff (\uc8051golden_1.IRAM[15] [5], _40550_);
  dff (\uc8051golden_1.IRAM[15] [6], _40551_);
  dff (\uc8051golden_1.IRAM[15] [7], _40322_);
  dff (\uc8051golden_1.IRAM[14] [0], _40532_);
  dff (\uc8051golden_1.IRAM[14] [1], _40533_);
  dff (\uc8051golden_1.IRAM[14] [2], _40535_);
  dff (\uc8051golden_1.IRAM[14] [3], _40536_);
  dff (\uc8051golden_1.IRAM[14] [4], _40537_);
  dff (\uc8051golden_1.IRAM[14] [5], _40538_);
  dff (\uc8051golden_1.IRAM[14] [6], _40539_);
  dff (\uc8051golden_1.IRAM[14] [7], _40541_);
  dff (\uc8051golden_1.IRAM[13] [0], _40520_);
  dff (\uc8051golden_1.IRAM[13] [1], _40521_);
  dff (\uc8051golden_1.IRAM[13] [2], _40523_);
  dff (\uc8051golden_1.IRAM[13] [3], _40524_);
  dff (\uc8051golden_1.IRAM[13] [4], _40525_);
  dff (\uc8051golden_1.IRAM[13] [5], _40526_);
  dff (\uc8051golden_1.IRAM[13] [6], _40527_);
  dff (\uc8051golden_1.IRAM[13] [7], _40528_);
  dff (\uc8051golden_1.IRAM[12] [0], _40508_);
  dff (\uc8051golden_1.IRAM[12] [1], _40509_);
  dff (\uc8051golden_1.IRAM[12] [2], _40510_);
  dff (\uc8051golden_1.IRAM[12] [3], _40512_);
  dff (\uc8051golden_1.IRAM[12] [4], _40513_);
  dff (\uc8051golden_1.IRAM[12] [5], _40514_);
  dff (\uc8051golden_1.IRAM[12] [6], _40515_);
  dff (\uc8051golden_1.IRAM[12] [7], _40516_);
  dff (\uc8051golden_1.IRAM[11] [0], _40495_);
  dff (\uc8051golden_1.IRAM[11] [1], _40496_);
  dff (\uc8051golden_1.IRAM[11] [2], _40497_);
  dff (\uc8051golden_1.IRAM[11] [3], _40498_);
  dff (\uc8051golden_1.IRAM[11] [4], _40501_);
  dff (\uc8051golden_1.IRAM[11] [5], _40502_);
  dff (\uc8051golden_1.IRAM[11] [6], _40503_);
  dff (\uc8051golden_1.IRAM[11] [7], _40504_);
  dff (\uc8051golden_1.IRAM[10] [0], _40484_);
  dff (\uc8051golden_1.IRAM[10] [1], _40485_);
  dff (\uc8051golden_1.IRAM[10] [2], _40486_);
  dff (\uc8051golden_1.IRAM[10] [3], _40487_);
  dff (\uc8051golden_1.IRAM[10] [4], _40488_);
  dff (\uc8051golden_1.IRAM[10] [5], _40490_);
  dff (\uc8051golden_1.IRAM[10] [6], _40491_);
  dff (\uc8051golden_1.IRAM[10] [7], _40492_);
  dff (\uc8051golden_1.IRAM[9] [0], _40472_);
  dff (\uc8051golden_1.IRAM[9] [1], _40473_);
  dff (\uc8051golden_1.IRAM[9] [2], _40474_);
  dff (\uc8051golden_1.IRAM[9] [3], _40475_);
  dff (\uc8051golden_1.IRAM[9] [4], _40476_);
  dff (\uc8051golden_1.IRAM[9] [5], _40478_);
  dff (\uc8051golden_1.IRAM[9] [6], _40479_);
  dff (\uc8051golden_1.IRAM[9] [7], _40480_);
  dff (\uc8051golden_1.IRAM[8] [0], _40458_);
  dff (\uc8051golden_1.IRAM[8] [1], _40461_);
  dff (\uc8051golden_1.IRAM[8] [2], _40462_);
  dff (\uc8051golden_1.IRAM[8] [3], _40463_);
  dff (\uc8051golden_1.IRAM[8] [4], _40464_);
  dff (\uc8051golden_1.IRAM[8] [5], _40465_);
  dff (\uc8051golden_1.IRAM[8] [6], _40467_);
  dff (\uc8051golden_1.IRAM[8] [7], _40468_);
  dff (\uc8051golden_1.IRAM[7] [0], _40446_);
  dff (\uc8051golden_1.IRAM[7] [1], _40447_);
  dff (\uc8051golden_1.IRAM[7] [2], _40448_);
  dff (\uc8051golden_1.IRAM[7] [3], _40449_);
  dff (\uc8051golden_1.IRAM[7] [4], _40452_);
  dff (\uc8051golden_1.IRAM[7] [5], _40453_);
  dff (\uc8051golden_1.IRAM[7] [6], _40454_);
  dff (\uc8051golden_1.IRAM[7] [7], _40455_);
  dff (\uc8051golden_1.IRAM[6] [0], _40435_);
  dff (\uc8051golden_1.IRAM[6] [1], _40436_);
  dff (\uc8051golden_1.IRAM[6] [2], _40437_);
  dff (\uc8051golden_1.IRAM[6] [3], _40438_);
  dff (\uc8051golden_1.IRAM[6] [4], _40439_);
  dff (\uc8051golden_1.IRAM[6] [5], _40441_);
  dff (\uc8051golden_1.IRAM[6] [6], _40442_);
  dff (\uc8051golden_1.IRAM[6] [7], _40443_);
  dff (\uc8051golden_1.IRAM[5] [0], _40423_);
  dff (\uc8051golden_1.IRAM[5] [1], _40424_);
  dff (\uc8051golden_1.IRAM[5] [2], _40425_);
  dff (\uc8051golden_1.IRAM[5] [3], _40426_);
  dff (\uc8051golden_1.IRAM[5] [4], _40427_);
  dff (\uc8051golden_1.IRAM[5] [5], _40429_);
  dff (\uc8051golden_1.IRAM[5] [6], _40430_);
  dff (\uc8051golden_1.IRAM[5] [7], _40431_);
  dff (\uc8051golden_1.IRAM[4] [0], _40410_);
  dff (\uc8051golden_1.IRAM[4] [1], _40412_);
  dff (\uc8051golden_1.IRAM[4] [2], _40413_);
  dff (\uc8051golden_1.IRAM[4] [3], _40414_);
  dff (\uc8051golden_1.IRAM[4] [4], _40415_);
  dff (\uc8051golden_1.IRAM[4] [5], _40416_);
  dff (\uc8051golden_1.IRAM[4] [6], _40418_);
  dff (\uc8051golden_1.IRAM[4] [7], _40419_);
  dff (\uc8051golden_1.IRAM[3] [0], _40398_);
  dff (\uc8051golden_1.IRAM[3] [1], _40399_);
  dff (\uc8051golden_1.IRAM[3] [2], _40400_);
  dff (\uc8051golden_1.IRAM[3] [3], _40401_);
  dff (\uc8051golden_1.IRAM[3] [4], _40403_);
  dff (\uc8051golden_1.IRAM[3] [5], _40404_);
  dff (\uc8051golden_1.IRAM[3] [6], _40405_);
  dff (\uc8051golden_1.IRAM[3] [7], _40406_);
  dff (\uc8051golden_1.IRAM[2] [0], _40387_);
  dff (\uc8051golden_1.IRAM[2] [1], _40388_);
  dff (\uc8051golden_1.IRAM[2] [2], _40389_);
  dff (\uc8051golden_1.IRAM[2] [3], _40390_);
  dff (\uc8051golden_1.IRAM[2] [4], _40391_);
  dff (\uc8051golden_1.IRAM[2] [5], _40392_);
  dff (\uc8051golden_1.IRAM[2] [6], _40393_);
  dff (\uc8051golden_1.IRAM[2] [7], _40394_);
  dff (\uc8051golden_1.IRAM[1] [0], _40374_);
  dff (\uc8051golden_1.IRAM[1] [1], _40375_);
  dff (\uc8051golden_1.IRAM[1] [2], _40376_);
  dff (\uc8051golden_1.IRAM[1] [3], _40378_);
  dff (\uc8051golden_1.IRAM[1] [4], _40379_);
  dff (\uc8051golden_1.IRAM[1] [5], _40380_);
  dff (\uc8051golden_1.IRAM[1] [6], _40381_);
  dff (\uc8051golden_1.IRAM[1] [7], _40382_);
  dff (\uc8051golden_1.IRAM[0] [0], _40361_);
  dff (\uc8051golden_1.IRAM[0] [1], _40362_);
  dff (\uc8051golden_1.IRAM[0] [2], _40363_);
  dff (\uc8051golden_1.IRAM[0] [3], _40364_);
  dff (\uc8051golden_1.IRAM[0] [4], _40366_);
  dff (\uc8051golden_1.IRAM[0] [5], _40367_);
  dff (\uc8051golden_1.IRAM[0] [6], _40368_);
  dff (\uc8051golden_1.IRAM[0] [7], _40370_);
  dff (\uc8051golden_1.B [0], _42889_);
  dff (\uc8051golden_1.B [1], _42890_);
  dff (\uc8051golden_1.B [2], _42891_);
  dff (\uc8051golden_1.B [3], _42892_);
  dff (\uc8051golden_1.B [4], _42893_);
  dff (\uc8051golden_1.B [5], _42894_);
  dff (\uc8051golden_1.B [6], _42895_);
  dff (\uc8051golden_1.B [7], _40323_);
  dff (\uc8051golden_1.ACC [0], _42896_);
  dff (\uc8051golden_1.ACC [1], _42898_);
  dff (\uc8051golden_1.ACC [2], _42899_);
  dff (\uc8051golden_1.ACC [3], _42900_);
  dff (\uc8051golden_1.ACC [4], _42901_);
  dff (\uc8051golden_1.ACC [5], _42902_);
  dff (\uc8051golden_1.ACC [6], _42903_);
  dff (\uc8051golden_1.ACC [7], _40324_);
  dff (\uc8051golden_1.PCON [0], _42905_);
  dff (\uc8051golden_1.PCON [1], _42906_);
  dff (\uc8051golden_1.PCON [2], _42907_);
  dff (\uc8051golden_1.PCON [3], _42908_);
  dff (\uc8051golden_1.PCON [4], _42909_);
  dff (\uc8051golden_1.PCON [5], _42910_);
  dff (\uc8051golden_1.PCON [6], _42911_);
  dff (\uc8051golden_1.PCON [7], _40325_);
  dff (\uc8051golden_1.TMOD [0], _42912_);
  dff (\uc8051golden_1.TMOD [1], _42913_);
  dff (\uc8051golden_1.TMOD [2], _42914_);
  dff (\uc8051golden_1.TMOD [3], _42916_);
  dff (\uc8051golden_1.TMOD [4], _42917_);
  dff (\uc8051golden_1.TMOD [5], _42918_);
  dff (\uc8051golden_1.TMOD [6], _42919_);
  dff (\uc8051golden_1.TMOD [7], _40326_);
  dff (\uc8051golden_1.DPL [0], _42921_);
  dff (\uc8051golden_1.DPL [1], _42922_);
  dff (\uc8051golden_1.DPL [2], _42923_);
  dff (\uc8051golden_1.DPL [3], _42924_);
  dff (\uc8051golden_1.DPL [4], _42925_);
  dff (\uc8051golden_1.DPL [5], _42926_);
  dff (\uc8051golden_1.DPL [6], _42927_);
  dff (\uc8051golden_1.DPL [7], _40328_);
  dff (\uc8051golden_1.DPH [0], _42928_);
  dff (\uc8051golden_1.DPH [1], _42929_);
  dff (\uc8051golden_1.DPH [2], _42930_);
  dff (\uc8051golden_1.DPH [3], _42931_);
  dff (\uc8051golden_1.DPH [4], _42932_);
  dff (\uc8051golden_1.DPH [5], _42934_);
  dff (\uc8051golden_1.DPH [6], _42935_);
  dff (\uc8051golden_1.DPH [7], _40329_);
  dff (\uc8051golden_1.TL1 [0], _42936_);
  dff (\uc8051golden_1.TL1 [1], _42938_);
  dff (\uc8051golden_1.TL1 [2], _42939_);
  dff (\uc8051golden_1.TL1 [3], _42940_);
  dff (\uc8051golden_1.TL1 [4], _42941_);
  dff (\uc8051golden_1.TL1 [5], _42942_);
  dff (\uc8051golden_1.TL1 [6], _42943_);
  dff (\uc8051golden_1.TL1 [7], _40330_);
  dff (\uc8051golden_1.TL0 [0], _42944_);
  dff (\uc8051golden_1.TL0 [1], _42945_);
  dff (\uc8051golden_1.TL0 [2], _42946_);
  dff (\uc8051golden_1.TL0 [3], _42947_);
  dff (\uc8051golden_1.TL0 [4], _42948_);
  dff (\uc8051golden_1.TL0 [5], _42949_);
  dff (\uc8051golden_1.TL0 [6], _42950_);
  dff (\uc8051golden_1.TL0 [7], _40331_);
  dff (\uc8051golden_1.TCON [0], _42952_);
  dff (\uc8051golden_1.TCON [1], _42953_);
  dff (\uc8051golden_1.TCON [2], _42954_);
  dff (\uc8051golden_1.TCON [3], _42956_);
  dff (\uc8051golden_1.TCON [4], _42957_);
  dff (\uc8051golden_1.TCON [5], _42958_);
  dff (\uc8051golden_1.TCON [6], _42959_);
  dff (\uc8051golden_1.TCON [7], _40332_);
  dff (\uc8051golden_1.TH1 [0], _42960_);
  dff (\uc8051golden_1.TH1 [1], _42961_);
  dff (\uc8051golden_1.TH1 [2], _42962_);
  dff (\uc8051golden_1.TH1 [3], _42963_);
  dff (\uc8051golden_1.TH1 [4], _42964_);
  dff (\uc8051golden_1.TH1 [5], _42965_);
  dff (\uc8051golden_1.TH1 [6], _42966_);
  dff (\uc8051golden_1.TH1 [7], _40334_);
  dff (\uc8051golden_1.TH0 [0], _42968_);
  dff (\uc8051golden_1.TH0 [1], _42969_);
  dff (\uc8051golden_1.TH0 [2], _42970_);
  dff (\uc8051golden_1.TH0 [3], _42971_);
  dff (\uc8051golden_1.TH0 [4], _42972_);
  dff (\uc8051golden_1.TH0 [5], _42974_);
  dff (\uc8051golden_1.TH0 [6], _42975_);
  dff (\uc8051golden_1.TH0 [7], _40335_);
  dff (\uc8051golden_1.PC [0], _42976_);
  dff (\uc8051golden_1.PC [1], _42977_);
  dff (\uc8051golden_1.PC [2], _42978_);
  dff (\uc8051golden_1.PC [3], _42980_);
  dff (\uc8051golden_1.PC [4], _42981_);
  dff (\uc8051golden_1.PC [5], _42982_);
  dff (\uc8051golden_1.PC [6], _42983_);
  dff (\uc8051golden_1.PC [7], _42984_);
  dff (\uc8051golden_1.PC [8], _42985_);
  dff (\uc8051golden_1.PC [9], _42986_);
  dff (\uc8051golden_1.PC [10], _42987_);
  dff (\uc8051golden_1.PC [11], _42988_);
  dff (\uc8051golden_1.PC [12], _42989_);
  dff (\uc8051golden_1.PC [13], _42991_);
  dff (\uc8051golden_1.PC [14], _42992_);
  dff (\uc8051golden_1.PC [15], _40336_);
  dff (\uc8051golden_1.P2 [0], _42993_);
  dff (\uc8051golden_1.P2 [1], _42994_);
  dff (\uc8051golden_1.P2 [2], _42995_);
  dff (\uc8051golden_1.P2 [3], _42996_);
  dff (\uc8051golden_1.P2 [4], _42997_);
  dff (\uc8051golden_1.P2 [5], _42998_);
  dff (\uc8051golden_1.P2 [6], _42999_);
  dff (\uc8051golden_1.P2 [7], _40337_);
  dff (\uc8051golden_1.P3 [0], _43001_);
  dff (\uc8051golden_1.P3 [1], _43002_);
  dff (\uc8051golden_1.P3 [2], _43003_);
  dff (\uc8051golden_1.P3 [3], _43004_);
  dff (\uc8051golden_1.P3 [4], _43005_);
  dff (\uc8051golden_1.P3 [5], _43006_);
  dff (\uc8051golden_1.P3 [6], _43007_);
  dff (\uc8051golden_1.P3 [7], _40338_);
  dff (\uc8051golden_1.P0 [0], _43009_);
  dff (\uc8051golden_1.P0 [1], _43010_);
  dff (\uc8051golden_1.P0 [2], _43011_);
  dff (\uc8051golden_1.P0 [3], _43012_);
  dff (\uc8051golden_1.P0 [4], _43013_);
  dff (\uc8051golden_1.P0 [5], _43014_);
  dff (\uc8051golden_1.P0 [6], _43015_);
  dff (\uc8051golden_1.P0 [7], _40339_);
  dff (\uc8051golden_1.P1 [0], _43017_);
  dff (\uc8051golden_1.P1 [1], _43018_);
  dff (\uc8051golden_1.P1 [2], _43019_);
  dff (\uc8051golden_1.P1 [3], _43020_);
  dff (\uc8051golden_1.P1 [4], _43021_);
  dff (\uc8051golden_1.P1 [5], _43022_);
  dff (\uc8051golden_1.P1 [6], _43023_);
  dff (\uc8051golden_1.P1 [7], _40340_);
  dff (\uc8051golden_1.IP [0], _43025_);
  dff (\uc8051golden_1.IP [1], _43026_);
  dff (\uc8051golden_1.IP [2], _43027_);
  dff (\uc8051golden_1.IP [3], _43028_);
  dff (\uc8051golden_1.IP [4], _43029_);
  dff (\uc8051golden_1.IP [5], _43030_);
  dff (\uc8051golden_1.IP [6], _43031_);
  dff (\uc8051golden_1.IP [7], _40341_);
  dff (\uc8051golden_1.IE [0], _43032_);
  dff (\uc8051golden_1.IE [1], _43034_);
  dff (\uc8051golden_1.IE [2], _43035_);
  dff (\uc8051golden_1.IE [3], _43036_);
  dff (\uc8051golden_1.IE [4], _43037_);
  dff (\uc8051golden_1.IE [5], _43038_);
  dff (\uc8051golden_1.IE [6], _43039_);
  dff (\uc8051golden_1.IE [7], _40342_);
  dff (\uc8051golden_1.SCON [0], _43041_);
  dff (\uc8051golden_1.SCON [1], _43042_);
  dff (\uc8051golden_1.SCON [2], _43043_);
  dff (\uc8051golden_1.SCON [3], _43044_);
  dff (\uc8051golden_1.SCON [4], _43045_);
  dff (\uc8051golden_1.SCON [5], _43046_);
  dff (\uc8051golden_1.SCON [6], _43047_);
  dff (\uc8051golden_1.SCON [7], _40343_);
  dff (\uc8051golden_1.SP [0], _43048_);
  dff (\uc8051golden_1.SP [1], _43049_);
  dff (\uc8051golden_1.SP [2], _43050_);
  dff (\uc8051golden_1.SP [3], _43052_);
  dff (\uc8051golden_1.SP [4], _43053_);
  dff (\uc8051golden_1.SP [5], _43054_);
  dff (\uc8051golden_1.SP [6], _43055_);
  dff (\uc8051golden_1.SP [7], _40345_);
  dff (\uc8051golden_1.SBUF [0], _43057_);
  dff (\uc8051golden_1.SBUF [1], _43058_);
  dff (\uc8051golden_1.SBUF [2], _43059_);
  dff (\uc8051golden_1.SBUF [3], _43060_);
  dff (\uc8051golden_1.SBUF [4], _43061_);
  dff (\uc8051golden_1.SBUF [5], _43062_);
  dff (\uc8051golden_1.SBUF [6], _43063_);
  dff (\uc8051golden_1.SBUF [7], _40346_);
  dff (\uc8051golden_1.PSW [0], _43065_);
  dff (\uc8051golden_1.PSW [1], _43066_);
  dff (\uc8051golden_1.PSW [2], _43067_);
  dff (\uc8051golden_1.PSW [3], _43068_);
  dff (\uc8051golden_1.PSW [4], _43069_);
  dff (\uc8051golden_1.PSW [5], _43071_);
  dff (\uc8051golden_1.PSW [6], _43072_);
  dff (\uc8051golden_1.PSW [7], _40347_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \uc8051golden_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \uc8051golden_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \uc8051golden_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \uc8051golden_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \uc8051golden_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \uc8051golden_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \uc8051golden_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \uc8051golden_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \uc8051golden_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \uc8051golden_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \uc8051golden_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \uc8051golden_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \uc8051golden_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \uc8051golden_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \uc8051golden_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \uc8051golden_1.PC [15]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [0], \uc8051golden_1.PC [0]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [1], \uc8051golden_1.PC [1]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [2], \uc8051golden_1.PC [2]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [3], \uc8051golden_1.PC [3]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [4], \uc8051golden_1.PC [4]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [5], \uc8051golden_1.PC [5]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [6], \uc8051golden_1.PC [6]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [7], \uc8051golden_1.PC [7]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [8], \uc8051golden_1.PC [8]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [9], \uc8051golden_1.PC [9]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [10], \uc8051golden_1.PC [10]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [11], \uc8051golden_1.PC [11]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [12], \uc8051golden_1.PC [12]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [13], \uc8051golden_1.PC [13]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [14], \uc8051golden_1.PC [14]);
  buf(\uc8051golden_1.RD_ROM_0_ADDR [15], \uc8051golden_1.PC [15]);
  buf(\uc8051golden_1.clk , clk);
  buf(\uc8051golden_1.rst , rst);
  buf(\uc8051golden_1.ACC_03 [0], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_03 [1], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_03 [2], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_03 [3], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_03 [4], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_03 [5], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_03 [6], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_03 [7], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.ACC_13 [0], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_13 [1], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_13 [2], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_13 [3], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_13 [4], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_13 [5], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_13 [6], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_13 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.ACC_23 [0], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_23 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.ACC_23 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_23 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_23 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_23 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_23 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_23 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_33 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.ACC_33 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.ACC_33 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_33 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_33 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_33 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_33 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_33 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_c4 [0], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_c4 [1], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_c4 [2], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_c4 [3], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_c4 [4], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.ACC_c4 [5], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_c4 [6], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_c4 [7], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_d6 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.ACC_d6 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.ACC_d6 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.ACC_d6 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.ACC_d6 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_d6 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_d6 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_d6 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_d7 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.ACC_d7 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.ACC_d7 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.ACC_d7 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.ACC_d7 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_d7 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_d7 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_d7 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_e4 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.ACC_e4 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.ACC_e4 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.ACC_e4 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.ACC_e4 [4], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.ACC_e4 [5], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.ACC_e4 [6], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.ACC_e4 [7], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.PC_22 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.PC_22 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.PC_22 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.PC_22 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.PC_22 [4], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.PC_22 [5], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.PC_22 [6], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.PC_22 [7], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.PC_22 [8], \uc8051golden_1.n1268 [0]);
  buf(\uc8051golden_1.PC_22 [9], \uc8051golden_1.n1268 [1]);
  buf(\uc8051golden_1.PC_22 [10], \uc8051golden_1.n1268 [2]);
  buf(\uc8051golden_1.PC_22 [11], \uc8051golden_1.n1268 [3]);
  buf(\uc8051golden_1.PC_22 [12], \uc8051golden_1.n1268 [4]);
  buf(\uc8051golden_1.PC_22 [13], \uc8051golden_1.n1268 [5]);
  buf(\uc8051golden_1.PC_22 [14], \uc8051golden_1.n1268 [6]);
  buf(\uc8051golden_1.PC_22 [15], \uc8051golden_1.n1268 [8]);
  buf(\uc8051golden_1.PC_32 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.PC_32 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.PC_32 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.PC_32 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.PC_32 [4], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.PC_32 [5], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.PC_32 [6], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.PC_32 [7], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.PC_32 [8], \uc8051golden_1.n1268 [0]);
  buf(\uc8051golden_1.PC_32 [9], \uc8051golden_1.n1268 [1]);
  buf(\uc8051golden_1.PC_32 [10], \uc8051golden_1.n1268 [2]);
  buf(\uc8051golden_1.PC_32 [11], \uc8051golden_1.n1268 [3]);
  buf(\uc8051golden_1.PC_32 [12], \uc8051golden_1.n1268 [4]);
  buf(\uc8051golden_1.PC_32 [13], \uc8051golden_1.n1268 [5]);
  buf(\uc8051golden_1.PC_32 [14], \uc8051golden_1.n1268 [6]);
  buf(\uc8051golden_1.PC_32 [15], \uc8051golden_1.n1268 [8]);
  buf(\uc8051golden_1.PSW_13 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_13 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_13 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_13 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_13 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_13 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_13 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_13 [7], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.PSW_24 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_24 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_24 [2], \uc8051golden_1.n1207 [2]);
  buf(\uc8051golden_1.PSW_24 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_24 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_24 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_24 [6], \uc8051golden_1.n1207 [6]);
  buf(\uc8051golden_1.PSW_24 [7], \uc8051golden_1.n1207 [7]);
  buf(\uc8051golden_1.PSW_25 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_25 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_25 [2], \uc8051golden_1.n1227 [2]);
  buf(\uc8051golden_1.PSW_25 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_25 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_25 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_25 [6], \uc8051golden_1.n1227 [6]);
  buf(\uc8051golden_1.PSW_25 [7], \uc8051golden_1.n1227 [7]);
  buf(\uc8051golden_1.PSW_26 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_26 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_26 [2], \uc8051golden_1.n1246 [2]);
  buf(\uc8051golden_1.PSW_26 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_26 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_26 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_26 [6], \uc8051golden_1.n1258 [6]);
  buf(\uc8051golden_1.PSW_26 [7], \uc8051golden_1.n1246 [7]);
  buf(\uc8051golden_1.PSW_27 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_27 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_27 [2], \uc8051golden_1.n1258 [2]);
  buf(\uc8051golden_1.PSW_27 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_27 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_27 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_27 [6], \uc8051golden_1.n1258 [6]);
  buf(\uc8051golden_1.PSW_27 [7], \uc8051golden_1.n1258 [7]);
  buf(\uc8051golden_1.PSW_28 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_28 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_28 [2], \uc8051golden_1.n1280 [2]);
  buf(\uc8051golden_1.PSW_28 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_28 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_28 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_28 [6], \uc8051golden_1.n1292 [6]);
  buf(\uc8051golden_1.PSW_28 [7], \uc8051golden_1.n1280 [7]);
  buf(\uc8051golden_1.PSW_29 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_29 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_29 [2], \uc8051golden_1.n1280 [2]);
  buf(\uc8051golden_1.PSW_29 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_29 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_29 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_29 [6], \uc8051golden_1.n1292 [6]);
  buf(\uc8051golden_1.PSW_29 [7], \uc8051golden_1.n1280 [7]);
  buf(\uc8051golden_1.PSW_2a [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2a [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2a [2], \uc8051golden_1.n1280 [2]);
  buf(\uc8051golden_1.PSW_2a [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2a [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2a [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2a [6], \uc8051golden_1.n1291 [6]);
  buf(\uc8051golden_1.PSW_2a [7], \uc8051golden_1.n1280 [7]);
  buf(\uc8051golden_1.PSW_2b [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2b [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2b [2], \uc8051golden_1.n1292 [2]);
  buf(\uc8051golden_1.PSW_2b [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2b [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2b [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2b [6], \uc8051golden_1.n1291 [6]);
  buf(\uc8051golden_1.PSW_2b [7], \uc8051golden_1.n1292 [7]);
  buf(\uc8051golden_1.PSW_2c [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2c [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2c [2], \uc8051golden_1.n1292 [2]);
  buf(\uc8051golden_1.PSW_2c [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2c [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2c [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2c [6], \uc8051golden_1.n1291 [6]);
  buf(\uc8051golden_1.PSW_2c [7], \uc8051golden_1.n1292 [7]);
  buf(\uc8051golden_1.PSW_2d [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2d [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2d [2], \uc8051golden_1.n1280 [2]);
  buf(\uc8051golden_1.PSW_2d [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2d [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2d [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2d [6], \uc8051golden_1.n1292 [6]);
  buf(\uc8051golden_1.PSW_2d [7], \uc8051golden_1.n1280 [7]);
  buf(\uc8051golden_1.PSW_2e [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2e [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2e [2], \uc8051golden_1.n1292 [2]);
  buf(\uc8051golden_1.PSW_2e [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2e [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2e [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2e [6], \uc8051golden_1.n1292 [6]);
  buf(\uc8051golden_1.PSW_2e [7], \uc8051golden_1.n1292 [7]);
  buf(\uc8051golden_1.PSW_2f [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2f [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2f [2], \uc8051golden_1.n1292 [2]);
  buf(\uc8051golden_1.PSW_2f [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2f [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2f [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2f [6], \uc8051golden_1.n1292 [6]);
  buf(\uc8051golden_1.PSW_2f [7], \uc8051golden_1.n1292 [7]);
  buf(\uc8051golden_1.PSW_33 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_33 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_33 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_33 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_33 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_33 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_33 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_33 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.PSW_34 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_34 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_34 [2], \uc8051golden_1.n1318 [2]);
  buf(\uc8051golden_1.PSW_34 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_34 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_34 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_34 [6], \uc8051golden_1.n1318 [6]);
  buf(\uc8051golden_1.PSW_34 [7], \uc8051golden_1.n1318 [7]);
  buf(\uc8051golden_1.PSW_35 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_35 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_35 [2], \uc8051golden_1.n1334 [2]);
  buf(\uc8051golden_1.PSW_35 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_35 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_35 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_35 [6], \uc8051golden_1.n1334 [6]);
  buf(\uc8051golden_1.PSW_35 [7], \uc8051golden_1.n1334 [7]);
  buf(\uc8051golden_1.PSW_36 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_36 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_36 [2], \uc8051golden_1.n1350 [2]);
  buf(\uc8051golden_1.PSW_36 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_36 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_36 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_36 [6], \uc8051golden_1.n1350 [6]);
  buf(\uc8051golden_1.PSW_36 [7], \uc8051golden_1.n1350 [7]);
  buf(\uc8051golden_1.PSW_37 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_37 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_37 [2], \uc8051golden_1.n1350 [2]);
  buf(\uc8051golden_1.PSW_37 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_37 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_37 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_37 [6], \uc8051golden_1.n1350 [6]);
  buf(\uc8051golden_1.PSW_37 [7], \uc8051golden_1.n1350 [7]);
  buf(\uc8051golden_1.PSW_38 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_38 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_38 [2], \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.PSW_38 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_38 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_38 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_38 [6], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.PSW_38 [7], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.PSW_39 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_39 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_39 [2], \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.PSW_39 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_39 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_39 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_39 [6], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.PSW_39 [7], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.PSW_3a [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3a [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3a [2], \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.PSW_3a [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3a [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3a [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3a [6], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.PSW_3a [7], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.PSW_3b [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3b [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3b [2], \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.PSW_3b [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3b [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3b [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3b [6], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.PSW_3b [7], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.PSW_3c [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3c [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3c [2], \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.PSW_3c [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3c [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3c [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3c [6], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.PSW_3c [7], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.PSW_3d [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3d [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3d [2], \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.PSW_3d [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3d [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3d [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3d [6], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.PSW_3d [7], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.PSW_3e [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3e [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3e [2], \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.PSW_3e [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3e [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3e [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3e [6], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.PSW_3e [7], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.PSW_3f [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3f [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3f [2], \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.PSW_3f [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3f [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3f [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3f [6], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.PSW_3f [7], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.PSW_72 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_72 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_72 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_72 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_72 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_72 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_72 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_72 [7], \uc8051golden_1.n1522 [7]);
  buf(\uc8051golden_1.PSW_82 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_82 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_82 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_82 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_82 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_82 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_82 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_82 [7], \uc8051golden_1.n1546 [7]);
  buf(\uc8051golden_1.PSW_84 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_84 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_84 [2], \uc8051golden_1.n1555 [2]);
  buf(\uc8051golden_1.PSW_84 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_84 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_84 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_84 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_84 [7], 1'b0);
  buf(\uc8051golden_1.PSW_94 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_94 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_94 [2], \uc8051golden_1.n1692 [2]);
  buf(\uc8051golden_1.PSW_94 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_94 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_94 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_94 [6], \uc8051golden_1.n1692 [6]);
  buf(\uc8051golden_1.PSW_94 [7], \uc8051golden_1.n1692 [7]);
  buf(\uc8051golden_1.PSW_95 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_95 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_95 [2], \uc8051golden_1.n1705 [2]);
  buf(\uc8051golden_1.PSW_95 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_95 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_95 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_95 [6], \uc8051golden_1.n1705 [6]);
  buf(\uc8051golden_1.PSW_95 [7], \uc8051golden_1.n1705 [7]);
  buf(\uc8051golden_1.PSW_96 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_96 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_96 [2], \uc8051golden_1.n1718 [2]);
  buf(\uc8051golden_1.PSW_96 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_96 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_96 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_96 [6], \uc8051golden_1.n1718 [6]);
  buf(\uc8051golden_1.PSW_96 [7], \uc8051golden_1.n1718 [7]);
  buf(\uc8051golden_1.PSW_97 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_97 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_97 [2], \uc8051golden_1.n1718 [2]);
  buf(\uc8051golden_1.PSW_97 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_97 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_97 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_97 [6], \uc8051golden_1.n1718 [6]);
  buf(\uc8051golden_1.PSW_97 [7], \uc8051golden_1.n1718 [7]);
  buf(\uc8051golden_1.PSW_98 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_98 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_98 [2], \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.PSW_98 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_98 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_98 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_98 [6], \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.PSW_98 [7], \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.PSW_99 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_99 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_99 [2], \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.PSW_99 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_99 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_99 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_99 [6], \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.PSW_99 [7], \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.PSW_9a [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9a [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9a [2], \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.PSW_9a [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9a [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9a [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9a [6], \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.PSW_9a [7], \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.PSW_9b [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9b [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9b [2], \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.PSW_9b [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9b [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9b [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9b [6], \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.PSW_9b [7], \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.PSW_9c [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9c [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9c [2], \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.PSW_9c [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9c [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9c [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9c [6], \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.PSW_9c [7], \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.PSW_9d [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9d [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9d [2], \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.PSW_9d [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9d [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9d [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9d [6], \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.PSW_9d [7], \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.PSW_9e [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9e [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9e [2], \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.PSW_9e [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9e [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9e [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9e [6], \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.PSW_9e [7], \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.PSW_9f [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9f [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9f [2], \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.PSW_9f [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9f [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9f [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9f [6], \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.PSW_9f [7], \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.PSW_a0 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_a0 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_a0 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_a0 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_a0 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_a0 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_a0 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_a0 [7], \uc8051golden_1.n1734 [7]);
  buf(\uc8051golden_1.PSW_a2 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_a2 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_a2 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_a2 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_a2 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_a2 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_a2 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_a2 [7], \uc8051golden_1.n1735 [7]);
  buf(\uc8051golden_1.PSW_a4 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_a4 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_a4 [2], \uc8051golden_1.n1746 [2]);
  buf(\uc8051golden_1.PSW_a4 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_a4 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_a4 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_a4 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_a4 [7], 1'b0);
  buf(\uc8051golden_1.PSW_b0 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b0 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b0 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b0 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b0 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b0 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b0 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b0 [7], \uc8051golden_1.n1750 [7]);
  buf(\uc8051golden_1.PSW_b3 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b3 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b3 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b3 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b3 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b3 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b3 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b3 [7], \uc8051golden_1.n1766 [7]);
  buf(\uc8051golden_1.PSW_b4 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b4 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b4 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b4 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b4 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b4 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b4 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b4 [7], \uc8051golden_1.n1772 [7]);
  buf(\uc8051golden_1.PSW_b5 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b5 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b5 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b5 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b5 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b5 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b5 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b5 [7], \uc8051golden_1.n1778 [7]);
  buf(\uc8051golden_1.PSW_b6 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b6 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b6 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b6 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b6 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b6 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b6 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b6 [7], \uc8051golden_1.n1784 [7]);
  buf(\uc8051golden_1.PSW_b7 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b7 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b7 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b7 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b7 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b7 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b7 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b7 [7], \uc8051golden_1.n1784 [7]);
  buf(\uc8051golden_1.PSW_b8 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b8 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b8 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b8 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b8 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b8 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b8 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b8 [7], \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.PSW_b9 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b9 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b9 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b9 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b9 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b9 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b9 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b9 [7], \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.PSW_ba [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_ba [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_ba [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_ba [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_ba [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_ba [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_ba [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_ba [7], \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.PSW_bb [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_bb [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_bb [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_bb [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_bb [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_bb [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_bb [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_bb [7], \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.PSW_bc [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_bc [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_bc [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_bc [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_bc [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_bc [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_bc [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_bc [7], \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.PSW_bd [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_bd [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_bd [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_bd [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_bd [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_bd [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_bd [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_bd [7], \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.PSW_be [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_be [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_be [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_be [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_be [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_be [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_be [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_be [7], \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.PSW_bf [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_bf [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_bf [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_bf [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_bf [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_bf [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_bf [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_bf [7], \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.PSW_c3 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_c3 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_c3 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_c3 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_c3 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_c3 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_c3 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_c3 [7], 1'b0);
  buf(\uc8051golden_1.PSW_d3 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_d3 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_d3 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_d3 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_d3 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_d3 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_d3 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_d3 [7], 1'b1);
  buf(\uc8051golden_1.PSW_d4 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_d4 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_d4 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_d4 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_d4 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_d4 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_d4 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_d4 [7], \uc8051golden_1.n1848 [7]);
  buf(\uc8051golden_1.RD_IRAM_0 [0], \uc8051golden_1.n1268 [0]);
  buf(\uc8051golden_1.RD_IRAM_0 [1], \uc8051golden_1.n1268 [1]);
  buf(\uc8051golden_1.RD_IRAM_0 [2], \uc8051golden_1.n1268 [2]);
  buf(\uc8051golden_1.RD_IRAM_0 [3], \uc8051golden_1.n1268 [3]);
  buf(\uc8051golden_1.RD_IRAM_0 [4], \uc8051golden_1.n1268 [4]);
  buf(\uc8051golden_1.RD_IRAM_0 [5], \uc8051golden_1.n1268 [5]);
  buf(\uc8051golden_1.RD_IRAM_0 [6], \uc8051golden_1.n1268 [6]);
  buf(\uc8051golden_1.RD_IRAM_0 [7], \uc8051golden_1.n1268 [8]);
  buf(\uc8051golden_1.RD_IRAM_1 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.RD_IRAM_1 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.RD_IRAM_1 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.RD_IRAM_1 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.RD_IRAM_1 [4], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.RD_IRAM_1 [5], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.RD_IRAM_1 [6], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.RD_IRAM_1 [7], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.n0006 [0], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0006 [1], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0007 [0], 1'b0);
  buf(\uc8051golden_1.n0007 [1], 1'b0);
  buf(\uc8051golden_1.n0007 [2], 1'b0);
  buf(\uc8051golden_1.n0007 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0007 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0007 [5], 1'b0);
  buf(\uc8051golden_1.n0007 [6], 1'b0);
  buf(\uc8051golden_1.n0007 [7], 1'b0);
  buf(\uc8051golden_1.n0011 [0], 1'b1);
  buf(\uc8051golden_1.n0011 [1], 1'b0);
  buf(\uc8051golden_1.n0011 [2], 1'b0);
  buf(\uc8051golden_1.n0011 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0011 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0011 [5], 1'b0);
  buf(\uc8051golden_1.n0011 [6], 1'b0);
  buf(\uc8051golden_1.n0011 [7], 1'b0);
  buf(\uc8051golden_1.n0019 [0], 1'b0);
  buf(\uc8051golden_1.n0019 [1], 1'b1);
  buf(\uc8051golden_1.n0019 [2], 1'b0);
  buf(\uc8051golden_1.n0019 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0019 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0019 [5], 1'b0);
  buf(\uc8051golden_1.n0019 [6], 1'b0);
  buf(\uc8051golden_1.n0019 [7], 1'b0);
  buf(\uc8051golden_1.n0023 [0], 1'b1);
  buf(\uc8051golden_1.n0023 [1], 1'b1);
  buf(\uc8051golden_1.n0023 [2], 1'b0);
  buf(\uc8051golden_1.n0023 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0023 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0023 [5], 1'b0);
  buf(\uc8051golden_1.n0023 [6], 1'b0);
  buf(\uc8051golden_1.n0023 [7], 1'b0);
  buf(\uc8051golden_1.n0027 [0], 1'b0);
  buf(\uc8051golden_1.n0027 [1], 1'b0);
  buf(\uc8051golden_1.n0027 [2], 1'b1);
  buf(\uc8051golden_1.n0027 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0027 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0027 [5], 1'b0);
  buf(\uc8051golden_1.n0027 [6], 1'b0);
  buf(\uc8051golden_1.n0027 [7], 1'b0);
  buf(\uc8051golden_1.n0031 [0], 1'b1);
  buf(\uc8051golden_1.n0031 [1], 1'b0);
  buf(\uc8051golden_1.n0031 [2], 1'b1);
  buf(\uc8051golden_1.n0031 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0031 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0031 [5], 1'b0);
  buf(\uc8051golden_1.n0031 [6], 1'b0);
  buf(\uc8051golden_1.n0031 [7], 1'b0);
  buf(\uc8051golden_1.n0035 [0], 1'b0);
  buf(\uc8051golden_1.n0035 [1], 1'b1);
  buf(\uc8051golden_1.n0035 [2], 1'b1);
  buf(\uc8051golden_1.n0035 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0035 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0035 [5], 1'b0);
  buf(\uc8051golden_1.n0035 [6], 1'b0);
  buf(\uc8051golden_1.n0035 [7], 1'b0);
  buf(\uc8051golden_1.n0039 [0], 1'b1);
  buf(\uc8051golden_1.n0039 [1], 1'b1);
  buf(\uc8051golden_1.n0039 [2], 1'b1);
  buf(\uc8051golden_1.n0039 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0039 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0039 [5], 1'b0);
  buf(\uc8051golden_1.n0039 [6], 1'b0);
  buf(\uc8051golden_1.n0039 [7], 1'b0);
  buf(\uc8051golden_1.n0561 [0], \uc8051golden_1.n1268 [0]);
  buf(\uc8051golden_1.n0561 [1], \uc8051golden_1.n1268 [1]);
  buf(\uc8051golden_1.n0561 [2], \uc8051golden_1.n1268 [2]);
  buf(\uc8051golden_1.n0561 [3], \uc8051golden_1.n1268 [3]);
  buf(\uc8051golden_1.n0561 [4], \uc8051golden_1.n1268 [4]);
  buf(\uc8051golden_1.n0561 [5], \uc8051golden_1.n1268 [5]);
  buf(\uc8051golden_1.n0561 [6], \uc8051golden_1.n1268 [6]);
  buf(\uc8051golden_1.n0561 [7], \uc8051golden_1.n1268 [8]);
  buf(\uc8051golden_1.n0594 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.n0594 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.n0594 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.n0594 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.n0594 [4], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.n0594 [5], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.n0594 [6], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.n0594 [7], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.n0701 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0701 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0701 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0701 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0701 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0701 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0701 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0701 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0701 [8], 1'b0);
  buf(\uc8051golden_1.n0701 [9], 1'b0);
  buf(\uc8051golden_1.n0701 [10], 1'b0);
  buf(\uc8051golden_1.n0701 [11], 1'b0);
  buf(\uc8051golden_1.n0701 [12], 1'b0);
  buf(\uc8051golden_1.n0701 [13], 1'b0);
  buf(\uc8051golden_1.n0701 [14], 1'b0);
  buf(\uc8051golden_1.n0701 [15], 1'b0);
  buf(\uc8051golden_1.n0733 [0], \uc8051golden_1.DPL [0]);
  buf(\uc8051golden_1.n0733 [1], \uc8051golden_1.DPL [1]);
  buf(\uc8051golden_1.n0733 [2], \uc8051golden_1.DPL [2]);
  buf(\uc8051golden_1.n0733 [3], \uc8051golden_1.DPL [3]);
  buf(\uc8051golden_1.n0733 [4], \uc8051golden_1.DPL [4]);
  buf(\uc8051golden_1.n0733 [5], \uc8051golden_1.DPL [5]);
  buf(\uc8051golden_1.n0733 [6], \uc8051golden_1.DPL [6]);
  buf(\uc8051golden_1.n0733 [7], \uc8051golden_1.DPL [7]);
  buf(\uc8051golden_1.n0733 [8], \uc8051golden_1.DPH [0]);
  buf(\uc8051golden_1.n0733 [9], \uc8051golden_1.DPH [1]);
  buf(\uc8051golden_1.n0733 [10], \uc8051golden_1.DPH [2]);
  buf(\uc8051golden_1.n0733 [11], \uc8051golden_1.DPH [3]);
  buf(\uc8051golden_1.n0733 [12], \uc8051golden_1.DPH [4]);
  buf(\uc8051golden_1.n0733 [13], \uc8051golden_1.DPH [5]);
  buf(\uc8051golden_1.n0733 [14], \uc8051golden_1.DPH [6]);
  buf(\uc8051golden_1.n0733 [15], \uc8051golden_1.DPH [7]);
  buf(\uc8051golden_1.n0994 [0], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0994 [1], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0994 [2], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0994 [3], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0994 [4], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0994 [5], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0994 [6], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0994 [7], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1071 [0], \uc8051golden_1.n1268 [0]);
  buf(\uc8051golden_1.n1071 [1], \uc8051golden_1.n1268 [1]);
  buf(\uc8051golden_1.n1071 [2], \uc8051golden_1.n1268 [2]);
  buf(\uc8051golden_1.n1071 [3], \uc8051golden_1.n1268 [3]);
  buf(\uc8051golden_1.n1073 [0], 1'b0);
  buf(\uc8051golden_1.n1073 [1], 1'b0);
  buf(\uc8051golden_1.n1073 [2], 1'b0);
  buf(\uc8051golden_1.n1073 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1075 [0], 1'b1);
  buf(\uc8051golden_1.n1075 [1], 1'b0);
  buf(\uc8051golden_1.n1075 [2], 1'b0);
  buf(\uc8051golden_1.n1075 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1076 [0], 1'b0);
  buf(\uc8051golden_1.n1076 [1], 1'b1);
  buf(\uc8051golden_1.n1076 [2], 1'b0);
  buf(\uc8051golden_1.n1076 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1077 [0], 1'b1);
  buf(\uc8051golden_1.n1077 [1], 1'b1);
  buf(\uc8051golden_1.n1077 [2], 1'b0);
  buf(\uc8051golden_1.n1077 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1078 [0], 1'b0);
  buf(\uc8051golden_1.n1078 [1], 1'b0);
  buf(\uc8051golden_1.n1078 [2], 1'b1);
  buf(\uc8051golden_1.n1078 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1079 [0], 1'b1);
  buf(\uc8051golden_1.n1079 [1], 1'b0);
  buf(\uc8051golden_1.n1079 [2], 1'b1);
  buf(\uc8051golden_1.n1079 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1080 [0], 1'b0);
  buf(\uc8051golden_1.n1080 [1], 1'b1);
  buf(\uc8051golden_1.n1080 [2], 1'b1);
  buf(\uc8051golden_1.n1080 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1081 [0], 1'b1);
  buf(\uc8051golden_1.n1081 [1], 1'b1);
  buf(\uc8051golden_1.n1081 [2], 1'b1);
  buf(\uc8051golden_1.n1081 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1118 , \uc8051golden_1.n1735 [7]);
  buf(\uc8051golden_1.n1146 , \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1147 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1147 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1147 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1147 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1147 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1147 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1147 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1147 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1147 [8], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1148 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1148 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1148 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1148 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1148 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1148 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1148 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1148 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1148 [8], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1149 [0], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1149 [1], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1149 [2], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1149 [3], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1149 [4], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1149 [5], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1149 [6], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1149 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1150 , \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1151 , \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1152 [0], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1152 [1], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1152 [2], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1153 , \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1154 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1154 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1155 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1155 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1155 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1155 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1155 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1155 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1155 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1155 [7], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1181 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.n1181 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.n1181 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.n1181 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.n1181 [4], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.n1181 [5], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.n1181 [6], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.n1181 [7], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.n1181 [8], \uc8051golden_1.n1268 [0]);
  buf(\uc8051golden_1.n1181 [9], \uc8051golden_1.n1268 [1]);
  buf(\uc8051golden_1.n1181 [10], \uc8051golden_1.n1268 [2]);
  buf(\uc8051golden_1.n1181 [11], \uc8051golden_1.n1268 [3]);
  buf(\uc8051golden_1.n1181 [12], \uc8051golden_1.n1268 [4]);
  buf(\uc8051golden_1.n1181 [13], \uc8051golden_1.n1268 [5]);
  buf(\uc8051golden_1.n1181 [14], \uc8051golden_1.n1268 [6]);
  buf(\uc8051golden_1.n1181 [15], \uc8051golden_1.n1268 [8]);
  buf(\uc8051golden_1.n1183 [0], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1183 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1183 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1183 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1183 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1183 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1183 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1183 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1185 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1185 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1185 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1185 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1185 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1185 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1185 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1185 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1185 [8], 1'b0);
  buf(\uc8051golden_1.n1189 [8], \uc8051golden_1.n1207 [7]);
  buf(\uc8051golden_1.n1190 , \uc8051golden_1.n1207 [7]);
  buf(\uc8051golden_1.n1191 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1191 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1191 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1191 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1192 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1192 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1192 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1192 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1192 [4], 1'b0);
  buf(\uc8051golden_1.n1196 [4], \uc8051golden_1.n1207 [6]);
  buf(\uc8051golden_1.n1197 , \uc8051golden_1.n1207 [6]);
  buf(\uc8051golden_1.n1198 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1198 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1198 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1198 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1198 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1198 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1198 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1198 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1198 [8], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1206 , \uc8051golden_1.n1207 [2]);
  buf(\uc8051golden_1.n1207 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1207 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1207 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1207 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1207 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1211 [8], \uc8051golden_1.n1227 [7]);
  buf(\uc8051golden_1.n1212 , \uc8051golden_1.n1227 [7]);
  buf(\uc8051golden_1.n1217 [4], \uc8051golden_1.n1227 [6]);
  buf(\uc8051golden_1.n1218 , \uc8051golden_1.n1227 [6]);
  buf(\uc8051golden_1.n1226 , \uc8051golden_1.n1227 [2]);
  buf(\uc8051golden_1.n1227 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1227 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1227 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1227 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1227 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1229 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.n1229 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.n1229 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.n1229 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.n1229 [4], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.n1229 [5], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.n1229 [6], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.n1229 [7], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.n1229 [8], 1'b0);
  buf(\uc8051golden_1.n1231 [8], \uc8051golden_1.n1246 [7]);
  buf(\uc8051golden_1.n1232 , \uc8051golden_1.n1246 [7]);
  buf(\uc8051golden_1.n1233 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.n1233 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.n1233 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.n1233 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.n1234 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.n1234 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.n1234 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.n1234 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.n1234 [4], 1'b0);
  buf(\uc8051golden_1.n1236 [4], \uc8051golden_1.n1258 [6]);
  buf(\uc8051golden_1.n1237 , \uc8051golden_1.n1258 [6]);
  buf(\uc8051golden_1.n1238 [0], \uc8051golden_1.n1852 [0]);
  buf(\uc8051golden_1.n1238 [1], \uc8051golden_1.n1852 [1]);
  buf(\uc8051golden_1.n1238 [2], \uc8051golden_1.n1852 [2]);
  buf(\uc8051golden_1.n1238 [3], \uc8051golden_1.n1852 [3]);
  buf(\uc8051golden_1.n1238 [4], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.n1238 [5], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.n1238 [6], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.n1238 [7], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.n1238 [8], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.n1245 , \uc8051golden_1.n1246 [2]);
  buf(\uc8051golden_1.n1246 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1246 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1246 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1246 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1246 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1246 [6], \uc8051golden_1.n1258 [6]);
  buf(\uc8051golden_1.n1249 [8], \uc8051golden_1.n1258 [7]);
  buf(\uc8051golden_1.n1250 , \uc8051golden_1.n1258 [7]);
  buf(\uc8051golden_1.n1257 , \uc8051golden_1.n1258 [2]);
  buf(\uc8051golden_1.n1258 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1258 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1258 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1258 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1258 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1260 [0], \uc8051golden_1.n1268 [0]);
  buf(\uc8051golden_1.n1260 [1], \uc8051golden_1.n1268 [1]);
  buf(\uc8051golden_1.n1260 [2], \uc8051golden_1.n1268 [2]);
  buf(\uc8051golden_1.n1260 [3], \uc8051golden_1.n1268 [3]);
  buf(\uc8051golden_1.n1260 [4], \uc8051golden_1.n1268 [4]);
  buf(\uc8051golden_1.n1260 [5], \uc8051golden_1.n1268 [5]);
  buf(\uc8051golden_1.n1260 [6], \uc8051golden_1.n1268 [6]);
  buf(\uc8051golden_1.n1260 [7], \uc8051golden_1.n1268 [8]);
  buf(\uc8051golden_1.n1260 [8], 1'b0);
  buf(\uc8051golden_1.n1262 [8], \uc8051golden_1.n1280 [7]);
  buf(\uc8051golden_1.n1263 , \uc8051golden_1.n1280 [7]);
  buf(\uc8051golden_1.n1264 [0], \uc8051golden_1.n1268 [0]);
  buf(\uc8051golden_1.n1264 [1], \uc8051golden_1.n1268 [1]);
  buf(\uc8051golden_1.n1264 [2], \uc8051golden_1.n1268 [2]);
  buf(\uc8051golden_1.n1264 [3], \uc8051golden_1.n1268 [3]);
  buf(\uc8051golden_1.n1264 [4], 1'b0);
  buf(\uc8051golden_1.n1266 [4], \uc8051golden_1.n1292 [6]);
  buf(\uc8051golden_1.n1267 , \uc8051golden_1.n1292 [6]);
  buf(\uc8051golden_1.n1268 [7], \uc8051golden_1.n1268 [8]);
  buf(\uc8051golden_1.n1275 , \uc8051golden_1.n1280 [2]);
  buf(\uc8051golden_1.n1276 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1276 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1276 [2], \uc8051golden_1.n1280 [2]);
  buf(\uc8051golden_1.n1276 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1276 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1276 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1276 [6], \uc8051golden_1.n1292 [6]);
  buf(\uc8051golden_1.n1276 [7], \uc8051golden_1.n1280 [7]);
  buf(\uc8051golden_1.n1278 [4], \uc8051golden_1.n1291 [6]);
  buf(\uc8051golden_1.n1279 , \uc8051golden_1.n1291 [6]);
  buf(\uc8051golden_1.n1280 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1280 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1280 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1280 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1280 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1280 [6], \uc8051golden_1.n1291 [6]);
  buf(\uc8051golden_1.n1282 [8], \uc8051golden_1.n1292 [7]);
  buf(\uc8051golden_1.n1283 , \uc8051golden_1.n1292 [7]);
  buf(\uc8051golden_1.n1290 , \uc8051golden_1.n1292 [2]);
  buf(\uc8051golden_1.n1291 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1291 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1291 [2], \uc8051golden_1.n1292 [2]);
  buf(\uc8051golden_1.n1291 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1291 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1291 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1291 [7], \uc8051golden_1.n1292 [7]);
  buf(\uc8051golden_1.n1292 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1292 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1292 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1292 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1292 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1295 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1295 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1295 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1295 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1295 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1295 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1295 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1295 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1295 [8], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1296 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1296 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1296 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1296 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1296 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1296 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1296 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1296 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1296 [8], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1297 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1297 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1297 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1297 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1297 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1297 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1297 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1297 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1298 , \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1299 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1299 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1299 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1299 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1299 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1299 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1299 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1299 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1300 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1300 [1], 1'b0);
  buf(\uc8051golden_1.n1300 [2], 1'b0);
  buf(\uc8051golden_1.n1300 [3], 1'b0);
  buf(\uc8051golden_1.n1300 [4], 1'b0);
  buf(\uc8051golden_1.n1300 [5], 1'b0);
  buf(\uc8051golden_1.n1300 [6], 1'b0);
  buf(\uc8051golden_1.n1300 [7], 1'b0);
  buf(\uc8051golden_1.n1303 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1303 [1], 1'b0);
  buf(\uc8051golden_1.n1303 [2], 1'b0);
  buf(\uc8051golden_1.n1303 [3], 1'b0);
  buf(\uc8051golden_1.n1303 [4], 1'b0);
  buf(\uc8051golden_1.n1303 [5], 1'b0);
  buf(\uc8051golden_1.n1303 [6], 1'b0);
  buf(\uc8051golden_1.n1303 [7], 1'b0);
  buf(\uc8051golden_1.n1303 [8], 1'b0);
  buf(\uc8051golden_1.n1305 [8], \uc8051golden_1.n1318 [7]);
  buf(\uc8051golden_1.n1306 , \uc8051golden_1.n1318 [7]);
  buf(\uc8051golden_1.n1307 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1307 [1], 1'b0);
  buf(\uc8051golden_1.n1307 [2], 1'b0);
  buf(\uc8051golden_1.n1307 [3], 1'b0);
  buf(\uc8051golden_1.n1307 [4], 1'b0);
  buf(\uc8051golden_1.n1309 [4], \uc8051golden_1.n1318 [6]);
  buf(\uc8051golden_1.n1310 , \uc8051golden_1.n1318 [6]);
  buf(\uc8051golden_1.n1317 , \uc8051golden_1.n1318 [2]);
  buf(\uc8051golden_1.n1318 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1318 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1318 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1318 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1318 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1322 [8], \uc8051golden_1.n1334 [7]);
  buf(\uc8051golden_1.n1323 , \uc8051golden_1.n1334 [7]);
  buf(\uc8051golden_1.n1325 [4], \uc8051golden_1.n1334 [6]);
  buf(\uc8051golden_1.n1326 , \uc8051golden_1.n1334 [6]);
  buf(\uc8051golden_1.n1333 , \uc8051golden_1.n1334 [2]);
  buf(\uc8051golden_1.n1334 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1334 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1334 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1334 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1334 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1338 [8], \uc8051golden_1.n1350 [7]);
  buf(\uc8051golden_1.n1339 , \uc8051golden_1.n1350 [7]);
  buf(\uc8051golden_1.n1341 [4], \uc8051golden_1.n1350 [6]);
  buf(\uc8051golden_1.n1342 , \uc8051golden_1.n1350 [6]);
  buf(\uc8051golden_1.n1349 , \uc8051golden_1.n1350 [2]);
  buf(\uc8051golden_1.n1350 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1350 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1350 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1350 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1350 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1354 [8], \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.n1355 , \uc8051golden_1.n1366 [7]);
  buf(\uc8051golden_1.n1357 [4], \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.n1358 , \uc8051golden_1.n1366 [6]);
  buf(\uc8051golden_1.n1365 , \uc8051golden_1.n1366 [2]);
  buf(\uc8051golden_1.n1366 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1366 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1366 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1366 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1366 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1520 , \uc8051golden_1.n1522 [7]);
  buf(\uc8051golden_1.n1521 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1521 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1521 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1521 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1521 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1521 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1521 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1522 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1522 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1522 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1522 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1522 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1522 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1522 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1545 , \uc8051golden_1.n1546 [7]);
  buf(\uc8051golden_1.n1546 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1546 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1546 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1546 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1546 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1546 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1546 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1553 [0], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1553 [1], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1553 [2], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1553 [3], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1554 , \uc8051golden_1.n1555 [2]);
  buf(\uc8051golden_1.n1555 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1555 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1555 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1555 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1555 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1555 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1555 [7], 1'b0);
  buf(\uc8051golden_1.n1680 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1680 [1], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1680 [2], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1680 [3], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1680 [4], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1680 [5], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1680 [6], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1680 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1683 , \uc8051golden_1.n1692 [7]);
  buf(\uc8051golden_1.n1685 , \uc8051golden_1.n1692 [6]);
  buf(\uc8051golden_1.n1691 , \uc8051golden_1.n1692 [2]);
  buf(\uc8051golden_1.n1692 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1692 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1692 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1692 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1692 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1696 , \uc8051golden_1.n1705 [7]);
  buf(\uc8051golden_1.n1698 , \uc8051golden_1.n1705 [6]);
  buf(\uc8051golden_1.n1704 , \uc8051golden_1.n1705 [2]);
  buf(\uc8051golden_1.n1705 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1705 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1705 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1705 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1705 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1709 , \uc8051golden_1.n1718 [7]);
  buf(\uc8051golden_1.n1711 , \uc8051golden_1.n1718 [6]);
  buf(\uc8051golden_1.n1717 , \uc8051golden_1.n1718 [2]);
  buf(\uc8051golden_1.n1718 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1718 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1718 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1718 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1718 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1722 , \uc8051golden_1.n1731 [7]);
  buf(\uc8051golden_1.n1724 , \uc8051golden_1.n1731 [6]);
  buf(\uc8051golden_1.n1730 , \uc8051golden_1.n1731 [2]);
  buf(\uc8051golden_1.n1731 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1731 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1731 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1731 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1731 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1733 , \uc8051golden_1.n1734 [7]);
  buf(\uc8051golden_1.n1734 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1734 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1734 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1734 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1734 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1734 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1734 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1735 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1735 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1735 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1735 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1735 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1735 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1735 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1739 [0], \uc8051golden_1.B [0]);
  buf(\uc8051golden_1.n1739 [1], \uc8051golden_1.B [1]);
  buf(\uc8051golden_1.n1739 [2], \uc8051golden_1.B [2]);
  buf(\uc8051golden_1.n1739 [3], \uc8051golden_1.B [3]);
  buf(\uc8051golden_1.n1739 [4], \uc8051golden_1.B [4]);
  buf(\uc8051golden_1.n1739 [5], \uc8051golden_1.B [5]);
  buf(\uc8051golden_1.n1739 [6], \uc8051golden_1.B [6]);
  buf(\uc8051golden_1.n1739 [7], \uc8051golden_1.B [7]);
  buf(\uc8051golden_1.n1739 [8], 1'b0);
  buf(\uc8051golden_1.n1739 [9], 1'b0);
  buf(\uc8051golden_1.n1739 [10], 1'b0);
  buf(\uc8051golden_1.n1739 [11], 1'b0);
  buf(\uc8051golden_1.n1739 [12], 1'b0);
  buf(\uc8051golden_1.n1739 [13], 1'b0);
  buf(\uc8051golden_1.n1739 [14], 1'b0);
  buf(\uc8051golden_1.n1739 [15], 1'b0);
  buf(\uc8051golden_1.n1745 , \uc8051golden_1.n1746 [2]);
  buf(\uc8051golden_1.n1746 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1746 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1746 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1746 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1746 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1746 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1746 [7], 1'b0);
  buf(\uc8051golden_1.n1749 , \uc8051golden_1.n1750 [7]);
  buf(\uc8051golden_1.n1750 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1750 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1750 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1750 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1750 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1750 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1750 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1765 , \uc8051golden_1.n1766 [7]);
  buf(\uc8051golden_1.n1766 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1766 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1766 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1766 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1766 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1766 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1766 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1771 , \uc8051golden_1.n1772 [7]);
  buf(\uc8051golden_1.n1772 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1772 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1772 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1772 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1772 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1772 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1772 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1777 , \uc8051golden_1.n1778 [7]);
  buf(\uc8051golden_1.n1778 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1778 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1778 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1778 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1778 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1778 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1778 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1783 , \uc8051golden_1.n1784 [7]);
  buf(\uc8051golden_1.n1784 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1784 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1784 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1784 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1784 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1784 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1784 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1789 , \uc8051golden_1.n1790 [7]);
  buf(\uc8051golden_1.n1790 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1790 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1790 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1790 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1790 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1790 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1790 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1791 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1791 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1791 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1791 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1791 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1791 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1791 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1791 [7], 1'b0);
  buf(\uc8051golden_1.n1792 [0], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1792 [1], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1792 [2], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1792 [3], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1793 [0], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1793 [1], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1793 [2], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1793 [3], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1793 [4], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1793 [5], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1793 [6], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1793 [7], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1828 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1828 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1828 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1828 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1828 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1828 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1828 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1828 [7], 1'b1);
  buf(\uc8051golden_1.n1847 , \uc8051golden_1.n1848 [7]);
  buf(\uc8051golden_1.n1848 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1848 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1848 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1848 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1848 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1848 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1848 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1852 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1852 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1852 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1852 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1853 [0], \uc8051golden_1.n1854 [4]);
  buf(\uc8051golden_1.n1853 [1], \uc8051golden_1.n1854 [5]);
  buf(\uc8051golden_1.n1853 [2], \uc8051golden_1.n1854 [6]);
  buf(\uc8051golden_1.n1853 [3], \uc8051golden_1.n1854 [7]);
  buf(\uc8051golden_1.n1854 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1854 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1854 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1854 [3], \uc8051golden_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_rom_0_addr[0], \uc8051golden_1.PC [0]);
  buf(rd_rom_0_addr[1], \uc8051golden_1.PC [1]);
  buf(rd_rom_0_addr[2], \uc8051golden_1.PC [2]);
  buf(rd_rom_0_addr[3], \uc8051golden_1.PC [3]);
  buf(rd_rom_0_addr[4], \uc8051golden_1.PC [4]);
  buf(rd_rom_0_addr[5], \uc8051golden_1.PC [5]);
  buf(rd_rom_0_addr[6], \uc8051golden_1.PC [6]);
  buf(rd_rom_0_addr[7], \uc8051golden_1.PC [7]);
  buf(rd_rom_0_addr[8], \uc8051golden_1.PC [8]);
  buf(rd_rom_0_addr[9], \uc8051golden_1.PC [9]);
  buf(rd_rom_0_addr[10], \uc8051golden_1.PC [10]);
  buf(rd_rom_0_addr[11], \uc8051golden_1.PC [11]);
  buf(rd_rom_0_addr[12], \uc8051golden_1.PC [12]);
  buf(rd_rom_0_addr[13], \uc8051golden_1.PC [13]);
  buf(rd_rom_0_addr[14], \uc8051golden_1.PC [14]);
  buf(rd_rom_0_addr[15], \uc8051golden_1.PC [15]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
