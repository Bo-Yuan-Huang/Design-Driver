/** This is a highly unoptimized implementation of SHA1 by Forrest Heller.
  * Source: http://www.forrestheller.com/verilog/
  *         http://www.forrestheller.com/verilog/sha1.v
  *
  */

/*** SHA1 By Forrest Heller (2009) ***/
/* This code is based on the C SHA1 implementation as described in RFC 3174 */
/* round constants */
`define kzero 32'h5A827999
`define kone 32'h6ED9EBA1
`define ktwo 32'h8F1BBCDC
`define kthree 32'hCA62C1D6
`define SHA1CircularShift(bits,word) (((word)<<(bits))|((word)>>(32-(bits))))
module sha1(input wire [511:0] block ,
 input wire [159:0] current_hash,
 output wire [159:0] new_hash);

/*temporary wire variable to help with W initialization*/
wire [31:0] Wt [63:0];
/*mirrors W in SHA1 RFC reference*/
wire [31:0] W [79:0];
/* These variables mirror those in the SHA1 RFC reference*/
wire [31:0] temp [79:0];
wire [31:0] A [80:0];
wire [31:0] B [80:0];
wire [31:0] C [80:0];
wire [31:0] D [80:0];
wire [31:0] E [80:0];

 /* intialize first 16 words of W with the contents of block*/
assign W[0] = (block[31:24]) | (block[23:16] << 8) | (block[15:8] << 16) |( block[7:0] << 24);
assign W[1] = (block[63:56]) | (block[55:48] << 8) | (block[47:40] << 16) |( block[39:32] << 24);
assign W[2] = (block[95:88]) | (block[87:80] << 8) | (block[79:72] << 16) |( block[71:64] << 24);
assign W[3] = (block[127:120]) | (block[119:112] << 8) | (block[111:104] << 16) |( block[103:96] << 24);
assign W[4] = (block[159:152]) | (block[151:144] << 8) | (block[143:136] << 16) |( block[135:128] << 24);
assign W[5] = (block[191:184]) | (block[183:176] << 8) | (block[175:168] << 16) |( block[167:160] << 24);
assign W[6] = (block[223:216]) | (block[215:208] << 8) | (block[207:200] << 16) |( block[199:192] << 24);
assign W[7] = (block[255:248]) | (block[247:240] << 8) | (block[239:232] << 16) |( block[231:224] << 24);
assign W[8] = (block[287:280]) | (block[279:272] << 8) | (block[271:264] << 16) |( block[263:256] << 24);
assign W[9] = (block[319:312]) | (block[311:304] << 8) | (block[303:296] << 16) |( block[295:288] << 24);
assign W[10] = (block[351:344]) | (block[343:336] << 8) | (block[335:328] << 16) |( block[327:320] << 24);
assign W[11] = (block[383:376]) | (block[375:368] << 8) | (block[367:360] << 16) |( block[359:352] << 24);
assign W[12] = (block[415:408]) | (block[407:400] << 8) | (block[399:392] << 16) |( block[391:384] << 24);
assign W[13] = (block[447:440]) | (block[439:432] << 8) | (block[431:424] << 16) |( block[423:416] << 24);
assign W[14] = (block[479:472]) | (block[471:464] << 8) | (block[463:456] << 16) |( block[455:448] << 24);
assign W[15] = (block[511:504]) | (block[503:496] << 8) | (block[495:488] << 16) |( block[487:480] << 24);
/* initialize rest of W */
assign Wt[0]= W[13] ^ W[8] ^ W[2] ^ W[0];
assign W[16] = `SHA1CircularShift(1,Wt[0]);
assign Wt[1]= W[14] ^ W[9] ^ W[3] ^ W[1];
assign W[17] = `SHA1CircularShift(1,Wt[1]);
assign Wt[2]= W[15] ^ W[10] ^ W[4] ^ W[2];
assign W[18] = `SHA1CircularShift(1,Wt[2]);
assign Wt[3]= W[16] ^ W[11] ^ W[5] ^ W[3];
assign W[19] = `SHA1CircularShift(1,Wt[3]);
assign Wt[4]= W[17] ^ W[12] ^ W[6] ^ W[4];
assign W[20] = `SHA1CircularShift(1,Wt[4]);
assign Wt[5]= W[18] ^ W[13] ^ W[7] ^ W[5];
assign W[21] = `SHA1CircularShift(1,Wt[5]);
assign Wt[6]= W[19] ^ W[14] ^ W[8] ^ W[6];
assign W[22] = `SHA1CircularShift(1,Wt[6]);
assign Wt[7]= W[20] ^ W[15] ^ W[9] ^ W[7];
assign W[23] = `SHA1CircularShift(1,Wt[7]);
assign Wt[8]= W[21] ^ W[16] ^ W[10] ^ W[8];
assign W[24] = `SHA1CircularShift(1,Wt[8]);
assign Wt[9]= W[22] ^ W[17] ^ W[11] ^ W[9];
assign W[25] = `SHA1CircularShift(1,Wt[9]);
assign Wt[10]= W[23] ^ W[18] ^ W[12] ^ W[10];
assign W[26] = `SHA1CircularShift(1,Wt[10]);
assign Wt[11]= W[24] ^ W[19] ^ W[13] ^ W[11];
assign W[27] = `SHA1CircularShift(1,Wt[11]);
assign Wt[12]= W[25] ^ W[20] ^ W[14] ^ W[12];
assign W[28] = `SHA1CircularShift(1,Wt[12]);
assign Wt[13]= W[26] ^ W[21] ^ W[15] ^ W[13];
assign W[29] = `SHA1CircularShift(1,Wt[13]);
assign Wt[14]= W[27] ^ W[22] ^ W[16] ^ W[14];
assign W[30] = `SHA1CircularShift(1,Wt[14]);
assign Wt[15]= W[28] ^ W[23] ^ W[17] ^ W[15];
assign W[31] = `SHA1CircularShift(1,Wt[15]);
assign Wt[16]= W[29] ^ W[24] ^ W[18] ^ W[16];
assign W[32] = `SHA1CircularShift(1,Wt[16]);
assign Wt[17]= W[30] ^ W[25] ^ W[19] ^ W[17];
assign W[33] = `SHA1CircularShift(1,Wt[17]);
assign Wt[18]= W[31] ^ W[26] ^ W[20] ^ W[18];
assign W[34] = `SHA1CircularShift(1,Wt[18]);
assign Wt[19]= W[32] ^ W[27] ^ W[21] ^ W[19];
assign W[35] = `SHA1CircularShift(1,Wt[19]);
assign Wt[20]= W[33] ^ W[28] ^ W[22] ^ W[20];
assign W[36] = `SHA1CircularShift(1,Wt[20]);
assign Wt[21]= W[34] ^ W[29] ^ W[23] ^ W[21];
assign W[37] = `SHA1CircularShift(1,Wt[21]);
assign Wt[22]= W[35] ^ W[30] ^ W[24] ^ W[22];
assign W[38] = `SHA1CircularShift(1,Wt[22]);
assign Wt[23]= W[36] ^ W[31] ^ W[25] ^ W[23];
assign W[39] = `SHA1CircularShift(1,Wt[23]);
assign Wt[24]= W[37] ^ W[32] ^ W[26] ^ W[24];
assign W[40] = `SHA1CircularShift(1,Wt[24]);
assign Wt[25]= W[38] ^ W[33] ^ W[27] ^ W[25];
assign W[41] = `SHA1CircularShift(1,Wt[25]);
assign Wt[26]= W[39] ^ W[34] ^ W[28] ^ W[26];
assign W[42] = `SHA1CircularShift(1,Wt[26]);
assign Wt[27]= W[40] ^ W[35] ^ W[29] ^ W[27];
assign W[43] = `SHA1CircularShift(1,Wt[27]);
assign Wt[28]= W[41] ^ W[36] ^ W[30] ^ W[28];
assign W[44] = `SHA1CircularShift(1,Wt[28]);
assign Wt[29]= W[42] ^ W[37] ^ W[31] ^ W[29];
assign W[45] = `SHA1CircularShift(1,Wt[29]);
assign Wt[30]= W[43] ^ W[38] ^ W[32] ^ W[30];
assign W[46] = `SHA1CircularShift(1,Wt[30]);
assign Wt[31]= W[44] ^ W[39] ^ W[33] ^ W[31];
assign W[47] = `SHA1CircularShift(1,Wt[31]);
assign Wt[32]= W[45] ^ W[40] ^ W[34] ^ W[32];
assign W[48] = `SHA1CircularShift(1,Wt[32]);
assign Wt[33]= W[46] ^ W[41] ^ W[35] ^ W[33];
assign W[49] = `SHA1CircularShift(1,Wt[33]);
assign Wt[34]= W[47] ^ W[42] ^ W[36] ^ W[34];
assign W[50] = `SHA1CircularShift(1,Wt[34]);
assign Wt[35]= W[48] ^ W[43] ^ W[37] ^ W[35];
assign W[51] = `SHA1CircularShift(1,Wt[35]);
assign Wt[36]= W[49] ^ W[44] ^ W[38] ^ W[36];
assign W[52] = `SHA1CircularShift(1,Wt[36]);
assign Wt[37]= W[50] ^ W[45] ^ W[39] ^ W[37];
assign W[53] = `SHA1CircularShift(1,Wt[37]);
assign Wt[38]= W[51] ^ W[46] ^ W[40] ^ W[38];
assign W[54] = `SHA1CircularShift(1,Wt[38]);
assign Wt[39]= W[52] ^ W[47] ^ W[41] ^ W[39];
assign W[55] = `SHA1CircularShift(1,Wt[39]);
assign Wt[40]= W[53] ^ W[48] ^ W[42] ^ W[40];
assign W[56] = `SHA1CircularShift(1,Wt[40]);
assign Wt[41]= W[54] ^ W[49] ^ W[43] ^ W[41];
assign W[57] = `SHA1CircularShift(1,Wt[41]);
assign Wt[42]= W[55] ^ W[50] ^ W[44] ^ W[42];
assign W[58] = `SHA1CircularShift(1,Wt[42]);
assign Wt[43]= W[56] ^ W[51] ^ W[45] ^ W[43];
assign W[59] = `SHA1CircularShift(1,Wt[43]);
assign Wt[44]= W[57] ^ W[52] ^ W[46] ^ W[44];
assign W[60] = `SHA1CircularShift(1,Wt[44]);
assign Wt[45]= W[58] ^ W[53] ^ W[47] ^ W[45];
assign W[61] = `SHA1CircularShift(1,Wt[45]);
assign Wt[46]= W[59] ^ W[54] ^ W[48] ^ W[46];
assign W[62] = `SHA1CircularShift(1,Wt[46]);
assign Wt[47]= W[60] ^ W[55] ^ W[49] ^ W[47];
assign W[63] = `SHA1CircularShift(1,Wt[47]);
assign Wt[48]= W[61] ^ W[56] ^ W[50] ^ W[48];
assign W[64] = `SHA1CircularShift(1,Wt[48]);
assign Wt[49]= W[62] ^ W[57] ^ W[51] ^ W[49];
assign W[65] = `SHA1CircularShift(1,Wt[49]);
assign Wt[50]= W[63] ^ W[58] ^ W[52] ^ W[50];
assign W[66] = `SHA1CircularShift(1,Wt[50]);
assign Wt[51]= W[64] ^ W[59] ^ W[53] ^ W[51];
assign W[67] = `SHA1CircularShift(1,Wt[51]);
assign Wt[52]= W[65] ^ W[60] ^ W[54] ^ W[52];
assign W[68] = `SHA1CircularShift(1,Wt[52]);
assign Wt[53]= W[66] ^ W[61] ^ W[55] ^ W[53];
assign W[69] = `SHA1CircularShift(1,Wt[53]);
assign Wt[54]= W[67] ^ W[62] ^ W[56] ^ W[54];
assign W[70] = `SHA1CircularShift(1,Wt[54]);
assign Wt[55]= W[68] ^ W[63] ^ W[57] ^ W[55];
assign W[71] = `SHA1CircularShift(1,Wt[55]);
assign Wt[56]= W[69] ^ W[64] ^ W[58] ^ W[56];
assign W[72] = `SHA1CircularShift(1,Wt[56]);
assign Wt[57]= W[70] ^ W[65] ^ W[59] ^ W[57];
assign W[73] = `SHA1CircularShift(1,Wt[57]);
assign Wt[58]= W[71] ^ W[66] ^ W[60] ^ W[58];
assign W[74] = `SHA1CircularShift(1,Wt[58]);
assign Wt[59]= W[72] ^ W[67] ^ W[61] ^ W[59];
assign W[75] = `SHA1CircularShift(1,Wt[59]);
assign Wt[60]= W[73] ^ W[68] ^ W[62] ^ W[60];
assign W[76] = `SHA1CircularShift(1,Wt[60]);
assign Wt[61]= W[74] ^ W[69] ^ W[63] ^ W[61];
assign W[77] = `SHA1CircularShift(1,Wt[61]);
assign Wt[62]= W[75] ^ W[70] ^ W[64] ^ W[62];
assign W[78] = `SHA1CircularShift(1,Wt[62]);
assign Wt[63]= W[76] ^ W[71] ^ W[65] ^ W[63];
assign W[79] = `SHA1CircularShift(1,Wt[63]);
/* assign initial hashes*/
assign A[0] = current_hash[31:0];
assign B[0] = current_hash[63:32];
assign C[0] = current_hash[95:64];
assign D[0] = current_hash[127:96];
assign E[0] = current_hash[159:128];

/* * * * * First Rounds [0-19] * * * * */
assign temp[0] = `SHA1CircularShift(5,A[0]) + ((B[0] & C[0]) | ((~B[0]) & D[0])) + E[0] + W[0] + `kzero;
assign E[0+1] = D[0];
assign D[0+1] = C[0];
assign C[0+1] = `SHA1CircularShift(30,B[0]);
assign B[0+1] = A[0];
assign A[0+1] = temp[0][31:0];
assign temp[1] = `SHA1CircularShift(5,A[1]) + ((B[1] & C[1]) | ((~B[1]) & D[1])) + E[1] + W[1] + `kzero;
assign E[1+1] = D[1];
assign D[1+1] = C[1];
assign C[1+1] = `SHA1CircularShift(30,B[1]);
assign B[1+1] = A[1];
assign A[1+1] = temp[1][31:0];
assign temp[2] = `SHA1CircularShift(5,A[2]) + ((B[2] & C[2]) | ((~B[2]) & D[2])) + E[2] + W[2] + `kzero;
assign E[2+1] = D[2];
assign D[2+1] = C[2];
assign C[2+1] = `SHA1CircularShift(30,B[2]);
assign B[2+1] = A[2];
assign A[2+1] = temp[2][31:0];
assign temp[3] = `SHA1CircularShift(5,A[3]) + ((B[3] & C[3]) | ((~B[3]) & D[3])) + E[3] + W[3] + `kzero;
assign E[3+1] = D[3];
assign D[3+1] = C[3];
assign C[3+1] = `SHA1CircularShift(30,B[3]);
assign B[3+1] = A[3];
assign A[3+1] = temp[3][31:0];
assign temp[4] = `SHA1CircularShift(5,A[4]) + ((B[4] & C[4]) | ((~B[4]) & D[4])) + E[4] + W[4] + `kzero;
assign E[4+1] = D[4];
assign D[4+1] = C[4];
assign C[4+1] = `SHA1CircularShift(30,B[4]);
assign B[4+1] = A[4];
assign A[4+1] = temp[4][31:0];
assign temp[5] = `SHA1CircularShift(5,A[5]) + ((B[5] & C[5]) | ((~B[5]) & D[5])) + E[5] + W[5] + `kzero;
assign E[5+1] = D[5];
assign D[5+1] = C[5];
assign C[5+1] = `SHA1CircularShift(30,B[5]);
assign B[5+1] = A[5];
assign A[5+1] = temp[5][31:0];
assign temp[6] = `SHA1CircularShift(5,A[6]) + ((B[6] & C[6]) | ((~B[6]) & D[6])) + E[6] + W[6] + `kzero;
assign E[6+1] = D[6];
assign D[6+1] = C[6];
assign C[6+1] = `SHA1CircularShift(30,B[6]);
assign B[6+1] = A[6];
assign A[6+1] = temp[6][31:0];
assign temp[7] = `SHA1CircularShift(5,A[7]) + ((B[7] & C[7]) | ((~B[7]) & D[7])) + E[7] + W[7] + `kzero;
assign E[7+1] = D[7];
assign D[7+1] = C[7];
assign C[7+1] = `SHA1CircularShift(30,B[7]);
assign B[7+1] = A[7];
assign A[7+1] = temp[7][31:0];
assign temp[8] = `SHA1CircularShift(5,A[8]) + ((B[8] & C[8]) | ((~B[8]) & D[8])) + E[8] + W[8] + `kzero;
assign E[8+1] = D[8];
assign D[8+1] = C[8];
assign C[8+1] = `SHA1CircularShift(30,B[8]);
assign B[8+1] = A[8];
assign A[8+1] = temp[8][31:0];
assign temp[9] = `SHA1CircularShift(5,A[9]) + ((B[9] & C[9]) | ((~B[9]) & D[9])) + E[9] + W[9] + `kzero;
assign E[9+1] = D[9];
assign D[9+1] = C[9];
assign C[9+1] = `SHA1CircularShift(30,B[9]);
assign B[9+1] = A[9];
assign A[9+1] = temp[9][31:0];
assign temp[10] = `SHA1CircularShift(5,A[10]) + ((B[10] & C[10]) | ((~B[10]) & D[10])) + E[10] + W[10] + `kzero;
assign E[10+1] = D[10];
assign D[10+1] = C[10];
assign C[10+1] = `SHA1CircularShift(30,B[10]);
assign B[10+1] = A[10];
assign A[10+1] = temp[10][31:0];
assign temp[11] = `SHA1CircularShift(5,A[11]) + ((B[11] & C[11]) | ((~B[11]) & D[11])) + E[11] + W[11] + `kzero;
assign E[11+1] = D[11];
assign D[11+1] = C[11];
assign C[11+1] = `SHA1CircularShift(30,B[11]);
assign B[11+1] = A[11];
assign A[11+1] = temp[11][31:0];
assign temp[12] = `SHA1CircularShift(5,A[12]) + ((B[12] & C[12]) | ((~B[12]) & D[12])) + E[12] + W[12] + `kzero;
assign E[12+1] = D[12];
assign D[12+1] = C[12];
assign C[12+1] = `SHA1CircularShift(30,B[12]);
assign B[12+1] = A[12];
assign A[12+1] = temp[12][31:0];
assign temp[13] = `SHA1CircularShift(5,A[13]) + ((B[13] & C[13]) | ((~B[13]) & D[13])) + E[13] + W[13] + `kzero;
assign E[13+1] = D[13];
assign D[13+1] = C[13];
assign C[13+1] = `SHA1CircularShift(30,B[13]);
assign B[13+1] = A[13];
assign A[13+1] = temp[13][31:0];
assign temp[14] = `SHA1CircularShift(5,A[14]) + ((B[14] & C[14]) | ((~B[14]) & D[14])) + E[14] + W[14] + `kzero;
assign E[14+1] = D[14];
assign D[14+1] = C[14];
assign C[14+1] = `SHA1CircularShift(30,B[14]);
assign B[14+1] = A[14];
assign A[14+1] = temp[14][31:0];
assign temp[15] = `SHA1CircularShift(5,A[15]) + ((B[15] & C[15]) | ((~B[15]) & D[15])) + E[15] + W[15] + `kzero;
assign E[15+1] = D[15];
assign D[15+1] = C[15];
assign C[15+1] = `SHA1CircularShift(30,B[15]);
assign B[15+1] = A[15];
assign A[15+1] = temp[15][31:0];
assign temp[16] = `SHA1CircularShift(5,A[16]) + ((B[16] & C[16]) | ((~B[16]) & D[16])) + E[16] + W[16] + `kzero;
assign E[16+1] = D[16];
assign D[16+1] = C[16];
assign C[16+1] = `SHA1CircularShift(30,B[16]);
assign B[16+1] = A[16];
assign A[16+1] = temp[16][31:0];
assign temp[17] = `SHA1CircularShift(5,A[17]) + ((B[17] & C[17]) | ((~B[17]) & D[17])) + E[17] + W[17] + `kzero;
assign E[17+1] = D[17];
assign D[17+1] = C[17];
assign C[17+1] = `SHA1CircularShift(30,B[17]);
assign B[17+1] = A[17];
assign A[17+1] = temp[17][31:0];
assign temp[18] = `SHA1CircularShift(5,A[18]) + ((B[18] & C[18]) | ((~B[18]) & D[18])) + E[18] + W[18] + `kzero;
assign E[18+1] = D[18];
assign D[18+1] = C[18];
assign C[18+1] = `SHA1CircularShift(30,B[18]);
assign B[18+1] = A[18];
assign A[18+1] = temp[18][31:0];
assign temp[19] = `SHA1CircularShift(5,A[19]) + ((B[19] & C[19]) | ((~B[19]) & D[19])) + E[19] + W[19] + `kzero;
assign E[19+1] = D[19];
assign D[19+1] = C[19];
assign C[19+1] = `SHA1CircularShift(30,B[19]);
assign B[19+1] = A[19];
assign A[19+1] = temp[19][31:0];

/* * * * * Second Rounds [20-39] * * * * */
assign temp[20] = `SHA1CircularShift(5,A[20]) + (B[20]^C[20]^D[20]) + E[20] + W[20] + `kone;
assign E[20+1] = D[20];
assign D[20+1] = C[20];
assign C[20+1] = `SHA1CircularShift(30,B[20]);
assign B[20+1] = A[20];
assign A[20+1] = temp[20][31:0];
assign temp[21] = `SHA1CircularShift(5,A[21]) + (B[21]^C[21]^D[21]) + E[21] + W[21] + `kone;
assign E[21+1] = D[21];
assign D[21+1] = C[21];
assign C[21+1] = `SHA1CircularShift(30,B[21]);
assign B[21+1] = A[21];
assign A[21+1] = temp[21][31:0];
assign temp[22] = `SHA1CircularShift(5,A[22]) + (B[22]^C[22]^D[22]) + E[22] + W[22] + `kone;
assign E[22+1] = D[22];
assign D[22+1] = C[22];
assign C[22+1] = `SHA1CircularShift(30,B[22]);
assign B[22+1] = A[22];
assign A[22+1] = temp[22][31:0];
assign temp[23] = `SHA1CircularShift(5,A[23]) + (B[23]^C[23]^D[23]) + E[23] + W[23] + `kone;
assign E[23+1] = D[23];
assign D[23+1] = C[23];
assign C[23+1] = `SHA1CircularShift(30,B[23]);
assign B[23+1] = A[23];
assign A[23+1] = temp[23][31:0];
assign temp[24] = `SHA1CircularShift(5,A[24]) + (B[24]^C[24]^D[24]) + E[24] + W[24] + `kone;
assign E[24+1] = D[24];
assign D[24+1] = C[24];
assign C[24+1] = `SHA1CircularShift(30,B[24]);
assign B[24+1] = A[24];
assign A[24+1] = temp[24][31:0];
assign temp[25] = `SHA1CircularShift(5,A[25]) + (B[25]^C[25]^D[25]) + E[25] + W[25] + `kone;
assign E[25+1] = D[25];
assign D[25+1] = C[25];
assign C[25+1] = `SHA1CircularShift(30,B[25]);
assign B[25+1] = A[25];
assign A[25+1] = temp[25][31:0];
assign temp[26] = `SHA1CircularShift(5,A[26]) + (B[26]^C[26]^D[26]) + E[26] + W[26] + `kone;
assign E[26+1] = D[26];
assign D[26+1] = C[26];
assign C[26+1] = `SHA1CircularShift(30,B[26]);
assign B[26+1] = A[26];
assign A[26+1] = temp[26][31:0];
assign temp[27] = `SHA1CircularShift(5,A[27]) + (B[27]^C[27]^D[27]) + E[27] + W[27] + `kone;
assign E[27+1] = D[27];
assign D[27+1] = C[27];
assign C[27+1] = `SHA1CircularShift(30,B[27]);
assign B[27+1] = A[27];
assign A[27+1] = temp[27][31:0];
assign temp[28] = `SHA1CircularShift(5,A[28]) + (B[28]^C[28]^D[28]) + E[28] + W[28] + `kone;
assign E[28+1] = D[28];
assign D[28+1] = C[28];
assign C[28+1] = `SHA1CircularShift(30,B[28]);
assign B[28+1] = A[28];
assign A[28+1] = temp[28][31:0];
assign temp[29] = `SHA1CircularShift(5,A[29]) + (B[29]^C[29]^D[29]) + E[29] + W[29] + `kone;
assign E[29+1] = D[29];
assign D[29+1] = C[29];
assign C[29+1] = `SHA1CircularShift(30,B[29]);
assign B[29+1] = A[29];
assign A[29+1] = temp[29][31:0];
assign temp[30] = `SHA1CircularShift(5,A[30]) + (B[30]^C[30]^D[30]) + E[30] + W[30] + `kone;
assign E[30+1] = D[30];
assign D[30+1] = C[30];
assign C[30+1] = `SHA1CircularShift(30,B[30]);
assign B[30+1] = A[30];
assign A[30+1] = temp[30][31:0];
assign temp[31] = `SHA1CircularShift(5,A[31]) + (B[31]^C[31]^D[31]) + E[31] + W[31] + `kone;
assign E[31+1] = D[31];
assign D[31+1] = C[31];
assign C[31+1] = `SHA1CircularShift(30,B[31]);
assign B[31+1] = A[31];
assign A[31+1] = temp[31][31:0];
assign temp[32] = `SHA1CircularShift(5,A[32]) + (B[32]^C[32]^D[32]) + E[32] + W[32] + `kone;
assign E[32+1] = D[32];
assign D[32+1] = C[32];
assign C[32+1] = `SHA1CircularShift(30,B[32]);
assign B[32+1] = A[32];
assign A[32+1] = temp[32][31:0];
assign temp[33] = `SHA1CircularShift(5,A[33]) + (B[33]^C[33]^D[33]) + E[33] + W[33] + `kone;
assign E[33+1] = D[33];
assign D[33+1] = C[33];
assign C[33+1] = `SHA1CircularShift(30,B[33]);
assign B[33+1] = A[33];
assign A[33+1] = temp[33][31:0];
assign temp[34] = `SHA1CircularShift(5,A[34]) + (B[34]^C[34]^D[34]) + E[34] + W[34] + `kone;
assign E[34+1] = D[34];
assign D[34+1] = C[34];
assign C[34+1] = `SHA1CircularShift(30,B[34]);
assign B[34+1] = A[34];
assign A[34+1] = temp[34][31:0];
assign temp[35] = `SHA1CircularShift(5,A[35]) + (B[35]^C[35]^D[35]) + E[35] + W[35] + `kone;
assign E[35+1] = D[35];
assign D[35+1] = C[35];
assign C[35+1] = `SHA1CircularShift(30,B[35]);
assign B[35+1] = A[35];
assign A[35+1] = temp[35][31:0];
assign temp[36] = `SHA1CircularShift(5,A[36]) + (B[36]^C[36]^D[36]) + E[36] + W[36] + `kone;
assign E[36+1] = D[36];
assign D[36+1] = C[36];
assign C[36+1] = `SHA1CircularShift(30,B[36]);
assign B[36+1] = A[36];
assign A[36+1] = temp[36][31:0];
assign temp[37] = `SHA1CircularShift(5,A[37]) + (B[37]^C[37]^D[37]) + E[37] + W[37] + `kone;
assign E[37+1] = D[37];
assign D[37+1] = C[37];
assign C[37+1] = `SHA1CircularShift(30,B[37]);
assign B[37+1] = A[37];
assign A[37+1] = temp[37][31:0];
assign temp[38] = `SHA1CircularShift(5,A[38]) + (B[38]^C[38]^D[38]) + E[38] + W[38] + `kone;
assign E[38+1] = D[38];
assign D[38+1] = C[38];
assign C[38+1] = `SHA1CircularShift(30,B[38]);
assign B[38+1] = A[38];
assign A[38+1] = temp[38][31:0];
assign temp[39] = `SHA1CircularShift(5,A[39]) + (B[39]^C[39]^D[39]) + E[39] + W[39] + `kone;
assign E[39+1] = D[39];
assign D[39+1] = C[39];
assign C[39+1] = `SHA1CircularShift(30,B[39]);
assign B[39+1] = A[39];
assign A[39+1] = temp[39][31:0];

/* * * * * Third Rounds [40-59] * * * * */
assign temp[40] = `SHA1CircularShift(5,A[40]) + ((B[40] & C[40]) | (B[40] & D[40]) | (C[40] & D[40])) + E[40] + W[40] + `ktwo;
assign E[40+1] = D[40];
assign D[40+1] = C[40];
assign C[40+1] = `SHA1CircularShift(30,B[40]);
assign B[40+1] = A[40];
assign A[40+1] = temp[40][31:0];
assign temp[41] = `SHA1CircularShift(5,A[41]) + ((B[41] & C[41]) | (B[41] & D[41]) | (C[41] & D[41])) + E[41] + W[41] + `ktwo;
assign E[41+1] = D[41];
assign D[41+1] = C[41];
assign C[41+1] = `SHA1CircularShift(30,B[41]);
assign B[41+1] = A[41];
assign A[41+1] = temp[41][31:0];
assign temp[42] = `SHA1CircularShift(5,A[42]) + ((B[42] & C[42]) | (B[42] & D[42]) | (C[42] & D[42])) + E[42] + W[42] + `ktwo;
assign E[42+1] = D[42];
assign D[42+1] = C[42];
assign C[42+1] = `SHA1CircularShift(30,B[42]);
assign B[42+1] = A[42];
assign A[42+1] = temp[42][31:0];
assign temp[43] = `SHA1CircularShift(5,A[43]) + ((B[43] & C[43]) | (B[43] & D[43]) | (C[43] & D[43])) + E[43] + W[43] + `ktwo;
assign E[43+1] = D[43];
assign D[43+1] = C[43];
assign C[43+1] = `SHA1CircularShift(30,B[43]);
assign B[43+1] = A[43];
assign A[43+1] = temp[43][31:0];
assign temp[44] = `SHA1CircularShift(5,A[44]) + ((B[44] & C[44]) | (B[44] & D[44]) | (C[44] & D[44])) + E[44] + W[44] + `ktwo;
assign E[44+1] = D[44];
assign D[44+1] = C[44];
assign C[44+1] = `SHA1CircularShift(30,B[44]);
assign B[44+1] = A[44];
assign A[44+1] = temp[44][31:0];
assign temp[45] = `SHA1CircularShift(5,A[45]) + ((B[45] & C[45]) | (B[45] & D[45]) | (C[45] & D[45])) + E[45] + W[45] + `ktwo;
assign E[45+1] = D[45];
assign D[45+1] = C[45];
assign C[45+1] = `SHA1CircularShift(30,B[45]);
assign B[45+1] = A[45];
assign A[45+1] = temp[45][31:0];
assign temp[46] = `SHA1CircularShift(5,A[46]) + ((B[46] & C[46]) | (B[46] & D[46]) | (C[46] & D[46])) + E[46] + W[46] + `ktwo;
assign E[46+1] = D[46];
assign D[46+1] = C[46];
assign C[46+1] = `SHA1CircularShift(30,B[46]);
assign B[46+1] = A[46];
assign A[46+1] = temp[46][31:0];
assign temp[47] = `SHA1CircularShift(5,A[47]) + ((B[47] & C[47]) | (B[47] & D[47]) | (C[47] & D[47])) + E[47] + W[47] + `ktwo;
assign E[47+1] = D[47];
assign D[47+1] = C[47];
assign C[47+1] = `SHA1CircularShift(30,B[47]);
assign B[47+1] = A[47];
assign A[47+1] = temp[47][31:0];
assign temp[48] = `SHA1CircularShift(5,A[48]) + ((B[48] & C[48]) | (B[48] & D[48]) | (C[48] & D[48])) + E[48] + W[48] + `ktwo;
assign E[48+1] = D[48];
assign D[48+1] = C[48];
assign C[48+1] = `SHA1CircularShift(30,B[48]);
assign B[48+1] = A[48];
assign A[48+1] = temp[48][31:0];
assign temp[49] = `SHA1CircularShift(5,A[49]) + ((B[49] & C[49]) | (B[49] & D[49]) | (C[49] & D[49])) + E[49] + W[49] + `ktwo;
assign E[49+1] = D[49];
assign D[49+1] = C[49];
assign C[49+1] = `SHA1CircularShift(30,B[49]);
assign B[49+1] = A[49];
assign A[49+1] = temp[49][31:0];
assign temp[50] = `SHA1CircularShift(5,A[50]) + ((B[50] & C[50]) | (B[50] & D[50]) | (C[50] & D[50])) + E[50] + W[50] + `ktwo;
assign E[50+1] = D[50];
assign D[50+1] = C[50];
assign C[50+1] = `SHA1CircularShift(30,B[50]);
assign B[50+1] = A[50];
assign A[50+1] = temp[50][31:0];
assign temp[51] = `SHA1CircularShift(5,A[51]) + ((B[51] & C[51]) | (B[51] & D[51]) | (C[51] & D[51])) + E[51] + W[51] + `ktwo;
assign E[51+1] = D[51];
assign D[51+1] = C[51];
assign C[51+1] = `SHA1CircularShift(30,B[51]);
assign B[51+1] = A[51];
assign A[51+1] = temp[51][31:0];
assign temp[52] = `SHA1CircularShift(5,A[52]) + ((B[52] & C[52]) | (B[52] & D[52]) | (C[52] & D[52])) + E[52] + W[52] + `ktwo;
assign E[52+1] = D[52];
assign D[52+1] = C[52];
assign C[52+1] = `SHA1CircularShift(30,B[52]);
assign B[52+1] = A[52];
assign A[52+1] = temp[52][31:0];
assign temp[53] = `SHA1CircularShift(5,A[53]) + ((B[53] & C[53]) | (B[53] & D[53]) | (C[53] & D[53])) + E[53] + W[53] + `ktwo;
assign E[53+1] = D[53];
assign D[53+1] = C[53];
assign C[53+1] = `SHA1CircularShift(30,B[53]);
assign B[53+1] = A[53];
assign A[53+1] = temp[53][31:0];
assign temp[54] = `SHA1CircularShift(5,A[54]) + ((B[54] & C[54]) | (B[54] & D[54]) | (C[54] & D[54])) + E[54] + W[54] + `ktwo;
assign E[54+1] = D[54];
assign D[54+1] = C[54];
assign C[54+1] = `SHA1CircularShift(30,B[54]);
assign B[54+1] = A[54];
assign A[54+1] = temp[54][31:0];
assign temp[55] = `SHA1CircularShift(5,A[55]) + ((B[55] & C[55]) | (B[55] & D[55]) | (C[55] & D[55])) + E[55] + W[55] + `ktwo;
assign E[55+1] = D[55];
assign D[55+1] = C[55];
assign C[55+1] = `SHA1CircularShift(30,B[55]);
assign B[55+1] = A[55];
assign A[55+1] = temp[55][31:0];
assign temp[56] = `SHA1CircularShift(5,A[56]) + ((B[56] & C[56]) | (B[56] & D[56]) | (C[56] & D[56])) + E[56] + W[56] + `ktwo;
assign E[56+1] = D[56];
assign D[56+1] = C[56];
assign C[56+1] = `SHA1CircularShift(30,B[56]);
assign B[56+1] = A[56];
assign A[56+1] = temp[56][31:0];
assign temp[57] = `SHA1CircularShift(5,A[57]) + ((B[57] & C[57]) | (B[57] & D[57]) | (C[57] & D[57])) + E[57] + W[57] + `ktwo;
assign E[57+1] = D[57];
assign D[57+1] = C[57];
assign C[57+1] = `SHA1CircularShift(30,B[57]);
assign B[57+1] = A[57];
assign A[57+1] = temp[57][31:0];
assign temp[58] = `SHA1CircularShift(5,A[58]) + ((B[58] & C[58]) | (B[58] & D[58]) | (C[58] & D[58])) + E[58] + W[58] + `ktwo;
assign E[58+1] = D[58];
assign D[58+1] = C[58];
assign C[58+1] = `SHA1CircularShift(30,B[58]);
assign B[58+1] = A[58];
assign A[58+1] = temp[58][31:0];
assign temp[59] = `SHA1CircularShift(5,A[59]) + ((B[59] & C[59]) | (B[59] & D[59]) | (C[59] & D[59])) + E[59] + W[59] + `ktwo;
assign E[59+1] = D[59];
assign D[59+1] = C[59];
assign C[59+1] = `SHA1CircularShift(30,B[59]);
assign B[59+1] = A[59];
assign A[59+1] = temp[59][31:0];

/* * * * * Fourth Rounds [60-79] * * * * */
assign temp[60] = `SHA1CircularShift(5,A[60]) + (B[60]^C[60]^D[60]) + E[60] + W[60] + `kthree;
assign E[60+1] = D[60];
assign D[60+1] = C[60];
assign C[60+1] = `SHA1CircularShift(30,B[60]);
assign B[60+1] = A[60];
assign A[60+1] = temp[60][31:0];
assign temp[61] = `SHA1CircularShift(5,A[61]) + (B[61]^C[61]^D[61]) + E[61] + W[61] + `kthree;
assign E[61+1] = D[61];
assign D[61+1] = C[61];
assign C[61+1] = `SHA1CircularShift(30,B[61]);
assign B[61+1] = A[61];
assign A[61+1] = temp[61][31:0];
assign temp[62] = `SHA1CircularShift(5,A[62]) + (B[62]^C[62]^D[62]) + E[62] + W[62] + `kthree;
assign E[62+1] = D[62];
assign D[62+1] = C[62];
assign C[62+1] = `SHA1CircularShift(30,B[62]);
assign B[62+1] = A[62];
assign A[62+1] = temp[62][31:0];
assign temp[63] = `SHA1CircularShift(5,A[63]) + (B[63]^C[63]^D[63]) + E[63] + W[63] + `kthree;
assign E[63+1] = D[63];
assign D[63+1] = C[63];
assign C[63+1] = `SHA1CircularShift(30,B[63]);
assign B[63+1] = A[63];
assign A[63+1] = temp[63][31:0];
assign temp[64] = `SHA1CircularShift(5,A[64]) + (B[64]^C[64]^D[64]) + E[64] + W[64] + `kthree;
assign E[64+1] = D[64];
assign D[64+1] = C[64];
assign C[64+1] = `SHA1CircularShift(30,B[64]);
assign B[64+1] = A[64];
assign A[64+1] = temp[64][31:0];
assign temp[65] = `SHA1CircularShift(5,A[65]) + (B[65]^C[65]^D[65]) + E[65] + W[65] + `kthree;
assign E[65+1] = D[65];
assign D[65+1] = C[65];
assign C[65+1] = `SHA1CircularShift(30,B[65]);
assign B[65+1] = A[65];
assign A[65+1] = temp[65][31:0];
assign temp[66] = `SHA1CircularShift(5,A[66]) + (B[66]^C[66]^D[66]) + E[66] + W[66] + `kthree;
assign E[66+1] = D[66];
assign D[66+1] = C[66];
assign C[66+1] = `SHA1CircularShift(30,B[66]);
assign B[66+1] = A[66];
assign A[66+1] = temp[66][31:0];
assign temp[67] = `SHA1CircularShift(5,A[67]) + (B[67]^C[67]^D[67]) + E[67] + W[67] + `kthree;
assign E[67+1] = D[67];
assign D[67+1] = C[67];
assign C[67+1] = `SHA1CircularShift(30,B[67]);
assign B[67+1] = A[67];
assign A[67+1] = temp[67][31:0];
assign temp[68] = `SHA1CircularShift(5,A[68]) + (B[68]^C[68]^D[68]) + E[68] + W[68] + `kthree;
assign E[68+1] = D[68];
assign D[68+1] = C[68];
assign C[68+1] = `SHA1CircularShift(30,B[68]);
assign B[68+1] = A[68];
assign A[68+1] = temp[68][31:0];
assign temp[69] = `SHA1CircularShift(5,A[69]) + (B[69]^C[69]^D[69]) + E[69] + W[69] + `kthree;
assign E[69+1] = D[69];
assign D[69+1] = C[69];
assign C[69+1] = `SHA1CircularShift(30,B[69]);
assign B[69+1] = A[69];
assign A[69+1] = temp[69][31:0];
assign temp[70] = `SHA1CircularShift(5,A[70]) + (B[70]^C[70]^D[70]) + E[70] + W[70] + `kthree;
assign E[70+1] = D[70];
assign D[70+1] = C[70];
assign C[70+1] = `SHA1CircularShift(30,B[70]);
assign B[70+1] = A[70];
assign A[70+1] = temp[70][31:0];
assign temp[71] = `SHA1CircularShift(5,A[71]) + (B[71]^C[71]^D[71]) + E[71] + W[71] + `kthree;
assign E[71+1] = D[71];
assign D[71+1] = C[71];
assign C[71+1] = `SHA1CircularShift(30,B[71]);
assign B[71+1] = A[71];
assign A[71+1] = temp[71][31:0];
assign temp[72] = `SHA1CircularShift(5,A[72]) + (B[72]^C[72]^D[72]) + E[72] + W[72] + `kthree;
assign E[72+1] = D[72];
assign D[72+1] = C[72];
assign C[72+1] = `SHA1CircularShift(30,B[72]);
assign B[72+1] = A[72];
assign A[72+1] = temp[72][31:0];
assign temp[73] = `SHA1CircularShift(5,A[73]) + (B[73]^C[73]^D[73]) + E[73] + W[73] + `kthree;
assign E[73+1] = D[73];
assign D[73+1] = C[73];
assign C[73+1] = `SHA1CircularShift(30,B[73]);
assign B[73+1] = A[73];
assign A[73+1] = temp[73][31:0];
assign temp[74] = `SHA1CircularShift(5,A[74]) + (B[74]^C[74]^D[74]) + E[74] + W[74] + `kthree;
assign E[74+1] = D[74];
assign D[74+1] = C[74];
assign C[74+1] = `SHA1CircularShift(30,B[74]);
assign B[74+1] = A[74];
assign A[74+1] = temp[74][31:0];
assign temp[75] = `SHA1CircularShift(5,A[75]) + (B[75]^C[75]^D[75]) + E[75] + W[75] + `kthree;
assign E[75+1] = D[75];
assign D[75+1] = C[75];
assign C[75+1] = `SHA1CircularShift(30,B[75]);
assign B[75+1] = A[75];
assign A[75+1] = temp[75][31:0];
assign temp[76] = `SHA1CircularShift(5,A[76]) + (B[76]^C[76]^D[76]) + E[76] + W[76] + `kthree;
assign E[76+1] = D[76];
assign D[76+1] = C[76];
assign C[76+1] = `SHA1CircularShift(30,B[76]);
assign B[76+1] = A[76];
assign A[76+1] = temp[76][31:0];
assign temp[77] = `SHA1CircularShift(5,A[77]) + (B[77]^C[77]^D[77]) + E[77] + W[77] + `kthree;
assign E[77+1] = D[77];
assign D[77+1] = C[77];
assign C[77+1] = `SHA1CircularShift(30,B[77]);
assign B[77+1] = A[77];
assign A[77+1] = temp[77][31:0];
assign temp[78] = `SHA1CircularShift(5,A[78]) + (B[78]^C[78]^D[78]) + E[78] + W[78] + `kthree;
assign E[78+1] = D[78];
assign D[78+1] = C[78];
assign C[78+1] = `SHA1CircularShift(30,B[78]);
assign B[78+1] = A[78];
assign A[78+1] = temp[78][31:0];
assign temp[79] = `SHA1CircularShift(5,A[79]) + (B[79]^C[79]^D[79]) + E[79] + W[79] + `kthree;
assign E[79+1] = D[79];
assign D[79+1] = C[79];
assign C[79+1] = `SHA1CircularShift(30,B[79]);
assign B[79+1] = A[79];
assign A[79+1] = temp[79][31:0];
assign new_hash[31:0] = current_hash[31:0] + A[80];
assign new_hash[63:32] = current_hash[63:32] + B[80];
assign new_hash[95:64] = current_hash[95:64] + C[80];
assign new_hash[127:96] = current_hash[127:96] + D[80];
assign new_hash[159:128] = current_hash[159:128] + E[80];
/* finally, add the new values to the current hash for a new hash
always @(A[80],B[80],C[80],D[80],E[80],current_hash) begin

	new_hash[31:0] <= current_hash[31:0] + A[80];
	new_hash[63:32] <= current_hash[63:32] + B[80];
	new_hash[95:64] <= current_hash[95:64] + C[80];
	new_hash[127:96] <= current_hash[127:96] + D[80];
	new_hash[159:128] <= current_hash[159:128] + E[80];
end*/
endmodule
