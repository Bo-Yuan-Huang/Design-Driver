
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1071 ;
  wire [3:0] \oc8051_golden_model_1.n1073 ;
  wire [3:0] \oc8051_golden_model_1.n1075 ;
  wire [3:0] \oc8051_golden_model_1.n1076 ;
  wire [3:0] \oc8051_golden_model_1.n1077 ;
  wire [3:0] \oc8051_golden_model_1.n1078 ;
  wire [3:0] \oc8051_golden_model_1.n1079 ;
  wire [3:0] \oc8051_golden_model_1.n1080 ;
  wire [3:0] \oc8051_golden_model_1.n1081 ;
  wire \oc8051_golden_model_1.n1118 ;
  wire \oc8051_golden_model_1.n1146 ;
  wire [8:0] \oc8051_golden_model_1.n1147 ;
  wire [8:0] \oc8051_golden_model_1.n1148 ;
  wire [7:0] \oc8051_golden_model_1.n1149 ;
  wire \oc8051_golden_model_1.n1150 ;
  wire \oc8051_golden_model_1.n1151 ;
  wire [2:0] \oc8051_golden_model_1.n1152 ;
  wire \oc8051_golden_model_1.n1153 ;
  wire [1:0] \oc8051_golden_model_1.n1154 ;
  wire [7:0] \oc8051_golden_model_1.n1155 ;
  wire [15:0] \oc8051_golden_model_1.n1181 ;
  wire [7:0] \oc8051_golden_model_1.n1183 ;
  wire [8:0] \oc8051_golden_model_1.n1185 ;
  wire [8:0] \oc8051_golden_model_1.n1189 ;
  wire \oc8051_golden_model_1.n1190 ;
  wire [3:0] \oc8051_golden_model_1.n1191 ;
  wire [4:0] \oc8051_golden_model_1.n1192 ;
  wire [4:0] \oc8051_golden_model_1.n1196 ;
  wire \oc8051_golden_model_1.n1197 ;
  wire [8:0] \oc8051_golden_model_1.n1198 ;
  wire \oc8051_golden_model_1.n1206 ;
  wire [7:0] \oc8051_golden_model_1.n1207 ;
  wire [8:0] \oc8051_golden_model_1.n1211 ;
  wire \oc8051_golden_model_1.n1212 ;
  wire [4:0] \oc8051_golden_model_1.n1217 ;
  wire \oc8051_golden_model_1.n1218 ;
  wire \oc8051_golden_model_1.n1226 ;
  wire [7:0] \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1229 ;
  wire [8:0] \oc8051_golden_model_1.n1231 ;
  wire \oc8051_golden_model_1.n1232 ;
  wire [3:0] \oc8051_golden_model_1.n1233 ;
  wire [4:0] \oc8051_golden_model_1.n1234 ;
  wire [4:0] \oc8051_golden_model_1.n1236 ;
  wire \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1238 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [7:0] \oc8051_golden_model_1.n1246 ;
  wire [8:0] \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1257 ;
  wire [7:0] \oc8051_golden_model_1.n1258 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [4:0] \oc8051_golden_model_1.n1278 ;
  wire \oc8051_golden_model_1.n1279 ;
  wire [7:0] \oc8051_golden_model_1.n1280 ;
  wire [8:0] \oc8051_golden_model_1.n1282 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire \oc8051_golden_model_1.n1290 ;
  wire [7:0] \oc8051_golden_model_1.n1291 ;
  wire [7:0] \oc8051_golden_model_1.n1292 ;
  wire [8:0] \oc8051_golden_model_1.n1295 ;
  wire [8:0] \oc8051_golden_model_1.n1296 ;
  wire [7:0] \oc8051_golden_model_1.n1297 ;
  wire \oc8051_golden_model_1.n1298 ;
  wire [7:0] \oc8051_golden_model_1.n1299 ;
  wire [7:0] \oc8051_golden_model_1.n1300 ;
  wire [8:0] \oc8051_golden_model_1.n1303 ;
  wire [8:0] \oc8051_golden_model_1.n1305 ;
  wire \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1307 ;
  wire [4:0] \oc8051_golden_model_1.n1309 ;
  wire \oc8051_golden_model_1.n1310 ;
  wire \oc8051_golden_model_1.n1317 ;
  wire [7:0] \oc8051_golden_model_1.n1318 ;
  wire [8:0] \oc8051_golden_model_1.n1322 ;
  wire \oc8051_golden_model_1.n1323 ;
  wire [4:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire [7:0] \oc8051_golden_model_1.n1334 ;
  wire [8:0] \oc8051_golden_model_1.n1338 ;
  wire \oc8051_golden_model_1.n1339 ;
  wire [4:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire [7:0] \oc8051_golden_model_1.n1350 ;
  wire [8:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [4:0] \oc8051_golden_model_1.n1357 ;
  wire \oc8051_golden_model_1.n1358 ;
  wire \oc8051_golden_model_1.n1365 ;
  wire [7:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1520 ;
  wire [6:0] \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [3:0] \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire [7:0] \oc8051_golden_model_1.n1555 ;
  wire [7:0] \oc8051_golden_model_1.n1680 ;
  wire \oc8051_golden_model_1.n1683 ;
  wire \oc8051_golden_model_1.n1685 ;
  wire \oc8051_golden_model_1.n1691 ;
  wire [7:0] \oc8051_golden_model_1.n1692 ;
  wire \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1698 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire \oc8051_golden_model_1.n1709 ;
  wire \oc8051_golden_model_1.n1711 ;
  wire \oc8051_golden_model_1.n1717 ;
  wire [7:0] \oc8051_golden_model_1.n1718 ;
  wire \oc8051_golden_model_1.n1722 ;
  wire \oc8051_golden_model_1.n1724 ;
  wire \oc8051_golden_model_1.n1730 ;
  wire [7:0] \oc8051_golden_model_1.n1731 ;
  wire \oc8051_golden_model_1.n1733 ;
  wire [7:0] \oc8051_golden_model_1.n1734 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire [15:0] \oc8051_golden_model_1.n1739 ;
  wire \oc8051_golden_model_1.n1745 ;
  wire [7:0] \oc8051_golden_model_1.n1746 ;
  wire \oc8051_golden_model_1.n1749 ;
  wire [7:0] \oc8051_golden_model_1.n1750 ;
  wire \oc8051_golden_model_1.n1765 ;
  wire [7:0] \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1771 ;
  wire [7:0] \oc8051_golden_model_1.n1772 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire [7:0] \oc8051_golden_model_1.n1778 ;
  wire \oc8051_golden_model_1.n1783 ;
  wire [7:0] \oc8051_golden_model_1.n1784 ;
  wire \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [7:0] \oc8051_golden_model_1.n1791 ;
  wire [3:0] \oc8051_golden_model_1.n1792 ;
  wire [7:0] \oc8051_golden_model_1.n1793 ;
  wire [7:0] \oc8051_golden_model_1.n1828 ;
  wire \oc8051_golden_model_1.n1847 ;
  wire [7:0] \oc8051_golden_model_1.n1848 ;
  wire [7:0] \oc8051_golden_model_1.n1852 ;
  wire [3:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1854 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not _43534_ (_42618_, rst);
  not _43535_ (_18751_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _43536_ (_18772_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _43537_ (_18773_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18772_);
  and _43538_ (_18784_, _18773_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _43539_ (_18795_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18772_);
  and _43540_ (_18806_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18772_);
  nor _43541_ (_18817_, _18806_, _18795_);
  and _43542_ (_18828_, _18817_, _18784_);
  nor _43543_ (_18839_, _18828_, _18751_);
  and _43544_ (_18850_, _18751_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _43545_ (_18861_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _43546_ (_18872_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18861_);
  nor _43547_ (_18883_, _18872_, _18850_);
  not _43548_ (_18894_, _18883_);
  and _43549_ (_18905_, _18894_, _18828_);
  or _43550_ (_18916_, _18905_, _18839_);
  and _43551_ (_22124_, _18916_, _42618_);
  nor _43552_ (_18937_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _43553_ (_18948_, _18937_);
  and _43554_ (_18959_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and _43555_ (_18970_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _43556_ (_18981_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _43557_ (_18992_, _18981_);
  not _43558_ (_19003_, _18872_);
  nor _43559_ (_19014_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not _43560_ (_19025_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _43561_ (_19036_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _19025_);
  nor _43562_ (_19047_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not _43563_ (_19058_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor _43564_ (_19069_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _19058_);
  nor _43565_ (_19080_, _19069_, _19047_);
  nor _43566_ (_19091_, _19080_, _19036_);
  not _43567_ (_19102_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _43568_ (_19112_, _19036_, _19102_);
  nor _43569_ (_19123_, _19112_, _19091_);
  and _43570_ (_19134_, _19123_, _19014_);
  not _43571_ (_19145_, _19134_);
  and _43572_ (_19156_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _43573_ (_19167_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _43574_ (_19178_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _43575_ (_19189_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _19178_);
  and _43576_ (_19200_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _43577_ (_19211_, _19200_, _19167_);
  and _43578_ (_19222_, _19211_, _19145_);
  nor _43579_ (_19233_, _19222_, _19003_);
  not _43580_ (_19244_, _18850_);
  nor _43581_ (_19255_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor _43582_ (_19266_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _19058_);
  nor _43583_ (_19277_, _19266_, _19255_);
  nor _43584_ (_19288_, _19277_, _19036_);
  not _43585_ (_19299_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _43586_ (_19310_, _19036_, _19299_);
  nor _43587_ (_19321_, _19310_, _19288_);
  and _43588_ (_19332_, _19321_, _19014_);
  not _43589_ (_19343_, _19332_);
  and _43590_ (_19354_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _43591_ (_19365_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _43592_ (_19376_, _19365_, _19354_);
  and _43593_ (_19387_, _19376_, _19343_);
  nor _43594_ (_19398_, _19387_, _19244_);
  nor _43595_ (_19409_, _19398_, _19233_);
  nor _43596_ (_19420_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor _43597_ (_19430_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _19058_);
  nor _43598_ (_19441_, _19430_, _19420_);
  nor _43599_ (_19452_, _19441_, _19036_);
  not _43600_ (_19463_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _43601_ (_19474_, _19036_, _19463_);
  nor _43602_ (_19485_, _19474_, _19452_);
  and _43603_ (_19496_, _19485_, _19014_);
  not _43604_ (_19507_, _19496_);
  and _43605_ (_19517_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _43606_ (_19528_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _43607_ (_19539_, _19528_, _19517_);
  and _43608_ (_19550_, _19539_, _19507_);
  nor _43609_ (_19561_, _19550_, _18894_);
  nor _43610_ (_19572_, _19561_, _18937_);
  and _43611_ (_19583_, _19572_, _19409_);
  nor _43612_ (_19594_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor _43613_ (_19604_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _19058_);
  nor _43614_ (_19615_, _19604_, _19594_);
  nor _43615_ (_19626_, _19615_, _19036_);
  not _43616_ (_19637_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _43617_ (_19648_, _19036_, _19637_);
  nor _43618_ (_19659_, _19648_, _19626_);
  and _43619_ (_19670_, _19659_, _19014_);
  not _43620_ (_19681_, _19670_);
  and _43621_ (_19691_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _43622_ (_19702_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _43623_ (_19713_, _19702_, _19691_);
  and _43624_ (_19724_, _19713_, _19681_);
  and _43625_ (_19735_, _19724_, _18937_);
  nor _43626_ (_19746_, _19735_, _19583_);
  not _43627_ (_19768_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _43628_ (_19779_, _19768_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _43629_ (_19791_, _19779_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43630_ (_19803_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _43631_ (_19815_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _43632_ (_19827_, _19815_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43633_ (_19839_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _43634_ (_19840_, _19839_, _19803_);
  not _43635_ (_19851_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43636_ (_19862_, _19779_, _19851_);
  and _43637_ (_19872_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _43638_ (_19883_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43639_ (_19894_, _19883_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _43640_ (_19905_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor _43641_ (_19916_, _19905_, _19872_);
  and _43642_ (_19927_, _19916_, _19840_);
  and _43643_ (_19938_, _19883_, _19768_);
  and _43644_ (_19948_, _19938_, _19659_);
  and _43645_ (_19959_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _43646_ (_19970_, _19959_, _19851_);
  and _43647_ (_19981_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _43648_ (_19992_, _19959_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43649_ (_20003_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor _43650_ (_20014_, _20003_, _19981_);
  not _43651_ (_20025_, _20014_);
  nor _43652_ (_20035_, _20025_, _19948_);
  and _43653_ (_20046_, _20035_, _19927_);
  not _43654_ (_20057_, _20046_);
  and _43655_ (_20068_, _20057_, _19746_);
  not _43656_ (_20079_, _20068_);
  nor _43657_ (_20090_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor _43658_ (_20101_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _19058_);
  nor _43659_ (_20112_, _20101_, _20090_);
  nor _43660_ (_20122_, _20112_, _19036_);
  not _43661_ (_20133_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _43662_ (_20144_, _19036_, _20133_);
  nor _43663_ (_20155_, _20144_, _20122_);
  and _43664_ (_20166_, _20155_, _19014_);
  not _43665_ (_20177_, _20166_);
  and _43666_ (_20188_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _43667_ (_20199_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _43668_ (_20209_, _20199_, _20188_);
  and _43669_ (_20220_, _20209_, _20177_);
  nor _43670_ (_20231_, _20220_, _19003_);
  nor _43671_ (_20242_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor _43672_ (_20253_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _19058_);
  nor _43673_ (_20264_, _20253_, _20242_);
  nor _43674_ (_20275_, _20264_, _19036_);
  not _43675_ (_20285_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _43676_ (_20296_, _19036_, _20285_);
  nor _43677_ (_20307_, _20296_, _20275_);
  and _43678_ (_20318_, _20307_, _19014_);
  not _43679_ (_20329_, _20318_);
  and _43680_ (_20340_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _43681_ (_20351_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _43682_ (_20362_, _20351_, _20340_);
  and _43683_ (_20372_, _20362_, _20329_);
  nor _43684_ (_20383_, _20372_, _19244_);
  nor _43685_ (_20394_, _20383_, _20231_);
  nor _43686_ (_20405_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor _43687_ (_20416_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _19058_);
  nor _43688_ (_20427_, _20416_, _20405_);
  nor _43689_ (_20438_, _20427_, _19036_);
  not _43690_ (_20449_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _43691_ (_20459_, _19036_, _20449_);
  nor _43692_ (_20470_, _20459_, _20438_);
  and _43693_ (_20481_, _20470_, _19014_);
  not _43694_ (_20492_, _20481_);
  and _43695_ (_20503_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _43696_ (_20514_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _43697_ (_20525_, _20514_, _20503_);
  and _43698_ (_20536_, _20525_, _20492_);
  nor _43699_ (_20546_, _20536_, _18894_);
  nor _43700_ (_20557_, _20546_, _18937_);
  and _43701_ (_20568_, _20557_, _20394_);
  nor _43702_ (_20579_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor _43703_ (_20590_, _19058_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor _43704_ (_20601_, _20590_, _20579_);
  nor _43705_ (_20612_, _20601_, _19036_);
  not _43706_ (_20623_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _43707_ (_20633_, _19036_, _20623_);
  nor _43708_ (_20644_, _20633_, _20612_);
  and _43709_ (_20655_, _20644_, _19014_);
  not _43710_ (_20676_, _20655_);
  and _43711_ (_20687_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _43712_ (_20688_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _43713_ (_20699_, _20688_, _20687_);
  and _43714_ (_20719_, _20699_, _20676_);
  and _43715_ (_20730_, _20719_, _18937_);
  nor _43716_ (_20731_, _20730_, _20568_);
  and _43717_ (_20752_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _43718_ (_20763_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _43719_ (_20764_, _20763_, _20752_);
  and _43720_ (_20775_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _43721_ (_20786_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _43722_ (_20797_, _20786_, _20775_);
  and _43723_ (_20817_, _20797_, _20764_);
  and _43724_ (_20818_, _20644_, _19938_);
  and _43725_ (_20829_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _43726_ (_20840_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _43727_ (_20851_, _20840_, _20829_);
  not _43728_ (_20862_, _20851_);
  nor _43729_ (_20873_, _20862_, _20818_);
  and _43730_ (_20884_, _20873_, _20817_);
  not _43731_ (_20895_, _20884_);
  and _43732_ (_20905_, _20895_, _20731_);
  and _43733_ (_20916_, _20905_, _20079_);
  not _43734_ (_20927_, _20916_);
  and _43735_ (_20948_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _43736_ (_20949_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _43737_ (_20960_, _20949_, _20948_);
  and _43738_ (_20971_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _43739_ (_20982_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _43740_ (_20993_, _20982_, _20971_);
  and _43741_ (_21003_, _20993_, _20960_);
  and _43742_ (_21014_, _20307_, _19938_);
  and _43743_ (_21025_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _43744_ (_21036_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _43745_ (_21047_, _21036_, _21025_);
  not _43746_ (_21058_, _21047_);
  nor _43747_ (_21069_, _21058_, _21014_);
  and _43748_ (_21080_, _21069_, _21003_);
  not _43749_ (_21090_, _21080_);
  and _43750_ (_21101_, _21090_, _20731_);
  and _43751_ (_21122_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _43752_ (_21123_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _43753_ (_21134_, _21123_, _21122_);
  and _43754_ (_21145_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _43755_ (_21156_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _43756_ (_21167_, _21156_, _21145_);
  and _43757_ (_21178_, _21167_, _21134_);
  and _43758_ (_21188_, _19938_, _19321_);
  and _43759_ (_21199_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _43760_ (_21210_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _43761_ (_21221_, _21210_, _21199_);
  not _43762_ (_21232_, _21221_);
  nor _43763_ (_21243_, _21232_, _21188_);
  and _43764_ (_21254_, _21243_, _21178_);
  not _43765_ (_21265_, _21254_);
  and _43766_ (_21276_, _21265_, _19746_);
  and _43767_ (_21286_, _21101_, _21276_);
  nor _43768_ (_21297_, _21286_, _20068_);
  and _43769_ (_21318_, _21286_, _20057_);
  nor _43770_ (_21319_, _21318_, _21297_);
  and _43771_ (_21330_, _21319_, _21101_);
  and _43772_ (_21341_, _20905_, _20068_);
  and _43773_ (_21352_, _20731_, _20057_);
  and _43774_ (_21363_, _20895_, _19746_);
  nor _43775_ (_21373_, _21363_, _21352_);
  nor _43776_ (_21384_, _21373_, _21341_);
  and _43777_ (_21395_, _21384_, _21330_);
  and _43778_ (_21406_, _21384_, _21318_);
  nor _43779_ (_21417_, _21406_, _21395_);
  nor _43780_ (_21428_, _21417_, _20927_);
  and _43781_ (_21439_, _21417_, _20927_);
  nor _43782_ (_21450_, _21439_, _21428_);
  not _43783_ (_21461_, _21450_);
  and _43784_ (_21471_, _21265_, _20731_);
  and _43785_ (_21482_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _43786_ (_21493_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _43787_ (_21504_, _21493_, _21482_);
  and _43788_ (_21515_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _43789_ (_21526_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _43790_ (_21537_, _21526_, _21515_);
  and _43791_ (_21548_, _21537_, _21504_);
  and _43792_ (_21558_, _20155_, _19938_);
  and _43793_ (_21569_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _43794_ (_21580_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor _43795_ (_21591_, _21580_, _21569_);
  not _43796_ (_21602_, _21591_);
  nor _43797_ (_21613_, _21602_, _21558_);
  and _43798_ (_21624_, _21613_, _21548_);
  not _43799_ (_21635_, _21624_);
  and _43800_ (_21646_, _21635_, _19746_);
  and _43801_ (_21666_, _21646_, _21471_);
  and _43802_ (_21667_, _21090_, _19746_);
  nor _43803_ (_21678_, _21667_, _21471_);
  nor _43804_ (_21689_, _21678_, _21286_);
  and _43805_ (_21700_, _21689_, _21666_);
  nor _43806_ (_21711_, _21101_, _20068_);
  nor _43807_ (_21722_, _21711_, _21330_);
  and _43808_ (_21733_, _21722_, _21700_);
  nor _43809_ (_21744_, _21384_, _21330_);
  nor _43810_ (_21754_, _21744_, _21395_);
  nor _43811_ (_21775_, _21754_, _21318_);
  nor _43812_ (_21776_, _21775_, _21406_);
  and _43813_ (_21787_, _21776_, _21733_);
  nor _43814_ (_21798_, _21776_, _21733_);
  nor _43815_ (_21809_, _21798_, _21787_);
  not _43816_ (_21820_, _21809_);
  and _43817_ (_21831_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _43818_ (_21841_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _43819_ (_21852_, _21841_, _21831_);
  and _43820_ (_21863_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and _43821_ (_21874_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor _43822_ (_21885_, _21874_, _21863_);
  and _43823_ (_21896_, _21885_, _21852_);
  and _43824_ (_21907_, _20470_, _19938_);
  and _43825_ (_21918_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _43826_ (_21929_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _43827_ (_21939_, _21929_, _21918_);
  not _43828_ (_21950_, _21939_);
  nor _43829_ (_21961_, _21950_, _21907_);
  and _43830_ (_21972_, _21961_, _21896_);
  not _43831_ (_21983_, _21972_);
  and _43832_ (_21994_, _21983_, _20731_);
  and _43833_ (_22005_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _43834_ (_22015_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _43835_ (_22026_, _22015_, _22005_);
  and _43836_ (_22037_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _43837_ (_22048_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor _43838_ (_22059_, _22048_, _22037_);
  and _43839_ (_22070_, _22059_, _22026_);
  and _43840_ (_22081_, _19938_, _19123_);
  and _43841_ (_22092_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _43842_ (_22102_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor _43843_ (_22113_, _22102_, _22092_);
  not _43844_ (_22125_, _22113_);
  nor _43845_ (_22136_, _22125_, _22081_);
  and _43846_ (_22147_, _22136_, _22070_);
  not _43847_ (_22158_, _22147_);
  and _43848_ (_22169_, _22158_, _19746_);
  and _43849_ (_22180_, _22169_, _21994_);
  and _43850_ (_22190_, _21983_, _19746_);
  not _43851_ (_22201_, _22190_);
  and _43852_ (_22222_, _22158_, _20731_);
  and _43853_ (_22223_, _22222_, _22201_);
  and _43854_ (_22234_, _22223_, _21646_);
  nor _43855_ (_22245_, _22234_, _22180_);
  and _43856_ (_22256_, _21635_, _20731_);
  nor _43857_ (_22267_, _22256_, _21276_);
  nor _43858_ (_22277_, _22267_, _21666_);
  not _43859_ (_22288_, _22277_);
  nor _43860_ (_22299_, _22288_, _22245_);
  nor _43861_ (_22310_, _21689_, _21666_);
  nor _43862_ (_22321_, _22310_, _21700_);
  and _43863_ (_22332_, _22321_, _22299_);
  nor _43864_ (_22343_, _21722_, _21700_);
  nor _43865_ (_22354_, _22343_, _21733_);
  and _43866_ (_22364_, _22354_, _22332_);
  and _43867_ (_22375_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _43868_ (_22386_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _43869_ (_22397_, _22386_, _22375_);
  and _43870_ (_22408_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _43871_ (_22419_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _43872_ (_22430_, _22419_, _22408_);
  and _43873_ (_22440_, _22430_, _22397_);
  and _43874_ (_22451_, _19938_, _19485_);
  and _43875_ (_22462_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and _43876_ (_22473_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _43877_ (_22484_, _22473_, _22462_);
  not _43878_ (_22495_, _22484_);
  nor _43879_ (_22516_, _22495_, _22451_);
  and _43880_ (_22517_, _22516_, _22440_);
  not _43881_ (_22527_, _22517_);
  and _43882_ (_22538_, _22527_, _20731_);
  and _43883_ (_22549_, _22538_, _22190_);
  nor _43884_ (_22560_, _22169_, _21994_);
  nor _43885_ (_22571_, _22560_, _22180_);
  and _43886_ (_22582_, _22571_, _22549_);
  nor _43887_ (_22593_, _22223_, _21646_);
  nor _43888_ (_22603_, _22593_, _22234_);
  and _43889_ (_22624_, _22603_, _22582_);
  and _43890_ (_22625_, _22288_, _22245_);
  nor _43891_ (_22636_, _22625_, _22299_);
  and _43892_ (_22647_, _22636_, _22624_);
  nor _43893_ (_22658_, _22321_, _22299_);
  nor _43894_ (_22669_, _22658_, _22332_);
  and _43895_ (_22680_, _22669_, _22647_);
  nor _43896_ (_22690_, _22354_, _22332_);
  nor _43897_ (_22701_, _22690_, _22364_);
  and _43898_ (_22712_, _22701_, _22680_);
  nor _43899_ (_22723_, _22712_, _22364_);
  nor _43900_ (_22734_, _22723_, _21820_);
  nor _43901_ (_22745_, _22734_, _21787_);
  nor _43902_ (_22756_, _22745_, _21461_);
  or _43903_ (_22767_, _22756_, _21341_);
  nor _43904_ (_22777_, _22767_, _21428_);
  nor _43905_ (_22788_, _22777_, _18992_);
  and _43906_ (_22799_, _22777_, _18992_);
  nor _43907_ (_22810_, _22799_, _22788_);
  not _43908_ (_22821_, _22810_);
  and _43909_ (_22842_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and _43910_ (_22843_, _22745_, _21461_);
  nor _43911_ (_22854_, _22843_, _22756_);
  and _43912_ (_22864_, _22854_, _22842_);
  and _43913_ (_22875_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and _43914_ (_22886_, _22723_, _21820_);
  nor _43915_ (_22897_, _22886_, _22734_);
  and _43916_ (_22908_, _22897_, _22875_);
  nor _43917_ (_22919_, _22897_, _22875_);
  nor _43918_ (_22930_, _22919_, _22908_);
  not _43919_ (_22941_, _22930_);
  and _43920_ (_22951_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor _43921_ (_22962_, _22701_, _22680_);
  nor _43922_ (_22973_, _22962_, _22712_);
  and _43923_ (_22984_, _22973_, _22951_);
  nor _43924_ (_22995_, _22973_, _22951_);
  nor _43925_ (_23006_, _22995_, _22984_);
  and _43926_ (_23017_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor _43927_ (_23028_, _22669_, _22647_);
  nor _43928_ (_23038_, _23028_, _22680_);
  and _43929_ (_23049_, _23038_, _23017_);
  nor _43930_ (_23060_, _23038_, _23017_);
  nor _43931_ (_23071_, _23060_, _23049_);
  not _43932_ (_23082_, _23071_);
  and _43933_ (_23103_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor _43934_ (_23104_, _22636_, _22624_);
  nor _43935_ (_23114_, _23104_, _22647_);
  and _43936_ (_23125_, _23114_, _23103_);
  and _43937_ (_23136_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor _43938_ (_23147_, _22603_, _22582_);
  nor _43939_ (_23158_, _23147_, _22624_);
  and _43940_ (_23169_, _23158_, _23136_);
  and _43941_ (_23180_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor _43942_ (_23191_, _22571_, _22549_);
  nor _43943_ (_23202_, _23191_, _22582_);
  and _43944_ (_23213_, _23202_, _23180_);
  nor _43945_ (_23223_, _23158_, _23136_);
  nor _43946_ (_23234_, _23223_, _23169_);
  and _43947_ (_23245_, _23234_, _23213_);
  nor _43948_ (_23256_, _23245_, _23169_);
  not _43949_ (_23267_, _23256_);
  nor _43950_ (_23278_, _23114_, _23103_);
  nor _43951_ (_23289_, _23278_, _23125_);
  and _43952_ (_23300_, _23289_, _23267_);
  nor _43953_ (_23311_, _23300_, _23125_);
  nor _43954_ (_23322_, _23311_, _23082_);
  nor _43955_ (_23332_, _23322_, _23049_);
  not _43956_ (_23343_, _23332_);
  and _43957_ (_23354_, _23343_, _23006_);
  nor _43958_ (_23365_, _23354_, _22984_);
  nor _43959_ (_23386_, _23365_, _22941_);
  nor _43960_ (_23387_, _23386_, _22908_);
  nor _43961_ (_23398_, _22854_, _22842_);
  nor _43962_ (_23409_, _23398_, _22864_);
  not _43963_ (_23420_, _23409_);
  nor _43964_ (_23431_, _23420_, _23387_);
  nor _43965_ (_23442_, _23431_, _22864_);
  nor _43966_ (_23452_, _23442_, _22821_);
  nor _43967_ (_23463_, _23452_, _22788_);
  not _43968_ (_23474_, _23463_);
  and _43969_ (_23485_, _23474_, _18970_);
  and _43970_ (_23496_, _23485_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _43971_ (_23507_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _43972_ (_23518_, _23507_, _23496_);
  and _43973_ (_23529_, _23518_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _43974_ (_23540_, _23529_, _18959_);
  not _43975_ (_23551_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _43976_ (_23561_, _18937_, _23551_);
  or _43977_ (_23572_, _23561_, _23540_);
  nand _43978_ (_23583_, _23540_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and _43979_ (_23594_, _23583_, _23572_);
  and _43980_ (_24283_, _23594_, _42618_);
  nor _43981_ (_23615_, _18828_, _18861_);
  and _43982_ (_23626_, _18828_, _18861_);
  or _43983_ (_23637_, _23626_, _23615_);
  and _43984_ (_02354_, _23637_, _42618_);
  and _43985_ (_23658_, _22527_, _19746_);
  and _43986_ (_02542_, _23658_, _42618_);
  nor _43987_ (_23678_, _22538_, _22190_);
  nor _43988_ (_23689_, _23678_, _22549_);
  and _43989_ (_02700_, _23689_, _42618_);
  nor _43990_ (_23710_, _23202_, _23180_);
  nor _43991_ (_23721_, _23710_, _23213_);
  and _43992_ (_02882_, _23721_, _42618_);
  nor _43993_ (_23742_, _23234_, _23213_);
  nor _43994_ (_23753_, _23742_, _23245_);
  and _43995_ (_03125_, _23753_, _42618_);
  nor _43996_ (_23773_, _23289_, _23267_);
  nor _43997_ (_23784_, _23773_, _23300_);
  and _43998_ (_03328_, _23784_, _42618_);
  and _43999_ (_23815_, _23311_, _23082_);
  nor _44000_ (_23816_, _23815_, _23322_);
  and _44001_ (_03527_, _23816_, _42618_);
  nor _44002_ (_23837_, _23343_, _23006_);
  nor _44003_ (_23848_, _23837_, _23354_);
  and _44004_ (_03728_, _23848_, _42618_);
  and _44005_ (_23869_, _23365_, _22941_);
  nor _44006_ (_23879_, _23869_, _23386_);
  and _44007_ (_03927_, _23879_, _42618_);
  and _44008_ (_23900_, _23420_, _23387_);
  nor _44009_ (_23911_, _23900_, _23431_);
  and _44010_ (_04023_, _23911_, _42618_);
  and _44011_ (_23932_, _23442_, _22821_);
  nor _44012_ (_23943_, _23932_, _23452_);
  and _44013_ (_04123_, _23943_, _42618_);
  nor _44014_ (_23963_, _23474_, _18970_);
  nor _44015_ (_23974_, _23963_, _23485_);
  and _44016_ (_04222_, _23974_, _42618_);
  and _44017_ (_23995_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor _44018_ (_24006_, _23995_, _23485_);
  nor _44019_ (_24017_, _24006_, _23496_);
  and _44020_ (_04321_, _24017_, _42618_);
  nor _44021_ (_24038_, _23507_, _23496_);
  nor _44022_ (_24048_, _24038_, _23518_);
  and _44023_ (_04414_, _24048_, _42618_);
  and _44024_ (_24069_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor _44025_ (_24080_, _24069_, _23518_);
  nor _44026_ (_24091_, _24080_, _23529_);
  and _44027_ (_04512_, _24091_, _42618_);
  nor _44028_ (_24112_, _23529_, _18959_);
  nor _44029_ (_24122_, _24112_, _23540_);
  and _44030_ (_04611_, _24122_, _42618_);
  and _44031_ (_24143_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18772_);
  nor _44032_ (_24154_, _24143_, _18773_);
  not _44033_ (_24165_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _44034_ (_24176_, _18795_, _24165_);
  and _44035_ (_24187_, _24176_, _24154_);
  and _44036_ (_24198_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _44037_ (_24208_, _24198_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44038_ (_24219_, _24198_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44039_ (_24230_, _24219_, _24208_);
  and _44040_ (_00925_, _24230_, _42618_);
  and _44041_ (_00951_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _42618_);
  not _44042_ (_24261_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _44043_ (_24272_, _20536_, _24261_);
  and _44044_ (_24284_, _20220_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44045_ (_24294_, _24284_, _24272_);
  nor _44046_ (_24305_, _24294_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44047_ (_24316_, _20372_, _24261_);
  and _44048_ (_24327_, _20719_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _44049_ (_24338_, _24327_, _24316_);
  and _44050_ (_24349_, _24338_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44051_ (_24360_, _24349_, _24305_);
  nor _44052_ (_24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _44053_ (_24381_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and _44054_ (_24392_, _24371_, _20884_);
  nor _44055_ (_24403_, _24392_, _24381_);
  not _44056_ (_24414_, _24403_);
  and _44057_ (_24425_, _19550_, _24261_);
  and _44058_ (_24436_, _19222_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44059_ (_24447_, _24436_, _24425_);
  nor _44060_ (_24458_, _24447_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44061_ (_24468_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44062_ (_24479_, _19387_, _24261_);
  and _44063_ (_24490_, _19724_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44064_ (_24501_, _24490_, _24479_);
  nor _44065_ (_24522_, _24501_, _24468_);
  nor _44066_ (_24523_, _24522_, _24458_);
  nor _44067_ (_24534_, _24523_, _24414_);
  and _44068_ (_24544_, _24523_, _24414_);
  nor _44069_ (_24555_, _24544_, _24534_);
  nor _44070_ (_24566_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and _44071_ (_24577_, _24371_, _20046_);
  nor _44072_ (_24588_, _24577_, _24566_);
  not _44073_ (_24599_, _24588_);
  nor _44074_ (_24610_, _20536_, _24261_);
  nor _44075_ (_24621_, _24610_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44076_ (_24631_, _20220_, _24261_);
  and _44077_ (_24642_, _20372_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44078_ (_24653_, _24642_, _24631_);
  nor _44079_ (_24664_, _24653_, _24468_);
  nor _44080_ (_24675_, _24664_, _24621_);
  nor _44081_ (_24686_, _24675_, _24599_);
  and _44082_ (_24697_, _24675_, _24599_);
  nor _44083_ (_24707_, _24697_, _24686_);
  not _44084_ (_24718_, _24707_);
  nor _44085_ (_24729_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and _44086_ (_24740_, _24371_, _21080_);
  nor _44087_ (_24751_, _24740_, _24729_);
  not _44088_ (_24762_, _24751_);
  nor _44089_ (_24773_, _19550_, _24261_);
  nor _44090_ (_24784_, _24773_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44091_ (_24794_, _19222_, _24261_);
  and _44092_ (_24805_, _19387_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44093_ (_24816_, _24805_, _24794_);
  nor _44094_ (_24827_, _24816_, _24468_);
  nor _44095_ (_24838_, _24827_, _24784_);
  nor _44096_ (_24849_, _24838_, _24762_);
  and _44097_ (_24860_, _24838_, _24762_);
  and _44098_ (_24871_, _24294_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44099_ (_24881_, _24871_);
  nor _44100_ (_24892_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and _44101_ (_24903_, _24371_, _21254_);
  nor _44102_ (_24914_, _24903_, _24892_);
  and _44103_ (_24925_, _24914_, _24881_);
  and _44104_ (_24936_, _24447_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44105_ (_24947_, _24936_);
  and _44106_ (_24958_, _24371_, _21624_);
  nor _44107_ (_24968_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor _44108_ (_24979_, _24968_, _24958_);
  and _44109_ (_24990_, _24979_, _24947_);
  nor _44110_ (_25001_, _24979_, _24947_);
  nor _44111_ (_25012_, _25001_, _24990_);
  not _44112_ (_25023_, _25012_);
  and _44113_ (_25034_, _24610_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44114_ (_25045_, _25034_);
  and _44115_ (_25065_, _24371_, _22147_);
  nor _44116_ (_25066_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor _44117_ (_25077_, _25066_, _25065_);
  and _44118_ (_25088_, _25077_, _25045_);
  and _44119_ (_25099_, _24773_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44120_ (_25110_, _25099_);
  nor _44121_ (_25121_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and _44122_ (_25132_, _24371_, _21972_);
  nor _44123_ (_25143_, _25132_, _25121_);
  nor _44124_ (_25154_, _25143_, _25110_);
  not _44125_ (_25165_, _25154_);
  nor _44126_ (_25176_, _25077_, _25045_);
  nor _44127_ (_25187_, _25176_, _25088_);
  and _44128_ (_25198_, _25187_, _25165_);
  nor _44129_ (_25209_, _25198_, _25088_);
  nor _44130_ (_25220_, _25209_, _25023_);
  nor _44131_ (_25231_, _25220_, _24990_);
  nor _44132_ (_25242_, _24914_, _24881_);
  nor _44133_ (_25253_, _25242_, _24925_);
  not _44134_ (_25264_, _25253_);
  nor _44135_ (_25275_, _25264_, _25231_);
  nor _44136_ (_25286_, _25275_, _24925_);
  nor _44137_ (_25297_, _25286_, _24860_);
  nor _44138_ (_25308_, _25297_, _24849_);
  nor _44139_ (_25328_, _25308_, _24718_);
  nor _44140_ (_25329_, _25328_, _24686_);
  not _44141_ (_25340_, _25329_);
  and _44142_ (_25351_, _25340_, _24555_);
  or _44143_ (_25362_, _25351_, _24534_);
  and _44144_ (_25373_, _20719_, _19724_);
  or _44145_ (_25384_, _25373_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _44146_ (_25395_, _24501_);
  and _44147_ (_25406_, _24338_, _25395_);
  nor _44148_ (_25417_, _24816_, _24653_);
  and _44149_ (_25428_, _25417_, _25406_);
  or _44150_ (_25439_, _25428_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44151_ (_25450_, _25439_, _25384_);
  and _44152_ (_25461_, _25450_, _25362_);
  and _44153_ (_25472_, _25461_, _24360_);
  nor _44154_ (_25483_, _25340_, _24555_);
  or _44155_ (_25494_, _25483_, _25351_);
  and _44156_ (_25505_, _25494_, _25472_);
  nor _44157_ (_25516_, _25472_, _24403_);
  nor _44158_ (_25527_, _25516_, _25505_);
  not _44159_ (_25538_, _25527_);
  and _44160_ (_25549_, _25527_, _24360_);
  not _44161_ (_25560_, _24523_);
  nor _44162_ (_25571_, _25472_, _24599_);
  and _44163_ (_25582_, _25308_, _24718_);
  nor _44164_ (_25593_, _25582_, _25328_);
  and _44165_ (_25604_, _25593_, _25472_);
  or _44166_ (_25615_, _25604_, _25571_);
  and _44167_ (_25636_, _25615_, _25560_);
  nor _44168_ (_25637_, _25615_, _25560_);
  nor _44169_ (_25648_, _25637_, _25636_);
  not _44170_ (_25659_, _25648_);
  not _44171_ (_25670_, _24675_);
  nor _44172_ (_25681_, _25472_, _24762_);
  nor _44173_ (_25692_, _24860_, _24849_);
  nor _44174_ (_25702_, _25692_, _25286_);
  and _44175_ (_25713_, _25692_, _25286_);
  or _44176_ (_25724_, _25713_, _25702_);
  and _44177_ (_25735_, _25724_, _25472_);
  or _44178_ (_25746_, _25735_, _25681_);
  and _44179_ (_25757_, _25746_, _25670_);
  nor _44180_ (_25768_, _25746_, _25670_);
  not _44181_ (_25779_, _24838_);
  and _44182_ (_25790_, _25264_, _25231_);
  or _44183_ (_25801_, _25790_, _25275_);
  and _44184_ (_25812_, _25801_, _25472_);
  nor _44185_ (_25823_, _25472_, _24914_);
  nor _44186_ (_25834_, _25823_, _25812_);
  and _44187_ (_25845_, _25834_, _25779_);
  and _44188_ (_25856_, _25209_, _25023_);
  nor _44189_ (_25867_, _25856_, _25220_);
  not _44190_ (_25878_, _25867_);
  and _44191_ (_25889_, _25878_, _25472_);
  nor _44192_ (_25900_, _25472_, _24979_);
  nor _44193_ (_25911_, _25900_, _25889_);
  and _44194_ (_25922_, _25911_, _24881_);
  nor _44195_ (_25933_, _25911_, _24881_);
  nor _44196_ (_25944_, _25933_, _25922_);
  not _44197_ (_25965_, _25944_);
  nor _44198_ (_25966_, _25187_, _25165_);
  nor _44199_ (_25977_, _25966_, _25198_);
  not _44200_ (_25988_, _25977_);
  and _44201_ (_25999_, _25988_, _25472_);
  nor _44202_ (_26010_, _25472_, _25077_);
  nor _44203_ (_26021_, _26010_, _25999_);
  and _44204_ (_26032_, _26021_, _24947_);
  and _44205_ (_26043_, _25472_, _25099_);
  nor _44206_ (_26054_, _26043_, _25143_);
  and _44207_ (_26064_, _26043_, _25143_);
  nor _44208_ (_26075_, _26064_, _26054_);
  and _44209_ (_26086_, _26075_, _25045_);
  nor _44210_ (_26097_, _26075_, _25045_);
  nor _44211_ (_26108_, _26097_, _26086_);
  and _44212_ (_26119_, _24371_, _22517_);
  nor _44213_ (_26130_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _44214_ (_26141_, _26130_, _26119_);
  nor _44215_ (_26152_, _26141_, _25110_);
  not _44216_ (_26163_, _26152_);
  and _44217_ (_26174_, _26163_, _26108_);
  nor _44218_ (_26185_, _26174_, _26086_);
  nor _44219_ (_26196_, _26021_, _24947_);
  nor _44220_ (_26207_, _26196_, _26032_);
  not _44221_ (_26218_, _26207_);
  nor _44222_ (_26229_, _26218_, _26185_);
  nor _44223_ (_26240_, _26229_, _26032_);
  nor _44224_ (_26251_, _26240_, _25965_);
  nor _44225_ (_26262_, _26251_, _25922_);
  nor _44226_ (_26273_, _25834_, _25779_);
  nor _44227_ (_26284_, _26273_, _25845_);
  not _44228_ (_26295_, _26284_);
  nor _44229_ (_26306_, _26295_, _26262_);
  nor _44230_ (_26317_, _26306_, _25845_);
  nor _44231_ (_26328_, _26317_, _25768_);
  nor _44232_ (_26339_, _26328_, _25757_);
  nor _44233_ (_26350_, _26339_, _25659_);
  or _44234_ (_26361_, _26350_, _25636_);
  or _44235_ (_26372_, _26361_, _25549_);
  and _44236_ (_26383_, _26372_, _25450_);
  nor _44237_ (_26394_, _26383_, _25538_);
  and _44238_ (_26405_, _25549_, _25450_);
  and _44239_ (_26415_, _26405_, _26361_);
  or _44240_ (_26426_, _26415_, _26394_);
  and _44241_ (_00971_, _26426_, _42618_);
  or _44242_ (_26447_, _25527_, _24360_);
  and _44243_ (_26458_, _26447_, _26383_);
  and _44244_ (_02836_, _26458_, _42618_);
  and _44245_ (_02848_, _25472_, _42618_);
  and _44246_ (_02870_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _42618_);
  and _44247_ (_02894_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _42618_);
  and _44248_ (_02916_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _42618_);
  or _44249_ (_26519_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44250_ (_26530_, _24198_, rst);
  and _44251_ (_02927_, _26530_, _26519_);
  and _44252_ (_26551_, _26458_, _25099_);
  or _44253_ (_26562_, _26551_, _26141_);
  nand _44254_ (_26573_, _26551_, _26141_);
  and _44255_ (_26584_, _26573_, _26562_);
  and _44256_ (_02940_, _26584_, _42618_);
  nor _44257_ (_26605_, _26163_, _26108_);
  or _44258_ (_26616_, _26605_, _26174_);
  nand _44259_ (_26627_, _26616_, _26458_);
  or _44260_ (_26638_, _26458_, _26075_);
  and _44261_ (_26649_, _26638_, _26627_);
  and _44262_ (_02954_, _26649_, _42618_);
  and _44263_ (_26670_, _26218_, _26185_);
  or _44264_ (_26681_, _26670_, _26229_);
  nand _44265_ (_26692_, _26681_, _26458_);
  or _44266_ (_26703_, _26458_, _26021_);
  and _44267_ (_26714_, _26703_, _26692_);
  and _44268_ (_02967_, _26714_, _42618_);
  and _44269_ (_26735_, _26240_, _25965_);
  or _44270_ (_26746_, _26735_, _26251_);
  nand _44271_ (_26756_, _26746_, _26458_);
  or _44272_ (_26767_, _26458_, _25911_);
  and _44273_ (_26778_, _26767_, _26756_);
  and _44274_ (_02981_, _26778_, _42618_);
  and _44275_ (_26799_, _26295_, _26262_);
  or _44276_ (_26810_, _26799_, _26306_);
  nand _44277_ (_26821_, _26810_, _26458_);
  or _44278_ (_26832_, _26458_, _25834_);
  and _44279_ (_26843_, _26832_, _26821_);
  and _44280_ (_02995_, _26843_, _42618_);
  or _44281_ (_26864_, _25768_, _25757_);
  and _44282_ (_26875_, _26864_, _26317_);
  nor _44283_ (_26886_, _26864_, _26317_);
  or _44284_ (_26897_, _26886_, _26875_);
  nand _44285_ (_26908_, _26897_, _26458_);
  or _44286_ (_26919_, _26458_, _25746_);
  and _44287_ (_26930_, _26919_, _26908_);
  and _44288_ (_03008_, _26930_, _42618_);
  and _44289_ (_26951_, _26339_, _25659_);
  or _44290_ (_26962_, _26951_, _26350_);
  nand _44291_ (_26973_, _26962_, _26458_);
  or _44292_ (_26984_, _26458_, _25615_);
  and _44293_ (_26995_, _26984_, _26973_);
  and _44294_ (_03022_, _26995_, _42618_);
  and _44295_ (_27016_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44296_ (_27027_, _27016_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _44297_ (_27038_, _27027_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _44298_ (_27049_, _27038_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _44299_ (_27060_, _27049_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _44300_ (_27071_, _27060_);
  not _44301_ (_27082_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44302_ (_27093_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18772_);
  and _44303_ (_27103_, _27093_, _27082_);
  and _44304_ (_27114_, _27103_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  not _44305_ (_27125_, _27114_);
  nor _44306_ (_27136_, _27049_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _44307_ (_27147_, _27136_, _27125_);
  and _44308_ (_27158_, _27147_, _27071_);
  not _44309_ (_27169_, _27158_);
  and _44310_ (_27180_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44311_ (_27191_, _27180_, _27093_);
  not _44312_ (_27202_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _44313_ (_27213_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18772_);
  and _44314_ (_27224_, _27213_, _27202_);
  and _44315_ (_27245_, _27224_, _27082_);
  and _44316_ (_27246_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _44317_ (_27257_, _27246_, _27191_);
  not _44318_ (_27268_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _44319_ (_27279_, _27103_, _27268_);
  and _44320_ (_27290_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _44321_ (_27301_, _27224_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44322_ (_27312_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _44323_ (_27323_, _27312_, _27290_);
  and _44324_ (_27334_, _27323_, _27257_);
  and _44325_ (_27345_, _27334_, _27169_);
  and _44326_ (_27356_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not _44327_ (_27367_, _27356_);
  and _44328_ (_27378_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _44329_ (_27389_, _27378_, _27191_);
  and _44330_ (_27400_, _27389_, _27367_);
  nor _44331_ (_27411_, _27038_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _44332_ (_27422_, _27411_);
  nor _44333_ (_27433_, _27125_, _27049_);
  and _44334_ (_27444_, _27433_, _27422_);
  or _44335_ (_27454_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44336_ (_27465_, _27454_, _18772_);
  nor _44337_ (_27476_, _27465_, _27213_);
  and _44338_ (_27487_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and _44339_ (_27498_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor _44340_ (_27509_, _27498_, _27487_);
  not _44341_ (_27520_, _27509_);
  nor _44342_ (_27531_, _27520_, _27444_);
  and _44343_ (_27542_, _27531_, _27400_);
  nor _44344_ (_27553_, _27542_, _27345_);
  nor _44345_ (_27564_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _44346_ (_27575_, _27564_, _27016_);
  and _44347_ (_27586_, _27575_, _27114_);
  and _44348_ (_27597_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _44349_ (_27608_, _27597_, _27586_);
  and _44350_ (_27619_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _44351_ (_27630_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and _44352_ (_27641_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or _44353_ (_27652_, _27641_, _27630_);
  nor _44354_ (_27663_, _27652_, _27619_);
  and _44355_ (_27674_, _27663_, _27608_);
  and _44356_ (_27685_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and _44357_ (_27696_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor _44358_ (_27707_, _27696_, _27685_);
  and _44359_ (_27718_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not _44360_ (_27729_, _27718_);
  not _44361_ (_27740_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44362_ (_27751_, _27114_, _27740_);
  and _44363_ (_27762_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _44364_ (_27773_, _27762_, _27751_);
  and _44365_ (_27784_, _27773_, _27729_);
  and _44366_ (_27795_, _27784_, _27707_);
  and _44367_ (_27806_, _27795_, _27674_);
  not _44368_ (_27816_, _27038_);
  nor _44369_ (_27827_, _27027_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _44370_ (_27838_, _27827_, _27125_);
  and _44371_ (_27849_, _27838_, _27816_);
  not _44372_ (_27860_, _27849_);
  and _44373_ (_27881_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _44374_ (_27882_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _44375_ (_27893_, _27882_, _27881_);
  and _44376_ (_27904_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _44377_ (_27915_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _44378_ (_27926_, _27915_, _27904_);
  and _44379_ (_27937_, _27926_, _27893_);
  and _44380_ (_27948_, _27937_, _27860_);
  nor _44381_ (_27959_, _27016_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44382_ (_27970_, _27959_, _27027_);
  and _44383_ (_27981_, _27970_, _27114_);
  and _44384_ (_27992_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _44385_ (_28003_, _27992_, _27981_);
  and _44386_ (_28014_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _44387_ (_28025_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and _44388_ (_28036_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _44389_ (_28047_, _28036_, _28025_);
  nor _44390_ (_28058_, _28047_, _28014_);
  and _44391_ (_28069_, _28058_, _28003_);
  and _44392_ (_28080_, _28069_, _27948_);
  and _44393_ (_28091_, _28080_, _27806_);
  not _44394_ (_28102_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and _44395_ (_28113_, _27060_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _44396_ (_28124_, _28113_, _28102_);
  and _44397_ (_28135_, _28113_, _28102_);
  nor _44398_ (_28145_, _28135_, _28124_);
  nor _44399_ (_28156_, _28145_, _27125_);
  not _44400_ (_28167_, _28156_);
  and _44401_ (_28188_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nor _44402_ (_28189_, _28188_, _27191_);
  and _44403_ (_28200_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and _44404_ (_28211_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor _44405_ (_28222_, _28211_, _28200_);
  and _44406_ (_28233_, _28222_, _28189_);
  and _44407_ (_28244_, _28233_, _28167_);
  not _44408_ (_28255_, _28113_);
  nor _44409_ (_28266_, _27060_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _44410_ (_28277_, _28266_, _27125_);
  and _44411_ (_28288_, _28277_, _28255_);
  not _44412_ (_28299_, _28288_);
  and _44413_ (_28310_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _44414_ (_28321_, _28310_, _27191_);
  and _44415_ (_28332_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _44416_ (_28343_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _44417_ (_28354_, _28343_, _28332_);
  and _44418_ (_28365_, _28354_, _28321_);
  and _44419_ (_28376_, _28365_, _28299_);
  nor _44420_ (_28387_, _28376_, _28244_);
  and _44421_ (_28398_, _28387_, _28091_);
  nand _44422_ (_28409_, _28398_, _27553_);
  and _44423_ (_28420_, _26426_, _24187_);
  not _44424_ (_28431_, _28420_);
  and _44425_ (_28442_, _23594_, _18828_);
  not _44426_ (_28453_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _44427_ (_28463_, _24143_, _28453_);
  and _44428_ (_28474_, _28463_, _18817_);
  nor _44429_ (_28485_, _20046_, _19724_);
  and _44430_ (_28496_, _20046_, _19724_);
  nor _44431_ (_28507_, _28496_, _28485_);
  not _44432_ (_28518_, _28507_);
  nor _44433_ (_28539_, _21080_, _20372_);
  nor _44434_ (_28540_, _21254_, _19387_);
  and _44435_ (_28551_, _21080_, _20372_);
  nor _44436_ (_28562_, _28551_, _28539_);
  and _44437_ (_28573_, _28562_, _28540_);
  nor _44438_ (_28584_, _28573_, _28539_);
  nor _44439_ (_28595_, _28584_, _28518_);
  and _44440_ (_28606_, _21254_, _19387_);
  nor _44441_ (_28617_, _28606_, _28540_);
  nor _44442_ (_28628_, _21624_, _20220_);
  and _44443_ (_28639_, _21624_, _20220_);
  nor _44444_ (_28650_, _28639_, _28628_);
  nor _44445_ (_28661_, _22147_, _19222_);
  and _44446_ (_28672_, _22147_, _19222_);
  nor _44447_ (_28683_, _28672_, _28661_);
  not _44448_ (_28694_, _28683_);
  nor _44449_ (_28705_, _21972_, _20536_);
  nor _44450_ (_28716_, _22517_, _19550_);
  and _44451_ (_28727_, _21972_, _20536_);
  nor _44452_ (_28738_, _28727_, _28705_);
  and _44453_ (_28749_, _28738_, _28716_);
  nor _44454_ (_28760_, _28749_, _28705_);
  nor _44455_ (_28770_, _28760_, _28694_);
  nor _44456_ (_28781_, _28770_, _28661_);
  nor _44457_ (_28792_, _28781_, _28650_);
  and _44458_ (_28803_, _28781_, _28650_);
  nor _44459_ (_28814_, _28803_, _28792_);
  not _44460_ (_28825_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _44461_ (_28836_, _19036_, _28825_);
  not _44462_ (_28847_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _44463_ (_28858_, _28847_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44464_ (_28869_, _28858_, _19080_);
  nor _44465_ (_28880_, _28869_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not _44466_ (_28891_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44467_ (_28912_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _28891_);
  and _44468_ (_28913_, _28912_, _20427_);
  not _44469_ (_28924_, _28913_);
  and _44470_ (_28935_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44471_ (_28946_, _28935_, _20112_);
  nor _44472_ (_28957_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44473_ (_28968_, _28957_, _19441_);
  nor _44474_ (_28979_, _28968_, _28946_);
  and _44475_ (_28990_, _28979_, _28924_);
  and _44476_ (_29001_, _28990_, _28880_);
  not _44477_ (_29012_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _44478_ (_29023_, _28858_, _19615_);
  nor _44479_ (_29034_, _29023_, _29012_);
  and _44480_ (_29045_, _28957_, _19277_);
  not _44481_ (_29056_, _29045_);
  and _44482_ (_29067_, _28935_, _20601_);
  and _44483_ (_29077_, _28912_, _20264_);
  nor _44484_ (_29088_, _29077_, _29067_);
  and _44485_ (_29099_, _29088_, _29056_);
  and _44486_ (_29110_, _29099_, _29034_);
  nor _44487_ (_29121_, _29110_, _29001_);
  nor _44488_ (_29132_, _29121_, _19036_);
  nor _44489_ (_29143_, _29132_, _28836_);
  and _44490_ (_29154_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _44491_ (_29165_, _29154_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _44492_ (_29176_, _29165_);
  and _44493_ (_29187_, _29176_, _29143_);
  and _44494_ (_29198_, _29176_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _44495_ (_29209_, _29198_, _29187_);
  and _44496_ (_29220_, _22517_, _19550_);
  nor _44497_ (_29231_, _29220_, _28716_);
  not _44498_ (_29242_, _29231_);
  nor _44499_ (_29253_, _29242_, _29209_);
  and _44500_ (_29264_, _29253_, _28738_);
  and _44501_ (_29275_, _28760_, _28694_);
  nor _44502_ (_29286_, _29275_, _28770_);
  and _44503_ (_29297_, _29286_, _29264_);
  not _44504_ (_29308_, _29297_);
  nor _44505_ (_29319_, _29308_, _28814_);
  nor _44506_ (_29330_, _28781_, _28639_);
  or _44507_ (_29341_, _29330_, _28628_);
  or _44508_ (_29352_, _29341_, _29319_);
  and _44509_ (_29363_, _29352_, _28617_);
  nor _44510_ (_29373_, _28562_, _28540_);
  nor _44511_ (_29384_, _29373_, _28573_);
  and _44512_ (_29395_, _29384_, _29363_);
  and _44513_ (_29406_, _28584_, _28518_);
  nor _44514_ (_29417_, _29406_, _28595_);
  and _44515_ (_29438_, _29417_, _29395_);
  or _44516_ (_29439_, _29438_, _28595_);
  nor _44517_ (_29450_, _29439_, _28485_);
  nor _44518_ (_29461_, _20884_, _20719_);
  and _44519_ (_29472_, _20884_, _20719_);
  nor _44520_ (_29483_, _29472_, _29461_);
  not _44521_ (_29494_, _29483_);
  nor _44522_ (_29505_, _29494_, _29450_);
  and _44523_ (_29516_, _29494_, _29450_);
  nor _44524_ (_29527_, _29516_, _29505_);
  and _44525_ (_29538_, _29527_, _28474_);
  not _44526_ (_29549_, _29538_);
  not _44527_ (_29560_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _44528_ (_29571_, _18773_, _29560_);
  and _44529_ (_29582_, _29571_, _18817_);
  not _44530_ (_29593_, _29582_);
  not _44531_ (_29604_, _19724_);
  nor _44532_ (_29615_, _20046_, _29604_);
  and _44533_ (_29626_, _21090_, _20372_);
  not _44534_ (_29637_, _19387_);
  and _44535_ (_29648_, _21254_, _29637_);
  nor _44536_ (_29659_, _29648_, _28562_);
  nor _44537_ (_29670_, _29659_, _29626_);
  nor _44538_ (_29680_, _29670_, _28507_);
  nor _44539_ (_29691_, _29680_, _29615_);
  and _44540_ (_29712_, _29670_, _28507_);
  nor _44541_ (_29713_, _29712_, _29680_);
  not _44542_ (_29724_, _29713_);
  and _44543_ (_29735_, _29648_, _28562_);
  nor _44544_ (_29746_, _29735_, _29659_);
  not _44545_ (_29757_, _29746_);
  not _44546_ (_29768_, _28617_);
  not _44547_ (_29779_, _28650_);
  not _44548_ (_29790_, _19550_);
  and _44549_ (_29801_, _22517_, _29790_);
  nor _44550_ (_29812_, _29801_, _28738_);
  not _44551_ (_29823_, _20536_);
  nor _44552_ (_29834_, _21972_, _29823_);
  nor _44553_ (_29845_, _29834_, _29812_);
  nor _44554_ (_29856_, _29845_, _28683_);
  not _44555_ (_29867_, _19222_);
  nor _44556_ (_29878_, _22147_, _29867_);
  nor _44557_ (_29889_, _29878_, _29856_);
  nor _44558_ (_29900_, _29889_, _29779_);
  and _44559_ (_29911_, _29889_, _29779_);
  nor _44560_ (_29922_, _29911_, _29900_);
  and _44561_ (_29933_, _29845_, _28683_);
  nor _44562_ (_29944_, _29933_, _29856_);
  not _44563_ (_29955_, _29944_);
  and _44564_ (_29966_, _29801_, _28738_);
  nor _44565_ (_29976_, _29966_, _29812_);
  not _44566_ (_29987_, _29976_);
  nor _44567_ (_29998_, _29231_, _29209_);
  and _44568_ (_30009_, _29998_, _29987_);
  and _44569_ (_30020_, _30009_, _29955_);
  and _44570_ (_30031_, _30020_, _29922_);
  not _44571_ (_30042_, _20220_);
  or _44572_ (_30053_, _21624_, _30042_);
  and _44573_ (_30064_, _21624_, _30042_);
  or _44574_ (_30075_, _29889_, _30064_);
  and _44575_ (_30085_, _30075_, _30053_);
  or _44576_ (_30096_, _30085_, _30031_);
  and _44577_ (_30107_, _30096_, _29768_);
  and _44578_ (_30118_, _30107_, _29757_);
  and _44579_ (_30129_, _30118_, _29724_);
  nor _44580_ (_30140_, _30129_, _29691_);
  nor _44581_ (_30151_, _30140_, _29483_);
  and _44582_ (_30162_, _30140_, _29483_);
  nor _44583_ (_30173_, _30162_, _30151_);
  nor _44584_ (_30184_, _30173_, _29593_);
  and _44585_ (_30194_, _18806_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _44586_ (_30205_, _30194_, _29571_);
  nor _44587_ (_30216_, _22517_, _21972_);
  and _44588_ (_30227_, _30216_, _22158_);
  and _44589_ (_30238_, _30227_, _21635_);
  and _44590_ (_30249_, _30238_, _21265_);
  and _44591_ (_30260_, _30249_, _21090_);
  and _44592_ (_30271_, _30260_, _20057_);
  and _44593_ (_30282_, _30271_, _29209_);
  not _44594_ (_30293_, _29209_);
  and _44595_ (_30303_, _21080_, _20046_);
  and _44596_ (_30314_, _22517_, _21972_);
  and _44597_ (_30335_, _30314_, _22147_);
  and _44598_ (_30336_, _30335_, _21624_);
  and _44599_ (_30347_, _30336_, _21254_);
  and _44600_ (_30358_, _30347_, _30303_);
  and _44601_ (_30369_, _30358_, _30293_);
  nor _44602_ (_30380_, _30369_, _30282_);
  and _44603_ (_30391_, _30380_, _20884_);
  nor _44604_ (_30402_, _30380_, _20884_);
  nor _44605_ (_30412_, _30402_, _30391_);
  and _44606_ (_30423_, _30412_, _30205_);
  not _44607_ (_30434_, _20719_);
  nor _44608_ (_30445_, _29209_, _30434_);
  not _44609_ (_30456_, _30445_);
  and _44610_ (_30467_, _29209_, _20884_);
  and _44611_ (_30478_, _30194_, _18784_);
  not _44612_ (_30489_, _30478_);
  nor _44613_ (_30500_, _30489_, _30467_);
  and _44614_ (_30511_, _30500_, _30456_);
  nor _44615_ (_30522_, _30511_, _30423_);
  and _44616_ (_30532_, _28463_, _24176_);
  not _44617_ (_30543_, _30532_);
  and _44618_ (_30554_, _22147_, _21972_);
  nor _44619_ (_30565_, _30554_, _21624_);
  and _44620_ (_30576_, _30565_, _30532_);
  and _44621_ (_30587_, _30576_, _21265_);
  nor _44622_ (_30598_, _30587_, _21090_);
  and _44623_ (_30609_, _30598_, _20046_);
  nor _44624_ (_30620_, _30303_, _20884_);
  nor _44625_ (_30631_, _30620_, _30576_);
  and _44626_ (_30641_, _30631_, _29209_);
  nor _44627_ (_30652_, _30641_, _30609_);
  and _44628_ (_30663_, _30652_, _20884_);
  nor _44629_ (_30674_, _30652_, _20884_);
  nor _44630_ (_30685_, _30674_, _30663_);
  nor _44631_ (_30696_, _30685_, _30543_);
  not _44632_ (_30707_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _44633_ (_30718_, _18806_, _30707_);
  and _44634_ (_30729_, _30718_, _28463_);
  not _44635_ (_30740_, _30729_);
  nor _44636_ (_30750_, _30740_, _29472_);
  and _44637_ (_30761_, _30718_, _24154_);
  and _44638_ (_30772_, _30761_, _29483_);
  nor _44639_ (_30783_, _30772_, _30750_);
  and _44640_ (_30794_, _30194_, _24154_);
  not _44641_ (_30805_, _30794_);
  nor _44642_ (_30816_, _30805_, _22517_);
  and _44643_ (_30827_, _30718_, _18773_);
  not _44644_ (_30838_, _30827_);
  nor _44645_ (_30849_, _30838_, _20046_);
  nor _44646_ (_30859_, _30849_, _30816_);
  and _44647_ (_30870_, _30194_, _28463_);
  not _44648_ (_30881_, _30870_);
  nor _44649_ (_30892_, _30881_, _29209_);
  and _44650_ (_30903_, _24176_, _18784_);
  and _44651_ (_30914_, _30903_, _29461_);
  and _44652_ (_30925_, _29571_, _24176_);
  and _44653_ (_30936_, _30925_, _20884_);
  nor _44654_ (_30947_, _30936_, _30914_);
  and _44655_ (_30958_, _24154_, _18817_);
  not _44656_ (_30968_, _30958_);
  nor _44657_ (_30979_, _30968_, _20884_);
  not _44658_ (_30990_, _30979_);
  nand _44659_ (_31001_, _30990_, _30947_);
  nor _44660_ (_31012_, _31001_, _30892_);
  and _44661_ (_31023_, _31012_, _30859_);
  and _44662_ (_31045_, _31023_, _30783_);
  not _44663_ (_31046_, _31045_);
  nor _44664_ (_31068_, _31046_, _30696_);
  and _44665_ (_31069_, _31068_, _30522_);
  not _44666_ (_31090_, _31069_);
  nor _44667_ (_31091_, _31090_, _30184_);
  and _44668_ (_31113_, _31091_, _29549_);
  not _44669_ (_31114_, _31113_);
  nor _44670_ (_31125_, _31114_, _28442_);
  and _44671_ (_31136_, _31125_, _28431_);
  not _44672_ (_31147_, _31136_);
  or _44673_ (_31168_, _31147_, _28409_);
  not _44674_ (_31169_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _44675_ (_31189_, \oc8051_top_1.oc8051_decoder1.wr , _18772_);
  not _44676_ (_31190_, _31189_);
  nor _44677_ (_31211_, _31190_, _27103_);
  and _44678_ (_31212_, _31211_, _31169_);
  not _44679_ (_31233_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _44680_ (_31234_, _28409_, _31233_);
  and _44681_ (_31255_, _31234_, _31212_);
  and _44682_ (_31256_, _31255_, _31168_);
  nor _44683_ (_31277_, _31211_, _31233_);
  not _44684_ (_31278_, _28474_);
  nor _44685_ (_31299_, _29505_, _29461_);
  nor _44686_ (_31300_, _31299_, _31278_);
  not _44687_ (_31320_, _31300_);
  and _44688_ (_31321_, _20884_, _30434_);
  nor _44689_ (_31342_, _31321_, _30151_);
  nor _44690_ (_31343_, _31342_, _29593_);
  and _44691_ (_31364_, _29209_, _20046_);
  and _44692_ (_31365_, _31364_, _30598_);
  nor _44693_ (_31386_, _31365_, _30467_);
  nor _44694_ (_31387_, _29209_, _20884_);
  not _44695_ (_31408_, _31387_);
  nor _44696_ (_31409_, _31408_, _30609_);
  nor _44697_ (_31429_, _31409_, _30543_);
  and _44698_ (_31430_, _31429_, _31386_);
  nor _44699_ (_31451_, _30925_, _30293_);
  and _44700_ (_31452_, _30805_, _29198_);
  nor _44701_ (_31473_, _31452_, _29187_);
  not _44702_ (_31474_, _31473_);
  nor _44703_ (_31495_, _31474_, _31451_);
  nor _44704_ (_31496_, _29198_, _29143_);
  not _44705_ (_31517_, _30761_);
  nor _44706_ (_31518_, _31517_, _29187_);
  nor _44707_ (_31538_, _31518_, _30729_);
  nor _44708_ (_31539_, _31538_, _31496_);
  and _44709_ (_31560_, _29165_, _29143_);
  and _44710_ (_31561_, _30718_, _29571_);
  and _44711_ (_31582_, _30903_, _29143_);
  nor _44712_ (_31583_, _31582_, _31561_);
  nor _44713_ (_31604_, _31583_, _31560_);
  nor _44714_ (_31605_, _30968_, _29209_);
  and _44715_ (_31626_, _30718_, _18784_);
  not _44716_ (_31627_, _31626_);
  nor _44717_ (_31647_, _31627_, _20884_);
  nor _44718_ (_31648_, _30881_, _22517_);
  or _44719_ (_31669_, _31648_, _30576_);
  or _44720_ (_31670_, _31669_, _31647_);
  or _44721_ (_31691_, _31670_, _31605_);
  or _44722_ (_31692_, _31691_, _31604_);
  or _44723_ (_31713_, _31692_, _31539_);
  or _44724_ (_31714_, _31713_, _31495_);
  nor _44725_ (_31735_, _31714_, _31430_);
  not _44726_ (_31736_, _31735_);
  nor _44727_ (_31756_, _31736_, _31343_);
  and _44728_ (_31757_, _31756_, _31320_);
  nor _44729_ (_31768_, _28376_, _27345_);
  not _44730_ (_31779_, _28244_);
  not _44731_ (_31790_, _27948_);
  nor _44732_ (_31801_, _31790_, _27542_);
  and _44733_ (_31812_, _31801_, _31779_);
  and _44734_ (_31823_, _31812_, _31768_);
  not _44735_ (_31834_, _28069_);
  nor _44736_ (_31845_, _27795_, _27674_);
  and _44737_ (_31855_, _31845_, _31834_);
  and _44738_ (_31866_, _31855_, _31823_);
  nand _44739_ (_31877_, _31866_, _31757_);
  or _44740_ (_31888_, _31866_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _44741_ (_31899_, _31211_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _44742_ (_31910_, _31899_, _31888_);
  and _44743_ (_31921_, _31910_, _31877_);
  or _44744_ (_31932_, _31921_, _31277_);
  or _44745_ (_31943_, _31932_, _31256_);
  and _44746_ (_06626_, _31943_, _42618_);
  and _44747_ (_31963_, _26584_, _24187_);
  not _44748_ (_31974_, _31963_);
  and _44749_ (_31985_, _29242_, _29209_);
  nor _44750_ (_31996_, _31985_, _29253_);
  nand _44751_ (_32007_, _31996_, _28474_);
  and _44752_ (_32018_, _30903_, _28716_);
  and _44753_ (_32029_, _30925_, _22517_);
  nor _44754_ (_32040_, _32029_, _32018_);
  nor _44755_ (_32051_, _31517_, _28716_);
  nor _44756_ (_32062_, _32051_, _30729_);
  or _44757_ (_32073_, _32062_, _29220_);
  and _44758_ (_32083_, _30194_, _28453_);
  not _44759_ (_32094_, _32083_);
  nor _44760_ (_32105_, _32094_, _21972_);
  and _44761_ (_32116_, _31561_, _20895_);
  nor _44762_ (_32127_, _32116_, _32105_);
  and _44763_ (_32138_, _32127_, _32073_);
  and _44764_ (_32149_, _32138_, _32040_);
  and _44765_ (_32160_, _23911_, _18828_);
  and _44766_ (_32171_, _31996_, _29582_);
  nor _44767_ (_32182_, _31627_, _29209_);
  nor _44768_ (_32192_, _30489_, _19550_);
  and _44769_ (_32203_, _30205_, _22517_);
  nor _44770_ (_32214_, _32203_, _32192_);
  nor _44771_ (_32225_, _30958_, _30532_);
  nor _44772_ (_32236_, _32225_, _22517_);
  not _44773_ (_32247_, _32236_);
  nand _44774_ (_32258_, _32247_, _32214_);
  or _44775_ (_32269_, _32258_, _32182_);
  or _44776_ (_32280_, _32269_, _32171_);
  nor _44777_ (_32291_, _32280_, _32160_);
  and _44778_ (_32301_, _32291_, _32149_);
  and _44779_ (_32312_, _32301_, _32007_);
  and _44780_ (_32323_, _32312_, _31974_);
  not _44781_ (_32334_, _32323_);
  or _44782_ (_32345_, _32334_, _28409_);
  not _44783_ (_32356_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _44784_ (_32367_, _28409_, _32356_);
  and _44785_ (_32378_, _32367_, _31212_);
  and _44786_ (_32389_, _32378_, _32345_);
  nor _44787_ (_32399_, _31211_, _32356_);
  not _44788_ (_32410_, _31757_);
  or _44789_ (_32421_, _32410_, _28409_);
  and _44790_ (_32432_, _32367_, _31899_);
  and _44791_ (_32443_, _32432_, _32421_);
  or _44792_ (_32454_, _32443_, _32399_);
  or _44793_ (_32465_, _32454_, _32389_);
  and _44794_ (_08867_, _32465_, _42618_);
  and _44795_ (_32486_, _23943_, _18828_);
  not _44796_ (_32497_, _32486_);
  and _44797_ (_32508_, _26649_, _24187_);
  nor _44798_ (_32518_, _28738_, _28716_);
  or _44799_ (_32529_, _32518_, _28749_);
  and _44800_ (_32540_, _32529_, _29253_);
  nor _44801_ (_32551_, _32529_, _29253_);
  or _44802_ (_32562_, _32551_, _32540_);
  and _44803_ (_32573_, _32562_, _28474_);
  not _44804_ (_32584_, _32573_);
  nor _44805_ (_32595_, _30565_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _44806_ (_32606_, _32595_, _21983_);
  nor _44807_ (_32617_, _32595_, _21983_);
  nor _44808_ (_32627_, _32617_, _32606_);
  nor _44809_ (_32638_, _32627_, _30543_);
  not _44810_ (_32649_, _32638_);
  and _44811_ (_32660_, _30761_, _28738_);
  nor _44812_ (_32671_, _30740_, _28727_);
  not _44813_ (_32682_, _32671_);
  and _44814_ (_32693_, _30903_, _28705_);
  and _44815_ (_32704_, _30925_, _21972_);
  nor _44816_ (_32715_, _32704_, _32693_);
  nand _44817_ (_32726_, _32715_, _32682_);
  nor _44818_ (_32736_, _32726_, _32660_);
  nor _44819_ (_32747_, _32094_, _22147_);
  not _44820_ (_32758_, _32747_);
  nor _44821_ (_32769_, _30968_, _21972_);
  nor _44822_ (_32780_, _30838_, _22517_);
  nor _44823_ (_32791_, _32780_, _32769_);
  and _44824_ (_32802_, _32791_, _32758_);
  and _44825_ (_32813_, _32802_, _32736_);
  and _44826_ (_32824_, _32813_, _32649_);
  and _44827_ (_32835_, _32824_, _32584_);
  nor _44828_ (_32845_, _30489_, _20536_);
  nor _44829_ (_32856_, _30314_, _30216_);
  not _44830_ (_32867_, _32856_);
  nor _44831_ (_32878_, _32867_, _29209_);
  and _44832_ (_32889_, _32867_, _29209_);
  nor _44833_ (_32900_, _32889_, _32878_);
  and _44834_ (_32911_, _32900_, _30205_);
  nor _44835_ (_32922_, _32911_, _32845_);
  not _44836_ (_32933_, _32922_);
  nor _44837_ (_32944_, _29998_, _29987_);
  nor _44838_ (_32955_, _32944_, _30009_);
  nor _44839_ (_32965_, _32955_, _29593_);
  nor _44840_ (_32976_, _32965_, _32933_);
  and _44841_ (_32987_, _32976_, _32835_);
  not _44842_ (_32998_, _32987_);
  nor _44843_ (_33009_, _32998_, _32508_);
  and _44844_ (_33020_, _33009_, _32497_);
  not _44845_ (_33031_, _33020_);
  or _44846_ (_33042_, _33031_, _28409_);
  not _44847_ (_33053_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _44848_ (_33064_, _28409_, _33053_);
  and _44849_ (_33074_, _33064_, _31212_);
  and _44850_ (_33085_, _33074_, _33042_);
  nor _44851_ (_33096_, _31211_, _33053_);
  not _44852_ (_33107_, _27674_);
  nor _44853_ (_33118_, _27795_, _33107_);
  and _44854_ (_33129_, _33118_, _28069_);
  and _44855_ (_33140_, _33129_, _31823_);
  nand _44856_ (_33151_, _33140_, _31757_);
  or _44857_ (_33162_, _33140_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _44858_ (_33172_, _33162_, _31899_);
  and _44859_ (_33183_, _33172_, _33151_);
  or _44860_ (_33194_, _33183_, _33096_);
  or _44861_ (_33205_, _33194_, _33085_);
  and _44862_ (_08878_, _33205_, _42618_);
  and _44863_ (_33226_, _26714_, _24187_);
  not _44864_ (_33237_, _33226_);
  and _44865_ (_33248_, _23974_, _18828_);
  nor _44866_ (_33259_, _30489_, _19222_);
  and _44867_ (_33270_, _30314_, _30293_);
  and _44868_ (_33281_, _30216_, _29209_);
  nor _44869_ (_33291_, _33281_, _33270_);
  nor _44870_ (_33302_, _33291_, _22147_);
  not _44871_ (_33313_, _30205_);
  and _44872_ (_33324_, _33291_, _22147_);
  or _44873_ (_33335_, _33324_, _33313_);
  nor _44874_ (_33346_, _33335_, _33302_);
  nor _44875_ (_33357_, _33346_, _33259_);
  nor _44876_ (_33368_, _30009_, _29955_);
  nor _44877_ (_33379_, _33368_, _30020_);
  nor _44878_ (_33390_, _33379_, _29593_);
  and _44879_ (_33400_, _30761_, _28683_);
  nor _44880_ (_33411_, _30740_, _28672_);
  not _44881_ (_33422_, _33411_);
  and _44882_ (_33433_, _30903_, _28661_);
  and _44883_ (_33444_, _30925_, _22147_);
  nor _44884_ (_33455_, _33444_, _33433_);
  nand _44885_ (_33466_, _33455_, _33422_);
  nor _44886_ (_33477_, _33466_, _33400_);
  nor _44887_ (_33488_, _30838_, _21972_);
  not _44888_ (_33499_, _33488_);
  nor _44889_ (_33509_, _30968_, _22147_);
  nor _44890_ (_33520_, _32094_, _21624_);
  nor _44891_ (_33531_, _33520_, _33509_);
  and _44892_ (_33542_, _33531_, _33499_);
  and _44893_ (_33553_, _33542_, _33477_);
  not _44894_ (_33564_, _33553_);
  nor _44895_ (_33575_, _33564_, _33390_);
  nor _44896_ (_33586_, _29286_, _29264_);
  nor _44897_ (_33597_, _33586_, _31278_);
  and _44898_ (_33608_, _33597_, _29308_);
  nor _44899_ (_33618_, _32617_, _22147_);
  and _44900_ (_33629_, _30554_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _44901_ (_33640_, _33629_, _33618_);
  nor _44902_ (_33651_, _33640_, _30543_);
  nor _44903_ (_33662_, _33651_, _33608_);
  and _44904_ (_33673_, _33662_, _33575_);
  and _44905_ (_33684_, _33673_, _33357_);
  not _44906_ (_33695_, _33684_);
  nor _44907_ (_33706_, _33695_, _33248_);
  and _44908_ (_33717_, _33706_, _33237_);
  not _44909_ (_33728_, _33717_);
  or _44910_ (_33738_, _33728_, _28409_);
  not _44911_ (_33749_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _44912_ (_33760_, _28409_, _33749_);
  and _44913_ (_33771_, _33760_, _31212_);
  and _44914_ (_33782_, _33771_, _33738_);
  nor _44915_ (_33793_, _31211_, _33749_);
  nand _44916_ (_33804_, _31823_, _28069_);
  or _44917_ (_33815_, _31845_, _33804_);
  and _44918_ (_33826_, _33815_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _44919_ (_33837_, _28069_, _27795_);
  and _44920_ (_33847_, _33837_, _33107_);
  not _44921_ (_33858_, _33847_);
  nor _44922_ (_33869_, _33858_, _31757_);
  and _44923_ (_33880_, _28069_, _27674_);
  and _44924_ (_33891_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _44925_ (_33902_, _33891_, _33869_);
  and _44926_ (_33913_, _33902_, _31823_);
  or _44927_ (_33924_, _33913_, _33826_);
  and _44928_ (_33935_, _33924_, _31899_);
  or _44929_ (_33945_, _33935_, _33793_);
  or _44930_ (_33956_, _33945_, _33782_);
  and _44931_ (_08889_, _33956_, _42618_);
  and _44932_ (_33977_, _24017_, _18828_);
  not _44933_ (_33988_, _33977_);
  and _44934_ (_33999_, _26778_, _24187_);
  and _44935_ (_34010_, _29308_, _28814_);
  or _44936_ (_34021_, _34010_, _31278_);
  nor _44937_ (_34032_, _34021_, _29319_);
  not _44938_ (_34043_, _34032_);
  nor _44939_ (_34054_, _30020_, _29922_);
  nor _44940_ (_34064_, _34054_, _30031_);
  nor _44941_ (_34075_, _34064_, _29593_);
  not _44942_ (_34086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _44943_ (_34097_, _30554_, _34086_);
  nor _44944_ (_34108_, _34097_, _21635_);
  or _44945_ (_34119_, _34108_, _30543_);
  nor _44946_ (_34130_, _34119_, _30565_);
  nor _44947_ (_34141_, _34130_, _34075_);
  nor _44948_ (_34152_, _30489_, _20220_);
  nor _44949_ (_34163_, _30335_, _29209_);
  nor _44950_ (_34173_, _30227_, _30293_);
  nor _44951_ (_34186_, _34173_, _34163_);
  and _44952_ (_34205_, _34186_, _21635_);
  not _44953_ (_34216_, _34205_);
  nor _44954_ (_34227_, _34186_, _21635_);
  nor _44955_ (_34238_, _34227_, _33313_);
  and _44956_ (_34249_, _34238_, _34216_);
  nor _44957_ (_34260_, _34249_, _34152_);
  and _44958_ (_34271_, _30903_, _28628_);
  and _44959_ (_34282_, _30925_, _21624_);
  nor _44960_ (_34292_, _34282_, _34271_);
  nor _44961_ (_34303_, _32094_, _21254_);
  not _44962_ (_34314_, _34303_);
  and _44963_ (_34325_, _34314_, _34292_);
  nor _44964_ (_34336_, _30740_, _28639_);
  and _44965_ (_34347_, _30761_, _28650_);
  nor _44966_ (_34358_, _34347_, _34336_);
  nor _44967_ (_34369_, _30968_, _21624_);
  nor _44968_ (_34380_, _30838_, _22147_);
  nor _44969_ (_34391_, _34380_, _34369_);
  and _44970_ (_34401_, _34391_, _34358_);
  and _44971_ (_34412_, _34401_, _34325_);
  and _44972_ (_34423_, _34412_, _34260_);
  and _44973_ (_34434_, _34423_, _34141_);
  and _44974_ (_34445_, _34434_, _34043_);
  not _44975_ (_34456_, _34445_);
  nor _44976_ (_34467_, _34456_, _33999_);
  and _44977_ (_34478_, _34467_, _33988_);
  not _44978_ (_34489_, _34478_);
  or _44979_ (_34500_, _34489_, _28409_);
  not _44980_ (_34510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _44981_ (_34521_, _28409_, _34510_);
  and _44982_ (_34532_, _34521_, _31212_);
  and _44983_ (_34543_, _34532_, _34500_);
  nor _44984_ (_34554_, _31211_, _34510_);
  and _44985_ (_34565_, _33804_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _44986_ (_34576_, _31845_, _28069_);
  not _44987_ (_34587_, _34576_);
  nor _44988_ (_34598_, _34587_, _31757_);
  nor _44989_ (_34609_, _33880_, _33837_);
  nor _44990_ (_34620_, _34609_, _34510_);
  or _44991_ (_34630_, _34620_, _34598_);
  and _44992_ (_34641_, _34630_, _31823_);
  or _44993_ (_34652_, _34641_, _34565_);
  and _44994_ (_34663_, _34652_, _31899_);
  or _44995_ (_34674_, _34663_, _34554_);
  or _44996_ (_34685_, _34674_, _34543_);
  and _44997_ (_08900_, _34685_, _42618_);
  and _44998_ (_34706_, _26843_, _24187_);
  not _44999_ (_34717_, _34706_);
  and _45000_ (_34727_, _24048_, _18828_);
  nor _45001_ (_34738_, _30096_, _28617_);
  and _45002_ (_34749_, _30096_, _28617_);
  nor _45003_ (_34760_, _34749_, _34738_);
  and _45004_ (_34771_, _34760_, _29582_);
  not _45005_ (_34782_, _34771_);
  nor _45006_ (_34793_, _29352_, _28617_);
  nor _45007_ (_34804_, _34793_, _29363_);
  and _45008_ (_34815_, _34804_, _28474_);
  and _45009_ (_34826_, _29209_, _21265_);
  nor _45010_ (_34837_, _29209_, _19387_);
  or _45011_ (_34847_, _34837_, _34826_);
  and _45012_ (_34858_, _34847_, _30478_);
  and _45013_ (_34869_, _30238_, _29209_);
  and _45014_ (_34880_, _30336_, _30293_);
  nor _45015_ (_34891_, _34880_, _34869_);
  nor _45016_ (_34902_, _34891_, _21254_);
  not _45017_ (_34913_, _34902_);
  and _45018_ (_34924_, _34891_, _21254_);
  nor _45019_ (_34935_, _34924_, _33313_);
  and _45020_ (_34946_, _34935_, _34913_);
  nor _45021_ (_34956_, _34946_, _34858_);
  nor _45022_ (_34967_, _30576_, _21265_);
  not _45023_ (_34978_, _34967_);
  nor _45024_ (_34989_, _30587_, _30543_);
  and _45025_ (_35000_, _34989_, _34978_);
  not _45026_ (_35011_, _35000_);
  and _45027_ (_35022_, _30761_, _28617_);
  and _45028_ (_35033_, _30903_, _28540_);
  nor _45029_ (_35044_, _30740_, _28606_);
  and _45030_ (_35055_, _30925_, _21254_);
  or _45031_ (_35065_, _35055_, _35044_);
  or _45032_ (_35076_, _35065_, _35033_);
  nor _45033_ (_35087_, _35076_, _35022_);
  nor _45034_ (_35098_, _30968_, _21254_);
  nor _45035_ (_35109_, _32094_, _21080_);
  nor _45036_ (_35120_, _30838_, _21624_);
  or _45037_ (_35131_, _35120_, _35109_);
  nor _45038_ (_35142_, _35131_, _35098_);
  and _45039_ (_35153_, _35142_, _35087_);
  and _45040_ (_35164_, _35153_, _35011_);
  and _45041_ (_35174_, _35164_, _34956_);
  not _45042_ (_35185_, _35174_);
  nor _45043_ (_35196_, _35185_, _34815_);
  and _45044_ (_35207_, _35196_, _34782_);
  not _45045_ (_35218_, _35207_);
  nor _45046_ (_35229_, _35218_, _34727_);
  and _45047_ (_35240_, _35229_, _34717_);
  not _45048_ (_35251_, _35240_);
  or _45049_ (_35262_, _35251_, _28409_);
  not _45050_ (_35273_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _45051_ (_35283_, _28409_, _35273_);
  and _45052_ (_35294_, _35283_, _31212_);
  and _45053_ (_35305_, _35294_, _35262_);
  nor _45054_ (_35316_, _31211_, _35273_);
  not _45055_ (_35327_, _31823_);
  and _45056_ (_35338_, _27806_, _31834_);
  nor _45057_ (_35349_, _27806_, _31834_);
  nor _45058_ (_35360_, _35349_, _35338_);
  or _45059_ (_35371_, _35360_, _35327_);
  and _45060_ (_35382_, _35371_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _45061_ (_35393_, _35338_, _32410_);
  and _45062_ (_35403_, _35349_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _45063_ (_35414_, _35403_, _35393_);
  and _45064_ (_35425_, _35414_, _31823_);
  or _45065_ (_35436_, _35425_, _35382_);
  and _45066_ (_35447_, _35436_, _31899_);
  or _45067_ (_35458_, _35447_, _35316_);
  or _45068_ (_35469_, _35458_, _35305_);
  and _45069_ (_08911_, _35469_, _42618_);
  and _45070_ (_35489_, _26930_, _24187_);
  not _45071_ (_35500_, _35489_);
  and _45072_ (_35511_, _24091_, _18828_);
  nor _45073_ (_35522_, _29384_, _29363_);
  nor _45074_ (_35533_, _35522_, _29395_);
  and _45075_ (_35544_, _35533_, _28474_);
  not _45076_ (_35555_, _35544_);
  nor _45077_ (_35566_, _30107_, _29757_);
  nor _45078_ (_35577_, _35566_, _30118_);
  nor _45079_ (_35588_, _35577_, _29593_);
  nor _45080_ (_35598_, _29209_, _20372_);
  and _45081_ (_35609_, _29209_, _21090_);
  nor _45082_ (_35620_, _35609_, _35598_);
  nor _45083_ (_35631_, _35620_, _30489_);
  nor _45084_ (_35642_, _30249_, _30293_);
  nor _45085_ (_35653_, _30347_, _29209_);
  nor _45086_ (_35664_, _35653_, _35642_);
  and _45087_ (_35675_, _35664_, _21090_);
  nor _45088_ (_35686_, _35664_, _21090_);
  or _45089_ (_35697_, _35686_, _33313_);
  nor _45090_ (_35707_, _35697_, _35675_);
  nor _45091_ (_35718_, _35707_, _35631_);
  not _45092_ (_35729_, _30641_);
  and _45093_ (_35740_, _35729_, _30598_);
  nor _45094_ (_35751_, _30641_, _30587_);
  nor _45095_ (_35762_, _35751_, _21080_);
  nor _45096_ (_35773_, _35762_, _35740_);
  nor _45097_ (_35784_, _35773_, _30543_);
  and _45098_ (_35795_, _30761_, _28562_);
  nor _45099_ (_35806_, _30740_, _28551_);
  not _45100_ (_35817_, _35806_);
  and _45101_ (_35827_, _30903_, _28539_);
  and _45102_ (_35838_, _30925_, _21080_);
  nor _45103_ (_35849_, _35838_, _35827_);
  nand _45104_ (_35860_, _35849_, _35817_);
  nor _45105_ (_35871_, _35860_, _35795_);
  nor _45106_ (_35882_, _32094_, _20046_);
  not _45107_ (_35893_, _35882_);
  nor _45108_ (_35904_, _30968_, _21080_);
  nor _45109_ (_35915_, _30838_, _21254_);
  nor _45110_ (_35926_, _35915_, _35904_);
  and _45111_ (_35937_, _35926_, _35893_);
  and _45112_ (_35948_, _35937_, _35871_);
  not _45113_ (_35958_, _35948_);
  nor _45114_ (_35969_, _35958_, _35784_);
  and _45115_ (_35980_, _35969_, _35718_);
  not _45116_ (_35991_, _35980_);
  nor _45117_ (_36002_, _35991_, _35588_);
  and _45118_ (_36013_, _36002_, _35555_);
  not _45119_ (_36024_, _36013_);
  nor _45120_ (_36035_, _36024_, _35511_);
  and _45121_ (_36046_, _36035_, _35500_);
  not _45122_ (_36057_, _36046_);
  or _45123_ (_36068_, _36057_, _28409_);
  not _45124_ (_36078_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _45125_ (_36089_, _28409_, _36078_);
  and _45126_ (_36100_, _36089_, _31212_);
  and _45127_ (_36111_, _36100_, _36068_);
  nor _45128_ (_36122_, _31211_, _36078_);
  and _45129_ (_36133_, _33118_, _31834_);
  and _45130_ (_36144_, _36133_, _31823_);
  nand _45131_ (_36155_, _36144_, _31757_);
  or _45132_ (_36166_, _36144_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _45133_ (_36177_, _36166_, _31899_);
  and _45134_ (_36188_, _36177_, _36155_);
  or _45135_ (_36199_, _36188_, _36122_);
  or _45136_ (_36209_, _36199_, _36111_);
  and _45137_ (_08922_, _36209_, _42618_);
  and _45138_ (_36230_, _26995_, _24187_);
  and _45139_ (_36241_, _24122_, _18828_);
  or _45140_ (_36252_, _29417_, _29395_);
  nor _45141_ (_36263_, _31278_, _29438_);
  and _45142_ (_36274_, _36263_, _36252_);
  nor _45143_ (_36284_, _30118_, _29724_);
  nor _45144_ (_36295_, _36284_, _30129_);
  nor _45145_ (_36306_, _36295_, _29593_);
  nor _45146_ (_36317_, _29209_, _29604_);
  or _45147_ (_36328_, _36317_, _30489_);
  nor _45148_ (_36339_, _36328_, _31364_);
  nor _45149_ (_36350_, _29209_, _21090_);
  nand _45150_ (_36361_, _36350_, _30347_);
  nand _45151_ (_36371_, _30260_, _29209_);
  and _45152_ (_36382_, _36371_, _36361_);
  and _45153_ (_36393_, _36382_, _20046_);
  nor _45154_ (_36404_, _36382_, _20046_);
  or _45155_ (_36415_, _36404_, _33313_);
  nor _45156_ (_36426_, _36415_, _36393_);
  nor _45157_ (_36437_, _36426_, _36339_);
  nor _45158_ (_36448_, _35740_, _20046_);
  and _45159_ (_36458_, _35740_, _20046_);
  or _45160_ (_36469_, _36458_, _36448_);
  and _45161_ (_36480_, _36469_, _30532_);
  and _45162_ (_36491_, _30761_, _28507_);
  nor _45163_ (_36502_, _30740_, _28496_);
  not _45164_ (_36513_, _36502_);
  and _45165_ (_36524_, _30903_, _28485_);
  and _45166_ (_36535_, _30925_, _20046_);
  nor _45167_ (_36545_, _36535_, _36524_);
  nand _45168_ (_36556_, _36545_, _36513_);
  nor _45169_ (_36567_, _36556_, _36491_);
  nor _45170_ (_36578_, _32094_, _20884_);
  nor _45171_ (_36589_, _30968_, _20046_);
  nor _45172_ (_36600_, _30838_, _21080_);
  or _45173_ (_36611_, _36600_, _36589_);
  nor _45174_ (_36621_, _36611_, _36578_);
  nand _45175_ (_36632_, _36621_, _36567_);
  nor _45176_ (_36643_, _36632_, _36480_);
  nand _45177_ (_36654_, _36643_, _36437_);
  or _45178_ (_36665_, _36654_, _36306_);
  or _45179_ (_36676_, _36665_, _36274_);
  or _45180_ (_36687_, _36676_, _36241_);
  or _45181_ (_36698_, _36687_, _36230_);
  or _45182_ (_36708_, _36698_, _28409_);
  not _45183_ (_36719_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _45184_ (_36730_, _28409_, _36719_);
  and _45185_ (_36741_, _36730_, _31212_);
  and _45186_ (_36752_, _36741_, _36708_);
  nor _45187_ (_36763_, _31211_, _36719_);
  nor _45188_ (_36774_, _28069_, _27674_);
  and _45189_ (_36785_, _36774_, _27795_);
  and _45190_ (_36795_, _36785_, _31823_);
  nand _45191_ (_36806_, _36795_, _31757_);
  or _45192_ (_36817_, _36795_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _45193_ (_36828_, _36817_, _31899_);
  and _45194_ (_36839_, _36828_, _36806_);
  or _45195_ (_36850_, _36839_, _36763_);
  or _45196_ (_36861_, _36850_, _36752_);
  and _45197_ (_08933_, _36861_, _42618_);
  and _45198_ (_36882_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45199_ (_36893_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or _45200_ (_36903_, _36893_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _45201_ (_36914_, _36903_);
  not _45202_ (_36925_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _45203_ (_36936_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _45204_ (_36947_, _36936_, _36925_);
  and _45205_ (_36958_, _36893_, _18772_);
  and _45206_ (_36969_, _36958_, _36947_);
  and _45207_ (_36980_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45208_ (_36991_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _45209_ (_37002_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45210_ (_37012_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _45211_ (_37023_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _45212_ (_37034_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45213_ (_37045_, _37034_, _37023_);
  and _45214_ (_37056_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _45215_ (_37067_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45216_ (_37078_, _37067_, _37023_);
  and _45217_ (_37089_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _45218_ (_37100_, _37089_, _37056_);
  not _45219_ (_37111_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45220_ (_37122_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _37111_);
  and _45221_ (_37133_, _37122_, _37023_);
  and _45222_ (_37144_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not _45223_ (_37155_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _45224_ (_37166_, _37155_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45225_ (_37177_, _37166_, _37023_);
  and _45226_ (_37188_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _45227_ (_37199_, _37188_, _37144_);
  nor _45228_ (_37210_, _37034_, _37023_);
  and _45229_ (_37221_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _45230_ (_37232_, _37034_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _45231_ (_37243_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _45232_ (_37253_, _37243_, _37221_);
  and _45233_ (_37264_, _37253_, _37199_);
  and _45234_ (_37275_, _37264_, _37100_);
  nor _45235_ (_37286_, _37275_, _37012_);
  and _45236_ (_37297_, _37286_, _37002_);
  nor _45237_ (_37308_, _37297_, _36991_);
  nor _45238_ (_37319_, _37308_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45239_ (_37330_, _37319_, _36980_);
  and _45240_ (_37341_, _37330_, _36969_);
  not _45241_ (_37352_, _37341_);
  not _45242_ (_37363_, _36947_);
  nor _45243_ (_37373_, _36958_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _45244_ (_37384_, _37373_, _37363_);
  and _45245_ (_37395_, _37384_, _37352_);
  not _45246_ (_37406_, _37395_);
  and _45247_ (_37417_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45248_ (_37428_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45249_ (_37439_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _45250_ (_37450_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _45251_ (_37461_, _37450_, _37439_);
  and _45252_ (_37472_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _45253_ (_37482_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _45254_ (_37493_, _37482_, _37472_);
  and _45255_ (_37504_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _45256_ (_37515_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _45257_ (_37526_, _37515_, _37504_);
  and _45258_ (_37537_, _37526_, _37493_);
  and _45259_ (_37548_, _37537_, _37461_);
  nor _45260_ (_37559_, _37548_, _37012_);
  and _45261_ (_37570_, _37559_, _37002_);
  nor _45262_ (_37581_, _37570_, _37428_);
  nor _45263_ (_37591_, _37581_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45264_ (_37602_, _37591_, _37417_);
  and _45265_ (_37613_, _37602_, _36969_);
  not _45266_ (_37624_, _37613_);
  nor _45267_ (_37635_, _36958_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _45268_ (_37646_, _37635_, _37363_);
  and _45269_ (_37657_, _37646_, _37624_);
  and _45270_ (_37668_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _45271_ (_37679_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45272_ (_37690_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or _45273_ (_37701_, _37012_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45274_ (_37712_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _45275_ (_37723_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _45276_ (_37734_, _37723_, _37712_);
  and _45277_ (_37745_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _45278_ (_37756_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _45279_ (_37765_, _37756_, _37745_);
  and _45280_ (_37776_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _45281_ (_37787_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _45282_ (_37798_, _37787_, _37776_);
  and _45283_ (_37809_, _37798_, _37765_);
  and _45284_ (_37820_, _37809_, _37734_);
  nor _45285_ (_37829_, _37820_, _37701_);
  or _45286_ (_37830_, _37829_, _37690_);
  and _45287_ (_37831_, _37830_, _37679_);
  nor _45288_ (_37832_, _37831_, _37668_);
  and _45289_ (_37833_, _37832_, _36969_);
  not _45290_ (_37834_, _37833_);
  nor _45291_ (_37835_, _36958_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _45292_ (_37836_, _37835_, _37363_);
  and _45293_ (_37837_, _37836_, _37834_);
  not _45294_ (_37838_, _37837_);
  not _45295_ (_37839_, _36969_);
  and _45296_ (_37840_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _45297_ (_37841_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _45298_ (_37842_, _37841_, _37840_);
  and _45299_ (_37843_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _45300_ (_37844_, _37843_, _37012_);
  and _45301_ (_37845_, _37844_, _37842_);
  and _45302_ (_37846_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not _45303_ (_37847_, _37846_);
  and _45304_ (_37848_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _45305_ (_37849_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _45306_ (_37850_, _37849_, _37848_);
  and _45307_ (_37851_, _37850_, _37847_);
  and _45308_ (_37852_, _37851_, _37845_);
  and _45309_ (_37853_, _37852_, _37002_);
  nor _45310_ (_37854_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _37002_);
  or _45311_ (_37855_, _37854_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45312_ (_37856_, _37855_, _37853_);
  and _45313_ (_37857_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _45314_ (_37858_, _37857_, _37856_);
  nor _45315_ (_37859_, _37858_, _37839_);
  not _45316_ (_37860_, _37859_);
  nor _45317_ (_37861_, _36958_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _45318_ (_37862_, _37861_, _37363_);
  and _45319_ (_37863_, _37862_, _37860_);
  and _45320_ (_37864_, _37863_, _37838_);
  and _45321_ (_37865_, _37864_, _37657_);
  and _45322_ (_37866_, _37865_, _37406_);
  and _45323_ (_37867_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _45324_ (_37868_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _45325_ (_37869_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _45326_ (_37870_, _37869_, _37868_);
  or _45327_ (_37871_, _37870_, _37867_);
  and _45328_ (_37872_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _45329_ (_37873_, _37872_, _37012_);
  and _45330_ (_37874_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _45331_ (_37875_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _45332_ (_37876_, _37875_, _37874_);
  nand _45333_ (_37877_, _37876_, _37873_);
  nor _45334_ (_37878_, _37877_, _37871_);
  and _45335_ (_37879_, _37878_, _37002_);
  nor _45336_ (_37880_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _37002_);
  or _45337_ (_37881_, _37880_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45338_ (_37882_, _37881_, _37879_);
  and _45339_ (_37883_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _45340_ (_37884_, _37883_, _37882_);
  nor _45341_ (_37885_, _37884_, _37839_);
  not _45342_ (_37886_, _37885_);
  nor _45343_ (_37887_, _36958_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _45344_ (_37888_, _37887_, _37363_);
  and _45345_ (_37889_, _37888_, _37886_);
  not _45346_ (_37890_, _37889_);
  and _45347_ (_37891_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45348_ (_37892_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45349_ (_37893_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and _45350_ (_37894_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _45351_ (_37895_, _37894_, _37893_);
  and _45352_ (_37896_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _45353_ (_37897_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _45354_ (_37898_, _37897_, _37896_);
  and _45355_ (_37899_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and _45356_ (_37900_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _45357_ (_37901_, _37900_, _37899_);
  and _45358_ (_37902_, _37901_, _37898_);
  and _45359_ (_37903_, _37902_, _37895_);
  nor _45360_ (_37904_, _37903_, _37012_);
  and _45361_ (_37905_, _37904_, _37002_);
  nor _45362_ (_37906_, _37905_, _37892_);
  nor _45363_ (_37907_, _37906_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45364_ (_37908_, _37907_, _37891_);
  and _45365_ (_37909_, _37908_, _36969_);
  not _45366_ (_37910_, _37909_);
  nor _45367_ (_37911_, _36958_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _45368_ (_37912_, _37911_, _37363_);
  and _45369_ (_37913_, _37912_, _37910_);
  and _45370_ (_37914_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and _45371_ (_37915_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _45372_ (_37916_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and _45373_ (_37917_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _45374_ (_37918_, _37917_, _37916_);
  and _45375_ (_37919_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _45376_ (_37920_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _45377_ (_37921_, _37920_, _37919_);
  and _45378_ (_37922_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _45379_ (_37923_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _45380_ (_37924_, _37923_, _37922_);
  and _45381_ (_37925_, _37924_, _37921_);
  and _45382_ (_37926_, _37925_, _37918_);
  nor _45383_ (_37927_, _37926_, _37012_);
  and _45384_ (_37928_, _37927_, _37002_);
  or _45385_ (_37929_, _37928_, _37915_);
  and _45386_ (_37930_, _37929_, _37679_);
  nor _45387_ (_37931_, _37930_, _37914_);
  and _45388_ (_37932_, _37931_, _36969_);
  not _45389_ (_37933_, _37932_);
  nor _45390_ (_37934_, _36958_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _45391_ (_37935_, _37934_, _37363_);
  and _45392_ (_37936_, _37935_, _37933_);
  not _45393_ (_37937_, _37936_);
  and _45394_ (_37938_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45395_ (_37939_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45396_ (_37940_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _45397_ (_37941_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _45398_ (_37942_, _37941_, _37940_);
  and _45399_ (_37943_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _45400_ (_37944_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _45401_ (_37945_, _37944_, _37943_);
  and _45402_ (_37946_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and _45403_ (_37947_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _45404_ (_37948_, _37947_, _37946_);
  and _45405_ (_37949_, _37948_, _37945_);
  and _45406_ (_37950_, _37949_, _37942_);
  nor _45407_ (_37951_, _37701_, _37950_);
  nor _45408_ (_37952_, _37951_, _37939_);
  nor _45409_ (_37953_, _37952_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45410_ (_37954_, _37953_, _37938_);
  and _45411_ (_37955_, _37954_, _36969_);
  not _45412_ (_37956_, _37955_);
  nor _45413_ (_37957_, _36958_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _45414_ (_37958_, _37957_, _37363_);
  and _45415_ (_37959_, _37958_, _37956_);
  nor _45416_ (_37960_, _37959_, _37937_);
  and _45417_ (_37961_, _37960_, _37913_);
  and _45418_ (_37962_, _37961_, _37890_);
  and _45419_ (_37963_, _37962_, _37866_);
  not _45420_ (_37964_, _37963_);
  and _45421_ (_37965_, _37959_, _37913_);
  and _45422_ (_37966_, _37965_, _37937_);
  and _45423_ (_37967_, _37966_, _37889_);
  and _45424_ (_37968_, _37866_, _37967_);
  not _45425_ (_37969_, _37913_);
  and _45426_ (_37970_, _37960_, _37969_);
  and _45427_ (_37971_, _37970_, _37889_);
  and _45428_ (_37972_, _37971_, _37866_);
  nor _45429_ (_37973_, _37972_, _37968_);
  and _45430_ (_37974_, _37973_, _37964_);
  and _45431_ (_37975_, _37970_, _37890_);
  nor _45432_ (_37976_, _37863_, _37657_);
  nor _45433_ (_37977_, _37838_, _37395_);
  and _45434_ (_37978_, _37977_, _37976_);
  and _45435_ (_37979_, _37978_, _37975_);
  and _45436_ (_37980_, _37978_, _37962_);
  nor _45437_ (_37981_, _37980_, _37979_);
  and _45438_ (_37982_, _37981_, _37974_);
  nor _45439_ (_37983_, _37982_, _36914_);
  not _45440_ (_37984_, _37983_);
  and _45441_ (_37985_, _37959_, _37937_);
  nor _45442_ (_37986_, _37837_, _37395_);
  and _45443_ (_37987_, _37976_, _37986_);
  not _45444_ (_37988_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _45445_ (_37989_, _18772_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _45446_ (_37990_, _37989_, _37988_);
  and _45447_ (_37991_, _37990_, _37987_);
  and _45448_ (_37992_, _37991_, _37985_);
  not _45449_ (_37993_, _36893_);
  nor _45450_ (_37994_, _37981_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _45451_ (_37995_, _37994_, _37993_);
  nor _45452_ (_37996_, _37995_, _37992_);
  and _45453_ (_37997_, _37996_, _37984_);
  nor _45454_ (_37998_, _37997_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45455_ (_37999_, _37998_, _36882_);
  and _45456_ (_38000_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _45457_ (_38001_, _37959_, _37969_);
  and _45458_ (_38002_, _38001_, _37936_);
  and _45459_ (_38003_, _38002_, _37890_);
  not _45460_ (_38004_, _37657_);
  and _45461_ (_38005_, _37864_, _37406_);
  and _45462_ (_38006_, _38005_, _38004_);
  and _45463_ (_38007_, _38006_, _38003_);
  and _45464_ (_38008_, _37961_, _37889_);
  and _45465_ (_38009_, _38008_, _38005_);
  and _45466_ (_38010_, _38009_, _38004_);
  nor _45467_ (_38011_, _38010_, _38007_);
  and _45468_ (_38012_, _37987_, _37961_);
  not _45469_ (_38013_, _37863_);
  and _45470_ (_38014_, _38013_, _37657_);
  and _45471_ (_38015_, _38014_, _37977_);
  and _45472_ (_38016_, _38001_, _37937_);
  and _45473_ (_38017_, _38016_, _37890_);
  and _45474_ (_38018_, _38017_, _38015_);
  nor _45475_ (_38019_, _38018_, _38012_);
  and _45476_ (_38020_, _38002_, _37889_);
  and _45477_ (_38021_, _38020_, _38015_);
  nor _45478_ (_38022_, _37959_, _37936_);
  and _45479_ (_38023_, _38022_, _37969_);
  and _45480_ (_38024_, _38023_, _37889_);
  and _45481_ (_38025_, _38024_, _38015_);
  nor _45482_ (_38026_, _38025_, _38021_);
  and _45483_ (_38027_, _37967_, _38006_);
  and _45484_ (_38028_, _38017_, _38005_);
  nor _45485_ (_38029_, _38028_, _38027_);
  and _45486_ (_38030_, _38029_, _38026_);
  and _45487_ (_38031_, _38030_, _38019_);
  and _45488_ (_38032_, _38031_, _38011_);
  and _45489_ (_38033_, _37962_, _38006_);
  and _45490_ (_38034_, _38020_, _38005_);
  and _45491_ (_38035_, _38034_, _38004_);
  nor _45492_ (_38036_, _38035_, _38033_);
  and _45493_ (_38037_, _38022_, _37913_);
  and _45494_ (_38038_, _38037_, _37889_);
  and _45495_ (_38039_, _38038_, _37987_);
  not _45496_ (_38040_, _38039_);
  and _45497_ (_38041_, _38037_, _37890_);
  and _45498_ (_38042_, _38041_, _37987_);
  and _45499_ (_38043_, _38024_, _37987_);
  nor _45500_ (_38044_, _38043_, _38042_);
  and _45501_ (_38045_, _38044_, _38040_);
  and _45502_ (_38046_, _38023_, _37890_);
  and _45503_ (_38047_, _38046_, _38015_);
  and _45504_ (_38048_, _37965_, _37936_);
  and _45505_ (_38049_, _38048_, _37890_);
  and _45506_ (_38050_, _38049_, _38015_);
  and _45507_ (_38051_, _37863_, _37837_);
  and _45508_ (_38052_, _38051_, _37406_);
  and _45509_ (_38053_, _38052_, _37890_);
  and _45510_ (_38054_, _38053_, _37961_);
  or _45511_ (_38055_, _38054_, _38050_);
  nor _45512_ (_38056_, _38055_, _38047_);
  and _45513_ (_38057_, _38056_, _38045_);
  and _45514_ (_38058_, _38057_, _38036_);
  not _45515_ (_38059_, _38015_);
  and _45516_ (_38060_, _38016_, _37889_);
  nor _45517_ (_38061_, _38060_, _38037_);
  nor _45518_ (_38062_, _38061_, _38059_);
  not _45519_ (_38063_, _38062_);
  and _45520_ (_38064_, _37966_, _37890_);
  and _45521_ (_38065_, _38064_, _38015_);
  and _45522_ (_38066_, _38015_, _38003_);
  nor _45523_ (_38067_, _38066_, _38065_);
  and _45524_ (_38068_, _37987_, _38002_);
  and _45525_ (_38069_, _38064_, _38005_);
  nor _45526_ (_38070_, _38069_, _38068_);
  and _45527_ (_38071_, _38070_, _38067_);
  and _45528_ (_38072_, _38071_, _38063_);
  and _45529_ (_38073_, _37975_, _38006_);
  and _45530_ (_38074_, _38060_, _38005_);
  nor _45531_ (_38075_, _38074_, _38073_);
  and _45532_ (_38076_, _38037_, _38006_);
  and _45533_ (_38077_, _37962_, _37395_);
  nor _45534_ (_38078_, _38077_, _38076_);
  and _45535_ (_38079_, _38078_, _38075_);
  and _45536_ (_38080_, _37971_, _38006_);
  and _45537_ (_38081_, _37975_, _38015_);
  nor _45538_ (_38082_, _38081_, _38080_);
  not _45539_ (_38083_, _38082_);
  nor _45540_ (_38084_, _37971_, _38008_);
  nor _45541_ (_38085_, _38084_, _38059_);
  nor _45542_ (_38086_, _38085_, _38083_);
  and _45543_ (_38087_, _38086_, _38079_);
  and _45544_ (_38088_, _38087_, _38072_);
  and _45545_ (_38089_, _38088_, _38058_);
  and _45546_ (_38090_, _38089_, _38032_);
  nor _45547_ (_38091_, _38090_, _36914_);
  and _45548_ (_38092_, \oc8051_top_1.oc8051_decoder1.state [0], _18772_);
  and _45549_ (_38093_, _38092_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _45550_ (_38094_, _38093_, _38076_);
  nor _45551_ (_38095_, _37992_, _38094_);
  not _45552_ (_38096_, _38095_);
  nor _45553_ (_38097_, _38096_, _38091_);
  nor _45554_ (_38098_, _38097_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45555_ (_38099_, _38098_, _38000_);
  and _45556_ (_38100_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45557_ (_38101_, _37395_, _37890_);
  and _45558_ (_38102_, _38101_, _38051_);
  and _45559_ (_38103_, _38102_, _37961_);
  and _45560_ (_38104_, _38052_, _38023_);
  nor _45561_ (_38105_, _38104_, _38103_);
  and _45562_ (_38106_, _37975_, _38052_);
  nor _45563_ (_38107_, _38106_, _38076_);
  and _45564_ (_38108_, _38107_, _38105_);
  and _45565_ (_38109_, _38102_, _38016_);
  and _45566_ (_38110_, _38052_, _38037_);
  or _45567_ (_38111_, _38110_, _38109_);
  and _45568_ (_38112_, _38052_, _38002_);
  and _45569_ (_38113_, _38102_, _37970_);
  nor _45570_ (_38114_, _38113_, _38112_);
  not _45571_ (_38115_, _38114_);
  nor _45572_ (_38116_, _38115_, _38111_);
  and _45573_ (_38117_, _38116_, _38108_);
  and _45574_ (_38118_, _38064_, _38052_);
  not _45575_ (_38119_, _38118_);
  and _45576_ (_38120_, _38020_, _37987_);
  not _45577_ (_38121_, _38053_);
  nor _45578_ (_38122_, _38048_, _38016_);
  nor _45579_ (_38123_, _38122_, _38121_);
  nor _45580_ (_38124_, _38123_, _38120_);
  and _45581_ (_38125_, _38124_, _38119_);
  and _45582_ (_38126_, _38125_, _37974_);
  and _45583_ (_38127_, _38126_, _38117_);
  nor _45584_ (_38128_, _38127_, _36914_);
  and _45585_ (_38129_, _37992_, _37913_);
  or _45586_ (_38130_, _38129_, _38094_);
  nor _45587_ (_38131_, _38130_, _38128_);
  nor _45588_ (_38132_, _38131_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45589_ (_38133_, _38132_, _38100_);
  nor _45590_ (_38134_, _38133_, _38099_);
  and _45591_ (_38135_, _38134_, _37999_);
  and _45592_ (_09484_, _38135_, _42618_);
  and _45593_ (_38136_, _31212_, _27948_);
  and _45594_ (_38137_, _27542_, _27345_);
  not _45595_ (_38138_, _28376_);
  nor _45596_ (_38139_, _38138_, _28244_);
  and _45597_ (_38140_, _38139_, _38137_);
  and _45598_ (_38141_, _38140_, _33118_);
  and _45599_ (_38142_, _38141_, _28069_);
  and _45600_ (_38143_, _38142_, _38136_);
  not _45601_ (_38144_, _38143_);
  and _45602_ (_38145_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _45603_ (_38146_, _24187_, _18828_);
  and _45604_ (_38147_, _28463_, _24165_);
  nor _45605_ (_38148_, _30958_, _38147_);
  and _45606_ (_38149_, _38148_, _38146_);
  nor _45607_ (_38150_, _30827_, _32083_);
  and _45608_ (_38151_, _38150_, _38149_);
  nor _45609_ (_38152_, _38151_, _20046_);
  not _45610_ (_38153_, _38152_);
  and _45611_ (_38154_, _38153_, _36567_);
  and _45612_ (_38155_, _38154_, _36437_);
  nor _45613_ (_38156_, _38155_, _38144_);
  nor _45614_ (_38157_, _38156_, _38145_);
  and _45615_ (_38158_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _45616_ (_38159_, _38151_, _21080_);
  not _45617_ (_38160_, _38159_);
  and _45618_ (_38161_, _38160_, _35871_);
  and _45619_ (_38162_, _38161_, _35718_);
  nor _45620_ (_38163_, _38162_, _38144_);
  nor _45621_ (_38164_, _38163_, _38158_);
  and _45622_ (_38165_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _45623_ (_38166_, _38151_, _21254_);
  not _45624_ (_38167_, _38166_);
  and _45625_ (_38168_, _38167_, _35087_);
  and _45626_ (_38169_, _38168_, _34956_);
  nor _45627_ (_38170_, _38169_, _38144_);
  nor _45628_ (_38171_, _38170_, _38165_);
  and _45629_ (_38172_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _45630_ (_38173_, _38151_, _21624_);
  not _45631_ (_38174_, _38173_);
  and _45632_ (_38175_, _38174_, _34292_);
  and _45633_ (_38176_, _38175_, _34358_);
  and _45634_ (_38177_, _38176_, _34260_);
  nor _45635_ (_38178_, _38177_, _38144_);
  nor _45636_ (_38179_, _38178_, _38172_);
  and _45637_ (_38180_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _45638_ (_38181_, _38151_, _22147_);
  not _45639_ (_38182_, _38181_);
  and _45640_ (_38183_, _38182_, _33477_);
  and _45641_ (_38184_, _38183_, _33357_);
  nor _45642_ (_38185_, _38184_, _38144_);
  nor _45643_ (_38186_, _38185_, _38180_);
  and _45644_ (_38187_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _45645_ (_38188_, _38151_, _21972_);
  not _45646_ (_38189_, _38188_);
  and _45647_ (_38190_, _38189_, _32736_);
  and _45648_ (_38191_, _38190_, _32922_);
  nor _45649_ (_38192_, _38191_, _38144_);
  nor _45650_ (_38193_, _38192_, _38187_);
  and _45651_ (_38194_, _38136_, _28069_);
  and _45652_ (_38195_, _38194_, _38141_);
  nor _45653_ (_38196_, _38195_, _27740_);
  nor _45654_ (_38197_, _31648_, _30816_);
  nor _45655_ (_38198_, _38149_, _22517_);
  nor _45656_ (_38199_, _38198_, _32780_);
  and _45657_ (_38200_, _38199_, _38197_);
  and _45658_ (_38201_, _38200_, _32214_);
  and _45659_ (_38202_, _38201_, _32040_);
  and _45660_ (_38203_, _38202_, _32073_);
  not _45661_ (_38204_, _38203_);
  and _45662_ (_38205_, _38204_, _38143_);
  nor _45663_ (_38206_, _38205_, _38196_);
  and _45664_ (_38207_, _38206_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _45665_ (_38208_, _38207_, _38193_);
  and _45666_ (_38209_, _38208_, _38186_);
  and _45667_ (_38210_, _38209_, _38179_);
  and _45668_ (_38211_, _38210_, _38171_);
  and _45669_ (_38212_, _38211_, _38164_);
  and _45670_ (_38213_, _38212_, _38157_);
  nor _45671_ (_38214_, _38195_, _28102_);
  nand _45672_ (_38215_, _38214_, _38213_);
  or _45673_ (_38216_, _38214_, _38213_);
  and _45674_ (_38217_, _38216_, _27125_);
  and _45675_ (_38218_, _38217_, _38215_);
  or _45676_ (_38219_, _38195_, _28156_);
  or _45677_ (_38220_, _38219_, _38218_);
  nor _45678_ (_38221_, _38151_, _20884_);
  not _45679_ (_38222_, _38221_);
  and _45680_ (_38223_, _38222_, _30947_);
  and _45681_ (_38224_, _38223_, _30783_);
  and _45682_ (_38225_, _38224_, _30522_);
  nand _45683_ (_38226_, _38225_, _38195_);
  and _45684_ (_38227_, _38226_, _38220_);
  and _45685_ (_09504_, _38227_, _42618_);
  not _45686_ (_38228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _45687_ (_38229_, _38206_, _38228_);
  nor _45688_ (_38230_, _38206_, _38228_);
  nor _45689_ (_38231_, _38230_, _38229_);
  and _45690_ (_38232_, _38231_, _27125_);
  nor _45691_ (_38233_, _38232_, _27751_);
  nor _45692_ (_38234_, _38233_, _38143_);
  nor _45693_ (_38235_, _38234_, _38205_);
  nand _45694_ (_10660_, _38235_, _42618_);
  nor _45695_ (_38236_, _38207_, _38193_);
  nor _45696_ (_38237_, _38236_, _38208_);
  nor _45697_ (_38238_, _38237_, _27114_);
  nor _45698_ (_38239_, _38238_, _27586_);
  nor _45699_ (_38240_, _38239_, _38143_);
  nor _45700_ (_38241_, _38240_, _38192_);
  nand _45701_ (_10671_, _38241_, _42618_);
  nor _45702_ (_38242_, _38208_, _38186_);
  nor _45703_ (_38243_, _38242_, _38209_);
  nor _45704_ (_38244_, _38243_, _27114_);
  nor _45705_ (_38245_, _38244_, _27981_);
  nor _45706_ (_38246_, _38245_, _38143_);
  nor _45707_ (_38247_, _38246_, _38185_);
  nand _45708_ (_10682_, _38247_, _42618_);
  nor _45709_ (_38248_, _38209_, _38179_);
  nor _45710_ (_38249_, _38248_, _38210_);
  nor _45711_ (_38250_, _38249_, _27114_);
  nor _45712_ (_38251_, _38250_, _27849_);
  nor _45713_ (_38252_, _38251_, _38143_);
  nor _45714_ (_38253_, _38252_, _38178_);
  nor _45715_ (_10693_, _38253_, rst);
  nor _45716_ (_38254_, _38210_, _38171_);
  nor _45717_ (_38255_, _38254_, _38211_);
  nor _45718_ (_38256_, _38255_, _27114_);
  nor _45719_ (_38257_, _38256_, _27444_);
  nor _45720_ (_38258_, _38257_, _38143_);
  nor _45721_ (_38259_, _38258_, _38170_);
  nor _45722_ (_10704_, _38259_, rst);
  nor _45723_ (_38260_, _38211_, _38164_);
  nor _45724_ (_38261_, _38260_, _38212_);
  nor _45725_ (_38262_, _38261_, _27114_);
  nor _45726_ (_38263_, _38262_, _27158_);
  nor _45727_ (_38264_, _38263_, _38143_);
  nor _45728_ (_38265_, _38264_, _38163_);
  nor _45729_ (_10715_, _38265_, rst);
  nor _45730_ (_38266_, _38212_, _38157_);
  nor _45731_ (_38267_, _38266_, _38213_);
  nor _45732_ (_38268_, _38267_, _27114_);
  nor _45733_ (_38269_, _38268_, _28288_);
  nor _45734_ (_38270_, _38269_, _38143_);
  nor _45735_ (_38271_, _38270_, _38156_);
  nor _45736_ (_10726_, _38271_, rst);
  and _45737_ (_38272_, _38140_, _34576_);
  nand _45738_ (_38273_, _38272_, _38136_);
  nor _45739_ (_38274_, _38273_, _31136_);
  and _45740_ (_38275_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18772_);
  and _45741_ (_38276_, _38275_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _45742_ (_38277_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _45743_ (_38278_, _38277_, _38276_);
  or _45744_ (_38279_, _38278_, _38274_);
  nor _45745_ (_38280_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not _45746_ (_38281_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _45747_ (_38282_, _38281_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _45748_ (_38283_, _38282_, _38280_);
  nor _45749_ (_38284_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _45750_ (_38285_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _45751_ (_38286_, _38285_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _45752_ (_38287_, _38286_, _38284_);
  not _45753_ (_38288_, _38287_);
  nor _45754_ (_38289_, _38288_, _31299_);
  nor _45755_ (_38290_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not _45756_ (_38291_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _45757_ (_38292_, _38291_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _45758_ (_38293_, _38292_, _38290_);
  and _45759_ (_38294_, _38293_, _38289_);
  nor _45760_ (_38295_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not _45761_ (_38296_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _45762_ (_38297_, _38296_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _45763_ (_38298_, _38297_, _38295_);
  and _45764_ (_38299_, _38298_, _38294_);
  and _45765_ (_38300_, _38299_, _38283_);
  nor _45766_ (_38301_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not _45767_ (_38302_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _45768_ (_38303_, _38302_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _45769_ (_38304_, _38303_, _38301_);
  and _45770_ (_38305_, _38304_, _38300_);
  nor _45771_ (_38306_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _45772_ (_38307_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _45773_ (_38308_, _38307_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _45774_ (_38309_, _38308_, _38306_);
  and _45775_ (_38310_, _38309_, _38305_);
  nor _45776_ (_38311_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _45777_ (_38312_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _45778_ (_38313_, _38312_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _45779_ (_38314_, _38313_, _38311_);
  and _45780_ (_38315_, _38314_, _38310_);
  nor _45781_ (_38316_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _45782_ (_38317_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _45783_ (_38318_, _38317_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _45784_ (_38319_, _38318_, _38316_);
  nand _45785_ (_38320_, _38319_, _38315_);
  or _45786_ (_38321_, _38319_, _38315_);
  and _45787_ (_38322_, _38321_, _28474_);
  and _45788_ (_38323_, _38322_, _38320_);
  not _45789_ (_38324_, _38323_);
  and _45790_ (_38325_, _23879_, _18828_);
  and _45791_ (_38326_, _29209_, _20372_);
  not _45792_ (_38327_, _38326_);
  and _45793_ (_38328_, _30271_, _20895_);
  and _45794_ (_38329_, _38328_, _29790_);
  and _45795_ (_38330_, _38329_, _29823_);
  and _45796_ (_38331_, _38330_, _29867_);
  and _45797_ (_38332_, _38331_, _30042_);
  nor _45798_ (_38333_, _38332_, _30293_);
  and _45799_ (_38334_, _29209_, _19387_);
  nor _45800_ (_38335_, _38334_, _38333_);
  and _45801_ (_38336_, _38335_, _38327_);
  and _45802_ (_38337_, _30358_, _20884_);
  and _45803_ (_38338_, _20220_, _19222_);
  and _45804_ (_38339_, _20536_, _19550_);
  and _45805_ (_38340_, _38339_, _38338_);
  and _45806_ (_38341_, _38340_, _38337_);
  and _45807_ (_38342_, _20372_, _19387_);
  and _45808_ (_38343_, _38342_, _38341_);
  nor _45809_ (_38344_, _38343_, _29209_);
  not _45810_ (_38345_, _38344_);
  and _45811_ (_38346_, _38345_, _38336_);
  nor _45812_ (_38347_, _29209_, _19724_);
  and _45813_ (_38348_, _29209_, _19724_);
  nor _45814_ (_38349_, _38348_, _38347_);
  and _45815_ (_38350_, _38349_, _38346_);
  and _45816_ (_38351_, _38350_, _30434_);
  nor _45817_ (_38352_, _38350_, _30434_);
  nor _45818_ (_38353_, _38352_, _38351_);
  and _45819_ (_38354_, _38353_, _30205_);
  and _45820_ (_38355_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and _45821_ (_38356_, _29209_, _30434_);
  nor _45822_ (_38357_, _38356_, _31387_);
  nor _45823_ (_38358_, _38357_, _30489_);
  nor _45824_ (_38359_, _31627_, _21624_);
  nor _45825_ (_38360_, _30968_, _20719_);
  or _45826_ (_38361_, _38360_, _38359_);
  or _45827_ (_38362_, _38361_, _38358_);
  nor _45828_ (_38363_, _38362_, _38355_);
  not _45829_ (_38364_, _38363_);
  nor _45830_ (_38365_, _38364_, _38354_);
  not _45831_ (_38366_, _38365_);
  nor _45832_ (_38367_, _38366_, _38325_);
  and _45833_ (_38368_, _38367_, _38324_);
  nand _45834_ (_38369_, _38368_, _38276_);
  and _45835_ (_38370_, _38369_, _42618_);
  and _45836_ (_12677_, _38370_, _38279_);
  and _45837_ (_38371_, _38140_, _33847_);
  and _45838_ (_38372_, _38371_, _38136_);
  nor _45839_ (_38373_, _38372_, _38276_);
  not _45840_ (_38374_, _38373_);
  nand _45841_ (_38375_, _38374_, _31136_);
  or _45842_ (_38376_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _45843_ (_38377_, _38376_, _42618_);
  and _45844_ (_12698_, _38377_, _38375_);
  nor _45845_ (_38378_, _38273_, _32323_);
  and _45846_ (_38379_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _45847_ (_38380_, _38379_, _38276_);
  or _45848_ (_38381_, _38380_, _38378_);
  and _45849_ (_38382_, _26458_, _24187_);
  not _45850_ (_38383_, _38382_);
  and _45851_ (_38384_, _38288_, _31299_);
  nor _45852_ (_38385_, _38384_, _38289_);
  and _45853_ (_38386_, _38385_, _28474_);
  nor _45854_ (_38387_, _31387_, _30467_);
  not _45855_ (_38388_, _38387_);
  nor _45856_ (_38389_, _38388_, _30380_);
  nor _45857_ (_38390_, _38389_, _29790_);
  and _45858_ (_38391_, _38389_, _29790_);
  or _45859_ (_38392_, _38391_, _33313_);
  nor _45860_ (_38393_, _38392_, _38390_);
  nor _45861_ (_38394_, _30968_, _19550_);
  and _45862_ (_38395_, _23658_, _18828_);
  nor _45863_ (_38396_, _31627_, _21254_);
  nor _45864_ (_38397_, _30489_, _22517_);
  or _45865_ (_38398_, _38397_, _38396_);
  or _45866_ (_38399_, _38398_, _38395_);
  nor _45867_ (_38400_, _38399_, _38394_);
  not _45868_ (_38401_, _38400_);
  nor _45869_ (_38402_, _38401_, _38393_);
  not _45870_ (_38403_, _38402_);
  nor _45871_ (_38404_, _38403_, _38386_);
  and _45872_ (_38405_, _38404_, _38383_);
  nand _45873_ (_38406_, _38405_, _38276_);
  and _45874_ (_38407_, _38406_, _42618_);
  and _45875_ (_13613_, _38407_, _38381_);
  nor _45876_ (_38408_, _38273_, _33020_);
  and _45877_ (_38409_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _45878_ (_38410_, _38409_, _38276_);
  or _45879_ (_38411_, _38410_, _38408_);
  nor _45880_ (_38412_, _38293_, _38289_);
  nor _45881_ (_38413_, _38412_, _38294_);
  and _45882_ (_38414_, _38413_, _28474_);
  not _45883_ (_38415_, _38414_);
  and _45884_ (_38416_, _25472_, _24187_);
  nor _45885_ (_38417_, _38329_, _30293_);
  and _45886_ (_38418_, _38337_, _19550_);
  nor _45887_ (_38419_, _38418_, _29209_);
  or _45888_ (_38420_, _38419_, _38417_);
  nor _45889_ (_38421_, _38420_, _29823_);
  and _45890_ (_38422_, _38420_, _29823_);
  or _45891_ (_38423_, _38422_, _38421_);
  and _45892_ (_38424_, _38423_, _30205_);
  nor _45893_ (_38425_, _30968_, _20536_);
  and _45894_ (_38426_, _23689_, _18828_);
  nor _45895_ (_38427_, _31627_, _21080_);
  nor _45896_ (_38428_, _30489_, _21972_);
  or _45897_ (_38429_, _38428_, _38427_);
  or _45898_ (_38430_, _38429_, _38426_);
  nor _45899_ (_38431_, _38430_, _38425_);
  not _45900_ (_38432_, _38431_);
  nor _45901_ (_38433_, _38432_, _38424_);
  not _45902_ (_38434_, _38433_);
  nor _45903_ (_38435_, _38434_, _38416_);
  and _45904_ (_38436_, _38435_, _38415_);
  nand _45905_ (_38437_, _38436_, _38276_);
  and _45906_ (_38438_, _38437_, _42618_);
  and _45907_ (_13624_, _38438_, _38411_);
  nor _45908_ (_38439_, _38273_, _33717_);
  and _45909_ (_38440_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _45910_ (_38441_, _38440_, _38276_);
  or _45911_ (_38442_, _38441_, _38439_);
  nor _45912_ (_38443_, _38298_, _38294_);
  nor _45913_ (_38444_, _38443_, _38299_);
  and _45914_ (_38445_, _38444_, _28474_);
  not _45915_ (_38446_, _38445_);
  and _45916_ (_38447_, _38418_, _20536_);
  and _45917_ (_38448_, _38447_, _30293_);
  and _45918_ (_38449_, _38330_, _29209_);
  nor _45919_ (_38450_, _38449_, _38448_);
  and _45920_ (_38451_, _38450_, _19222_);
  nor _45921_ (_38452_, _38450_, _19222_);
  nor _45922_ (_38453_, _38452_, _38451_);
  and _45923_ (_38454_, _38453_, _30205_);
  not _45924_ (_38455_, _38454_);
  nor _45925_ (_38456_, _30489_, _22147_);
  and _45926_ (_38457_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _45927_ (_38458_, _38457_, _38456_);
  and _45928_ (_38459_, _23721_, _18828_);
  nor _45929_ (_38460_, _31627_, _20046_);
  nor _45930_ (_38461_, _30968_, _19222_);
  or _45931_ (_38462_, _38461_, _38460_);
  nor _45932_ (_38463_, _38462_, _38459_);
  and _45933_ (_38464_, _38463_, _38458_);
  and _45934_ (_38465_, _38464_, _38455_);
  and _45935_ (_38466_, _38465_, _38446_);
  nand _45936_ (_38467_, _38466_, _38276_);
  and _45937_ (_38468_, _38467_, _42618_);
  and _45938_ (_13635_, _38468_, _38442_);
  nor _45939_ (_38469_, _38273_, _34478_);
  and _45940_ (_38470_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _45941_ (_38471_, _38470_, _38276_);
  or _45942_ (_38472_, _38471_, _38469_);
  nor _45943_ (_38473_, _38299_, _38283_);
  nor _45944_ (_38474_, _38473_, _38300_);
  and _45945_ (_38475_, _38474_, _28474_);
  not _45946_ (_38476_, _38475_);
  and _45947_ (_38477_, _23753_, _18828_);
  not _45948_ (_38478_, _38477_);
  nor _45949_ (_38479_, _38331_, _30042_);
  not _45950_ (_38480_, _38479_);
  and _45951_ (_38481_, _38480_, _38333_);
  and _45952_ (_38482_, _38447_, _19222_);
  nor _45953_ (_38483_, _38482_, _20220_);
  nor _45954_ (_38484_, _38483_, _38341_);
  nor _45955_ (_38485_, _38484_, _29209_);
  nor _45956_ (_38486_, _38485_, _38481_);
  nor _45957_ (_38487_, _38486_, _33313_);
  nor _45958_ (_38488_, _30968_, _20220_);
  nor _45959_ (_38489_, _30489_, _21624_);
  and _45960_ (_38490_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _45961_ (_38491_, _38490_, _38489_);
  or _45962_ (_38492_, _38491_, _31647_);
  nor _45963_ (_38493_, _38492_, _38488_);
  not _45964_ (_38494_, _38493_);
  nor _45965_ (_38495_, _38494_, _38487_);
  and _45966_ (_38496_, _38495_, _38478_);
  and _45967_ (_38497_, _38496_, _38476_);
  nand _45968_ (_38498_, _38497_, _38276_);
  and _45969_ (_38499_, _38498_, _42618_);
  and _45970_ (_13646_, _38499_, _38472_);
  nor _45971_ (_38500_, _38273_, _35240_);
  and _45972_ (_38501_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _45973_ (_38502_, _38501_, _38276_);
  or _45974_ (_38503_, _38502_, _38500_);
  nor _45975_ (_38504_, _38304_, _38300_);
  nor _45976_ (_38505_, _38504_, _38305_);
  and _45977_ (_38506_, _38505_, _28474_);
  not _45978_ (_38507_, _38506_);
  and _45979_ (_38508_, _23784_, _18828_);
  nor _45980_ (_38509_, _38341_, _29209_);
  nor _45981_ (_38510_, _38509_, _38333_);
  nor _45982_ (_38511_, _38510_, _29637_);
  and _45983_ (_38512_, _38510_, _29637_);
  nor _45984_ (_38513_, _38512_, _38511_);
  and _45985_ (_38514_, _38513_, _30205_);
  and _45986_ (_38515_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _45987_ (_38516_, _29209_, _21265_);
  or _45988_ (_38517_, _38516_, _30489_);
  nor _45989_ (_38518_, _38517_, _38334_);
  nor _45990_ (_38519_, _31627_, _22517_);
  nor _45991_ (_38520_, _30968_, _19387_);
  or _45992_ (_38521_, _38520_, _38519_);
  or _45993_ (_38522_, _38521_, _38518_);
  nor _45994_ (_38523_, _38522_, _38515_);
  not _45995_ (_38524_, _38523_);
  nor _45996_ (_38525_, _38524_, _38514_);
  not _45997_ (_38526_, _38525_);
  nor _45998_ (_38527_, _38526_, _38508_);
  and _45999_ (_38528_, _38527_, _38507_);
  nand _46000_ (_38529_, _38528_, _38276_);
  and _46001_ (_38530_, _38529_, _42618_);
  and _46002_ (_13657_, _38530_, _38503_);
  nor _46003_ (_38531_, _38273_, _36046_);
  and _46004_ (_38532_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _46005_ (_38533_, _38532_, _38276_);
  or _46006_ (_38534_, _38533_, _38531_);
  nor _46007_ (_38535_, _38309_, _38305_);
  not _46008_ (_38536_, _38535_);
  nor _46009_ (_38537_, _38310_, _31278_);
  and _46010_ (_38538_, _38537_, _38536_);
  not _46011_ (_38539_, _38538_);
  and _46012_ (_38540_, _23816_, _18828_);
  and _46013_ (_38541_, _38341_, _19387_);
  nor _46014_ (_38542_, _38541_, _29209_);
  not _46015_ (_38543_, _38542_);
  and _46016_ (_38544_, _38543_, _38335_);
  and _46017_ (_38545_, _38544_, _20372_);
  nor _46018_ (_38546_, _38544_, _20372_);
  nor _46019_ (_38547_, _38546_, _38545_);
  nor _46020_ (_38548_, _38547_, _33313_);
  and _46021_ (_38549_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _46022_ (_38550_, _36350_, _30489_);
  and _46023_ (_38551_, _38550_, _38327_);
  nor _46024_ (_38552_, _31627_, _21972_);
  nor _46025_ (_38553_, _30968_, _20372_);
  or _46026_ (_38554_, _38553_, _38552_);
  or _46027_ (_38555_, _38554_, _38551_);
  nor _46028_ (_38556_, _38555_, _38549_);
  not _46029_ (_38557_, _38556_);
  nor _46030_ (_38558_, _38557_, _38548_);
  not _46031_ (_38559_, _38558_);
  nor _46032_ (_38560_, _38559_, _38540_);
  and _46033_ (_38561_, _38560_, _38539_);
  nand _46034_ (_38562_, _38561_, _38276_);
  and _46035_ (_38563_, _38562_, _42618_);
  and _46036_ (_13668_, _38563_, _38534_);
  or _46037_ (_38564_, _38273_, _36698_);
  not _46038_ (_38565_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand _46039_ (_38566_, _38273_, _38565_);
  and _46040_ (_38567_, _38566_, _38564_);
  or _46041_ (_38568_, _38567_, _38276_);
  not _46042_ (_38569_, _38276_);
  nor _46043_ (_38570_, _38314_, _38310_);
  nor _46044_ (_38571_, _38570_, _38315_);
  and _46045_ (_38572_, _38571_, _28474_);
  and _46046_ (_38573_, _23848_, _18828_);
  and _46047_ (_38574_, _38346_, _19724_);
  nor _46048_ (_38575_, _38346_, _19724_);
  or _46049_ (_38576_, _38575_, _38574_);
  and _46050_ (_38577_, _38576_, _30205_);
  or _46051_ (_38578_, _29209_, _20057_);
  nor _46052_ (_38579_, _38348_, _30489_);
  and _46053_ (_38580_, _38579_, _38578_);
  nor _46054_ (_38581_, _31627_, _22147_);
  nor _46055_ (_38582_, _30968_, _19724_);
  and _46056_ (_38583_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or _46057_ (_38584_, _38583_, _38582_);
  or _46058_ (_38585_, _38584_, _38581_);
  or _46059_ (_38586_, _38585_, _38580_);
  or _46060_ (_38587_, _38586_, _38577_);
  or _46061_ (_38588_, _38587_, _38573_);
  or _46062_ (_38589_, _38588_, _38572_);
  or _46063_ (_38590_, _38589_, _38569_);
  and _46064_ (_38591_, _38590_, _42618_);
  and _46065_ (_13679_, _38591_, _38568_);
  nand _46066_ (_38592_, _38374_, _32323_);
  or _46067_ (_38593_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _46068_ (_38594_, _38593_, _42618_);
  and _46069_ (_13690_, _38594_, _38592_);
  nand _46070_ (_38595_, _38374_, _33020_);
  or _46071_ (_38596_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _46072_ (_38597_, _38596_, _42618_);
  and _46073_ (_13701_, _38597_, _38595_);
  nand _46074_ (_38598_, _38374_, _33717_);
  or _46075_ (_38599_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _46076_ (_38600_, _38599_, _42618_);
  and _46077_ (_13711_, _38600_, _38598_);
  nand _46078_ (_38601_, _38374_, _34478_);
  or _46079_ (_38602_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _46080_ (_38603_, _38602_, _42618_);
  and _46081_ (_13722_, _38603_, _38601_);
  nand _46082_ (_38604_, _38374_, _35240_);
  or _46083_ (_38605_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _46084_ (_38606_, _38605_, _42618_);
  and _46085_ (_13733_, _38606_, _38604_);
  nand _46086_ (_38607_, _38374_, _36046_);
  or _46087_ (_38608_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _46088_ (_38609_, _38608_, _42618_);
  and _46089_ (_13744_, _38609_, _38607_);
  or _46090_ (_38610_, _38373_, _36698_);
  or _46091_ (_38611_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _46092_ (_38612_, _38611_, _42618_);
  and _46093_ (_13755_, _38612_, _38610_);
  not _46094_ (_38613_, _27345_);
  nor _46095_ (_38614_, _28376_, _38613_);
  and _46096_ (_38615_, _38614_, _31899_);
  and _46097_ (_38616_, _38615_, _31812_);
  not _46098_ (_38617_, _31855_);
  nor _46099_ (_38618_, _38617_, _31757_);
  not _46100_ (_38619_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _46101_ (_38620_, _31855_, _38619_);
  or _46102_ (_38621_, _38620_, _38618_);
  and _46103_ (_38622_, _38621_, _38616_);
  nor _46104_ (_38623_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _46105_ (_38624_, _38623_);
  nand _46106_ (_38625_, _38624_, _31757_);
  and _46107_ (_38626_, _38623_, _38619_);
  nor _46108_ (_38627_, _38626_, _38616_);
  and _46109_ (_38628_, _38627_, _38625_);
  nor _46110_ (_38629_, _27542_, _38613_);
  and _46111_ (_38630_, _31212_, _28398_);
  and _46112_ (_38631_, _38630_, _38629_);
  or _46113_ (_38632_, _38631_, _38628_);
  or _46114_ (_38633_, _38632_, _38622_);
  nand _46115_ (_38634_, _38631_, _38225_);
  and _46116_ (_38635_, _38634_, _42618_);
  and _46117_ (_15158_, _38635_, _38633_);
  and _46118_ (_38636_, _38616_, _33129_);
  nand _46119_ (_38637_, _38636_, _31757_);
  not _46120_ (_38638_, _38631_);
  or _46121_ (_38639_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _46122_ (_38640_, _38639_, _38638_);
  and _46123_ (_38641_, _38640_, _38637_);
  nor _46124_ (_38642_, _38638_, _38191_);
  or _46125_ (_38645_, _38642_, _38641_);
  and _46126_ (_17339_, _38645_, _42618_);
  or _46127_ (_38647_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _46128_ (_38648_, _23943_, _23911_);
  or _46129_ (_38649_, _38648_, _23974_);
  or _46130_ (_38650_, _38649_, _24017_);
  or _46131_ (_38651_, _38650_, _24048_);
  or _46132_ (_38652_, _38651_, _24091_);
  or _46133_ (_38653_, _38652_, _24122_);
  or _46134_ (_38654_, _38653_, _23594_);
  and _46135_ (_38655_, _38654_, _18828_);
  or _46136_ (_38657_, _31342_, _30140_);
  not _46137_ (_38666_, _31321_);
  nand _46138_ (_38672_, _38666_, _30140_);
  and _46139_ (_38678_, _38672_, _29582_);
  and _46140_ (_38681_, _38678_, _38657_);
  not _46141_ (_38682_, _29461_);
  nand _46142_ (_38683_, _29450_, _38682_);
  or _46143_ (_38684_, _29472_, _29450_);
  and _46144_ (_38685_, _28474_, _38684_);
  and _46145_ (_38686_, _38685_, _38683_);
  and _46146_ (_38687_, _38342_, _25373_);
  and _46147_ (_38688_, _38340_, _24187_);
  nand _46148_ (_38689_, _38688_, _38687_);
  nand _46149_ (_38690_, _38689_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _46150_ (_38691_, _38690_, _38686_);
  or _46151_ (_38692_, _38691_, _38681_);
  or _46152_ (_38693_, _38692_, _38655_);
  and _46153_ (_38694_, _38693_, _38647_);
  or _46154_ (_38695_, _38694_, _38616_);
  not _46155_ (_38696_, _38616_);
  and _46156_ (_38697_, _33858_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _46157_ (_38698_, _38697_, _33869_);
  or _46158_ (_38699_, _38698_, _38696_);
  and _46159_ (_38700_, _38699_, _38695_);
  or _46160_ (_38701_, _38700_, _38631_);
  nand _46161_ (_38702_, _38631_, _38184_);
  and _46162_ (_38703_, _38702_, _42618_);
  and _46163_ (_17350_, _38703_, _38701_);
  and _46164_ (_38704_, _38616_, _34576_);
  nand _46165_ (_38707_, _38704_, _31757_);
  or _46166_ (_38708_, _38704_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _46167_ (_38709_, _38708_, _38638_);
  and _46168_ (_38710_, _38709_, _38707_);
  nor _46169_ (_38711_, _38638_, _38177_);
  or _46170_ (_38712_, _38711_, _38710_);
  and _46171_ (_17361_, _38712_, _42618_);
  or _46172_ (_38713_, _38696_, _35360_);
  nor _46173_ (_38714_, _38638_, _38169_);
  and _46174_ (_38715_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _46175_ (_38716_, _38715_, _38714_);
  nor _46176_ (_38743_, _38716_, rst);
  and _46177_ (_38717_, _38743_, _38713_);
  and _46178_ (_38718_, _35349_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _46179_ (_38719_, _38718_, _35393_);
  and _46180_ (_38720_, _38616_, _42618_);
  and _46181_ (_38721_, _38720_, _38719_);
  or _46182_ (_17372_, _38721_, _38717_);
  and _46183_ (_38722_, _38616_, _36133_);
  nand _46184_ (_38723_, _38722_, _31757_);
  or _46185_ (_38724_, _38722_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _46186_ (_38725_, _38724_, _38638_);
  and _46187_ (_38726_, _38725_, _38723_);
  nor _46188_ (_38727_, _38638_, _38162_);
  or _46189_ (_38728_, _38727_, _38726_);
  and _46190_ (_17383_, _38728_, _42618_);
  and _46191_ (_38729_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _46192_ (_38730_, _38729_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _46193_ (_38731_, _30096_, _29582_);
  and _46194_ (_38732_, _28474_, _29352_);
  nand _46195_ (_38733_, _30958_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _46196_ (_38734_, _38733_, _38729_);
  or _46197_ (_38735_, _38734_, _38732_);
  or _46198_ (_38736_, _38735_, _38731_);
  and _46199_ (_38737_, _38736_, _38730_);
  or _46200_ (_38738_, _38737_, _38616_);
  not _46201_ (_38739_, _36785_);
  nor _46202_ (_38740_, _38739_, _31757_);
  or _46203_ (_38742_, _36785_, _34086_);
  nand _46204_ (_38746_, _38742_, _38616_);
  or _46205_ (_38752_, _38746_, _38740_);
  and _46206_ (_38757_, _38752_, _38738_);
  or _46207_ (_38764_, _38757_, _38631_);
  nand _46208_ (_38772_, _38631_, _38155_);
  and _46209_ (_38780_, _38772_, _42618_);
  and _46210_ (_17394_, _38780_, _38764_);
  not _46211_ (_38781_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46212_ (_38782_, _38275_, _38781_);
  and _46213_ (_38783_, _38782_, _38368_);
  nor _46214_ (_38784_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _46215_ (_38785_, _38784_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46216_ (_38786_, _27542_, _38613_);
  and _46217_ (_38787_, _38786_, _28387_);
  and _46218_ (_38788_, _38787_, _28091_);
  and _46219_ (_38789_, _38788_, _31212_);
  nor _46220_ (_38790_, _38789_, _38785_);
  nor _46221_ (_38791_, _38790_, _31136_);
  and _46222_ (_38792_, _27948_, _27542_);
  and _46223_ (_38793_, _38792_, _31768_);
  not _46224_ (_38794_, _31899_);
  nor _46225_ (_38795_, _38794_, _28244_);
  and _46226_ (_38796_, _38795_, _38793_);
  and _46227_ (_38797_, _38796_, _31855_);
  and _46228_ (_38798_, _38797_, _31757_);
  nor _46229_ (_38799_, _38797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _46230_ (_38800_, _38799_);
  not _46231_ (_38801_, _38782_);
  and _46232_ (_38802_, _38790_, _38801_);
  and _46233_ (_38803_, _38802_, _38800_);
  not _46234_ (_38804_, _38803_);
  nor _46235_ (_38805_, _38804_, _38798_);
  nor _46236_ (_38806_, _38805_, _38782_);
  not _46237_ (_38807_, _38806_);
  nor _46238_ (_38808_, _38807_, _38791_);
  nor _46239_ (_38809_, _38808_, _38783_);
  and _46240_ (_17963_, _38809_, _42618_);
  nor _46241_ (_38810_, _38801_, _38405_);
  not _46242_ (_38811_, _38790_);
  and _46243_ (_38812_, _38811_, _32323_);
  and _46244_ (_38813_, _27806_, _28069_);
  and _46245_ (_38814_, _32410_, _38813_);
  not _46246_ (_38815_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _46247_ (_38821_, _38813_, _38815_);
  nor _46248_ (_38832_, _38821_, _38814_);
  and _46249_ (_38833_, _38796_, _38801_);
  not _46250_ (_38834_, _38833_);
  nor _46251_ (_38835_, _38834_, _38832_);
  nor _46252_ (_38846_, _38796_, _38815_);
  nor _46253_ (_38852_, _38846_, _38811_);
  nor _46254_ (_38853_, _38852_, _38782_);
  or _46255_ (_38854_, _38853_, _38835_);
  not _46256_ (_38855_, _38854_);
  nor _46257_ (_38856_, _38855_, _38812_);
  nor _46258_ (_38857_, _38856_, _38810_);
  nor _46259_ (_19757_, _38857_, rst);
  nor _46260_ (_38858_, _38801_, _38436_);
  and _46261_ (_38859_, _38811_, _33020_);
  not _46262_ (_38860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _46263_ (_38861_, _38796_, _38860_);
  nor _46264_ (_38862_, _38861_, _38811_);
  not _46265_ (_38863_, _33129_);
  nor _46266_ (_38864_, _38863_, _31757_);
  nor _46267_ (_38865_, _33129_, _38860_);
  nor _46268_ (_38866_, _38865_, _38864_);
  nand _46269_ (_38867_, _38802_, _38796_);
  or _46270_ (_38868_, _38867_, _38866_);
  and _46271_ (_38869_, _38868_, _38862_);
  or _46272_ (_38870_, _38869_, _38782_);
  nor _46273_ (_38871_, _38870_, _38859_);
  nor _46274_ (_38872_, _38871_, _38858_);
  nor _46275_ (_19769_, _38872_, rst);
  nor _46276_ (_38873_, _38801_, _38466_);
  and _46277_ (_38874_, _38811_, _33717_);
  not _46278_ (_38875_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _46279_ (_38876_, _38796_, _38875_);
  nor _46280_ (_38877_, _38876_, _38811_);
  not _46281_ (_38878_, _38877_);
  not _46282_ (_38879_, _38796_);
  nor _46283_ (_38880_, _33847_, _38875_);
  nor _46284_ (_38881_, _38880_, _33869_);
  nor _46285_ (_38882_, _38881_, _38879_);
  nor _46286_ (_38883_, _38882_, _38878_);
  nor _46287_ (_38884_, _38883_, _38782_);
  not _46288_ (_38885_, _38884_);
  nor _46289_ (_38886_, _38885_, _38874_);
  nor _46290_ (_38887_, _38886_, _38873_);
  nor _46291_ (_19780_, _38887_, rst);
  nor _46292_ (_38888_, _38790_, _34478_);
  and _46293_ (_38889_, _38802_, _38879_);
  and _46294_ (_38890_, _38889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _46295_ (_38891_, _38890_, _38888_);
  and _46296_ (_38892_, _34587_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _46297_ (_38893_, _38892_, _34598_);
  nor _46298_ (_38894_, _38893_, _38834_);
  and _46299_ (_38895_, _38894_, _38790_);
  nor _46300_ (_38896_, _38895_, _38782_);
  and _46301_ (_38897_, _38896_, _38891_);
  and _46302_ (_38898_, _38782_, _38497_);
  or _46303_ (_38899_, _38898_, _38897_);
  nor _46304_ (_19792_, _38899_, rst);
  nor _46305_ (_38900_, _38790_, _35240_);
  and _46306_ (_38901_, _38796_, _35338_);
  and _46307_ (_38902_, _38901_, _31757_);
  nor _46308_ (_38903_, _38901_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not _46309_ (_38904_, _38903_);
  and _46310_ (_38905_, _38904_, _38802_);
  not _46311_ (_38906_, _38905_);
  nor _46312_ (_38907_, _38906_, _38902_);
  or _46313_ (_38908_, _38907_, _38900_);
  and _46314_ (_38909_, _38908_, _38801_);
  nor _46315_ (_38910_, _38801_, _38528_);
  or _46316_ (_38911_, _38910_, _38909_);
  and _46317_ (_19804_, _38911_, _42618_);
  nor _46318_ (_38912_, _38790_, _36046_);
  and _46319_ (_38913_, _38796_, _36133_);
  nor _46320_ (_38914_, _38913_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not _46321_ (_38915_, _38914_);
  not _46322_ (_38916_, _38802_);
  and _46323_ (_38917_, _38913_, _31757_);
  nor _46324_ (_38918_, _38917_, _38916_);
  and _46325_ (_38919_, _38918_, _38915_);
  or _46326_ (_38920_, _38919_, _38912_);
  and _46327_ (_38921_, _38920_, _38801_);
  nor _46328_ (_38922_, _38801_, _38561_);
  or _46329_ (_38923_, _38922_, _38921_);
  and _46330_ (_19816_, _38923_, _42618_);
  or _46331_ (_38924_, _38801_, _38589_);
  and _46332_ (_38925_, _38811_, _36698_);
  and _46333_ (_38926_, _38796_, _36785_);
  or _46334_ (_38927_, _38926_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _46335_ (_38928_, _38926_, _31757_);
  and _46336_ (_38929_, _38928_, _38802_);
  and _46337_ (_38930_, _38929_, _38927_);
  or _46338_ (_38931_, _38930_, _38782_);
  or _46339_ (_38932_, _38931_, _38925_);
  and _46340_ (_38933_, _38932_, _38924_);
  and _46341_ (_19828_, _38933_, _42618_);
  and _46342_ (_38934_, _28376_, _27345_);
  and _46343_ (_38935_, _38792_, _31779_);
  and _46344_ (_38936_, _38935_, _38934_);
  and _46345_ (_38937_, _38936_, _31855_);
  nand _46346_ (_38938_, _38937_, _31757_);
  or _46347_ (_38939_, _38937_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46348_ (_38940_, _38939_, _31899_);
  and _46349_ (_38941_, _38940_, _38938_);
  and _46350_ (_38942_, _38140_, _28091_);
  nand _46351_ (_38943_, _38942_, _38225_);
  or _46352_ (_38944_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46353_ (_38945_, _38944_, _31212_);
  and _46354_ (_38946_, _38945_, _38943_);
  not _46355_ (_38947_, _31211_);
  and _46356_ (_38948_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _46357_ (_38949_, _38948_, rst);
  or _46358_ (_38950_, _38949_, _38946_);
  or _46359_ (_31034_, _38950_, _38941_);
  and _46360_ (_38951_, _38934_, _31812_);
  and _46361_ (_38952_, _38951_, _31855_);
  nand _46362_ (_38953_, _38952_, _31757_);
  or _46363_ (_38954_, _38952_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _46364_ (_38955_, _38954_, _31899_);
  and _46365_ (_38956_, _38955_, _38953_);
  and _46366_ (_38957_, _38629_, _38139_);
  and _46367_ (_38958_, _38957_, _28091_);
  nand _46368_ (_38959_, _38958_, _38225_);
  or _46369_ (_38960_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _46370_ (_38961_, _38960_, _31212_);
  and _46371_ (_38962_, _38961_, _38959_);
  and _46372_ (_38963_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _46373_ (_38964_, _38963_, rst);
  or _46374_ (_38965_, _38964_, _38962_);
  or _46375_ (_31057_, _38965_, _38956_);
  and _46376_ (_38966_, _28376_, _38613_);
  and _46377_ (_38967_, _38966_, _38935_);
  and _46378_ (_38968_, _38967_, _31855_);
  nand _46379_ (_38969_, _38968_, _31757_);
  or _46380_ (_38970_, _38968_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _46381_ (_38971_, _38970_, _31899_);
  and _46382_ (_38972_, _38971_, _38969_);
  and _46383_ (_38973_, _38786_, _38139_);
  and _46384_ (_38974_, _38973_, _28091_);
  not _46385_ (_38975_, _38974_);
  nor _46386_ (_38976_, _38975_, _38225_);
  and _46387_ (_38977_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _46388_ (_38978_, _38977_, _38976_);
  and _46389_ (_38979_, _38978_, _31212_);
  and _46390_ (_38980_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _46391_ (_38981_, _38980_, rst);
  or _46392_ (_38982_, _38981_, _38979_);
  or _46393_ (_31079_, _38982_, _38972_);
  and _46394_ (_38983_, _38966_, _31812_);
  and _46395_ (_38984_, _38983_, _31855_);
  nand _46396_ (_38985_, _38984_, _31757_);
  or _46397_ (_38986_, _38984_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _46398_ (_38987_, _38986_, _31899_);
  and _46399_ (_38988_, _38987_, _38985_);
  and _46400_ (_38989_, _38139_, _27553_);
  and _46401_ (_38990_, _38989_, _28091_);
  not _46402_ (_38991_, _38990_);
  nor _46403_ (_38992_, _38991_, _38225_);
  and _46404_ (_38993_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _46405_ (_38994_, _38993_, _38992_);
  and _46406_ (_38995_, _38994_, _31212_);
  and _46407_ (_38996_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _46408_ (_38997_, _38996_, rst);
  or _46409_ (_38998_, _38997_, _38995_);
  or _46410_ (_31102_, _38998_, _38988_);
  or _46411_ (_38999_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _46412_ (_39000_, _38999_, _31899_);
  and _46413_ (_39001_, _38936_, _38813_);
  nand _46414_ (_39002_, _39001_, _31757_);
  and _46415_ (_39003_, _39002_, _39000_);
  nand _46416_ (_39004_, _38942_, _38203_);
  and _46417_ (_39005_, _39004_, _31212_);
  and _46418_ (_39006_, _39005_, _38999_);
  not _46419_ (_39007_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _46420_ (_39008_, _31211_, _39007_);
  or _46421_ (_39009_, _39008_, rst);
  or _46422_ (_39010_, _39009_, _39006_);
  or _46423_ (_40308_, _39010_, _39003_);
  and _46424_ (_39011_, _33118_, _28080_);
  and _46425_ (_39012_, _39011_, _38140_);
  nand _46426_ (_39013_, _39012_, _31757_);
  or _46427_ (_39014_, _39012_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46428_ (_39015_, _39014_, _31899_);
  and _46429_ (_39016_, _39015_, _39013_);
  nand _46430_ (_39017_, _38942_, _38191_);
  or _46431_ (_39018_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46432_ (_39019_, _39018_, _31212_);
  and _46433_ (_39020_, _39019_, _39017_);
  and _46434_ (_39021_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _46435_ (_39022_, _39021_, rst);
  or _46436_ (_39023_, _39022_, _39020_);
  or _46437_ (_40310_, _39023_, _39016_);
  not _46438_ (_39024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  not _46439_ (_39025_, _34609_);
  and _46440_ (_39026_, _38936_, _39025_);
  nor _46441_ (_39035_, _39026_, _39024_);
  and _46442_ (_39046_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _46443_ (_39057_, _39046_, _33869_);
  and _46444_ (_39066_, _39057_, _38936_);
  or _46445_ (_39072_, _39066_, _39035_);
  and _46446_ (_39083_, _39072_, _31899_);
  nand _46447_ (_39094_, _38942_, _38184_);
  or _46448_ (_39105_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _46449_ (_39116_, _39105_, _31212_);
  and _46450_ (_39127_, _39116_, _39094_);
  nor _46451_ (_39138_, _31211_, _39024_);
  or _46452_ (_39149_, _39138_, rst);
  or _46453_ (_39160_, _39149_, _39127_);
  or _46454_ (_40312_, _39160_, _39083_);
  and _46455_ (_39181_, _38936_, _34576_);
  nand _46456_ (_39192_, _39181_, _31757_);
  or _46457_ (_39203_, _39181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _46458_ (_39214_, _39203_, _31899_);
  and _46459_ (_39225_, _39214_, _39192_);
  nand _46460_ (_39236_, _38942_, _38177_);
  or _46461_ (_39240_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _46462_ (_39241_, _39240_, _31212_);
  and _46463_ (_39242_, _39241_, _39236_);
  and _46464_ (_39243_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _46465_ (_39244_, _39243_, rst);
  or _46466_ (_39245_, _39244_, _39242_);
  or _46467_ (_40314_, _39245_, _39225_);
  not _46468_ (_39246_, _38936_);
  or _46469_ (_39247_, _39246_, _35360_);
  and _46470_ (_39248_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46471_ (_39249_, _35349_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _46472_ (_39250_, _39249_, _35393_);
  and _46473_ (_39251_, _39250_, _38936_);
  or _46474_ (_39252_, _39251_, _39248_);
  and _46475_ (_39253_, _39252_, _31899_);
  nand _46476_ (_39254_, _38942_, _38169_);
  or _46477_ (_39255_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46478_ (_39256_, _39255_, _31212_);
  and _46479_ (_39257_, _39256_, _39254_);
  not _46480_ (_39258_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor _46481_ (_39259_, _31211_, _39258_);
  or _46482_ (_39260_, _39259_, rst);
  or _46483_ (_39261_, _39260_, _39257_);
  or _46484_ (_40316_, _39261_, _39253_);
  and _46485_ (_39262_, _38936_, _36133_);
  nand _46486_ (_39263_, _39262_, _31757_);
  or _46487_ (_39264_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _46488_ (_39265_, _39264_, _31899_);
  and _46489_ (_39266_, _39265_, _39263_);
  nand _46490_ (_39267_, _38942_, _38162_);
  or _46491_ (_39268_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _46492_ (_39269_, _39268_, _31212_);
  and _46493_ (_39270_, _39269_, _39267_);
  and _46494_ (_39271_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _46495_ (_39272_, _39271_, rst);
  or _46496_ (_39273_, _39272_, _39270_);
  or _46497_ (_40318_, _39273_, _39266_);
  and _46498_ (_39274_, _38936_, _36785_);
  nand _46499_ (_39275_, _39274_, _31757_);
  or _46500_ (_39276_, _39274_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _46501_ (_39277_, _39276_, _31899_);
  and _46502_ (_39278_, _39277_, _39275_);
  nand _46503_ (_39279_, _38942_, _38155_);
  or _46504_ (_39280_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _46505_ (_39281_, _39280_, _31212_);
  and _46506_ (_39282_, _39281_, _39279_);
  and _46507_ (_39283_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _46508_ (_39284_, _39283_, rst);
  or _46509_ (_39285_, _39284_, _39282_);
  or _46510_ (_40320_, _39285_, _39278_);
  and _46511_ (_39286_, _38951_, _38813_);
  nand _46512_ (_39287_, _39286_, _31757_);
  or _46513_ (_39288_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _46514_ (_39289_, _39288_, _31899_);
  and _46515_ (_39290_, _39289_, _39287_);
  nand _46516_ (_39291_, _38958_, _38203_);
  and _46517_ (_39292_, _39291_, _31212_);
  and _46518_ (_39293_, _39292_, _39288_);
  not _46519_ (_39294_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _46520_ (_39295_, _31211_, _39294_);
  or _46521_ (_39296_, _39295_, rst);
  or _46522_ (_39297_, _39296_, _39293_);
  or _46523_ (_40322_, _39297_, _39290_);
  and _46524_ (_39298_, _38951_, _33129_);
  nand _46525_ (_39299_, _39298_, _31757_);
  or _46526_ (_39300_, _39298_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _46527_ (_39301_, _39300_, _31899_);
  and _46528_ (_39302_, _39301_, _39299_);
  nand _46529_ (_39303_, _38958_, _38191_);
  or _46530_ (_39304_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _46531_ (_39305_, _39304_, _31212_);
  and _46532_ (_39306_, _39305_, _39303_);
  and _46533_ (_39307_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _46534_ (_39308_, _39307_, rst);
  or _46535_ (_39309_, _39308_, _39306_);
  or _46536_ (_40324_, _39309_, _39302_);
  and _46537_ (_39310_, _38951_, _33847_);
  nand _46538_ (_39311_, _39310_, _31757_);
  or _46539_ (_39312_, _39310_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _46540_ (_39313_, _39312_, _31899_);
  and _46541_ (_39314_, _39313_, _39311_);
  nand _46542_ (_39315_, _38958_, _38184_);
  or _46543_ (_39316_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _46544_ (_39317_, _39316_, _31212_);
  and _46545_ (_39318_, _39317_, _39315_);
  and _46546_ (_39319_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _46547_ (_39320_, _39319_, rst);
  or _46548_ (_39321_, _39320_, _39318_);
  or _46549_ (_40326_, _39321_, _39314_);
  and _46550_ (_39322_, _38951_, _34576_);
  nand _46551_ (_39323_, _39322_, _31757_);
  or _46552_ (_39324_, _39322_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _46553_ (_39325_, _39324_, _31899_);
  and _46554_ (_39326_, _39325_, _39323_);
  nand _46555_ (_39327_, _38958_, _38177_);
  or _46556_ (_39328_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _46557_ (_39329_, _39328_, _31212_);
  and _46558_ (_39330_, _39329_, _39327_);
  and _46559_ (_39331_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _46560_ (_39332_, _39331_, rst);
  or _46561_ (_39333_, _39332_, _39330_);
  or _46562_ (_40327_, _39333_, _39326_);
  and _46563_ (_39334_, _38951_, _35338_);
  nand _46564_ (_39335_, _39334_, _31757_);
  or _46565_ (_39336_, _39334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _46566_ (_39337_, _39336_, _31899_);
  and _46567_ (_39338_, _39337_, _39335_);
  nand _46568_ (_39339_, _38958_, _38169_);
  or _46569_ (_39340_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _46570_ (_39341_, _39340_, _31212_);
  and _46571_ (_39342_, _39341_, _39339_);
  not _46572_ (_39343_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor _46573_ (_39344_, _31211_, _39343_);
  or _46574_ (_39345_, _39344_, rst);
  or _46575_ (_39346_, _39345_, _39342_);
  or _46576_ (_40329_, _39346_, _39338_);
  and _46577_ (_39347_, _38951_, _36133_);
  nand _46578_ (_39348_, _39347_, _31757_);
  or _46579_ (_39349_, _39347_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _46580_ (_39350_, _39349_, _31899_);
  and _46581_ (_39351_, _39350_, _39348_);
  nand _46582_ (_39352_, _38958_, _38162_);
  or _46583_ (_39353_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _46584_ (_39354_, _39353_, _31212_);
  and _46585_ (_39355_, _39354_, _39352_);
  and _46586_ (_39356_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _46587_ (_39357_, _39356_, rst);
  or _46588_ (_39358_, _39357_, _39355_);
  or _46589_ (_40331_, _39358_, _39351_);
  and _46590_ (_39359_, _38951_, _36785_);
  nand _46591_ (_39360_, _39359_, _31757_);
  or _46592_ (_39361_, _39359_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _46593_ (_39362_, _39361_, _31899_);
  and _46594_ (_39363_, _39362_, _39360_);
  nand _46595_ (_39364_, _38958_, _38155_);
  or _46596_ (_39365_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _46597_ (_39366_, _39365_, _31212_);
  and _46598_ (_39367_, _39366_, _39364_);
  and _46599_ (_39368_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _46600_ (_39369_, _39368_, rst);
  or _46601_ (_39370_, _39369_, _39367_);
  or _46602_ (_40333_, _39370_, _39363_);
  nand _46603_ (_39371_, _38974_, _31757_);
  or _46604_ (_39372_, _38974_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _46605_ (_39373_, _39372_, _31899_);
  and _46606_ (_39374_, _39373_, _39371_);
  nor _46607_ (_39375_, _38975_, _38203_);
  not _46608_ (_39376_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _46609_ (_39377_, _38974_, _39376_);
  or _46610_ (_39378_, _39377_, _39375_);
  and _46611_ (_39379_, _39378_, _31212_);
  nor _46612_ (_39380_, _31211_, _39376_);
  or _46613_ (_39381_, _39380_, rst);
  or _46614_ (_39382_, _39381_, _39379_);
  or _46615_ (_40335_, _39382_, _39374_);
  and _46616_ (_39383_, _38967_, _33129_);
  nand _46617_ (_39384_, _39383_, _31757_);
  or _46618_ (_39385_, _39383_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _46619_ (_39386_, _39385_, _31899_);
  and _46620_ (_39387_, _39386_, _39384_);
  nor _46621_ (_39388_, _38975_, _38191_);
  and _46622_ (_39389_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _46623_ (_39390_, _39389_, _39388_);
  and _46624_ (_39391_, _39390_, _31212_);
  and _46625_ (_39392_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _46626_ (_39393_, _39392_, rst);
  or _46627_ (_39394_, _39393_, _39391_);
  or _46628_ (_40337_, _39394_, _39387_);
  and _46629_ (_39395_, _38967_, _33847_);
  nand _46630_ (_39396_, _39395_, _31757_);
  or _46631_ (_39397_, _39395_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _46632_ (_39398_, _39397_, _31899_);
  and _46633_ (_39399_, _39398_, _39396_);
  nor _46634_ (_39400_, _38975_, _38184_);
  and _46635_ (_39401_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _46636_ (_39402_, _39401_, _39400_);
  and _46637_ (_39403_, _39402_, _31212_);
  and _46638_ (_39404_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _46639_ (_39405_, _39404_, rst);
  or _46640_ (_39406_, _39405_, _39403_);
  or _46641_ (_40339_, _39406_, _39399_);
  and _46642_ (_39407_, _38967_, _34576_);
  nand _46643_ (_39408_, _39407_, _31757_);
  or _46644_ (_39409_, _39407_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _46645_ (_39410_, _39409_, _31899_);
  and _46646_ (_39411_, _39410_, _39408_);
  nor _46647_ (_39412_, _38975_, _38177_);
  and _46648_ (_39413_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _46649_ (_39414_, _39413_, _39412_);
  and _46650_ (_39415_, _39414_, _31212_);
  and _46651_ (_39416_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _46652_ (_39417_, _39416_, rst);
  or _46653_ (_39418_, _39417_, _39415_);
  or _46654_ (_40341_, _39418_, _39411_);
  and _46655_ (_39419_, _38967_, _35338_);
  nand _46656_ (_39420_, _39419_, _31757_);
  or _46657_ (_39421_, _39419_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _46658_ (_39422_, _39421_, _31899_);
  and _46659_ (_39423_, _39422_, _39420_);
  nor _46660_ (_39424_, _38975_, _38169_);
  not _46661_ (_39425_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor _46662_ (_39426_, _38974_, _39425_);
  or _46663_ (_39427_, _39426_, _39424_);
  and _46664_ (_39428_, _39427_, _31212_);
  nor _46665_ (_39429_, _31211_, _39425_);
  or _46666_ (_39430_, _39429_, rst);
  or _46667_ (_39431_, _39430_, _39428_);
  or _46668_ (_40343_, _39431_, _39423_);
  and _46669_ (_39432_, _38967_, _36133_);
  nand _46670_ (_39433_, _39432_, _31757_);
  or _46671_ (_39434_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _46672_ (_39435_, _39434_, _31899_);
  and _46673_ (_39436_, _39435_, _39433_);
  nor _46674_ (_39437_, _38975_, _38162_);
  and _46675_ (_39438_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _46676_ (_39439_, _39438_, _39437_);
  and _46677_ (_39440_, _39439_, _31212_);
  and _46678_ (_39441_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _46679_ (_39442_, _39441_, rst);
  or _46680_ (_39443_, _39442_, _39440_);
  or _46681_ (_40345_, _39443_, _39436_);
  and _46682_ (_39444_, _38967_, _36785_);
  nand _46683_ (_39445_, _39444_, _31757_);
  or _46684_ (_39446_, _39444_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _46685_ (_39447_, _39446_, _31899_);
  and _46686_ (_39448_, _39447_, _39445_);
  nor _46687_ (_39449_, _38975_, _38155_);
  and _46688_ (_39450_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _46689_ (_39451_, _39450_, _39449_);
  and _46690_ (_39452_, _39451_, _31212_);
  and _46691_ (_39453_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _46692_ (_39454_, _39453_, rst);
  or _46693_ (_39455_, _39454_, _39452_);
  or _46694_ (_40347_, _39455_, _39448_);
  and _46695_ (_39456_, _38983_, _38813_);
  nand _46696_ (_39461_, _39456_, _31757_);
  or _46697_ (_39467_, _39456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _46698_ (_39468_, _39467_, _31899_);
  and _46699_ (_39469_, _39468_, _39461_);
  nor _46700_ (_39470_, _38991_, _38203_);
  not _46701_ (_39471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _46702_ (_39472_, _38990_, _39471_);
  or _46703_ (_39473_, _39472_, _39470_);
  and _46704_ (_39474_, _39473_, _31212_);
  nor _46705_ (_39475_, _31211_, _39471_);
  or _46706_ (_39476_, _39475_, rst);
  or _46707_ (_39477_, _39476_, _39474_);
  or _46708_ (_40349_, _39477_, _39469_);
  and _46709_ (_39478_, _38983_, _33129_);
  nand _46710_ (_39479_, _39478_, _31757_);
  or _46711_ (_39480_, _39478_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _46712_ (_39481_, _39480_, _31899_);
  and _46713_ (_39482_, _39481_, _39479_);
  nor _46714_ (_39483_, _38991_, _38191_);
  and _46715_ (_39484_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _46716_ (_39485_, _39484_, _39483_);
  and _46717_ (_39486_, _39485_, _31212_);
  and _46718_ (_39487_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _46719_ (_39488_, _39487_, rst);
  or _46720_ (_39489_, _39488_, _39486_);
  or _46721_ (_40351_, _39489_, _39482_);
  and _46722_ (_39490_, _38983_, _33847_);
  nand _46723_ (_39491_, _39490_, _31757_);
  or _46724_ (_39492_, _39490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _46725_ (_39493_, _39492_, _31899_);
  and _46726_ (_39494_, _39493_, _39491_);
  nor _46727_ (_39495_, _38991_, _38184_);
  and _46728_ (_39496_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _46729_ (_39497_, _39496_, _39495_);
  and _46730_ (_39498_, _39497_, _31212_);
  and _46731_ (_39499_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _46732_ (_39500_, _39499_, rst);
  or _46733_ (_39501_, _39500_, _39498_);
  or _46734_ (_40353_, _39501_, _39494_);
  and _46735_ (_39502_, _38983_, _34576_);
  nand _46736_ (_39503_, _39502_, _31757_);
  or _46737_ (_39504_, _39502_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _46738_ (_39505_, _39504_, _31899_);
  and _46739_ (_39506_, _39505_, _39503_);
  nor _46740_ (_39507_, _38991_, _38177_);
  and _46741_ (_39508_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _46742_ (_39509_, _39508_, _39507_);
  and _46743_ (_39510_, _39509_, _31212_);
  and _46744_ (_39511_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _46745_ (_39512_, _39511_, rst);
  or _46746_ (_39513_, _39512_, _39510_);
  or _46747_ (_40355_, _39513_, _39506_);
  and _46748_ (_39514_, _38983_, _35338_);
  nand _46749_ (_39515_, _39514_, _31757_);
  or _46750_ (_39516_, _39514_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _46751_ (_39517_, _39516_, _31899_);
  and _46752_ (_39518_, _39517_, _39515_);
  nor _46753_ (_39519_, _38991_, _38169_);
  not _46754_ (_39520_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor _46755_ (_39521_, _38990_, _39520_);
  or _46756_ (_39522_, _39521_, _39519_);
  and _46757_ (_39523_, _39522_, _31212_);
  nor _46758_ (_39524_, _31211_, _39520_);
  or _46759_ (_39525_, _39524_, rst);
  or _46760_ (_39526_, _39525_, _39523_);
  or _46761_ (_40356_, _39526_, _39518_);
  and _46762_ (_39527_, _38983_, _36133_);
  nand _46763_ (_39528_, _39527_, _31757_);
  or _46764_ (_39529_, _39527_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _46765_ (_39530_, _39529_, _31899_);
  and _46766_ (_39531_, _39530_, _39528_);
  nor _46767_ (_39532_, _38991_, _38162_);
  and _46768_ (_39533_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _46769_ (_39534_, _39533_, _39532_);
  and _46770_ (_39535_, _39534_, _31212_);
  and _46771_ (_39536_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _46772_ (_39537_, _39536_, rst);
  or _46773_ (_39538_, _39537_, _39535_);
  or _46774_ (_40358_, _39538_, _39531_);
  and _46775_ (_39539_, _38983_, _36785_);
  nand _46776_ (_39540_, _39539_, _31757_);
  or _46777_ (_39541_, _39539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _46778_ (_39542_, _39541_, _31899_);
  and _46779_ (_39543_, _39542_, _39540_);
  nor _46780_ (_39544_, _38991_, _38155_);
  and _46781_ (_39545_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _46782_ (_39546_, _39545_, _39544_);
  and _46783_ (_39547_, _39546_, _31212_);
  and _46784_ (_39548_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _46785_ (_39549_, _39548_, rst);
  or _46786_ (_39550_, _39549_, _39547_);
  or _46787_ (_40360_, _39550_, _39543_);
  and _46788_ (_40810_, t0_i, _42618_);
  and _46789_ (_40813_, t1_i, _42618_);
  not _46790_ (_39551_, _31212_);
  nor _46791_ (_39552_, _39551_, _27948_);
  and _46792_ (_39553_, _39552_, _34576_);
  and _46793_ (_39554_, _39553_, _38140_);
  nand _46794_ (_39565_, _39554_, _38225_);
  nor _46795_ (_39576_, _28069_, _27948_);
  and _46796_ (_39587_, _39576_, _38141_);
  and _46797_ (_39598_, _39587_, _31212_);
  not _46798_ (_39609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _46799_ (_39616_, _39609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _46800_ (_39617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _46801_ (_39618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _39617_);
  nor _46802_ (_39619_, _39618_, _39616_);
  or _46803_ (_39620_, _39619_, _39598_);
  and _46804_ (_39621_, _39620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _46805_ (_39622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _46806_ (_39623_, t1_i);
  and _46807_ (_39624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _39623_);
  nor _46808_ (_39625_, _39624_, _39622_);
  not _46809_ (_39626_, _39625_);
  not _46810_ (_39627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _46811_ (_39628_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39627_);
  nor _46812_ (_39629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _46813_ (_39630_, _39629_);
  and _46814_ (_39631_, _39630_, _39628_);
  and _46815_ (_39632_, _39631_, _39626_);
  not _46816_ (_39633_, _39632_);
  nand _46817_ (_39634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _46818_ (_39635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or _46819_ (_39636_, _39635_, _39634_);
  nor _46820_ (_39637_, _39636_, _39633_);
  and _46821_ (_39638_, _39637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _46822_ (_39639_, _39638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _46823_ (_39640_, _39639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _46824_ (_39641_, _39640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _46825_ (_39642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _46826_ (_39643_, _39636_, _39642_);
  and _46827_ (_39644_, _39643_, _39632_);
  and _46828_ (_39645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _46829_ (_39646_, _39645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _46830_ (_39647_, _39646_, _39644_);
  nor _46831_ (_39648_, _39647_, _39619_);
  and _46832_ (_39649_, _39648_, _39641_);
  and _46833_ (_39650_, _39647_, _39616_);
  and _46834_ (_39651_, _39650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _46835_ (_39652_, _39651_, _39649_);
  nor _46836_ (_39653_, _39652_, _39598_);
  or _46837_ (_39654_, _39653_, _39621_);
  or _46838_ (_39655_, _39554_, _39654_);
  and _46839_ (_39656_, _39655_, _42618_);
  and _46840_ (_40816_, _39656_, _39565_);
  and _46841_ (_39657_, _39552_, _38272_);
  and _46842_ (_39658_, _39657_, _42618_);
  and _46843_ (_39659_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _46844_ (_39660_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _46845_ (_39661_, _39660_);
  and _46846_ (_39662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _46847_ (_39663_, _39662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _46848_ (_39664_, _39663_, _39644_);
  and _46849_ (_39665_, _39664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _46850_ (_39666_, _39665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _46851_ (_39667_, _39666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _46852_ (_39668_, _39667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _46853_ (_39669_, _39668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _46854_ (_39670_, _39669_, _39661_);
  and _46855_ (_39671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not _46856_ (_39672_, _39618_);
  and _46857_ (_39673_, _39669_, _39646_);
  nor _46858_ (_39674_, _39673_, _39672_);
  or _46859_ (_39675_, _39674_, _39671_);
  or _46860_ (_39676_, _39646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _46861_ (_39677_, _39676_, _39675_);
  or _46862_ (_39678_, _39677_, _39670_);
  nor _46863_ (_39680_, _39668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _46864_ (_39686_, _39680_, _39598_);
  and _46865_ (_39687_, _39686_, _39678_);
  not _46866_ (_39688_, _39598_);
  nor _46867_ (_39689_, _39688_, _38225_);
  or _46868_ (_39690_, _39689_, _39687_);
  nor _46869_ (_39691_, _39554_, rst);
  and _46870_ (_39692_, _39691_, _39690_);
  or _46871_ (_40819_, _39692_, _39659_);
  and _46872_ (_39693_, _39633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or _46873_ (_39694_, _39693_, _39673_);
  and _46874_ (_39695_, _39694_, _39618_);
  or _46875_ (_39696_, _39693_, _39669_);
  and _46876_ (_39697_, _39696_, _39660_);
  nand _46877_ (_39698_, _39632_, _39609_);
  and _46878_ (_39699_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _46879_ (_39700_, _39699_, _39698_);
  or _46880_ (_39701_, _39700_, _39650_);
  or _46881_ (_39702_, _39701_, _39697_);
  nor _46882_ (_39703_, _39702_, _39695_);
  nor _46883_ (_39704_, _39703_, _39598_);
  and _46884_ (_40822_, _39704_, _39691_);
  and _46885_ (_39705_, _39552_, _35338_);
  and _46886_ (_39706_, _39705_, _38140_);
  nor _46887_ (_39707_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _46888_ (_39708_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _46889_ (_39709_, t0_i);
  and _46890_ (_39710_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _39709_);
  nor _46891_ (_39711_, _39710_, _39708_);
  not _46892_ (_39712_, _39711_);
  not _46893_ (_39713_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _46894_ (_39714_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _46895_ (_39715_, _39714_, _39713_);
  and _46896_ (_39716_, _39715_, _39712_);
  not _46897_ (_39717_, _39716_);
  and _46898_ (_39718_, _39717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and _46899_ (_39719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _46900_ (_39720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _46901_ (_39721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _46902_ (_39722_, _39721_, _39720_);
  and _46903_ (_39723_, _39722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _46904_ (_39724_, _39723_, _39716_);
  and _46905_ (_39725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _46906_ (_39726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _46907_ (_39727_, _39726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _46908_ (_39728_, _39727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _46909_ (_39729_, _39728_, _39725_);
  and _46910_ (_39730_, _39729_, _39724_);
  and _46911_ (_39731_, _39730_, _39719_);
  or _46912_ (_39732_, _39731_, _39718_);
  and _46913_ (_39733_, _39732_, _39707_);
  and _46914_ (_39734_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _46915_ (_39735_, _39734_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _46916_ (_39736_, _39735_, _39723_);
  and _46917_ (_39737_, _39736_, _39716_);
  or _46918_ (_39738_, _39737_, _39718_);
  not _46919_ (_39739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _46920_ (_39740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _39739_);
  and _46921_ (_39741_, _39729_, _39719_);
  or _46922_ (_39742_, _39741_, _39718_);
  and _46923_ (_39743_, _39742_, _39740_);
  or _46924_ (_39744_, _39743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _46925_ (_39745_, _39744_, _39738_);
  or _46926_ (_39746_, _39745_, _39733_);
  nand _46927_ (_39747_, _39746_, _42618_);
  nor _46928_ (_39748_, _39747_, _39706_);
  and _46929_ (_39749_, _39552_, _33847_);
  and _46930_ (_39750_, _39749_, _38140_);
  not _46931_ (_39751_, _39750_);
  and _46932_ (_40825_, _39751_, _39748_);
  and _46933_ (_39752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _46934_ (_39753_, _39752_, _39724_);
  or _46935_ (_39754_, _39753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _46936_ (_39755_, _39707_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _46937_ (_39756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _46938_ (_39757_, _39756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _46939_ (_39758_, _39757_, _39740_);
  and _46940_ (_39759_, _39735_, _39724_);
  not _46941_ (_39760_, _39759_);
  and _46942_ (_39761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _46943_ (_39762_, _39761_, _39760_);
  or _46944_ (_39763_, _39762_, _39758_);
  nand _46945_ (_39767_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _46946_ (_39775_, _39767_, _39759_);
  and _46947_ (_39776_, _39775_, _39763_);
  or _46948_ (_39777_, _39776_, _39755_);
  and _46949_ (_39778_, _39777_, _39754_);
  or _46950_ (_39779_, _39778_, _39706_);
  and _46951_ (_39780_, _39552_, _38371_);
  not _46952_ (_39781_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _46953_ (_39782_, _39706_, _39781_);
  nor _46954_ (_39783_, _39782_, _39780_);
  and _46955_ (_39784_, _39783_, _39779_);
  nor _46956_ (_39785_, _39751_, _38225_);
  or _46957_ (_39786_, _39785_, _39784_);
  and _46958_ (_40828_, _39786_, _42618_);
  not _46959_ (_39787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _46960_ (_39788_, _39716_, _39739_);
  and _46961_ (_39789_, _39788_, _39736_);
  and _46962_ (_39790_, _39789_, _39729_);
  and _46963_ (_39791_, _39790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _46964_ (_39792_, _39791_, _39787_);
  and _46965_ (_39793_, _39791_, _39787_);
  or _46966_ (_39794_, _39793_, _39792_);
  and _46967_ (_39795_, _39794_, _39758_);
  and _46968_ (_39796_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _46969_ (_39797_, _39796_, _39728_);
  and _46970_ (_39798_, _39797_, _39725_);
  and _46971_ (_39799_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _46972_ (_39800_, _39799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _46973_ (_39801_, _39796_, _39741_);
  and _46974_ (_39802_, _39801_, _39800_);
  and _46975_ (_39803_, _39802_, _39761_);
  and _46976_ (_39804_, _39730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _46977_ (_39805_, _39804_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not _46978_ (_39806_, _39707_);
  nor _46979_ (_39807_, _39731_, _39806_);
  and _46980_ (_39808_, _39807_, _39805_);
  or _46981_ (_39809_, _39808_, _39803_);
  or _46982_ (_39810_, _39809_, _39795_);
  or _46983_ (_39811_, _39810_, _39706_);
  nand _46984_ (_39812_, _39706_, _38225_);
  and _46985_ (_39813_, _39812_, _39811_);
  or _46986_ (_39814_, _39813_, _39750_);
  nand _46987_ (_39815_, _39750_, _39787_);
  and _46988_ (_39816_, _39815_, _42618_);
  and _46989_ (_40831_, _39816_, _39814_);
  not _46990_ (_39817_, _39796_);
  or _46991_ (_39818_, _39817_, _39741_);
  or _46992_ (_39819_, _39796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _46993_ (_39820_, _39761_, _42618_);
  and _46994_ (_39821_, _39820_, _39819_);
  nand _46995_ (_39822_, _39821_, _39818_);
  nor _46996_ (_39823_, _39822_, _39706_);
  and _46997_ (_40834_, _39823_, _39751_);
  and _46998_ (_39824_, _39552_, _38142_);
  or _46999_ (_39825_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _47000_ (_39826_, _39825_, _42618_);
  nand _47001_ (_39827_, _39824_, _38225_);
  and _47002_ (_40837_, _39827_, _39826_);
  not _47003_ (_39828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _47004_ (_39829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _47005_ (_39830_, _39829_, _39598_);
  and _47006_ (_39831_, _39830_, _39632_);
  nor _47007_ (_39832_, _39831_, _39828_);
  and _47008_ (_39833_, _39831_, _39828_);
  or _47009_ (_39834_, _39833_, _39832_);
  and _47010_ (_39835_, _39646_, _39643_);
  and _47011_ (_39836_, _39835_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _47012_ (_39837_, _39836_, _39616_);
  nor _47013_ (_39838_, _39837_, _39598_);
  or _47014_ (_39839_, _39838_, _39554_);
  or _47015_ (_39840_, _39839_, _39834_);
  nand _47016_ (_39841_, _39554_, _38203_);
  and _47017_ (_39842_, _39841_, _42618_);
  and _47018_ (_41323_, _39842_, _39840_);
  not _47019_ (_39847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _47020_ (_39848_, _39830_, _39847_);
  not _47021_ (_39849_, _39829_);
  and _47022_ (_39850_, _39632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _47023_ (_39851_, _39850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _47024_ (_39852_, _39850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _47025_ (_39853_, _39852_, _39851_);
  and _47026_ (_39854_, _39853_, _39849_);
  and _47027_ (_39855_, _39640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _47028_ (_39856_, _39855_, _39616_);
  and _47029_ (_39857_, _39856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _47030_ (_39858_, _39857_, _39854_);
  nor _47031_ (_39859_, _39858_, _39598_);
  or _47032_ (_39860_, _39859_, _39554_);
  or _47033_ (_39861_, _39860_, _39848_);
  nand _47034_ (_39862_, _39554_, _38191_);
  and _47035_ (_39863_, _39862_, _42618_);
  and _47036_ (_41325_, _39863_, _39861_);
  not _47037_ (_39873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _47038_ (_39874_, _39830_, _39873_);
  nor _47039_ (_39875_, _39851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _47040_ (_39876_, _39851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _47041_ (_39877_, _39876_, _39875_);
  and _47042_ (_39878_, _39877_, _39849_);
  and _47043_ (_39879_, _39650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _47044_ (_39880_, _39879_, _39878_);
  nor _47045_ (_39881_, _39880_, _39598_);
  or _47046_ (_39882_, _39881_, _39874_);
  and _47047_ (_39883_, _39882_, _39691_);
  not _47048_ (_39884_, _38184_);
  and _47049_ (_39885_, _39658_, _39884_);
  or _47050_ (_41327_, _39885_, _39883_);
  not _47051_ (_39886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _47052_ (_39887_, _39830_, _39886_);
  or _47053_ (_39888_, _39876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _47054_ (_39889_, _39829_, _39637_);
  and _47055_ (_39890_, _39889_, _39888_);
  and _47056_ (_39891_, _39650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _47057_ (_39892_, _39891_, _39890_);
  nor _47058_ (_39893_, _39892_, _39598_);
  or _47059_ (_39894_, _39893_, _39887_);
  and _47060_ (_39895_, _39894_, _39691_);
  not _47061_ (_39896_, _38177_);
  and _47062_ (_39897_, _39658_, _39896_);
  or _47063_ (_41328_, _39897_, _39895_);
  nor _47064_ (_39898_, _39830_, _39642_);
  and _47065_ (_39899_, _39856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _47066_ (_39900_, _39637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _47067_ (_39901_, _39900_, _39644_);
  and _47068_ (_39902_, _39901_, _39849_);
  nor _47069_ (_39903_, _39902_, _39899_);
  nor _47070_ (_39904_, _39903_, _39598_);
  or _47071_ (_39905_, _39904_, _39898_);
  and _47072_ (_39906_, _39905_, _39691_);
  not _47073_ (_39907_, _38169_);
  and _47074_ (_39908_, _39658_, _39907_);
  or _47075_ (_41330_, _39908_, _39906_);
  and _47076_ (_39909_, _39620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _47077_ (_39910_, _39856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _47078_ (_39911_, _39619_);
  and _47079_ (_39912_, _39644_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _47080_ (_39913_, _39644_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _47081_ (_39914_, _39913_, _39912_);
  and _47082_ (_39915_, _39914_, _39911_);
  nor _47083_ (_39916_, _39915_, _39910_);
  nor _47084_ (_39917_, _39916_, _39598_);
  or _47085_ (_39918_, _39917_, _39909_);
  and _47086_ (_39919_, _39918_, _39691_);
  not _47087_ (_39920_, _38162_);
  and _47088_ (_39921_, _39658_, _39920_);
  or _47089_ (_41332_, _39921_, _39919_);
  and _47090_ (_39922_, _39620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _47091_ (_39923_, _39616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47092_ (_39924_, _39923_, _39632_);
  and _47093_ (_39925_, _39924_, _39835_);
  or _47094_ (_39926_, _39912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _47095_ (_39927_, _39926_, _39911_);
  nor _47096_ (_39928_, _39927_, _39640_);
  nor _47097_ (_39929_, _39928_, _39925_);
  nor _47098_ (_39930_, _39929_, _39598_);
  or _47099_ (_39931_, _39930_, _39922_);
  and _47100_ (_39932_, _39931_, _39691_);
  not _47101_ (_39933_, _38155_);
  and _47102_ (_39934_, _39658_, _39933_);
  or _47103_ (_41334_, _39934_, _39932_);
  and _47104_ (_39935_, _39644_, _39617_);
  nor _47105_ (_39936_, _39646_, _39609_);
  not _47106_ (_39937_, _39936_);
  and _47107_ (_39938_, _39937_, _39935_);
  nand _47108_ (_39939_, _39938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or _47109_ (_39940_, _39938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47110_ (_39941_, _39940_, _39939_);
  or _47111_ (_39942_, _39941_, _39598_);
  nand _47112_ (_39943_, _39598_, _38203_);
  and _47113_ (_39944_, _39943_, _39691_);
  and _47114_ (_39945_, _39944_, _39942_);
  and _47115_ (_39946_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or _47116_ (_41336_, _39946_, _39945_);
  nand _47117_ (_39947_, _39598_, _38191_);
  nor _47118_ (_39948_, _39647_, _39672_);
  not _47119_ (_39949_, _39948_);
  not _47120_ (_39950_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _47121_ (_39951_, _39935_, _39618_);
  nor _47122_ (_39952_, _39951_, _39950_);
  and _47123_ (_39953_, _39952_, _39949_);
  or _47124_ (_39954_, _39953_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _47125_ (_39955_, _39953_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _47126_ (_39956_, _39955_, _39954_);
  or _47127_ (_39957_, _39956_, _39598_);
  and _47128_ (_39958_, _39957_, _39691_);
  and _47129_ (_39959_, _39958_, _39947_);
  and _47130_ (_39960_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _47131_ (_41338_, _39960_, _39959_);
  nand _47132_ (_39961_, _39598_, _38184_);
  or _47133_ (_39962_, _39936_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _47134_ (_39963_, _39962_);
  and _47135_ (_39964_, _39662_, _39644_);
  and _47136_ (_39965_, _39964_, _39963_);
  or _47137_ (_39966_, _39965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _47138_ (_39967_, _39664_, _39617_);
  nand _47139_ (_39968_, _39937_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _47140_ (_39969_, _39968_, _39967_);
  and _47141_ (_39970_, _39969_, _39966_);
  or _47142_ (_39971_, _39970_, _39598_);
  and _47143_ (_39972_, _39971_, _39691_);
  and _47144_ (_39973_, _39972_, _39961_);
  and _47145_ (_39974_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _47146_ (_41340_, _39974_, _39973_);
  nand _47147_ (_39975_, _39598_, _38177_);
  and _47148_ (_39976_, _39665_, _39646_);
  and _47149_ (_39977_, _39664_, _39646_);
  or _47150_ (_39978_, _39977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _47151_ (_39979_, _39978_, _39618_);
  nor _47152_ (_39980_, _39979_, _39976_);
  and _47153_ (_39981_, _39967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _47154_ (_39982_, _39967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _47155_ (_39983_, _39982_, _39981_);
  and _47156_ (_39984_, _39983_, _39672_);
  or _47157_ (_39985_, _39984_, _39980_);
  or _47158_ (_39986_, _39985_, _39598_);
  and _47159_ (_39987_, _39986_, _39691_);
  and _47160_ (_39988_, _39987_, _39975_);
  and _47161_ (_39989_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _47162_ (_41342_, _39989_, _39988_);
  nand _47163_ (_39990_, _39598_, _38169_);
  or _47164_ (_39991_, _39976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _47165_ (_39992_, _39991_, _39618_);
  and _47166_ (_39993_, _39976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _47167_ (_39994_, _39993_, _39992_);
  and _47168_ (_39995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47169_ (_39996_, _39662_, _39643_);
  and _47170_ (_39997_, _39996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47171_ (_39998_, _39997_, _39632_);
  and _47172_ (_39999_, _39998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _47173_ (_40000_, _39999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _47174_ (_40001_, _39999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47175_ (_40002_, _40001_, _40000_);
  and _47176_ (_40003_, _40002_, _39660_);
  or _47177_ (_40004_, _40003_, _39995_);
  or _47178_ (_40005_, _40004_, _39994_);
  or _47179_ (_40006_, _40005_, _39598_);
  and _47180_ (_40007_, _40006_, _39691_);
  and _47181_ (_40008_, _40007_, _39990_);
  and _47182_ (_40009_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _47183_ (_41344_, _40009_, _40008_);
  nand _47184_ (_40010_, _39598_, _38162_);
  not _47185_ (_40011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47186_ (_40012_, _39666_, _39660_);
  and _47187_ (_40013_, _39993_, _39618_);
  nor _47188_ (_40014_, _40013_, _40012_);
  nand _47189_ (_40015_, _40014_, _40011_);
  or _47190_ (_40016_, _40014_, _40011_);
  and _47191_ (_40017_, _40016_, _40015_);
  or _47192_ (_40018_, _40017_, _39598_);
  and _47193_ (_40019_, _40018_, _39691_);
  and _47194_ (_40020_, _40019_, _40010_);
  and _47195_ (_40021_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _47196_ (_41345_, _40021_, _40020_);
  nand _47197_ (_40022_, _39598_, _38155_);
  and _47198_ (_40023_, _39963_, _39667_);
  or _47199_ (_40024_, _40023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _47200_ (_40025_, _40023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47201_ (_40026_, _40025_, _40024_);
  or _47202_ (_40027_, _40026_, _39598_);
  and _47203_ (_40028_, _40027_, _39691_);
  and _47204_ (_40029_, _40028_, _40022_);
  and _47205_ (_40030_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _47206_ (_41347_, _40030_, _40029_);
  nor _47207_ (_40031_, _39717_, _39706_);
  or _47208_ (_40032_, _40031_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47209_ (_40033_, _39716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47210_ (_40034_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47211_ (_40035_, _40034_, _39736_);
  nand _47212_ (_40036_, _40035_, _40033_);
  or _47213_ (_40037_, _40036_, _39706_);
  and _47214_ (_40038_, _40037_, _40032_);
  or _47215_ (_40039_, _40038_, _39750_);
  nand _47216_ (_40040_, _39750_, _38203_);
  and _47217_ (_40041_, _40040_, _42618_);
  and _47218_ (_41349_, _40041_, _40039_);
  nor _47219_ (_40042_, _40033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _47220_ (_40043_, _40033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _47221_ (_40044_, _40043_, _40042_);
  and _47222_ (_40045_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _47223_ (_40046_, _40045_, _39759_);
  nor _47224_ (_40047_, _40046_, _40044_);
  nor _47225_ (_40048_, _40047_, _39706_);
  and _47226_ (_40049_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _47227_ (_40050_, _40049_, _40048_);
  and _47228_ (_40051_, _40050_, _39751_);
  nor _47229_ (_40052_, _39751_, _38191_);
  or _47230_ (_40053_, _40052_, _40051_);
  and _47231_ (_41351_, _40053_, _42618_);
  nand _47232_ (_40054_, _39780_, _38184_);
  and _47233_ (_40055_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _47234_ (_40056_, _40043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _47235_ (_40057_, _40033_, _39720_);
  nor _47236_ (_40058_, _40057_, _40056_);
  and _47237_ (_40059_, _39757_, _39759_);
  and _47238_ (_40060_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _47239_ (_40061_, _40060_, _40058_);
  nor _47240_ (_40062_, _40061_, _39706_);
  or _47241_ (_40063_, _40062_, _40055_);
  or _47242_ (_40064_, _40063_, _39780_);
  and _47243_ (_40065_, _40064_, _42618_);
  and _47244_ (_41353_, _40065_, _40054_);
  nand _47245_ (_40066_, _39780_, _38177_);
  and _47246_ (_40067_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _47247_ (_40068_, _39722_, _39716_);
  nor _47248_ (_40069_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _47249_ (_40070_, _40069_, _40068_);
  and _47250_ (_40071_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _47251_ (_40072_, _40071_, _40070_);
  nor _47252_ (_40073_, _40072_, _39706_);
  or _47253_ (_40074_, _40073_, _40067_);
  or _47254_ (_40075_, _40074_, _39780_);
  and _47255_ (_40076_, _40075_, _42618_);
  and _47256_ (_41355_, _40076_, _40066_);
  nand _47257_ (_40077_, _39780_, _38169_);
  and _47258_ (_40078_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _47259_ (_40079_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _47260_ (_40080_, _40079_, _39724_);
  and _47261_ (_40081_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _47262_ (_40082_, _40081_, _40080_);
  nor _47263_ (_40083_, _40082_, _39706_);
  or _47264_ (_40084_, _40083_, _40078_);
  or _47265_ (_40085_, _40084_, _39780_);
  and _47266_ (_40086_, _40085_, _42618_);
  and _47267_ (_41357_, _40086_, _40077_);
  and _47268_ (_40087_, _39724_, _39806_);
  and _47269_ (_40088_, _40087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _47270_ (_40089_, _40087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _47271_ (_40090_, _40089_, _40088_);
  and _47272_ (_40091_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _47273_ (_40092_, _40091_, _40090_);
  nor _47274_ (_40093_, _40092_, _39706_);
  and _47275_ (_40094_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _47276_ (_40095_, _40094_, _40093_);
  and _47277_ (_40096_, _40095_, _39751_);
  nor _47278_ (_40097_, _39751_, _38162_);
  or _47279_ (_40098_, _40097_, _40096_);
  and _47280_ (_41359_, _40098_, _42618_);
  not _47281_ (_40099_, _40088_);
  nor _47282_ (_40100_, _40099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _47283_ (_40101_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _47284_ (_40102_, _40101_, _39716_);
  and _47285_ (_40103_, _40102_, _39736_);
  nor _47286_ (_40104_, _40103_, _40100_);
  nor _47287_ (_40105_, _40104_, _39706_);
  or _47288_ (_40106_, _40099_, _39706_);
  and _47289_ (_40107_, _40106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _47290_ (_40108_, _40107_, _40105_);
  and _47291_ (_40109_, _40108_, _39751_);
  nor _47292_ (_40110_, _39751_, _38155_);
  or _47293_ (_40111_, _40110_, _40109_);
  and _47294_ (_41361_, _40111_, _42618_);
  or _47295_ (_40112_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47296_ (_40113_, _40112_, _39758_);
  and _47297_ (_40114_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _47298_ (_40115_, _40114_, _40113_);
  and _47299_ (_40116_, _39796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _47300_ (_40117_, _39796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47301_ (_40118_, _40117_, _39761_);
  nor _47302_ (_40119_, _40118_, _40116_);
  and _47303_ (_40120_, _39724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _47304_ (_40121_, _39724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47305_ (_40122_, _40121_, _39707_);
  nor _47306_ (_40123_, _40122_, _40120_);
  or _47307_ (_40124_, _40123_, _40119_);
  or _47308_ (_40125_, _40124_, _40115_);
  or _47309_ (_40126_, _40125_, _39706_);
  nand _47310_ (_40127_, _39706_, _38203_);
  and _47311_ (_40128_, _40127_, _40126_);
  or _47312_ (_40129_, _40128_, _39750_);
  or _47313_ (_40130_, _39751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _47314_ (_40131_, _40130_, _42618_);
  and _47315_ (_41362_, _40131_, _40129_);
  nand _47316_ (_40132_, _39706_, _38191_);
  or _47317_ (_40133_, _40114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _47318_ (_40134_, _39737_, _39726_);
  not _47319_ (_40135_, _40134_);
  or _47320_ (_40136_, _40135_, _39757_);
  and _47321_ (_40137_, _40136_, _39758_);
  and _47322_ (_40138_, _40137_, _40133_);
  not _47323_ (_40139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _47324_ (_40140_, _40116_, _40139_);
  and _47325_ (_40141_, _40116_, _40139_);
  or _47326_ (_40142_, _40141_, _40140_);
  and _47327_ (_40143_, _40142_, _39761_);
  or _47328_ (_40144_, _40120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _47329_ (_40145_, _40120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _47330_ (_40146_, _40145_, _39806_);
  and _47331_ (_40147_, _40146_, _40144_);
  or _47332_ (_40148_, _40147_, _40143_);
  or _47333_ (_40149_, _40148_, _40138_);
  or _47334_ (_40150_, _40149_, _39706_);
  and _47335_ (_40151_, _40150_, _40132_);
  or _47336_ (_40152_, _40151_, _39750_);
  nand _47337_ (_40153_, _39750_, _40139_);
  and _47338_ (_40154_, _40153_, _42618_);
  and _47339_ (_41364_, _40154_, _40152_);
  nand _47340_ (_40155_, _39706_, _38184_);
  and _47341_ (_40156_, _39726_, _39716_);
  and _47342_ (_40157_, _40156_, _39723_);
  or _47343_ (_40158_, _40157_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47344_ (_40159_, _39727_, _39724_);
  nor _47345_ (_40160_, _40159_, _39806_);
  and _47346_ (_40161_, _40160_, _40158_);
  or _47347_ (_40162_, _40134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47348_ (_40163_, _39737_, _39727_);
  not _47349_ (_40164_, _40163_);
  and _47350_ (_40165_, _40164_, _39740_);
  and _47351_ (_40166_, _40165_, _40162_);
  and _47352_ (_40167_, _39726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47353_ (_40168_, _40167_, _39796_);
  or _47354_ (_40169_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47355_ (_40170_, _39796_, _39727_);
  nand _47356_ (_40171_, _40170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47357_ (_40172_, _40171_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47358_ (_40173_, _40172_, _40169_);
  or _47359_ (_40174_, _40173_, _40166_);
  or _47360_ (_40175_, _40174_, _40161_);
  or _47361_ (_40176_, _40175_, _39706_);
  and _47362_ (_40177_, _40176_, _40155_);
  or _47363_ (_40178_, _40177_, _39750_);
  or _47364_ (_40179_, _39751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47365_ (_40180_, _40179_, _42618_);
  and _47366_ (_41366_, _40180_, _40178_);
  nand _47367_ (_40181_, _39706_, _38177_);
  not _47368_ (_40182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47369_ (_40183_, _40163_, _39739_);
  nor _47370_ (_40184_, _40183_, _40182_);
  and _47371_ (_40185_, _40183_, _40182_);
  or _47372_ (_40186_, _40185_, _40184_);
  and _47373_ (_40187_, _40186_, _39758_);
  or _47374_ (_40188_, _40170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _47375_ (_40189_, _39797_);
  and _47376_ (_40190_, _40189_, _39761_);
  and _47377_ (_40191_, _40190_, _40188_);
  or _47378_ (_40192_, _40159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47379_ (_40193_, _39728_, _39724_);
  nor _47380_ (_40194_, _40193_, _39806_);
  and _47381_ (_40195_, _40194_, _40192_);
  or _47382_ (_40196_, _40195_, _40191_);
  or _47383_ (_40197_, _40196_, _40187_);
  or _47384_ (_40198_, _40197_, _39706_);
  and _47385_ (_40199_, _40198_, _40181_);
  or _47386_ (_40200_, _40199_, _39750_);
  nand _47387_ (_40201_, _39750_, _40182_);
  and _47388_ (_40202_, _40201_, _42618_);
  and _47389_ (_41368_, _40202_, _40200_);
  nand _47390_ (_40203_, _39706_, _38169_);
  or _47391_ (_40204_, _40193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47392_ (_40205_, _40157_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47393_ (_40206_, _40205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47394_ (_40207_, _40206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _47395_ (_40208_, _40207_, _39806_);
  and _47396_ (_40209_, _40208_, _40204_);
  and _47397_ (_40210_, _39737_, _39728_);
  nand _47398_ (_40211_, _40210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _47399_ (_40212_, _40210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47400_ (_40213_, _40212_, _39740_);
  and _47401_ (_40214_, _40213_, _40211_);
  and _47402_ (_40215_, _39797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _47403_ (_40216_, _40215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47404_ (_40217_, _40216_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47405_ (_40218_, _39797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _47406_ (_40219_, _40218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47407_ (_40220_, _40219_, _40217_);
  or _47408_ (_40221_, _40220_, _40214_);
  or _47409_ (_40222_, _40221_, _40209_);
  or _47410_ (_40223_, _40222_, _39706_);
  and _47411_ (_40224_, _40223_, _40203_);
  or _47412_ (_40225_, _40224_, _39750_);
  or _47413_ (_40226_, _39751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47414_ (_40227_, _40226_, _42618_);
  and _47415_ (_41370_, _40227_, _40225_);
  nand _47416_ (_40228_, _39706_, _38162_);
  not _47417_ (_40229_, _40207_);
  nor _47418_ (_40230_, _40229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47419_ (_40231_, _40229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _47420_ (_40232_, _40231_, _40230_);
  and _47421_ (_40233_, _40232_, _39707_);
  nor _47422_ (_40234_, _40211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _47423_ (_40235_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _47424_ (_40236_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47425_ (_40237_, _40236_, _39758_);
  and _47426_ (_40238_, _40237_, _40235_);
  not _47427_ (_40239_, _39798_);
  and _47428_ (_40240_, _40239_, _39761_);
  or _47429_ (_40241_, _40218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47430_ (_40242_, _40241_, _40240_);
  or _47431_ (_40243_, _40242_, _40238_);
  or _47432_ (_40244_, _40243_, _40233_);
  nor _47433_ (_40245_, _40244_, _39706_);
  nor _47434_ (_40246_, _40245_, _39780_);
  and _47435_ (_40247_, _40246_, _40228_);
  and _47436_ (_40248_, _39750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _47437_ (_40249_, _40248_, _40247_);
  and _47438_ (_41372_, _40249_, _42618_);
  or _47439_ (_40250_, _39790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _47440_ (_40251_, _40250_, _39758_);
  nor _47441_ (_40252_, _40251_, _39791_);
  or _47442_ (_40253_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _47443_ (_40254_, _39799_);
  and _47444_ (_40255_, _40254_, _39761_);
  and _47445_ (_40256_, _40255_, _40253_);
  or _47446_ (_40257_, _39730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _47447_ (_40258_, _39804_, _39806_);
  and _47448_ (_40259_, _40258_, _40257_);
  or _47449_ (_40260_, _40259_, _40256_);
  nor _47450_ (_40261_, _40260_, _40252_);
  nor _47451_ (_40262_, _40261_, _39706_);
  and _47452_ (_40263_, _39706_, _39933_);
  or _47453_ (_40264_, _40263_, _40262_);
  and _47454_ (_40265_, _40264_, _39751_);
  and _47455_ (_40266_, _39750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _47456_ (_40267_, _40266_, _40265_);
  and _47457_ (_41374_, _40267_, _42618_);
  nor _47458_ (_40268_, _39824_, _39756_);
  and _47459_ (_40269_, _39824_, _38204_);
  or _47460_ (_40270_, _40269_, _40268_);
  and _47461_ (_41376_, _40270_, _42618_);
  or _47462_ (_40271_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47463_ (_40272_, _40271_, _42618_);
  nand _47464_ (_40273_, _39824_, _38191_);
  and _47465_ (_41378_, _40273_, _40272_);
  or _47466_ (_40274_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _47467_ (_40275_, _40274_, _42618_);
  nand _47468_ (_40276_, _39824_, _38184_);
  and _47469_ (_41379_, _40276_, _40275_);
  or _47470_ (_40277_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _47471_ (_40278_, _40277_, _42618_);
  nand _47472_ (_40279_, _39824_, _38177_);
  and _47473_ (_41381_, _40279_, _40278_);
  or _47474_ (_40280_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _47475_ (_40281_, _40280_, _42618_);
  nand _47476_ (_40282_, _39824_, _38169_);
  and _47477_ (_41383_, _40282_, _40281_);
  or _47478_ (_40283_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _47479_ (_40284_, _40283_, _42618_);
  nand _47480_ (_40285_, _39824_, _38162_);
  and _47481_ (_41385_, _40285_, _40284_);
  or _47482_ (_40286_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _47483_ (_40287_, _40286_, _42618_);
  nand _47484_ (_40288_, _39824_, _38155_);
  and _47485_ (_41387_, _40288_, _40287_);
  not _47486_ (_40289_, _27542_);
  nor _47487_ (_40290_, _38794_, _27948_);
  nand _47488_ (_40291_, _40290_, _40289_);
  nor _47489_ (_40292_, _40291_, _28244_);
  and _47490_ (_40293_, _40292_, _38966_);
  and _47491_ (_40294_, _40293_, _31855_);
  nand _47492_ (_40295_, _40294_, _31757_);
  and _47493_ (_40296_, _38136_, _31855_);
  and _47494_ (_40297_, _40296_, _38989_);
  not _47495_ (_40298_, _40297_);
  or _47496_ (_40299_, _40294_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _47497_ (_40300_, _40299_, _40298_);
  and _47498_ (_40301_, _40300_, _40295_);
  nor _47499_ (_40302_, _40298_, _38225_);
  or _47500_ (_40303_, _40302_, _40301_);
  and _47501_ (_42556_, _40303_, _42618_);
  and _47502_ (_40304_, _39552_, _38813_);
  and _47503_ (_40305_, _40304_, _38973_);
  not _47504_ (_40306_, _40305_);
  and _47505_ (_40307_, _31790_, _27542_);
  and _47506_ (_40309_, _40307_, _38795_);
  and _47507_ (_40311_, _40309_, _38966_);
  and _47508_ (_40313_, _40311_, _31855_);
  or _47509_ (_40315_, _40313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _47510_ (_40317_, _40315_, _40306_);
  nand _47511_ (_40319_, _40313_, _31757_);
  and _47512_ (_40321_, _40319_, _40317_);
  nor _47513_ (_40323_, _40306_, _38225_);
  or _47514_ (_40325_, _40323_, _40321_);
  and _47515_ (_42559_, _40325_, _42618_);
  and _47516_ (_40328_, _40304_, _38140_);
  and _47517_ (_40330_, _40290_, _27542_);
  and _47518_ (_40332_, _40330_, _31779_);
  and _47519_ (_40334_, _40332_, _38934_);
  nand _47520_ (_40336_, _40334_, _27795_);
  and _47521_ (_40338_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _47522_ (_40340_, _40338_, _40328_);
  or _47523_ (_40342_, _27806_, _33837_);
  and _47524_ (_40344_, _40342_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _47525_ (_40346_, _40344_, _38740_);
  and _47526_ (_40348_, _40346_, _40334_);
  or _47527_ (_40350_, _40348_, _40340_);
  nand _47528_ (_40352_, _40328_, _38155_);
  and _47529_ (_40354_, _40352_, _42618_);
  and _47530_ (_42561_, _40354_, _40350_);
  not _47531_ (_40357_, _40328_);
  nor _47532_ (_40359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _47533_ (_40361_, _40359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _47534_ (_40362_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _47535_ (_40363_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _47536_ (_40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _47537_ (_40365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40364_);
  and _47538_ (_40366_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47539_ (_40367_, _40366_, _40365_);
  nor _47540_ (_40368_, _40367_, _40363_);
  or _47541_ (_40369_, _40368_, _40362_);
  and _47542_ (_40370_, _40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _47543_ (_40371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _47544_ (_40372_, _40371_, _40370_);
  nor _47545_ (_40373_, _40372_, _40363_);
  and _47546_ (_40374_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40364_);
  and _47547_ (_40375_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47548_ (_40376_, _40375_, _40374_);
  nand _47549_ (_40377_, _40376_, _40373_);
  or _47550_ (_40378_, _40377_, _40369_);
  and _47551_ (_40379_, _40378_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _47552_ (_40380_, _40379_, _40361_);
  and _47553_ (_40381_, _38140_, _31855_);
  and _47554_ (_40382_, _40381_, _40290_);
  or _47555_ (_40383_, _40382_, _40380_);
  and _47556_ (_40384_, _40383_, _40357_);
  nand _47557_ (_40385_, _40382_, _31757_);
  and _47558_ (_40386_, _40385_, _40384_);
  nor _47559_ (_40387_, _40357_, _38225_);
  or _47560_ (_40388_, _40387_, _40386_);
  and _47561_ (_42564_, _40388_, _42618_);
  and _47562_ (_40389_, _39587_, _31899_);
  nand _47563_ (_40390_, _40389_, _31757_);
  not _47564_ (_40391_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _47565_ (_40392_, _40391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _47566_ (_40393_, _40376_, _40363_);
  not _47567_ (_40394_, _40393_);
  or _47568_ (_40395_, _40394_, _40373_);
  or _47569_ (_40396_, _40395_, _40369_);
  and _47570_ (_40397_, _40396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _47571_ (_40398_, _40397_, _40392_);
  or _47572_ (_40399_, _40398_, _40389_);
  and _47573_ (_40400_, _40399_, _40357_);
  and _47574_ (_40401_, _40400_, _40390_);
  nor _47575_ (_40402_, _40357_, _38162_);
  or _47576_ (_40403_, _40402_, _40401_);
  and _47577_ (_42566_, _40403_, _42618_);
  not _47578_ (_40404_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _47579_ (_40405_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40404_);
  nand _47580_ (_40406_, _40368_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _47581_ (_40407_, _40393_, _40373_);
  or _47582_ (_40408_, _40407_, _40406_);
  and _47583_ (_40409_, _40408_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _47584_ (_40410_, _40409_, _40405_);
  and _47585_ (_40411_, _40290_, _38142_);
  or _47586_ (_40412_, _40411_, _40410_);
  and _47587_ (_40413_, _40412_, _40357_);
  nand _47588_ (_40414_, _40411_, _31757_);
  and _47589_ (_40415_, _40414_, _40413_);
  nor _47590_ (_40416_, _40357_, _38191_);
  or _47591_ (_40417_, _40416_, _40415_);
  and _47592_ (_42568_, _40417_, _42618_);
  and _47593_ (_40418_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _47594_ (_40419_, _40406_, _40395_);
  and _47595_ (_40420_, _40419_, _40418_);
  and _47596_ (_40421_, _40290_, _38272_);
  or _47597_ (_40422_, _40421_, _40420_);
  and _47598_ (_40423_, _40422_, _40357_);
  nand _47599_ (_40424_, _40421_, _31757_);
  and _47600_ (_40425_, _40424_, _40423_);
  nor _47601_ (_40426_, _40357_, _38177_);
  or _47602_ (_40427_, _40426_, _40425_);
  and _47603_ (_42570_, _40427_, _42618_);
  nand _47604_ (_40428_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _47605_ (_40429_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40364_);
  and _47606_ (_40430_, _40429_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _47607_ (_40431_, _40430_, _40428_);
  or _47608_ (_40432_, _40431_, _40363_);
  and _47609_ (_40433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _47610_ (_40434_, _40433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _47611_ (_40435_, _40434_);
  and _47612_ (_40436_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _47613_ (_40437_, _40436_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _47614_ (_40438_, _40437_);
  and _47615_ (_40439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _47616_ (_40440_, _40439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47617_ (_40441_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _47618_ (_40442_, _40441_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _47619_ (_40443_, _40442_, _40440_);
  and _47620_ (_40444_, _40443_, _40438_);
  and _47621_ (_40445_, _40444_, _40435_);
  not _47622_ (_40446_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _47623_ (_40447_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _47624_ (_40448_, _40447_, _40446_);
  nand _47625_ (_40449_, _40448_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _47626_ (_40450_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _47627_ (_40451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _47628_ (_40452_, _40451_, _40450_);
  and _47629_ (_40453_, _40452_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _47630_ (_40454_, _40453_);
  and _47631_ (_40455_, _40454_, _40449_);
  nand _47632_ (_40456_, _40455_, _40445_);
  and _47633_ (_40457_, _40456_, _40432_);
  and _47634_ (_40458_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _47635_ (_40459_, _40458_, _40364_);
  and _47636_ (_40460_, _40459_, _40457_);
  not _47637_ (_40461_, _40460_);
  not _47638_ (_40462_, _40459_);
  and _47639_ (_40463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40363_);
  not _47640_ (_40464_, _40463_);
  not _47641_ (_40465_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _47642_ (_40466_, _40448_, _40465_);
  not _47643_ (_40467_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _47644_ (_40468_, _40452_, _40467_);
  nor _47645_ (_40469_, _40468_, _40466_);
  not _47646_ (_40470_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _47647_ (_40471_, _40433_, _40470_);
  not _47648_ (_40472_, _40471_);
  and _47649_ (_40473_, _40472_, _40469_);
  nor _47650_ (_40474_, _40473_, _40464_);
  not _47651_ (_40475_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47652_ (_40476_, _40436_, _40475_);
  not _47653_ (_40477_, _40476_);
  not _47654_ (_40478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47655_ (_40479_, _40439_, _40478_);
  not _47656_ (_40480_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _47657_ (_40481_, _40441_, _40480_);
  nor _47658_ (_40482_, _40481_, _40479_);
  and _47659_ (_40483_, _40482_, _40477_);
  nor _47660_ (_40484_, _40483_, _40464_);
  nor _47661_ (_40485_, _40484_, _40474_);
  or _47662_ (_40486_, _40485_, _40462_);
  and _47663_ (_40487_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42618_);
  and _47664_ (_40488_, _40487_, _40486_);
  and _47665_ (_42605_, _40488_, _40461_);
  nor _47666_ (_40489_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _47667_ (_40490_, _40489_);
  not _47668_ (_40491_, _40457_);
  and _47669_ (_40492_, _40485_, _40491_);
  nor _47670_ (_40493_, _40492_, _40490_);
  nand _47671_ (_40494_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42618_);
  nor _47672_ (_42607_, _40494_, _40493_);
  and _47673_ (_40495_, _40455_, _40435_);
  nand _47674_ (_40496_, _40495_, _40457_);
  or _47675_ (_40497_, _40474_, _40457_);
  and _47676_ (_40498_, _40497_, _40459_);
  and _47677_ (_40499_, _40498_, _40496_);
  or _47678_ (_40500_, _40499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor _47679_ (_40501_, _40462_, _40457_);
  nand _47680_ (_40502_, _40501_, _40484_);
  or _47681_ (_40503_, _40461_, _40444_);
  and _47682_ (_40504_, _40503_, _42618_);
  and _47683_ (_40505_, _40504_, _40502_);
  and _47684_ (_42609_, _40505_, _40500_);
  and _47685_ (_40506_, _40496_, _40489_);
  or _47686_ (_40507_, _40506_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _47687_ (_40508_, _40489_, _40457_);
  not _47688_ (_40509_, _40508_);
  or _47689_ (_40510_, _40509_, _40444_);
  or _47690_ (_40511_, _40474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand _47691_ (_40512_, _40489_, _40484_);
  and _47692_ (_40513_, _40512_, _40511_);
  or _47693_ (_40514_, _40513_, _40457_);
  and _47694_ (_40515_, _40514_, _42618_);
  and _47695_ (_40516_, _40515_, _40510_);
  and _47696_ (_42611_, _40516_, _40507_);
  nand _47697_ (_40517_, _40492_, _40363_);
  nor _47698_ (_40518_, _40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _47699_ (_40519_, _40518_, _40458_);
  and _47700_ (_40520_, _40519_, _42618_);
  and _47701_ (_42613_, _40520_, _40517_);
  and _47702_ (_40521_, _40492_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _47703_ (_40522_, _40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _47704_ (_40523_, _40522_, _40518_);
  nor _47705_ (_40524_, _40523_, _40491_);
  or _47706_ (_40525_, _40524_, _40458_);
  or _47707_ (_40526_, _40525_, _40521_);
  not _47708_ (_40527_, _40458_);
  or _47709_ (_40528_, _40523_, _40527_);
  and _47710_ (_40529_, _40528_, _42618_);
  and _47711_ (_42615_, _40529_, _40526_);
  and _47712_ (_40530_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42618_);
  and _47713_ (_42616_, _40530_, _40458_);
  nor _47714_ (_42621_, _40359_, rst);
  and _47715_ (_42623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _42618_);
  nor _47716_ (_40531_, _40492_, _40458_);
  and _47717_ (_40532_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _47718_ (_40533_, _40532_, _40531_);
  and _47719_ (_00130_, _40533_, _42618_);
  and _47720_ (_40534_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _47721_ (_40535_, _40534_, _40531_);
  and _47722_ (_00132_, _40535_, _42618_);
  and _47723_ (_40536_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42618_);
  and _47724_ (_00134_, _40536_, _40458_);
  not _47725_ (_40537_, _40481_);
  nor _47726_ (_40538_, _40468_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _47727_ (_40539_, _40538_, _40466_);
  or _47728_ (_40540_, _40539_, _40471_);
  and _47729_ (_40541_, _40540_, _40537_);
  or _47730_ (_40542_, _40541_, _40479_);
  nor _47731_ (_40543_, _40485_, _40457_);
  and _47732_ (_40544_, _40543_, _40477_);
  and _47733_ (_40545_, _40544_, _40542_);
  not _47734_ (_40546_, _40442_);
  or _47735_ (_40547_, _40453_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _47736_ (_40548_, _40547_, _40449_);
  or _47737_ (_40549_, _40548_, _40434_);
  and _47738_ (_40550_, _40549_, _40546_);
  or _47739_ (_40551_, _40550_, _40440_);
  and _47740_ (_40552_, _40457_, _40438_);
  and _47741_ (_40553_, _40552_, _40551_);
  or _47742_ (_40554_, _40553_, _40458_);
  or _47743_ (_40555_, _40554_, _40545_);
  or _47744_ (_40556_, _40527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _47745_ (_40557_, _40556_, _42618_);
  and _47746_ (_00136_, _40557_, _40555_);
  not _47747_ (_40558_, _40440_);
  or _47748_ (_40559_, _40442_, _40434_);
  and _47749_ (_40560_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _47750_ (_40561_, _40560_, _40559_);
  and _47751_ (_40562_, _40561_, _40558_);
  and _47752_ (_40563_, _40562_, _40552_);
  nor _47753_ (_40564_, _40479_, _40476_);
  or _47754_ (_40565_, _40481_, _40471_);
  and _47755_ (_40566_, _40469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _47756_ (_40567_, _40566_, _40565_);
  and _47757_ (_40568_, _40567_, _40564_);
  and _47758_ (_40569_, _40568_, _40543_);
  or _47759_ (_40570_, _40569_, _40458_);
  or _47760_ (_40571_, _40570_, _40563_);
  or _47761_ (_40578_, _40527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _47762_ (_40579_, _40578_, _42618_);
  and _47763_ (_00138_, _40579_, _40571_);
  or _47764_ (_40590_, _40471_, _40464_);
  nor _47765_ (_40596_, _40590_, _40469_);
  nand _47766_ (_40599_, _40596_, _40483_);
  nor _47767_ (_40600_, _40599_, _40457_);
  not _47768_ (_40601_, _40455_);
  and _47769_ (_40602_, _40601_, _40445_);
  and _47770_ (_40603_, _40602_, _40432_);
  or _47771_ (_40604_, _40603_, _40458_);
  or _47772_ (_40605_, _40604_, _40600_);
  or _47773_ (_40606_, _40527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _47774_ (_40607_, _40606_, _42618_);
  and _47775_ (_00139_, _40607_, _40605_);
  and _47776_ (_40608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42618_);
  and _47777_ (_00141_, _40608_, _40458_);
  and _47778_ (_40609_, _40458_, _40364_);
  or _47779_ (_40610_, _40609_, _40493_);
  or _47780_ (_40611_, _40610_, _40501_);
  and _47781_ (_00143_, _40611_, _42618_);
  not _47782_ (_40617_, _40531_);
  and _47783_ (_40621_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _47784_ (_40622_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _47785_ (_40624_, _40453_, _40364_);
  or _47786_ (_40625_, _40624_, _40622_);
  nor _47787_ (_40631_, _40449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47788_ (_40634_, _40631_, _40434_);
  nand _47789_ (_40635_, _40634_, _40625_);
  or _47790_ (_40636_, _40435_, _40366_);
  and _47791_ (_40639_, _40636_, _40635_);
  or _47792_ (_40645_, _40639_, _40442_);
  or _47793_ (_40647_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40364_);
  or _47794_ (_40648_, _40647_, _40546_);
  and _47795_ (_40650_, _40648_, _40558_);
  and _47796_ (_40656_, _40650_, _40645_);
  and _47797_ (_40659_, _40440_, _40366_);
  or _47798_ (_40660_, _40659_, _40437_);
  or _47799_ (_40661_, _40660_, _40656_);
  or _47800_ (_40664_, _40647_, _40438_);
  and _47801_ (_40670_, _40664_, _40457_);
  and _47802_ (_40672_, _40670_, _40661_);
  and _47803_ (_40675_, _40468_, _40364_);
  or _47804_ (_40676_, _40675_, _40622_);
  and _47805_ (_40682_, _40466_, _40364_);
  nor _47806_ (_40684_, _40682_, _40471_);
  nand _47807_ (_40686_, _40684_, _40676_);
  or _47808_ (_40687_, _40472_, _40366_);
  and _47809_ (_40693_, _40687_, _40686_);
  or _47810_ (_40696_, _40693_, _40481_);
  not _47811_ (_40697_, _40479_);
  or _47812_ (_40699_, _40647_, _40537_);
  and _47813_ (_40705_, _40699_, _40697_);
  and _47814_ (_40708_, _40705_, _40696_);
  and _47815_ (_40709_, _40479_, _40366_);
  or _47816_ (_40710_, _40709_, _40476_);
  or _47817_ (_40713_, _40710_, _40708_);
  and _47818_ (_40719_, _40647_, _40543_);
  or _47819_ (_40721_, _40719_, _40544_);
  and _47820_ (_40722_, _40721_, _40713_);
  or _47821_ (_40725_, _40722_, _40672_);
  and _47822_ (_40731_, _40725_, _40527_);
  or _47823_ (_40733_, _40731_, _40621_);
  and _47824_ (_00145_, _40733_, _42618_);
  and _47825_ (_40735_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _47826_ (_40741_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40364_);
  and _47827_ (_40744_, _40741_, _40438_);
  or _47828_ (_40745_, _40744_, _40444_);
  or _47829_ (_40747_, _40624_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _47830_ (_40753_, _40747_, _40634_);
  nand _47831_ (_40756_, _40434_, _40375_);
  nand _47832_ (_40757_, _40756_, _40443_);
  or _47833_ (_40758_, _40757_, _40753_);
  and _47834_ (_40763_, _40758_, _40745_);
  and _47835_ (_40768_, _40437_, _40375_);
  or _47836_ (_40769_, _40768_, _40763_);
  and _47837_ (_40770_, _40769_, _40457_);
  and _47838_ (_40775_, _40482_, _40471_);
  or _47839_ (_40780_, _40775_, _40476_);
  and _47840_ (_40781_, _40780_, _40375_);
  or _47841_ (_40782_, _40675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _47842_ (_40786_, _40684_, _40482_);
  and _47843_ (_40792_, _40786_, _40782_);
  not _47844_ (_40793_, _40482_);
  and _47845_ (_40794_, _40741_, _40793_);
  or _47846_ (_40798_, _40794_, _40792_);
  and _47847_ (_40803_, _40798_, _40477_);
  or _47848_ (_40804_, _40803_, _40781_);
  and _47849_ (_40805_, _40804_, _40543_);
  or _47850_ (_40806_, _40805_, _40770_);
  and _47851_ (_40807_, _40806_, _40527_);
  or _47852_ (_40808_, _40807_, _40735_);
  and _47853_ (_00147_, _40808_, _42618_);
  and _47854_ (_40809_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not _47855_ (_40811_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _47856_ (_40812_, _40453_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47857_ (_40814_, _40812_, _40811_);
  nor _47858_ (_40815_, _40449_, _40364_);
  nor _47859_ (_40817_, _40815_, _40434_);
  nand _47860_ (_40818_, _40817_, _40814_);
  or _47861_ (_40820_, _40435_, _40365_);
  and _47862_ (_40821_, _40820_, _40818_);
  or _47863_ (_40823_, _40821_, _40442_);
  or _47864_ (_40824_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47865_ (_40826_, _40824_, _40546_);
  and _47866_ (_40827_, _40826_, _40558_);
  and _47867_ (_40829_, _40827_, _40823_);
  and _47868_ (_40830_, _40440_, _40365_);
  or _47869_ (_40832_, _40830_, _40437_);
  or _47870_ (_40833_, _40832_, _40829_);
  or _47871_ (_40835_, _40824_, _40438_);
  and _47872_ (_40836_, _40835_, _40457_);
  and _47873_ (_40838_, _40836_, _40833_);
  and _47874_ (_40839_, _40468_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47875_ (_40840_, _40839_, _40811_);
  and _47876_ (_40841_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47877_ (_40842_, _40841_, _40471_);
  nand _47878_ (_40843_, _40842_, _40840_);
  or _47879_ (_40844_, _40472_, _40365_);
  and _47880_ (_40845_, _40844_, _40843_);
  or _47881_ (_40846_, _40845_, _40481_);
  or _47882_ (_40847_, _40824_, _40537_);
  and _47883_ (_40848_, _40847_, _40697_);
  and _47884_ (_40849_, _40848_, _40846_);
  and _47885_ (_40850_, _40479_, _40365_);
  or _47886_ (_40851_, _40850_, _40476_);
  or _47887_ (_40852_, _40851_, _40849_);
  and _47888_ (_40853_, _40824_, _40543_);
  or _47889_ (_40854_, _40853_, _40544_);
  and _47890_ (_40855_, _40854_, _40852_);
  or _47891_ (_40856_, _40855_, _40838_);
  and _47892_ (_40857_, _40856_, _40527_);
  or _47893_ (_40858_, _40857_, _40809_);
  and _47894_ (_00149_, _40858_, _42618_);
  and _47895_ (_40859_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _47896_ (_40860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _47897_ (_40861_, _40860_, _40438_);
  or _47898_ (_40862_, _40861_, _40444_);
  or _47899_ (_40863_, _40812_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _47900_ (_40864_, _40863_, _40817_);
  nand _47901_ (_40865_, _40434_, _40374_);
  nand _47902_ (_40866_, _40865_, _40443_);
  or _47903_ (_40867_, _40866_, _40864_);
  and _47904_ (_40868_, _40867_, _40862_);
  and _47905_ (_40869_, _40437_, _40374_);
  or _47906_ (_40870_, _40869_, _40868_);
  and _47907_ (_40871_, _40870_, _40457_);
  and _47908_ (_40872_, _40780_, _40374_);
  or _47909_ (_40873_, _40839_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _47910_ (_40874_, _40842_, _40482_);
  and _47911_ (_40875_, _40874_, _40873_);
  and _47912_ (_40876_, _40860_, _40793_);
  or _47913_ (_40877_, _40876_, _40875_);
  and _47914_ (_40878_, _40877_, _40477_);
  or _47915_ (_40879_, _40878_, _40872_);
  and _47916_ (_40880_, _40879_, _40543_);
  or _47917_ (_40881_, _40880_, _40871_);
  and _47918_ (_40882_, _40881_, _40527_);
  or _47919_ (_40883_, _40882_, _40859_);
  and _47920_ (_00150_, _40883_, _42618_);
  or _47921_ (_40884_, _40490_, _40485_);
  and _47922_ (_40885_, _40884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _47923_ (_40886_, _40885_, _40508_);
  and _47924_ (_00152_, _40886_, _42618_);
  and _47925_ (_40887_, _40486_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _47926_ (_40888_, _40887_, _40460_);
  and _47927_ (_00154_, _40888_, _42618_);
  and _47928_ (_40889_, _40334_, _38813_);
  or _47929_ (_40890_, _40889_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _47930_ (_40891_, _40890_, _40357_);
  nand _47931_ (_40892_, _40889_, _31757_);
  and _47932_ (_40893_, _40892_, _40891_);
  nor _47933_ (_40894_, _40357_, _38203_);
  or _47934_ (_40895_, _40894_, _40893_);
  and _47935_ (_00156_, _40895_, _42618_);
  not _47936_ (_40896_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _47937_ (_40897_, _40334_, _33847_);
  nand _47938_ (_40898_, _40897_, _40896_);
  and _47939_ (_40899_, _40898_, _40357_);
  or _47940_ (_40900_, _40897_, _32410_);
  and _47941_ (_40901_, _40900_, _40899_);
  nor _47942_ (_40902_, _40357_, _38184_);
  or _47943_ (_40903_, _40902_, _40901_);
  and _47944_ (_00158_, _40903_, _42618_);
  nand _47945_ (_40904_, _40334_, _35338_);
  nor _47946_ (_40905_, _40904_, _31757_);
  and _47947_ (_40906_, _40904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or _47948_ (_40907_, _40906_, _40328_);
  or _47949_ (_40908_, _40907_, _40905_);
  nand _47950_ (_40909_, _40328_, _38169_);
  and _47951_ (_40910_, _40909_, _42618_);
  and _47952_ (_00160_, _40910_, _40908_);
  and _47953_ (_40911_, _40311_, _38813_);
  or _47954_ (_40912_, _40911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _47955_ (_40913_, _40912_, _40306_);
  nand _47956_ (_40914_, _40911_, _31757_);
  and _47957_ (_40915_, _40914_, _40913_);
  nor _47958_ (_40916_, _40306_, _38203_);
  or _47959_ (_40917_, _40916_, _40915_);
  and _47960_ (_00161_, _40917_, _42618_);
  and _47961_ (_40918_, _40311_, _33129_);
  or _47962_ (_40919_, _40918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _47963_ (_40920_, _40919_, _40306_);
  nand _47964_ (_40921_, _40918_, _31757_);
  and _47965_ (_40922_, _40921_, _40920_);
  nor _47966_ (_40923_, _40306_, _38191_);
  or _47967_ (_40924_, _40923_, _40922_);
  and _47968_ (_00163_, _40924_, _42618_);
  nand _47969_ (_40925_, _40311_, _39025_);
  and _47970_ (_40926_, _40925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _47971_ (_40927_, _40926_, _40305_);
  and _47972_ (_40928_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _47973_ (_40929_, _40928_, _33869_);
  and _47974_ (_40930_, _40929_, _40311_);
  or _47975_ (_40931_, _40930_, _40927_);
  nand _47976_ (_40932_, _40305_, _38184_);
  and _47977_ (_40933_, _40932_, _42618_);
  and _47978_ (_00165_, _40933_, _40931_);
  and _47979_ (_40934_, _40311_, _34576_);
  or _47980_ (_40935_, _40934_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _47981_ (_40936_, _40935_, _40306_);
  nand _47982_ (_40937_, _40934_, _31757_);
  and _47983_ (_40938_, _40937_, _40936_);
  nor _47984_ (_40939_, _40306_, _38177_);
  or _47985_ (_40940_, _40939_, _40938_);
  and _47986_ (_00167_, _40940_, _42618_);
  and _47987_ (_40941_, _40311_, _35338_);
  or _47988_ (_40942_, _40941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _47989_ (_40943_, _40942_, _40306_);
  nand _47990_ (_40944_, _40941_, _31757_);
  and _47991_ (_40945_, _40944_, _40943_);
  nor _47992_ (_40946_, _40306_, _38169_);
  or _47993_ (_40947_, _40946_, _40945_);
  and _47994_ (_00169_, _40947_, _42618_);
  and _47995_ (_40948_, _40311_, _36133_);
  or _47996_ (_40949_, _40948_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _47997_ (_40950_, _40949_, _40306_);
  nand _47998_ (_40951_, _40948_, _31757_);
  and _47999_ (_40952_, _40951_, _40950_);
  nor _48000_ (_40953_, _40306_, _38162_);
  or _48001_ (_40954_, _40953_, _40952_);
  and _48002_ (_00171_, _40954_, _42618_);
  and _48003_ (_40955_, _40311_, _36785_);
  or _48004_ (_40956_, _40955_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _48005_ (_40957_, _40956_, _40306_);
  nand _48006_ (_40958_, _40955_, _31757_);
  and _48007_ (_40959_, _40958_, _40957_);
  nor _48008_ (_40960_, _40306_, _38155_);
  or _48009_ (_40961_, _40960_, _40959_);
  and _48010_ (_00173_, _40961_, _42618_);
  and _48011_ (_40962_, _40293_, _38813_);
  nand _48012_ (_40963_, _40962_, _31757_);
  or _48013_ (_40964_, _40962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _48014_ (_40965_, _40964_, _40298_);
  and _48015_ (_40966_, _40965_, _40963_);
  nor _48016_ (_40967_, _40298_, _38203_);
  or _48017_ (_40968_, _40967_, _40966_);
  and _48018_ (_00174_, _40968_, _42618_);
  and _48019_ (_40969_, _40293_, _33129_);
  nand _48020_ (_40970_, _40969_, _31757_);
  or _48021_ (_40971_, _40969_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _48022_ (_40972_, _40971_, _40298_);
  and _48023_ (_40973_, _40972_, _40970_);
  nor _48024_ (_40974_, _40298_, _38191_);
  or _48025_ (_40975_, _40974_, _40973_);
  and _48026_ (_00176_, _40975_, _42618_);
  and _48027_ (_40976_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _48028_ (_40977_, _40976_, _33869_);
  and _48029_ (_40978_, _40977_, _40293_);
  nand _48030_ (_40979_, _40293_, _39025_);
  and _48031_ (_40980_, _40979_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _48032_ (_40981_, _40980_, _40297_);
  or _48033_ (_40982_, _40981_, _40978_);
  nand _48034_ (_40983_, _40297_, _38184_);
  and _48035_ (_40984_, _40983_, _42618_);
  and _48036_ (_00178_, _40984_, _40982_);
  and _48037_ (_40985_, _40293_, _34576_);
  nand _48038_ (_40986_, _40985_, _31757_);
  or _48039_ (_40987_, _40985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _48040_ (_40988_, _40987_, _40986_);
  or _48041_ (_40989_, _40988_, _40297_);
  nand _48042_ (_40990_, _40297_, _38177_);
  and _48043_ (_40991_, _40990_, _42618_);
  and _48044_ (_00180_, _40991_, _40989_);
  and _48045_ (_40992_, _40293_, _35338_);
  nand _48046_ (_40993_, _40992_, _31757_);
  or _48047_ (_40994_, _40992_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _48048_ (_40995_, _40994_, _40298_);
  and _48049_ (_40996_, _40995_, _40993_);
  nor _48050_ (_40997_, _40298_, _38169_);
  or _48051_ (_40998_, _40997_, _40996_);
  and _48052_ (_00182_, _40998_, _42618_);
  and _48053_ (_40999_, _40293_, _36133_);
  nand _48054_ (_41000_, _40999_, _31757_);
  or _48055_ (_41001_, _40999_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _48056_ (_41002_, _41001_, _41000_);
  or _48057_ (_41003_, _41002_, _40297_);
  nand _48058_ (_41004_, _40297_, _38162_);
  and _48059_ (_41005_, _41004_, _42618_);
  and _48060_ (_00184_, _41005_, _41003_);
  and _48061_ (_41006_, _40293_, _36785_);
  nand _48062_ (_41007_, _41006_, _31757_);
  or _48063_ (_41008_, _41006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _48064_ (_41009_, _41008_, _41007_);
  or _48065_ (_41010_, _41009_, _40297_);
  nand _48066_ (_41011_, _40297_, _38155_);
  and _48067_ (_41012_, _41011_, _42618_);
  and _48068_ (_00185_, _41012_, _41010_);
  and _48069_ (_41013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _48070_ (_41014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _48071_ (_41015_, _40359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _48072_ (_41016_, _41015_, _41014_);
  not _48073_ (_41017_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _48074_ (_41018_, _41017_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _48075_ (_41019_, _41018_, _41016_);
  nor _48076_ (_41020_, _41019_, _41013_);
  or _48077_ (_41021_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _48078_ (_41022_, _41021_, _42618_);
  nor _48079_ (_00545_, _41022_, _41020_);
  nor _48080_ (_41023_, _41020_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _48081_ (_41024_, _41023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _48082_ (_41025_, _41023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _48083_ (_41026_, _41025_, _42618_);
  and _48084_ (_00548_, _41026_, _41024_);
  not _48085_ (_41027_, rxd_i);
  and _48086_ (_41028_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _41027_);
  nor _48087_ (_41029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _48088_ (_41030_, _41029_);
  and _48089_ (_41031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _48090_ (_41032_, _41031_, _41030_);
  and _48091_ (_41033_, _41032_, _41028_);
  not _48092_ (_41034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _48093_ (_41035_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _41034_);
  and _48094_ (_41036_, _41035_, _41029_);
  or _48095_ (_41037_, _41036_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or _48096_ (_41038_, _41037_, _41033_);
  and _48097_ (_41039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _42618_);
  and _48098_ (_00551_, _41039_, _41038_);
  and _48099_ (_41040_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _48100_ (_41041_, _41040_, _41030_);
  not _48101_ (_41042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _48102_ (_41043_, _41029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48103_ (_41044_, _41043_, _41042_);
  nor _48104_ (_41045_, _41044_, _41041_);
  not _48105_ (_41046_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _48106_ (_41047_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _41046_);
  not _48107_ (_41048_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _48108_ (_41049_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _41048_);
  and _48109_ (_41050_, _41049_, _41047_);
  not _48110_ (_41051_, _41050_);
  or _48111_ (_41052_, _41051_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and _48112_ (_41053_, _41050_, _41041_);
  and _48113_ (_41054_, _41041_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48114_ (_41055_, _41054_, _41053_);
  and _48115_ (_41056_, _41055_, _41052_);
  or _48116_ (_41057_, _41056_, _41045_);
  not _48117_ (_41058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand _48118_ (_41059_, _41029_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor _48119_ (_41060_, _41059_, _41058_);
  not _48120_ (_41061_, _41060_);
  or _48121_ (_41062_, _41061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _48122_ (_41063_, _41062_, _41057_);
  nand _48123_ (_00554_, _41063_, _41039_);
  not _48124_ (_41064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _48125_ (_41065_, _41041_);
  nor _48126_ (_41066_, _41042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _48127_ (_41067_, _41066_);
  not _48128_ (_41068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48129_ (_41069_, _41029_, _41068_);
  and _48130_ (_41070_, _41069_, _41067_);
  and _48131_ (_41071_, _41070_, _41065_);
  nor _48132_ (_41072_, _41071_, _41064_);
  and _48133_ (_41073_, _41071_, rxd_i);
  or _48134_ (_41074_, _41073_, rst);
  or _48135_ (_00556_, _41074_, _41072_);
  nor _48136_ (_41075_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48137_ (_41076_, _41075_, _41047_);
  and _48138_ (_41077_, _41076_, _41054_);
  nand _48139_ (_41078_, _41077_, _41027_);
  or _48140_ (_41079_, _41077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _48141_ (_41080_, _41079_, _42618_);
  and _48142_ (_00559_, _41080_, _41078_);
  and _48143_ (_41081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48144_ (_41082_, _41081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _48145_ (_41083_, _41082_, _41046_);
  and _48146_ (_41084_, _41083_, _41054_);
  and _48147_ (_41085_, _41032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48148_ (_41086_, _41085_, _41054_);
  nor _48149_ (_41087_, _41082_, _41065_);
  or _48150_ (_41088_, _41087_, _41086_);
  and _48151_ (_41089_, _41088_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _48152_ (_41090_, _41089_, _41084_);
  and _48153_ (_00562_, _41090_, _42618_);
  and _48154_ (_41091_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _42618_);
  nand _48155_ (_41092_, _41091_, _41068_);
  nand _48156_ (_41093_, _41039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _48157_ (_00564_, _41093_, _41092_);
  and _48158_ (_41094_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41068_);
  not _48159_ (_41095_, _41032_);
  nand _48160_ (_41096_, _41036_, _41058_);
  and _48161_ (_41097_, _41096_, _41095_);
  and _48162_ (_41098_, _41097_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _48163_ (_41099_, _41098_, _41041_);
  or _48164_ (_41100_, _41050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor _48165_ (_41101_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _48166_ (_41102_, _41101_, _41053_);
  and _48167_ (_41103_, _41102_, _41100_);
  and _48168_ (_41104_, _41103_, _41099_);
  or _48169_ (_41105_, _41104_, _41060_);
  nand _48170_ (_41106_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _48171_ (_41107_, _41106_, _41041_);
  or _48172_ (_41108_, _41107_, _41051_);
  and _48173_ (_41109_, _41108_, _41061_);
  or _48174_ (_41110_, _41109_, rxd_i);
  and _48175_ (_41111_, _41110_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48176_ (_41112_, _41111_, _41105_);
  or _48177_ (_41113_, _41112_, _41094_);
  and _48178_ (_00567_, _41113_, _42618_);
  and _48179_ (_41114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _48180_ (_41115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _48181_ (_41116_, _41015_, _41115_);
  or _48182_ (_41117_, _41116_, _41018_);
  nor _48183_ (_41118_, _41117_, _41114_);
  or _48184_ (_41119_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _48185_ (_41120_, _41119_, _42618_);
  nor _48186_ (_00570_, _41120_, _41118_);
  nor _48187_ (_41121_, _41118_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _48188_ (_41122_, _41121_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _48189_ (_41123_, _41121_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _48190_ (_41124_, _41123_, _42618_);
  and _48191_ (_00572_, _41124_, _41122_);
  not _48192_ (_41125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  nor _48193_ (_41126_, _31834_, _27948_);
  and _48194_ (_41127_, _41126_, _33118_);
  and _48195_ (_41128_, _41127_, _31212_);
  and _48196_ (_41129_, _41128_, _38957_);
  and _48197_ (_41130_, _41129_, _42618_);
  nand _48198_ (_41131_, _41130_, _41125_);
  nor _48199_ (_41132_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not _48200_ (_41133_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _48201_ (_41134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _48202_ (_41135_, _41134_, _41133_);
  and _48203_ (_41136_, _41135_, _41132_);
  not _48204_ (_41137_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _48205_ (_41138_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _48206_ (_41139_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _48207_ (_41140_, _41139_, _41138_);
  and _48208_ (_41141_, _41140_, _41137_);
  and _48209_ (_41142_, _41141_, _41136_);
  not _48210_ (_41143_, _41142_);
  or _48211_ (_41144_, _41143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  or _48212_ (_41145_, _41142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not _48213_ (_41146_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _48214_ (_41147_, _41059_, _41146_);
  and _48215_ (_41148_, _41147_, _41145_);
  and _48216_ (_41149_, _41148_, _41144_);
  nor _48217_ (_41150_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _48218_ (_41151_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _48219_ (_41152_, _41151_, _41150_);
  and _48220_ (_41153_, _41030_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _48221_ (_41154_, _41153_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _48222_ (_41155_, _41154_, _41152_);
  not _48223_ (_41156_, _41155_);
  or _48224_ (_41157_, _41156_, _41145_);
  and _48225_ (_41158_, _41152_, _41153_);
  or _48226_ (_41159_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _41146_);
  nor _48227_ (_41160_, _41159_, _41158_);
  nor _48228_ (_41161_, _41160_, _41147_);
  and _48229_ (_41162_, _41161_, _41157_);
  nor _48230_ (_41163_, _41162_, _41149_);
  nor _48231_ (_41164_, _41129_, rst);
  nand _48232_ (_41165_, _41164_, _41163_);
  and _48233_ (_00575_, _41165_, _41131_);
  nor _48234_ (_41166_, _41143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _48235_ (_41167_, _41158_, _41166_);
  and _48236_ (_41168_, _41147_, _41142_);
  or _48237_ (_41169_, _41146_, rst);
  nor _48238_ (_41170_, _41169_, _41168_);
  and _48239_ (_41171_, _41170_, _41167_);
  or _48240_ (_00578_, _41171_, _41130_);
  or _48241_ (_41172_, _41156_, _41166_);
  or _48242_ (_41173_, _41158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _48243_ (_41174_, _41059_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _48244_ (_41175_, _41174_, _41173_);
  and _48245_ (_41176_, _41175_, _41172_);
  or _48246_ (_41177_, _41176_, _41168_);
  and _48247_ (_00580_, _41177_, _41164_);
  and _48248_ (_41178_, _41154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _48249_ (_41179_, _41178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _48250_ (_41180_, _41179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nand _48251_ (_41181_, _41180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or _48252_ (_41182_, _41180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _48253_ (_41183_, _41182_, _41181_);
  and _48254_ (_00583_, _41183_, _41164_);
  nor _48255_ (_41184_, _41155_, _41147_);
  and _48256_ (_41185_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _48257_ (_41186_, _41185_, _41164_);
  and _48258_ (_41187_, _41130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _48259_ (_00586_, _41187_, _41186_);
  and _48260_ (_41188_, _40296_, _38140_);
  or _48261_ (_41189_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _48262_ (_41190_, _41189_, _42618_);
  nand _48263_ (_41191_, _41188_, _38225_);
  and _48264_ (_00588_, _41191_, _41190_);
  and _48265_ (_41192_, _40292_, _38934_);
  and _48266_ (_41193_, _41192_, _31855_);
  nand _48267_ (_41194_, _41193_, _31757_);
  and _48268_ (_41195_, _40304_, _38957_);
  not _48269_ (_41196_, _41195_);
  or _48270_ (_41197_, _41193_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _48271_ (_41198_, _41197_, _41196_);
  and _48272_ (_41199_, _41198_, _41194_);
  nor _48273_ (_41200_, _41196_, _38225_);
  or _48274_ (_41201_, _41200_, _41199_);
  and _48275_ (_00591_, _41201_, _42618_);
  nor _48276_ (_41202_, _41060_, _41053_);
  not _48277_ (_41203_, _41202_);
  nor _48278_ (_41204_, _41097_, _41041_);
  nor _48279_ (_41205_, _41204_, _41203_);
  nor _48280_ (_41206_, _41205_, _41068_);
  or _48281_ (_41207_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _48282_ (_41208_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _41068_);
  or _48283_ (_41209_, _41208_, _41202_);
  and _48284_ (_41210_, _41209_, _42618_);
  and _48285_ (_01206_, _41210_, _41207_);
  or _48286_ (_41211_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _48287_ (_41212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _41068_);
  or _48288_ (_41213_, _41212_, _41202_);
  and _48289_ (_41214_, _41213_, _42618_);
  and _48290_ (_01208_, _41214_, _41211_);
  or _48291_ (_41215_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _48292_ (_41216_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41068_);
  or _48293_ (_41217_, _41216_, _41202_);
  and _48294_ (_41218_, _41217_, _42618_);
  and _48295_ (_01210_, _41218_, _41215_);
  or _48296_ (_41219_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _48297_ (_41220_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41068_);
  or _48298_ (_41221_, _41220_, _41202_);
  and _48299_ (_41222_, _41221_, _42618_);
  and _48300_ (_01212_, _41222_, _41219_);
  or _48301_ (_41223_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _48302_ (_41224_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41068_);
  or _48303_ (_41225_, _41224_, _41202_);
  and _48304_ (_41226_, _41225_, _42618_);
  and _48305_ (_01214_, _41226_, _41223_);
  or _48306_ (_41227_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _48307_ (_41228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41068_);
  or _48308_ (_41229_, _41228_, _41202_);
  and _48309_ (_41230_, _41229_, _42618_);
  and _48310_ (_01216_, _41230_, _41227_);
  or _48311_ (_41231_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _48312_ (_41232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41068_);
  or _48313_ (_41233_, _41232_, _41202_);
  and _48314_ (_41234_, _41233_, _42618_);
  and _48315_ (_01218_, _41234_, _41231_);
  or _48316_ (_41235_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _48317_ (_41236_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _41068_);
  or _48318_ (_41237_, _41236_, _41202_);
  and _48319_ (_41238_, _41237_, _42618_);
  and _48320_ (_01220_, _41238_, _41235_);
  nor _48321_ (_41239_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _48322_ (_41240_, _41239_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _48323_ (_41241_, _41051_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or _48324_ (_41242_, _41050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _48325_ (_41243_, _41242_, _41041_);
  and _48326_ (_41244_, _41243_, _41241_);
  or _48327_ (_41245_, _41032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _48328_ (_41246_, _41245_, _41096_);
  and _48329_ (_41247_, _41246_, _41065_);
  or _48330_ (_41248_, _41247_, _41244_);
  or _48331_ (_41249_, _41248_, _41060_);
  or _48332_ (_41250_, _41061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _48333_ (_41251_, _41250_, _41039_);
  and _48334_ (_41252_, _41251_, _41249_);
  or _48335_ (_01221_, _41252_, _41240_);
  and _48336_ (_41253_, _41050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _48337_ (_41254_, _41253_, _41097_);
  or _48338_ (_41255_, _41254_, _41205_);
  and _48339_ (_41256_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _48340_ (_41257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _41068_);
  nand _48341_ (_41258_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48342_ (_41259_, _41258_, _41202_);
  or _48343_ (_41260_, _41259_, _41257_);
  or _48344_ (_41261_, _41260_, _41256_);
  and _48345_ (_01223_, _41261_, _42618_);
  not _48346_ (_41262_, _41206_);
  and _48347_ (_41263_, _41262_, _41091_);
  or _48348_ (_41264_, _41254_, _41203_);
  and _48349_ (_41265_, _41039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _48350_ (_41266_, _41265_, _41264_);
  or _48351_ (_01225_, _41266_, _41263_);
  or _48352_ (_41267_, _41084_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _48353_ (_41268_, _41084_, _41027_);
  and _48354_ (_41269_, _41268_, _42618_);
  and _48355_ (_01227_, _41269_, _41267_);
  or _48356_ (_41270_, _41086_, _41048_);
  or _48357_ (_41271_, _41054_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48358_ (_41272_, _41271_, _42618_);
  and _48359_ (_01229_, _41272_, _41270_);
  and _48360_ (_41273_, _41086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _48361_ (_41274_, _41075_, _41081_);
  and _48362_ (_41275_, _41274_, _41054_);
  or _48363_ (_41276_, _41275_, _41273_);
  and _48364_ (_01231_, _41276_, _42618_);
  and _48365_ (_41277_, _41088_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _48366_ (_41278_, _41081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48367_ (_41279_, _41278_, _41087_);
  or _48368_ (_41280_, _41279_, _41277_);
  and _48369_ (_01233_, _41280_, _42618_);
  and _48370_ (_41281_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41068_);
  and _48371_ (_41282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48372_ (_41283_, _41282_, _41281_);
  and _48373_ (_01235_, _41283_, _42618_);
  and _48374_ (_41284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41068_);
  and _48375_ (_41285_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48376_ (_41286_, _41285_, _41284_);
  and _48377_ (_01237_, _41286_, _42618_);
  and _48378_ (_41287_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41068_);
  and _48379_ (_41288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48380_ (_41289_, _41288_, _41287_);
  and _48381_ (_01239_, _41289_, _42618_);
  and _48382_ (_41290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41068_);
  and _48383_ (_41291_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48384_ (_41292_, _41291_, _41290_);
  and _48385_ (_01241_, _41292_, _42618_);
  and _48386_ (_41293_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41068_);
  and _48387_ (_41294_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48388_ (_41295_, _41294_, _41293_);
  and _48389_ (_01243_, _41295_, _42618_);
  and _48390_ (_41296_, _41039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _48391_ (_01245_, _41296_, _41240_);
  and _48392_ (_41297_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48393_ (_41298_, _41297_, _41257_);
  and _48394_ (_01247_, _41298_, _42618_);
  nor _48395_ (_41299_, _41154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _48396_ (_41300_, _41299_, _41178_);
  and _48397_ (_01249_, _41300_, _41164_);
  nor _48398_ (_41301_, _41178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _48399_ (_41302_, _41301_, _41179_);
  and _48400_ (_01251_, _41302_, _41164_);
  nor _48401_ (_41303_, _41179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _48402_ (_41304_, _41303_, _41180_);
  and _48403_ (_01253_, _41304_, _41164_);
  and _48404_ (_41305_, _41142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _48405_ (_41306_, _41305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _48406_ (_41307_, _41306_, _41147_);
  or _48407_ (_41308_, _41155_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _48408_ (_41309_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _48409_ (_41310_, _41309_, _41308_);
  nor _48410_ (_41311_, _41310_, _41307_);
  nor _48411_ (_41312_, _41311_, _41129_);
  nor _48412_ (_41313_, _41030_, _38203_);
  and _48413_ (_41314_, _41313_, _41129_);
  or _48414_ (_41315_, _41314_, _41312_);
  and _48415_ (_01255_, _41315_, _42618_);
  not _48416_ (_41316_, _41184_);
  and _48417_ (_41317_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _48418_ (_41318_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _48419_ (_41319_, _41318_, _41317_);
  and _48420_ (_41320_, _41319_, _41164_);
  nand _48421_ (_41321_, _41029_, _38191_);
  nand _48422_ (_41322_, _41030_, _38203_);
  and _48423_ (_41324_, _41322_, _41130_);
  and _48424_ (_41326_, _41324_, _41321_);
  or _48425_ (_01256_, _41326_, _41320_);
  nor _48426_ (_41329_, _41184_, _41137_);
  and _48427_ (_41331_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or _48428_ (_41333_, _41331_, _41329_);
  and _48429_ (_41335_, _41333_, _41164_);
  nand _48430_ (_41337_, _41029_, _38184_);
  nand _48431_ (_41339_, _41030_, _38191_);
  and _48432_ (_41341_, _41339_, _41130_);
  and _48433_ (_41343_, _41341_, _41337_);
  or _48434_ (_01258_, _41343_, _41335_);
  nand _48435_ (_41346_, _41184_, _41137_);
  or _48436_ (_41348_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _48437_ (_41350_, _41348_, _41346_);
  and _48438_ (_41352_, _41350_, _41164_);
  nand _48439_ (_41354_, _41030_, _38184_);
  nand _48440_ (_41356_, _41029_, _38177_);
  and _48441_ (_41358_, _41356_, _41130_);
  and _48442_ (_41360_, _41358_, _41354_);
  or _48443_ (_01260_, _41360_, _41352_);
  nand _48444_ (_41363_, _41184_, _41133_);
  or _48445_ (_41365_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _48446_ (_41367_, _41365_, _41363_);
  and _48447_ (_41369_, _41367_, _41164_);
  nand _48448_ (_41371_, _41030_, _38177_);
  nand _48449_ (_41373_, _41029_, _38169_);
  and _48450_ (_41375_, _41373_, _41130_);
  and _48451_ (_41377_, _41375_, _41371_);
  or _48452_ (_01262_, _41377_, _41369_);
  or _48453_ (_41380_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _48454_ (_41382_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _48455_ (_41384_, _41382_, _41380_);
  and _48456_ (_41386_, _41384_, _41164_);
  nand _48457_ (_41388_, _41029_, _38162_);
  nand _48458_ (_41389_, _41030_, _38169_);
  and _48459_ (_41390_, _41389_, _41130_);
  and _48460_ (_41391_, _41390_, _41388_);
  or _48461_ (_01264_, _41391_, _41386_);
  or _48462_ (_41392_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or _48463_ (_41393_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _48464_ (_41394_, _41393_, _41392_);
  and _48465_ (_41395_, _41394_, _41164_);
  nand _48466_ (_41396_, _41029_, _38155_);
  nand _48467_ (_41397_, _41030_, _38162_);
  and _48468_ (_41398_, _41397_, _41130_);
  and _48469_ (_41399_, _41398_, _41396_);
  or _48470_ (_01266_, _41399_, _41395_);
  or _48471_ (_41400_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _48472_ (_41401_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _48473_ (_41402_, _41401_, _41400_);
  and _48474_ (_41403_, _41402_, _41164_);
  nand _48475_ (_41404_, _41029_, _38225_);
  nand _48476_ (_41405_, _41030_, _38155_);
  and _48477_ (_41406_, _41405_, _41130_);
  and _48478_ (_41407_, _41406_, _41404_);
  or _48479_ (_01268_, _41407_, _41403_);
  and _48480_ (_41408_, _41129_, _41030_);
  nand _48481_ (_41409_, _41408_, _38225_);
  and _48482_ (_41410_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _48483_ (_41411_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _48484_ (_41412_, _41411_, _41410_);
  or _48485_ (_41413_, _41412_, _41129_);
  and _48486_ (_41414_, _41413_, _42618_);
  and _48487_ (_01270_, _41414_, _41409_);
  or _48488_ (_41415_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _48489_ (_41416_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _48490_ (_41417_, _41416_, _41415_);
  and _48491_ (_41418_, _41417_, _41164_);
  or _48492_ (_41419_, _41017_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _48493_ (_41420_, _41419_, _41030_);
  and _48494_ (_41421_, _41420_, _41130_);
  or _48495_ (_01272_, _41421_, _41418_);
  nand _48496_ (_41422_, _41188_, _38203_);
  or _48497_ (_41423_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _48498_ (_41424_, _41423_, _42618_);
  and _48499_ (_01274_, _41424_, _41422_);
  or _48500_ (_41425_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _48501_ (_41426_, _41425_, _42618_);
  nand _48502_ (_41427_, _41188_, _38191_);
  and _48503_ (_01276_, _41427_, _41426_);
  or _48504_ (_41428_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _48505_ (_41429_, _41428_, _42618_);
  nand _48506_ (_41430_, _41188_, _38184_);
  and _48507_ (_01278_, _41430_, _41429_);
  or _48508_ (_41431_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _48509_ (_41432_, _41431_, _42618_);
  nand _48510_ (_41433_, _41188_, _38177_);
  and _48511_ (_01280_, _41433_, _41432_);
  or _48512_ (_41434_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _48513_ (_41435_, _41434_, _42618_);
  nand _48514_ (_41436_, _41188_, _38169_);
  and _48515_ (_01282_, _41436_, _41435_);
  or _48516_ (_41437_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _48517_ (_41438_, _41437_, _42618_);
  nand _48518_ (_41439_, _41188_, _38162_);
  and _48519_ (_01284_, _41439_, _41438_);
  or _48520_ (_41440_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _48521_ (_41441_, _41440_, _42618_);
  nand _48522_ (_41442_, _41188_, _38155_);
  and _48523_ (_01286_, _41442_, _41441_);
  not _48524_ (_41443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _48525_ (_41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41443_);
  or _48526_ (_41445_, _41444_, _41029_);
  nor _48527_ (_41446_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48528_ (_41447_, _41446_, _41445_);
  or _48529_ (_41448_, _41447_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _48530_ (_41449_, _41448_, _41192_);
  or _48531_ (_41450_, _38813_, _41034_);
  nand _48532_ (_41451_, _41450_, _41192_);
  or _48533_ (_41452_, _41451_, _38814_);
  and _48534_ (_41453_, _41452_, _41449_);
  or _48535_ (_41454_, _41453_, _41195_);
  nand _48536_ (_41455_, _41195_, _38203_);
  and _48537_ (_41456_, _41455_, _42618_);
  and _48538_ (_01288_, _41456_, _41454_);
  or _48539_ (_41457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _48540_ (_41458_, _41457_, _41192_);
  nand _48541_ (_41459_, _38863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _48542_ (_41460_, _41459_, _41192_);
  or _48543_ (_41461_, _41460_, _38864_);
  and _48544_ (_41462_, _41461_, _41458_);
  or _48545_ (_41463_, _41462_, _41195_);
  nand _48546_ (_41464_, _41195_, _38191_);
  and _48547_ (_41465_, _41464_, _42618_);
  and _48548_ (_01290_, _41465_, _41463_);
  not _48549_ (_41466_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _48550_ (_41467_, _41043_, _41466_);
  and _48551_ (_41468_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _48552_ (_41469_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _48553_ (_41470_, _41467_, _41469_);
  or _48554_ (_41471_, _41470_, _41468_);
  or _48555_ (_41472_, _41471_, _41192_);
  or _48556_ (_41473_, _33847_, _41469_);
  nand _48557_ (_41474_, _41473_, _41192_);
  or _48558_ (_41475_, _41474_, _33869_);
  and _48559_ (_41476_, _41475_, _41472_);
  or _48560_ (_41477_, _41476_, _41195_);
  nand _48561_ (_41478_, _41195_, _38184_);
  and _48562_ (_41479_, _41478_, _42618_);
  and _48563_ (_01291_, _41479_, _41477_);
  and _48564_ (_41480_, _41192_, _34576_);
  nand _48565_ (_41481_, _41480_, _31757_);
  or _48566_ (_41482_, _41480_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _48567_ (_41483_, _41482_, _41196_);
  and _48568_ (_41484_, _41483_, _41481_);
  nor _48569_ (_41485_, _41196_, _38177_);
  or _48570_ (_41486_, _41485_, _41484_);
  and _48571_ (_01293_, _41486_, _42618_);
  and _48572_ (_41487_, _41192_, _35338_);
  nand _48573_ (_41488_, _41487_, _31757_);
  or _48574_ (_41489_, _41487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _48575_ (_41490_, _41489_, _41196_);
  and _48576_ (_41491_, _41490_, _41488_);
  nor _48577_ (_41492_, _41196_, _38169_);
  or _48578_ (_41493_, _41492_, _41491_);
  and _48579_ (_01295_, _41493_, _42618_);
  and _48580_ (_41494_, _41192_, _36133_);
  nand _48581_ (_41495_, _41494_, _31757_);
  or _48582_ (_41496_, _41494_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _48583_ (_41497_, _41496_, _41196_);
  and _48584_ (_41498_, _41497_, _41495_);
  nor _48585_ (_41499_, _41196_, _38162_);
  or _48586_ (_41500_, _41499_, _41498_);
  and _48587_ (_01297_, _41500_, _42618_);
  and _48588_ (_41501_, _41192_, _36785_);
  nand _48589_ (_41502_, _41501_, _31757_);
  or _48590_ (_41503_, _41501_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _48591_ (_41504_, _41503_, _41196_);
  and _48592_ (_41505_, _41504_, _41502_);
  nor _48593_ (_41506_, _41196_, _38155_);
  or _48594_ (_41507_, _41506_, _41505_);
  and _48595_ (_01299_, _41507_, _42618_);
  and _48596_ (_01626_, t2_i, _42618_);
  nor _48597_ (_41508_, t2_i, rst);
  and _48598_ (_01628_, _41508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand _48599_ (_41509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _42618_);
  nor _48600_ (_01631_, _41509_, t2ex_i);
  and _48601_ (_01634_, t2ex_i, _42618_);
  and _48602_ (_41510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _48603_ (_41511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _48604_ (_41512_, _41511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _48605_ (_41513_, _41512_, _41510_);
  not _48606_ (_41514_, _41513_);
  and _48607_ (_41515_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _48608_ (_41516_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor _48609_ (_41517_, _41516_, _41515_);
  and _48610_ (_41518_, _38137_, _28387_);
  and _48611_ (_41519_, _41518_, _39749_);
  nor _48612_ (_41520_, _41519_, _41517_);
  and _48613_ (_41521_, _27795_, _33107_);
  and _48614_ (_41522_, _41126_, _41521_);
  and _48615_ (_41523_, _41518_, _41522_);
  and _48616_ (_41524_, _41523_, _31212_);
  not _48617_ (_41525_, _41524_);
  nor _48618_ (_41526_, _41525_, _38225_);
  or _48619_ (_41527_, _41526_, _41520_);
  and _48620_ (_41528_, _41518_, _39553_);
  not _48621_ (_41529_, _41528_);
  and _48622_ (_41530_, _41529_, _41527_);
  and _48623_ (_41531_, _41528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _48624_ (_41532_, _41531_, _41530_);
  and _48625_ (_01637_, _41532_, _42618_);
  nand _48626_ (_41533_, _41528_, _38225_);
  nor _48627_ (_41534_, _41519_, _41514_);
  or _48628_ (_41535_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not _48629_ (_41536_, _41534_);
  or _48630_ (_41537_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _48631_ (_41538_, _41537_, _41535_);
  or _48632_ (_41539_, _41538_, _41528_);
  and _48633_ (_41540_, _41539_, _42618_);
  and _48634_ (_01640_, _41540_, _41533_);
  and _48635_ (_41541_, _41518_, _39705_);
  and _48636_ (_41542_, _39552_, _36133_);
  and _48637_ (_41543_, _41542_, _41518_);
  nor _48638_ (_41544_, _41543_, _41541_);
  not _48639_ (_41545_, _41511_);
  or _48640_ (_41546_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _48641_ (_41547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _48642_ (_41548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _41547_);
  and _48643_ (_41549_, _41548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _48644_ (_41550_, _41549_, _41546_);
  and _48645_ (_41551_, _41550_, _41545_);
  and _48646_ (_41552_, _41551_, _41544_);
  and _48647_ (_41553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _48648_ (_41554_, _41553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _48649_ (_41555_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _48650_ (_41556_, _41555_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _48651_ (_41557_, _41556_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _48652_ (_41558_, _41557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _48653_ (_41559_, _41558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _48654_ (_41560_, _41559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _48655_ (_41561_, _41560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _48656_ (_41562_, _41561_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _48657_ (_41563_, _41562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _48658_ (_41564_, _41563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _48659_ (_41565_, _41564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _48660_ (_41566_, _41565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _48661_ (_41567_, _41566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not _48662_ (_41568_, _41567_);
  nand _48663_ (_41569_, _41568_, _41552_);
  or _48664_ (_41570_, _41552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _48665_ (_41571_, _41570_, _42618_);
  and _48666_ (_01643_, _41571_, _41569_);
  nand _48667_ (_41572_, _41541_, _38225_);
  and _48668_ (_41573_, _41518_, _36133_);
  and _48669_ (_41574_, _41573_, _39552_);
  not _48670_ (_41575_, _41574_);
  not _48671_ (_41576_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _48672_ (_41577_, _41510_, _41576_);
  and _48673_ (_41578_, _41577_, _41511_);
  and _48674_ (_41579_, _41578_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not _48675_ (_41580_, _41578_);
  not _48676_ (_41581_, _41512_);
  and _48677_ (_41582_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _48678_ (_41583_, _41567_, _41550_);
  and _48679_ (_41584_, _41583_, _41582_);
  and _48680_ (_41585_, _41558_, _41550_);
  or _48681_ (_41586_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _48682_ (_41587_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _48683_ (_41588_, _41587_, _41586_);
  or _48684_ (_41589_, _41588_, _41584_);
  and _48685_ (_41590_, _41589_, _41580_);
  or _48686_ (_41591_, _41590_, _41579_);
  or _48687_ (_41592_, _41591_, _41541_);
  and _48688_ (_41593_, _41592_, _41575_);
  and _48689_ (_41594_, _41593_, _41572_);
  and _48690_ (_41595_, _41574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _48691_ (_41596_, _41595_, _41594_);
  and _48692_ (_01646_, _41596_, _42618_);
  and _48693_ (_41597_, _41566_, _41550_);
  or _48694_ (_41598_, _41597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _48695_ (_41599_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _48696_ (_41600_, _41599_, _41583_);
  and _48697_ (_41601_, _41600_, _41598_);
  or _48698_ (_41602_, _41601_, _41578_);
  or _48699_ (_41603_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _48700_ (_41604_, _41603_, _41544_);
  and _48701_ (_41605_, _41604_, _41602_);
  and _48702_ (_41606_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _48703_ (_41607_, _41606_, _41605_);
  not _48704_ (_41608_, _38225_);
  and _48705_ (_41609_, _41543_, _41608_);
  or _48706_ (_41610_, _41609_, _41607_);
  and _48707_ (_01649_, _41610_, _42618_);
  and _48708_ (_41611_, _41580_, _41550_);
  and _48709_ (_41612_, _41611_, _41511_);
  nand _48710_ (_41613_, _41612_, _41567_);
  nand _48711_ (_41614_, _41613_, _41544_);
  or _48712_ (_41615_, _41544_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _48713_ (_41616_, _41615_, _42618_);
  and _48714_ (_01652_, _41616_, _41614_);
  or _48715_ (_41617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _48716_ (_41618_, _40309_, _38614_);
  or _48717_ (_41619_, _41618_, _41617_);
  nand _48718_ (_41620_, _38617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _48719_ (_41621_, _41620_, _41618_);
  or _48720_ (_41622_, _41621_, _38618_);
  and _48721_ (_41623_, _41622_, _41619_);
  and _48722_ (_41624_, _41518_, _40304_);
  or _48723_ (_41625_, _41624_, _41623_);
  nand _48724_ (_41626_, _41624_, _38225_);
  and _48725_ (_41627_, _41626_, _42618_);
  and _48726_ (_01655_, _41627_, _41625_);
  or _48727_ (_41628_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not _48728_ (_41629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _48729_ (_41630_, _41513_, _41629_);
  and _48730_ (_41631_, _41630_, _41628_);
  or _48731_ (_41632_, _41631_, _41519_);
  nand _48732_ (_41633_, _41519_, _38203_);
  and _48733_ (_41634_, _41633_, _41632_);
  or _48734_ (_41635_, _41634_, _41528_);
  not _48735_ (_41636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _48736_ (_41637_, _41528_, _41636_);
  and _48737_ (_41638_, _41637_, _42618_);
  and _48738_ (_02111_, _41638_, _41635_);
  nand _48739_ (_41639_, _41519_, _38191_);
  and _48740_ (_41640_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _48741_ (_41641_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _48742_ (_41642_, _41641_, _41640_);
  or _48743_ (_41643_, _41642_, _41519_);
  and _48744_ (_41644_, _41643_, _41639_);
  or _48745_ (_41645_, _41644_, _41528_);
  or _48746_ (_41646_, _41529_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _48747_ (_41647_, _41646_, _42618_);
  and _48748_ (_02113_, _41647_, _41645_);
  nand _48749_ (_41648_, _41519_, _38184_);
  and _48750_ (_41649_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48751_ (_41650_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _48752_ (_41651_, _41650_, _41649_);
  or _48753_ (_41652_, _41651_, _41519_);
  and _48754_ (_41653_, _41652_, _41648_);
  or _48755_ (_41654_, _41653_, _41528_);
  or _48756_ (_41655_, _41529_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48757_ (_41656_, _41655_, _42618_);
  and _48758_ (_02115_, _41656_, _41654_);
  nand _48759_ (_41657_, _41519_, _38177_);
  and _48760_ (_41658_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _48761_ (_41659_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _48762_ (_41660_, _41659_, _41658_);
  or _48763_ (_41661_, _41660_, _41519_);
  and _48764_ (_41662_, _41661_, _41657_);
  or _48765_ (_41663_, _41662_, _41528_);
  or _48766_ (_41664_, _41529_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _48767_ (_41665_, _41664_, _42618_);
  and _48768_ (_02117_, _41665_, _41663_);
  nand _48769_ (_41666_, _41519_, _38169_);
  not _48770_ (_41667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor _48771_ (_41668_, _41513_, _41667_);
  and _48772_ (_41669_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _48773_ (_41670_, _41669_, _41668_);
  or _48774_ (_41671_, _41670_, _41519_);
  and _48775_ (_41672_, _41671_, _41666_);
  or _48776_ (_41673_, _41672_, _41528_);
  nand _48777_ (_41674_, _41528_, _41667_);
  and _48778_ (_41675_, _41674_, _42618_);
  and _48779_ (_02118_, _41675_, _41673_);
  and _48780_ (_41676_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48781_ (_41677_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _48782_ (_41678_, _41677_, _41676_);
  nor _48783_ (_41679_, _41678_, _41519_);
  nor _48784_ (_41680_, _41525_, _38162_);
  or _48785_ (_41681_, _41680_, _41679_);
  and _48786_ (_41682_, _41681_, _41529_);
  and _48787_ (_41683_, _41528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _48788_ (_41684_, _41683_, _41682_);
  and _48789_ (_02120_, _41684_, _42618_);
  and _48790_ (_41685_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _48791_ (_41686_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _48792_ (_41687_, _41686_, _41685_);
  nor _48793_ (_41688_, _41687_, _41519_);
  nor _48794_ (_41689_, _41525_, _38155_);
  or _48795_ (_41690_, _41689_, _41688_);
  and _48796_ (_41691_, _41690_, _41529_);
  and _48797_ (_41692_, _41528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _48798_ (_41693_, _41692_, _41691_);
  and _48799_ (_02122_, _41693_, _42618_);
  or _48800_ (_41694_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not _48801_ (_41695_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _48802_ (_41696_, _41534_, _41695_);
  and _48803_ (_41697_, _41696_, _41694_);
  or _48804_ (_41698_, _41697_, _41528_);
  nand _48805_ (_41699_, _41528_, _38203_);
  and _48806_ (_41700_, _41699_, _42618_);
  and _48807_ (_02124_, _41700_, _41698_);
  and _48808_ (_41701_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _48809_ (_41702_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _48810_ (_41703_, _41702_, _41701_);
  or _48811_ (_41704_, _41703_, _41528_);
  nand _48812_ (_41705_, _41528_, _38191_);
  and _48813_ (_41706_, _41705_, _42618_);
  and _48814_ (_02125_, _41706_, _41704_);
  nand _48815_ (_41707_, _41528_, _38184_);
  and _48816_ (_41708_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _48817_ (_41709_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _48818_ (_41710_, _41709_, _41708_);
  or _48819_ (_41711_, _41710_, _41528_);
  and _48820_ (_41712_, _41711_, _42618_);
  and _48821_ (_02127_, _41712_, _41707_);
  nand _48822_ (_41713_, _41528_, _38177_);
  and _48823_ (_41714_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _48824_ (_41715_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _48825_ (_41716_, _41715_, _41714_);
  or _48826_ (_41717_, _41716_, _41528_);
  and _48827_ (_41718_, _41717_, _42618_);
  and _48828_ (_02129_, _41718_, _41713_);
  nand _48829_ (_41719_, _41528_, _38169_);
  not _48830_ (_41720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _48831_ (_41721_, _41534_, _41720_);
  and _48832_ (_41722_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _48833_ (_41723_, _41722_, _41721_);
  or _48834_ (_41724_, _41723_, _41528_);
  and _48835_ (_41725_, _41724_, _42618_);
  and _48836_ (_02131_, _41725_, _41719_);
  nand _48837_ (_41726_, _41528_, _38162_);
  and _48838_ (_41727_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _48839_ (_41728_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _48840_ (_41729_, _41728_, _41727_);
  or _48841_ (_41730_, _41729_, _41528_);
  and _48842_ (_41731_, _41730_, _42618_);
  and _48843_ (_02132_, _41731_, _41726_);
  nand _48844_ (_41732_, _41528_, _38155_);
  and _48845_ (_41733_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _48846_ (_41734_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _48847_ (_41735_, _41734_, _41733_);
  or _48848_ (_41736_, _41735_, _41528_);
  and _48849_ (_41737_, _41736_, _42618_);
  and _48850_ (_02134_, _41737_, _41732_);
  or _48851_ (_41738_, _41550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _48852_ (_41739_, _41550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _48853_ (_41740_, _41512_, _41636_);
  nand _48854_ (_41741_, _41740_, _41567_);
  nand _48855_ (_41742_, _41741_, _41739_);
  and _48856_ (_41743_, _41742_, _41738_);
  or _48857_ (_41744_, _41743_, _41578_);
  and _48858_ (_41745_, _41578_, _41636_);
  nor _48859_ (_41746_, _41745_, _41541_);
  and _48860_ (_41747_, _41746_, _41744_);
  not _48861_ (_41748_, _41541_);
  nor _48862_ (_41749_, _41748_, _38203_);
  or _48863_ (_41750_, _41749_, _41574_);
  or _48864_ (_41751_, _41750_, _41747_);
  nand _48865_ (_41752_, _41543_, _41629_);
  and _48866_ (_41753_, _41752_, _42618_);
  and _48867_ (_02136_, _41753_, _41751_);
  and _48868_ (_41754_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _48869_ (_41755_, _41754_, _41611_);
  and _48870_ (_41756_, _41755_, _41567_);
  and _48871_ (_41757_, _41578_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _48872_ (_41758_, _41739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand _48873_ (_41759_, _41553_, _41550_);
  and _48874_ (_41760_, _41759_, _41580_);
  and _48875_ (_41761_, _41760_, _41758_);
  nor _48876_ (_41762_, _41761_, _41757_);
  nand _48877_ (_41763_, _41762_, _41544_);
  or _48878_ (_41764_, _41763_, _41756_);
  nand _48879_ (_41765_, _41541_, _38191_);
  or _48880_ (_41766_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _48881_ (_41767_, _41766_, _42618_);
  and _48882_ (_41768_, _41767_, _41765_);
  and _48883_ (_02138_, _41768_, _41764_);
  and _48884_ (_41769_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48885_ (_41770_, _41769_, _41583_);
  and _48886_ (_41771_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _48887_ (_41772_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _48888_ (_41773_, _41772_, _41578_);
  or _48889_ (_41774_, _41773_, _41771_);
  or _48890_ (_41775_, _41774_, _41770_);
  nor _48891_ (_41776_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor _48892_ (_41777_, _41776_, _41541_);
  and _48893_ (_41778_, _41777_, _41775_);
  nor _48894_ (_41779_, _41748_, _38184_);
  or _48895_ (_41780_, _41779_, _41778_);
  or _48896_ (_41781_, _41780_, _41574_);
  or _48897_ (_41782_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _48898_ (_41783_, _41782_, _42618_);
  and _48899_ (_02139_, _41783_, _41781_);
  and _48900_ (_41784_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _48901_ (_41785_, _41784_, _41583_);
  nand _48902_ (_41786_, _41554_, _41550_);
  and _48903_ (_41787_, _41786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _48904_ (_41788_, _41786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _48905_ (_41789_, _41788_, _41578_);
  or _48906_ (_41790_, _41789_, _41787_);
  or _48907_ (_41791_, _41790_, _41785_);
  nor _48908_ (_41792_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor _48909_ (_41793_, _41792_, _41541_);
  and _48910_ (_41794_, _41793_, _41791_);
  nor _48911_ (_41795_, _41748_, _38177_);
  or _48912_ (_41796_, _41795_, _41794_);
  or _48913_ (_41797_, _41796_, _41574_);
  or _48914_ (_41798_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _48915_ (_41799_, _41798_, _42618_);
  and _48916_ (_02141_, _41799_, _41797_);
  nor _48917_ (_41800_, _41512_, _41667_);
  and _48918_ (_41801_, _41800_, _41583_);
  not _48919_ (_41802_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _48920_ (_41803_, _41555_, _41550_);
  nor _48921_ (_41804_, _41803_, _41802_);
  and _48922_ (_41805_, _41803_, _41802_);
  or _48923_ (_41806_, _41805_, _41578_);
  or _48924_ (_41807_, _41806_, _41804_);
  or _48925_ (_41808_, _41807_, _41801_);
  and _48926_ (_41809_, _41578_, _41667_);
  nor _48927_ (_41810_, _41809_, _41541_);
  and _48928_ (_41811_, _41810_, _41808_);
  nor _48929_ (_41812_, _41748_, _38169_);
  or _48930_ (_41813_, _41812_, _41811_);
  or _48931_ (_41814_, _41813_, _41574_);
  nand _48932_ (_41815_, _41543_, _41802_);
  and _48933_ (_41816_, _41815_, _42618_);
  and _48934_ (_02143_, _41816_, _41814_);
  and _48935_ (_41817_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48936_ (_41818_, _41817_, _41583_);
  nand _48937_ (_41819_, _41556_, _41550_);
  and _48938_ (_41820_, _41819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _48939_ (_41821_, _41819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _48940_ (_41822_, _41821_, _41578_);
  or _48941_ (_41823_, _41822_, _41820_);
  or _48942_ (_41824_, _41823_, _41818_);
  nor _48943_ (_41825_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor _48944_ (_41826_, _41825_, _41541_);
  and _48945_ (_41827_, _41826_, _41824_);
  nor _48946_ (_41828_, _41748_, _38162_);
  or _48947_ (_41829_, _41828_, _41827_);
  or _48948_ (_41830_, _41829_, _41574_);
  or _48949_ (_41831_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _48950_ (_41832_, _41831_, _42618_);
  and _48951_ (_02145_, _41832_, _41830_);
  nor _48952_ (_41833_, _41748_, _38155_);
  and _48953_ (_41834_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _48954_ (_41835_, _41834_, _41583_);
  and _48955_ (_41836_, _41557_, _41550_);
  nor _48956_ (_41837_, _41836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _48957_ (_41838_, _41837_, _41585_);
  or _48958_ (_41839_, _41838_, _41578_);
  or _48959_ (_41840_, _41839_, _41835_);
  nor _48960_ (_41841_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _48961_ (_41842_, _41841_, _41541_);
  and _48962_ (_41843_, _41842_, _41840_);
  or _48963_ (_41844_, _41843_, _41574_);
  or _48964_ (_41845_, _41844_, _41833_);
  or _48965_ (_41846_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _48966_ (_41847_, _41846_, _42618_);
  and _48967_ (_02146_, _41847_, _41845_);
  not _48968_ (_41848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _48969_ (_41849_, _41512_, _41848_);
  and _48970_ (_41850_, _41849_, _41583_);
  and _48971_ (_41851_, _41559_, _41550_);
  or _48972_ (_41852_, _41851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _48973_ (_41853_, _41851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _48974_ (_41854_, _41853_, _41852_);
  or _48975_ (_41855_, _41854_, _41578_);
  or _48976_ (_41856_, _41855_, _41850_);
  and _48977_ (_41857_, _41578_, _41848_);
  nor _48978_ (_41858_, _41857_, _41541_);
  and _48979_ (_41859_, _41858_, _41856_);
  and _48980_ (_41860_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _48981_ (_41861_, _41860_, _41574_);
  or _48982_ (_41862_, _41861_, _41859_);
  nand _48983_ (_41863_, _41543_, _38203_);
  and _48984_ (_41864_, _41863_, _42618_);
  and _48985_ (_02148_, _41864_, _41862_);
  and _48986_ (_41865_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _48987_ (_41866_, _41865_, _41583_);
  and _48988_ (_41867_, _41560_, _41550_);
  or _48989_ (_41868_, _41867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _48990_ (_41869_, _41867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _48991_ (_41870_, _41869_, _41868_);
  or _48992_ (_41871_, _41870_, _41578_);
  or _48993_ (_41872_, _41871_, _41866_);
  nor _48994_ (_41873_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _48995_ (_41874_, _41873_, _41541_);
  and _48996_ (_41875_, _41874_, _41872_);
  and _48997_ (_41876_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _48998_ (_41877_, _41876_, _41574_);
  or _48999_ (_41878_, _41877_, _41875_);
  nand _49000_ (_41879_, _41574_, _38191_);
  and _49001_ (_41880_, _41879_, _42618_);
  and _49002_ (_02150_, _41880_, _41878_);
  and _49003_ (_41881_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _49004_ (_41882_, _41881_, _41583_);
  nand _49005_ (_41883_, _41561_, _41550_);
  and _49006_ (_41884_, _41883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _49007_ (_41885_, _41883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _49008_ (_41886_, _41885_, _41578_);
  or _49009_ (_41887_, _41886_, _41884_);
  or _49010_ (_41888_, _41887_, _41882_);
  nor _49011_ (_41889_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _49012_ (_41890_, _41889_, _41541_);
  and _49013_ (_41891_, _41890_, _41888_);
  and _49014_ (_41892_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _49015_ (_41893_, _41892_, _41574_);
  or _49016_ (_41894_, _41893_, _41891_);
  nand _49017_ (_41895_, _41574_, _38184_);
  and _49018_ (_41896_, _41895_, _42618_);
  and _49019_ (_02152_, _41896_, _41894_);
  and _49020_ (_41897_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _49021_ (_41898_, _41897_, _41583_);
  nand _49022_ (_41899_, _41562_, _41550_);
  and _49023_ (_41900_, _41899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor _49024_ (_41901_, _41899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49025_ (_41902_, _41901_, _41578_);
  or _49026_ (_41903_, _41902_, _41900_);
  or _49027_ (_41904_, _41903_, _41898_);
  nor _49028_ (_41905_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _49029_ (_41906_, _41905_, _41541_);
  and _49030_ (_41907_, _41906_, _41904_);
  and _49031_ (_41908_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49032_ (_41909_, _41908_, _41574_);
  or _49033_ (_41910_, _41909_, _41907_);
  nand _49034_ (_41911_, _41574_, _38177_);
  and _49035_ (_41912_, _41911_, _42618_);
  and _49036_ (_02153_, _41912_, _41910_);
  nor _49037_ (_41913_, _41512_, _41720_);
  and _49038_ (_41914_, _41913_, _41583_);
  not _49039_ (_41915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _49040_ (_41916_, _41563_, _41550_);
  nor _49041_ (_41917_, _41916_, _41915_);
  and _49042_ (_41918_, _41916_, _41915_);
  or _49043_ (_41919_, _41918_, _41578_);
  or _49044_ (_41920_, _41919_, _41917_);
  or _49045_ (_41921_, _41920_, _41914_);
  and _49046_ (_41922_, _41578_, _41720_);
  nor _49047_ (_41923_, _41922_, _41541_);
  and _49048_ (_41924_, _41923_, _41921_);
  and _49049_ (_41925_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _49050_ (_41926_, _41925_, _41574_);
  or _49051_ (_41927_, _41926_, _41924_);
  nand _49052_ (_41928_, _41574_, _38169_);
  and _49053_ (_41929_, _41928_, _42618_);
  and _49054_ (_02155_, _41929_, _41927_);
  and _49055_ (_41930_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _49056_ (_41931_, _41930_, _41583_);
  nand _49057_ (_41932_, _41564_, _41550_);
  and _49058_ (_41933_, _41932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _49059_ (_41934_, _41932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _49060_ (_41935_, _41934_, _41578_);
  or _49061_ (_41936_, _41935_, _41933_);
  or _49062_ (_41937_, _41936_, _41931_);
  nor _49063_ (_41938_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor _49064_ (_41939_, _41938_, _41541_);
  and _49065_ (_41940_, _41939_, _41937_);
  and _49066_ (_41941_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _49067_ (_41942_, _41941_, _41574_);
  or _49068_ (_41943_, _41942_, _41940_);
  nand _49069_ (_41944_, _41574_, _38162_);
  and _49070_ (_41945_, _41944_, _42618_);
  and _49071_ (_02157_, _41945_, _41943_);
  and _49072_ (_41946_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _49073_ (_41947_, _41946_, _41583_);
  and _49074_ (_41948_, _41565_, _41550_);
  nor _49075_ (_41949_, _41948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _49076_ (_41950_, _41949_, _41597_);
  or _49077_ (_41951_, _41950_, _41578_);
  or _49078_ (_41952_, _41951_, _41947_);
  nor _49079_ (_41953_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _49080_ (_41954_, _41953_, _41541_);
  and _49081_ (_41955_, _41954_, _41952_);
  and _49082_ (_41956_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _49083_ (_41957_, _41956_, _41574_);
  or _49084_ (_41958_, _41957_, _41955_);
  nand _49085_ (_41959_, _41574_, _38155_);
  and _49086_ (_41960_, _41959_, _42618_);
  and _49087_ (_02159_, _41960_, _41958_);
  not _49088_ (_41961_, _41624_);
  and _49089_ (_41962_, _41618_, _38813_);
  or _49090_ (_41963_, _41962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _49091_ (_41964_, _41963_, _41961_);
  nand _49092_ (_41965_, _41962_, _31757_);
  and _49093_ (_41966_, _41965_, _41964_);
  nor _49094_ (_41967_, _41961_, _38203_);
  or _49095_ (_41968_, _41967_, _41966_);
  and _49096_ (_02160_, _41968_, _42618_);
  and _49097_ (_41969_, _41618_, _33129_);
  or _49098_ (_41970_, _41969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _49099_ (_41971_, _41970_, _41961_);
  nand _49100_ (_41972_, _41969_, _31757_);
  and _49101_ (_41973_, _41972_, _41971_);
  nor _49102_ (_41974_, _41961_, _38191_);
  or _49103_ (_41975_, _41974_, _41973_);
  and _49104_ (_02162_, _41975_, _42618_);
  nand _49105_ (_41976_, _41618_, _39025_);
  and _49106_ (_41977_, _41976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _49107_ (_41978_, _41977_, _41624_);
  and _49108_ (_41979_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _49109_ (_41980_, _41979_, _33869_);
  and _49110_ (_41981_, _41980_, _41618_);
  or _49111_ (_41982_, _41981_, _41978_);
  nand _49112_ (_41983_, _41624_, _38184_);
  and _49113_ (_41984_, _41983_, _42618_);
  and _49114_ (_02164_, _41984_, _41982_);
  and _49115_ (_41985_, _41618_, _34576_);
  or _49116_ (_41986_, _41985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _49117_ (_41987_, _41986_, _41961_);
  nand _49118_ (_41988_, _41985_, _31757_);
  and _49119_ (_41989_, _41988_, _41987_);
  nor _49120_ (_41990_, _41961_, _38177_);
  or _49121_ (_41991_, _41990_, _41989_);
  and _49122_ (_02166_, _41991_, _42618_);
  and _49123_ (_41992_, _41618_, _35338_);
  or _49124_ (_41993_, _41992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _49125_ (_41994_, _41993_, _41961_);
  nand _49126_ (_41995_, _41992_, _31757_);
  and _49127_ (_41996_, _41995_, _41994_);
  nor _49128_ (_41997_, _41961_, _38169_);
  or _49129_ (_41998_, _41997_, _41996_);
  and _49130_ (_02167_, _41998_, _42618_);
  and _49131_ (_41999_, _41618_, _36133_);
  or _49132_ (_42000_, _41999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _49133_ (_42001_, _42000_, _41961_);
  nand _49134_ (_42002_, _41999_, _31757_);
  and _49135_ (_42003_, _42002_, _42001_);
  nor _49136_ (_42004_, _41961_, _38162_);
  or _49137_ (_42005_, _42004_, _42003_);
  and _49138_ (_02169_, _42005_, _42618_);
  not _49139_ (_42006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49140_ (_42007_, _41510_, _42006_);
  or _49141_ (_42008_, _42007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _49142_ (_42009_, _42008_, _41618_);
  nand _49143_ (_42010_, _38739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _49144_ (_42011_, _42010_, _41618_);
  or _49145_ (_42012_, _42011_, _38740_);
  and _49146_ (_42013_, _42012_, _42009_);
  or _49147_ (_42014_, _42013_, _41624_);
  nand _49148_ (_42015_, _41624_, _38155_);
  and _49149_ (_42016_, _42015_, _42618_);
  and _49150_ (_02171_, _42016_, _42014_);
  and _49151_ (_42017_, _38227_, _38135_);
  not _49152_ (_42018_, _42017_);
  not _49153_ (_42019_, _38133_);
  and _49154_ (_42020_, _42019_, _38099_);
  and _49155_ (_42021_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _49156_ (_42022_, _42021_, _38711_);
  nor _49157_ (_42023_, _42022_, _31790_);
  and _49158_ (_42024_, _42022_, _31790_);
  or _49159_ (_42025_, _42024_, _42023_);
  not _49160_ (_42026_, _42025_);
  and _49161_ (_42027_, _37657_, _27795_);
  nor _49162_ (_42028_, _37657_, _27795_);
  nor _49163_ (_42029_, _42028_, _42027_);
  and _49164_ (_42030_, _28376_, _28244_);
  not _49165_ (_42031_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _49166_ (_42032_, _31189_, _42031_);
  and _49167_ (_42033_, _42032_, _33880_);
  and _49168_ (_42034_, _42033_, _42030_);
  and _49169_ (_42035_, _42034_, _42029_);
  and _49170_ (_42036_, _42035_, _27345_);
  and _49171_ (_42037_, _38716_, _40289_);
  nor _49172_ (_42038_, _38716_, _40289_);
  nor _49173_ (_42039_, _42038_, _42037_);
  and _49174_ (_42040_, _42039_, _42036_);
  and _49175_ (_42041_, _42040_, _42026_);
  not _49176_ (_42042_, _38716_);
  nor _49177_ (_42043_, _42022_, _38004_);
  and _49178_ (_42044_, _42043_, _42042_);
  and _49179_ (_42045_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor _49180_ (_42046_, _42022_, _37657_);
  and _49181_ (_42047_, _42046_, _42042_);
  and _49182_ (_42048_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor _49183_ (_42049_, _42048_, _42045_);
  and _49184_ (_42050_, _42022_, _37657_);
  and _49185_ (_42051_, _42050_, _42042_);
  and _49186_ (_42052_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _49187_ (_42053_, _42022_, _38004_);
  and _49188_ (_42054_, _42053_, _38716_);
  and _49189_ (_42055_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor _49190_ (_42056_, _42055_, _42052_);
  and _49191_ (_42057_, _42056_, _42049_);
  and _49192_ (_42058_, _42050_, _38716_);
  and _49193_ (_42059_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _49194_ (_42060_, _42043_, _38716_);
  and _49195_ (_42061_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor _49196_ (_42062_, _42061_, _42059_);
  and _49197_ (_42063_, _42046_, _38716_);
  and _49198_ (_42064_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _49199_ (_42065_, _42053_, _42042_);
  and _49200_ (_42066_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor _49201_ (_42067_, _42066_, _42064_);
  and _49202_ (_42068_, _42067_, _42062_);
  and _49203_ (_42069_, _42068_, _42057_);
  nor _49204_ (_42070_, _42069_, _42041_);
  and _49205_ (_42071_, _42041_, _41608_);
  nor _49206_ (_42072_, _42071_, _42070_);
  not _49207_ (_42073_, _42072_);
  and _49208_ (_42074_, _42073_, _42020_);
  not _49209_ (_42075_, _42074_);
  not _49210_ (_42076_, _37999_);
  nor _49211_ (_42077_, _42019_, _38099_);
  and _49212_ (_42078_, _42077_, _37999_);
  not _49213_ (_42079_, _36958_);
  and _49214_ (_42080_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and _49215_ (_42081_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _49216_ (_42082_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _49217_ (_42083_, _42082_, _42081_);
  and _49218_ (_42084_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _49219_ (_42085_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _49220_ (_42086_, _42085_, _42084_);
  and _49221_ (_42087_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _49222_ (_42088_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _49223_ (_42089_, _42088_, _42087_);
  and _49224_ (_42090_, _42089_, _42086_);
  and _49225_ (_42091_, _42090_, _42083_);
  nor _49226_ (_42092_, _37012_, _42079_);
  not _49227_ (_42093_, _42092_);
  nor _49228_ (_42094_, _42093_, _42091_);
  nor _49229_ (_42095_, _42094_, _42080_);
  not _49230_ (_42096_, _42095_);
  and _49231_ (_42097_, _42096_, _42078_);
  nor _49232_ (_42098_, _42097_, _42076_);
  and _49233_ (_42099_, _42098_, _42075_);
  and _49234_ (_42100_, _42099_, _42018_);
  and _49235_ (_42101_, _37987_, _38008_);
  nor _49236_ (_42102_, _42101_, _38073_);
  and _49237_ (_42103_, _37962_, _37987_);
  nor _49238_ (_42104_, _42103_, _38027_);
  not _49239_ (_42105_, _42104_);
  nor _49240_ (_42106_, _42105_, _38080_);
  and _49241_ (_42107_, _42106_, _42102_);
  and _49242_ (_42108_, _38045_, _38011_);
  and _49243_ (_42109_, _42108_, _38036_);
  and _49244_ (_42110_, _42109_, _42107_);
  nor _49245_ (_42111_, _42110_, _36914_);
  nor _49246_ (_42112_, _38043_, _38039_);
  not _49247_ (_42113_, _37990_);
  nor _49248_ (_42114_, _42113_, _42112_);
  nor _49249_ (_42115_, _42114_, _42111_);
  not _49250_ (_42116_, _42115_);
  and _49251_ (_42117_, _42116_, _42100_);
  and _49252_ (_42118_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and _49253_ (_42119_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _49254_ (_42120_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _49255_ (_42121_, _42120_, _42119_);
  and _49256_ (_42122_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _49257_ (_42123_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _49258_ (_42124_, _42123_, _42122_);
  and _49259_ (_42125_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _49260_ (_42126_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _49261_ (_42127_, _42126_, _42125_);
  and _49262_ (_42128_, _42127_, _42124_);
  and _49263_ (_42129_, _42128_, _42121_);
  nor _49264_ (_42130_, _42129_, _42093_);
  nor _49265_ (_42131_, _42130_, _42118_);
  not _49266_ (_42132_, _42131_);
  and _49267_ (_42133_, _42132_, _42078_);
  not _49268_ (_42134_, _42133_);
  and _49269_ (_42135_, _42076_, _38133_);
  and _49270_ (_42136_, _42135_, _38099_);
  not _49271_ (_42137_, _38265_);
  and _49272_ (_42138_, _42137_, _38135_);
  nor _49273_ (_42139_, _42138_, _42136_);
  and _49274_ (_42140_, _42139_, _42134_);
  and _49275_ (_42141_, _38134_, _42076_);
  and _49276_ (_42142_, _42020_, _37999_);
  and _49277_ (_42143_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _49278_ (_42144_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _49279_ (_42145_, _42144_, _42143_);
  and _49280_ (_42146_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _49281_ (_42147_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _49282_ (_42148_, _42147_, _42146_);
  and _49283_ (_42149_, _42148_, _42145_);
  and _49284_ (_42150_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _49285_ (_42151_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor _49286_ (_42152_, _42151_, _42150_);
  and _49287_ (_42153_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _49288_ (_42154_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _49289_ (_42155_, _42154_, _42153_);
  and _49290_ (_42156_, _42155_, _42152_);
  and _49291_ (_42157_, _42156_, _42149_);
  nor _49292_ (_42158_, _42157_, _42041_);
  and _49293_ (_42159_, _42041_, _39920_);
  nor _49294_ (_42160_, _42159_, _42158_);
  not _49295_ (_42161_, _42160_);
  and _49296_ (_42162_, _42161_, _42142_);
  nor _49297_ (_42163_, _42162_, _42141_);
  and _49298_ (_42164_, _42163_, _42140_);
  not _49299_ (_42165_, _42164_);
  and _49300_ (_42166_, _42165_, _42117_);
  and _49301_ (_42167_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _49302_ (_42168_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _49303_ (_42169_, _42168_, _42167_);
  and _49304_ (_42170_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and _49305_ (_42171_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _49306_ (_42172_, _42171_, _42170_);
  and _49307_ (_42173_, _42172_, _42169_);
  and _49308_ (_42174_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _49309_ (_42175_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor _49310_ (_42176_, _42175_, _42174_);
  and _49311_ (_42177_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _49312_ (_42178_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _49313_ (_42179_, _42178_, _42177_);
  and _49314_ (_42180_, _42179_, _42176_);
  and _49315_ (_42181_, _42180_, _42173_);
  nor _49316_ (_42182_, _42181_, _42041_);
  and _49317_ (_42183_, _42041_, _39884_);
  nor _49318_ (_42184_, _42183_, _42182_);
  not _49319_ (_42185_, _42184_);
  and _49320_ (_42186_, _42185_, _42142_);
  not _49321_ (_42187_, _42186_);
  and _49322_ (_42188_, _37999_, _38133_);
  and _49323_ (_42189_, _42188_, _38099_);
  and _49324_ (_42190_, _42189_, _37837_);
  not _49325_ (_42191_, _42190_);
  not _49326_ (_42192_, _38247_);
  and _49327_ (_42193_, _42192_, _38135_);
  and _49328_ (_42194_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _49329_ (_42195_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _49330_ (_42196_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _49331_ (_42197_, _42196_, _42195_);
  and _49332_ (_42198_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _49333_ (_42199_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _49334_ (_42200_, _42199_, _42198_);
  and _49335_ (_42201_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _49336_ (_42202_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _49337_ (_42203_, _42202_, _42201_);
  and _49338_ (_42204_, _42203_, _42200_);
  and _49339_ (_42205_, _42204_, _42197_);
  nor _49340_ (_42206_, _42205_, _42093_);
  nor _49341_ (_42207_, _42206_, _42194_);
  not _49342_ (_42208_, _42207_);
  and _49343_ (_42209_, _42208_, _42078_);
  nor _49344_ (_42210_, _42209_, _42193_);
  and _49345_ (_42211_, _42210_, _42191_);
  and _49346_ (_42212_, _42211_, _42187_);
  nor _49347_ (_42213_, _42212_, _42116_);
  nor _49348_ (_42214_, _42213_, _42166_);
  not _49349_ (_42215_, _42214_);
  and _49350_ (_42216_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _49351_ (_42217_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _49352_ (_42218_, _42217_, _42216_);
  and _49353_ (_42219_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _49354_ (_42220_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _49355_ (_42221_, _42220_, _42219_);
  and _49356_ (_42222_, _42221_, _42218_);
  and _49357_ (_42223_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _49358_ (_42224_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _49359_ (_42225_, _42224_, _42223_);
  and _49360_ (_42226_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _49361_ (_42227_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor _49362_ (_42228_, _42227_, _42226_);
  and _49363_ (_42229_, _42228_, _42225_);
  and _49364_ (_42230_, _42229_, _42222_);
  nor _49365_ (_42231_, _42230_, _42041_);
  and _49366_ (_42232_, _42041_, _39907_);
  nor _49367_ (_42233_, _42232_, _42231_);
  not _49368_ (_42234_, _42233_);
  and _49369_ (_42235_, _42234_, _42142_);
  not _49370_ (_42236_, _42235_);
  not _49371_ (_42237_, _38259_);
  and _49372_ (_42238_, _42237_, _38135_);
  nor _49373_ (_42239_, _42238_, _42135_);
  and _49374_ (_42240_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and _49375_ (_42241_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _49376_ (_42242_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _49377_ (_42243_, _42242_, _42241_);
  and _49378_ (_42244_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _49379_ (_42245_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _49380_ (_42246_, _42245_, _42244_);
  and _49381_ (_42247_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _49382_ (_42248_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _49383_ (_42249_, _42248_, _42247_);
  and _49384_ (_42250_, _42249_, _42246_);
  and _49385_ (_42251_, _42250_, _42243_);
  nor _49386_ (_42252_, _42251_, _42093_);
  nor _49387_ (_42253_, _42252_, _42240_);
  not _49388_ (_42254_, _42253_);
  and _49389_ (_42255_, _42254_, _42078_);
  and _49390_ (_42256_, _42189_, _42042_);
  nor _49391_ (_42257_, _42256_, _42255_);
  and _49392_ (_42258_, _42257_, _42239_);
  and _49393_ (_42259_, _42258_, _42236_);
  not _49394_ (_42260_, _42259_);
  and _49395_ (_42261_, _42260_, _42117_);
  and _49396_ (_42262_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _49397_ (_42263_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _49398_ (_42264_, _42263_, _42262_);
  and _49399_ (_42265_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _49400_ (_42266_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _49401_ (_42267_, _42266_, _42265_);
  and _49402_ (_42268_, _42267_, _42264_);
  and _49403_ (_42269_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _49404_ (_42270_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _49405_ (_42271_, _42270_, _42269_);
  and _49406_ (_42272_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _49407_ (_42273_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _49408_ (_42274_, _42273_, _42272_);
  and _49409_ (_42275_, _42274_, _42271_);
  and _49410_ (_42276_, _42275_, _42268_);
  nor _49411_ (_42277_, _42276_, _42041_);
  not _49412_ (_42278_, _38191_);
  and _49413_ (_42279_, _42041_, _42278_);
  nor _49414_ (_42280_, _42279_, _42277_);
  not _49415_ (_42281_, _42280_);
  and _49416_ (_42282_, _42281_, _42142_);
  not _49417_ (_42283_, _42282_);
  and _49418_ (_42284_, _42020_, _42076_);
  and _49419_ (_42285_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _49420_ (_42286_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _49421_ (_42287_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _49422_ (_42288_, _42287_, _42286_);
  and _49423_ (_42289_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _49424_ (_42290_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _49425_ (_42291_, _42290_, _42289_);
  and _49426_ (_42292_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _49427_ (_42293_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _49428_ (_42294_, _42293_, _42292_);
  and _49429_ (_42295_, _42294_, _42291_);
  and _49430_ (_42296_, _42295_, _42288_);
  nor _49431_ (_42297_, _42296_, _42093_);
  nor _49432_ (_42298_, _42297_, _42285_);
  not _49433_ (_42299_, _42298_);
  and _49434_ (_42300_, _42299_, _42078_);
  nor _49435_ (_42301_, _42300_, _42284_);
  not _49436_ (_42302_, _38241_);
  and _49437_ (_42303_, _42302_, _38135_);
  and _49438_ (_42304_, _42189_, _37863_);
  nor _49439_ (_42305_, _42304_, _42303_);
  and _49440_ (_42306_, _42305_, _42301_);
  and _49441_ (_42307_, _42306_, _42283_);
  nor _49442_ (_42308_, _42307_, _42116_);
  nor _49443_ (_42309_, _42308_, _42261_);
  and _49444_ (_42310_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _49445_ (_42311_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _49446_ (_42312_, _42311_, _42310_);
  and _49447_ (_42313_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _49448_ (_42314_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _49449_ (_42315_, _42314_, _42313_);
  and _49450_ (_42316_, _42315_, _42312_);
  and _49451_ (_42317_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _49452_ (_42318_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor _49453_ (_42319_, _42318_, _42317_);
  and _49454_ (_42320_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _49455_ (_42321_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _49456_ (_42322_, _42321_, _42320_);
  and _49457_ (_42323_, _42322_, _42319_);
  and _49458_ (_42324_, _42323_, _42316_);
  nor _49459_ (_42325_, _42324_, _42041_);
  and _49460_ (_42326_, _42041_, _39896_);
  nor _49461_ (_42327_, _42326_, _42325_);
  not _49462_ (_42328_, _42327_);
  and _49463_ (_42329_, _42328_, _42142_);
  not _49464_ (_42330_, _42329_);
  not _49465_ (_42331_, _38253_);
  and _49466_ (_42332_, _42331_, _38135_);
  not _49467_ (_42333_, _42332_);
  not _49468_ (_42334_, _42022_);
  and _49469_ (_42335_, _42189_, _42334_);
  and _49470_ (_42336_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _49471_ (_42337_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _49472_ (_42338_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _49473_ (_42339_, _42338_, _42337_);
  and _49474_ (_42340_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _49475_ (_42341_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _49476_ (_42342_, _42341_, _42340_);
  and _49477_ (_42343_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _49478_ (_42344_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _49479_ (_42345_, _42344_, _42343_);
  and _49480_ (_42346_, _42345_, _42342_);
  and _49481_ (_42347_, _42346_, _42339_);
  nor _49482_ (_42348_, _42347_, _42093_);
  nor _49483_ (_42349_, _42348_, _42336_);
  not _49484_ (_42350_, _42349_);
  and _49485_ (_42351_, _42350_, _42078_);
  nor _49486_ (_42352_, _42351_, _42335_);
  and _49487_ (_42353_, _42352_, _42333_);
  and _49488_ (_42354_, _42353_, _42330_);
  not _49489_ (_42355_, _42354_);
  and _49490_ (_42356_, _42355_, _42117_);
  and _49491_ (_42357_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _49492_ (_42358_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor _49493_ (_42359_, _42358_, _42357_);
  and _49494_ (_42360_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _49495_ (_42361_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _49496_ (_42362_, _42361_, _42360_);
  and _49497_ (_42363_, _42362_, _42359_);
  and _49498_ (_42364_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _49499_ (_42365_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _49500_ (_42366_, _42365_, _42364_);
  and _49501_ (_42367_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _49502_ (_42368_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor _49503_ (_42369_, _42368_, _42367_);
  and _49504_ (_42370_, _42369_, _42366_);
  and _49505_ (_42371_, _42370_, _42363_);
  nor _49506_ (_42372_, _42371_, _42041_);
  and _49507_ (_42373_, _42041_, _38204_);
  nor _49508_ (_42374_, _42373_, _42372_);
  not _49509_ (_42375_, _42374_);
  and _49510_ (_42376_, _42375_, _42142_);
  not _49511_ (_42377_, _42376_);
  and _49512_ (_42378_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _49513_ (_42379_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _49514_ (_42380_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _49515_ (_42381_, _42380_, _42379_);
  and _49516_ (_42382_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _49517_ (_42383_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _49518_ (_42384_, _42383_, _42382_);
  and _49519_ (_42385_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _49520_ (_42386_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _49521_ (_42387_, _42386_, _42385_);
  and _49522_ (_42388_, _42387_, _42384_);
  and _49523_ (_42389_, _42388_, _42381_);
  nor _49524_ (_42390_, _42389_, _42093_);
  nor _49525_ (_42391_, _42390_, _42378_);
  not _49526_ (_42392_, _42391_);
  and _49527_ (_42393_, _42392_, _42078_);
  not _49528_ (_42394_, _42393_);
  not _49529_ (_42395_, _38235_);
  and _49530_ (_42396_, _42395_, _38135_);
  and _49531_ (_42397_, _42189_, _37657_);
  nor _49532_ (_42398_, _42397_, _42396_);
  and _49533_ (_42399_, _42398_, _42394_);
  and _49534_ (_42400_, _42399_, _42377_);
  nor _49535_ (_42401_, _42400_, _42116_);
  nor _49536_ (_42402_, _42401_, _42356_);
  or _49537_ (_42403_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not _49538_ (_42404_, _42402_);
  or _49539_ (_42405_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _49540_ (_42406_, _42405_, _42403_);
  or _49541_ (_42407_, _42406_, _42309_);
  not _49542_ (_42408_, _38271_);
  and _49543_ (_42409_, _42408_, _38135_);
  not _49544_ (_42410_, _42409_);
  and _49545_ (_42411_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _49546_ (_42412_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor _49547_ (_42413_, _42412_, _42411_);
  and _49548_ (_42414_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _49549_ (_42415_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor _49550_ (_42416_, _42415_, _42414_);
  and _49551_ (_42417_, _42416_, _42413_);
  and _49552_ (_42418_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _49553_ (_42419_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor _49554_ (_42420_, _42419_, _42418_);
  and _49555_ (_42421_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _49556_ (_42422_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _49557_ (_42423_, _42422_, _42421_);
  and _49558_ (_42424_, _42423_, _42420_);
  and _49559_ (_42425_, _42424_, _42417_);
  nor _49560_ (_42426_, _42425_, _42041_);
  and _49561_ (_42427_, _42041_, _39933_);
  nor _49562_ (_42428_, _42427_, _42426_);
  not _49563_ (_42429_, _42428_);
  and _49564_ (_42430_, _42429_, _42142_);
  not _49565_ (_42431_, _42430_);
  nor _49566_ (_42432_, _42020_, _37999_);
  and _49567_ (_42433_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _49568_ (_42434_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _49569_ (_42435_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _49570_ (_42436_, _42435_, _42434_);
  and _49571_ (_42437_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _49572_ (_42438_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _49573_ (_42439_, _42438_, _42437_);
  and _49574_ (_42440_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _49575_ (_42441_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _49576_ (_42442_, _42441_, _42440_);
  and _49577_ (_42443_, _42442_, _42439_);
  and _49578_ (_42444_, _42443_, _42436_);
  nor _49579_ (_42445_, _42444_, _42093_);
  nor _49580_ (_42446_, _42445_, _42433_);
  not _49581_ (_42447_, _42446_);
  and _49582_ (_42448_, _42447_, _42077_);
  nor _49583_ (_42449_, _42448_, _42432_);
  and _49584_ (_42450_, _42449_, _42431_);
  and _49585_ (_42451_, _42450_, _42410_);
  and _49586_ (_42452_, _42451_, _42117_);
  nor _49587_ (_42453_, _42355_, _42117_);
  nor _49588_ (_42454_, _42453_, _42452_);
  not _49589_ (_42455_, _42309_);
  or _49590_ (_42456_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _49591_ (_42457_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _49592_ (_42458_, _42457_, _42456_);
  or _49593_ (_42459_, _42458_, _42455_);
  and _49594_ (_42460_, _42459_, _42454_);
  and _49595_ (_42461_, _42460_, _42407_);
  and _49596_ (_42462_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and _49597_ (_42463_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _49598_ (_42464_, _42463_, _42455_);
  or _49599_ (_42465_, _42464_, _42462_);
  not _49600_ (_42466_, _42454_);
  and _49601_ (_42467_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and _49602_ (_42468_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _49603_ (_42469_, _42468_, _42309_);
  or _49604_ (_42470_, _42469_, _42467_);
  and _49605_ (_42471_, _42470_, _42466_);
  and _49606_ (_42472_, _42471_, _42465_);
  or _49607_ (_42473_, _42472_, _42461_);
  and _49608_ (_42474_, _42473_, _42215_);
  nor _49609_ (_42475_, _28244_, _27103_);
  nor _49610_ (_42476_, _42475_, _31190_);
  and _49611_ (_42477_, _28244_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49612_ (_42478_, _42477_, _40289_);
  nor _49613_ (_42479_, _27674_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _49614_ (_42480_, _42479_, _42478_);
  nand _49615_ (_42481_, _42480_, _42309_);
  or _49616_ (_42482_, _42480_, _42309_);
  and _49617_ (_42483_, _42482_, _42481_);
  not _49618_ (_42484_, _42483_);
  and _49619_ (_42485_, _42477_, _31790_);
  nor _49620_ (_42486_, _27795_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _49621_ (_42487_, _42486_, _42485_);
  not _49622_ (_42488_, _42487_);
  and _49623_ (_42489_, _42488_, _42402_);
  nor _49624_ (_42490_, _42488_, _42402_);
  nor _49625_ (_42491_, _42490_, _42489_);
  and _49626_ (_42492_, _42491_, _42484_);
  and _49627_ (_42493_, _42477_, _38138_);
  nor _49628_ (_42494_, _42477_, _27948_);
  nor _49629_ (_42495_, _42494_, _42493_);
  nor _49630_ (_42496_, _42495_, _42454_);
  and _49631_ (_42497_, _42495_, _42454_);
  nor _49632_ (_42498_, _42497_, _42496_);
  and _49633_ (_42499_, _42477_, _38613_);
  nor _49634_ (_42500_, _28069_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _49635_ (_42501_, _42500_, _42499_);
  not _49636_ (_42502_, _42501_);
  nor _49637_ (_42503_, _42502_, _42214_);
  and _49638_ (_42504_, _42502_, _42214_);
  nor _49639_ (_42505_, _42504_, _42503_);
  and _49640_ (_42506_, _42505_, _42498_);
  and _49641_ (_42507_, _42506_, _42492_);
  and _49642_ (_42508_, _42507_, _42476_);
  or _49643_ (_42509_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _49644_ (_42510_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and _49645_ (_42511_, _42510_, _42509_);
  or _49646_ (_42512_, _42511_, _42309_);
  or _49647_ (_42513_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _49648_ (_42514_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _49649_ (_42515_, _42514_, _42513_);
  or _49650_ (_42516_, _42515_, _42455_);
  and _49651_ (_42517_, _42516_, _42454_);
  and _49652_ (_42518_, _42517_, _42512_);
  and _49653_ (_42519_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and _49654_ (_42520_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _49655_ (_42521_, _42520_, _42455_);
  or _49656_ (_42522_, _42521_, _42519_);
  and _49657_ (_42523_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and _49658_ (_42524_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _49659_ (_42525_, _42524_, _42309_);
  or _49660_ (_42526_, _42525_, _42523_);
  and _49661_ (_42527_, _42526_, _42466_);
  and _49662_ (_42528_, _42527_, _42522_);
  or _49663_ (_42529_, _42528_, _42518_);
  and _49664_ (_42530_, _42529_, _42214_);
  or _49665_ (_42531_, _42530_, _42508_);
  or _49666_ (_42532_, _42531_, _42474_);
  nor _49667_ (_42533_, _42259_, _42117_);
  nor _49668_ (_42534_, _42477_, _27542_);
  not _49669_ (_42535_, _42534_);
  and _49670_ (_42536_, _42535_, _42533_);
  nor _49671_ (_42537_, _42535_, _42533_);
  nor _49672_ (_42538_, _42537_, _42536_);
  nor _49673_ (_42539_, _42165_, _42117_);
  nor _49674_ (_42540_, _42477_, _38613_);
  not _49675_ (_42541_, _42540_);
  nor _49676_ (_42542_, _42541_, _42539_);
  and _49677_ (_42543_, _42541_, _42539_);
  nor _49678_ (_42544_, _42543_, _42542_);
  and _49679_ (_42545_, _42544_, _42538_);
  nor _49680_ (_42546_, _42100_, _31779_);
  and _49681_ (_42547_, _42100_, _31779_);
  nor _49682_ (_42548_, _42547_, _42546_);
  nor _49683_ (_42549_, _42451_, _42117_);
  nor _49684_ (_42550_, _42477_, _28376_);
  not _49685_ (_42551_, _42550_);
  and _49686_ (_42552_, _42551_, _42549_);
  nor _49687_ (_42553_, _42551_, _42549_);
  nor _49688_ (_42554_, _42553_, _42552_);
  and _49689_ (_42555_, _42554_, _42548_);
  and _49690_ (_42557_, _42555_, _42545_);
  and _49691_ (_42558_, _42557_, _42508_);
  not _49692_ (_42560_, _42558_);
  or _49693_ (_42562_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not _49694_ (_42563_, _42508_);
  nor _49695_ (_42565_, _42558_, _42563_);
  nor _49696_ (_42567_, _42565_, rst);
  and _49697_ (_42569_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _49698_ (_42571_, _42569_, _28935_);
  nor _49699_ (_42572_, _42571_, _31757_);
  nand _49700_ (_42573_, _28935_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _49701_ (_42574_, _20601_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49702_ (_42575_, _42574_, _42573_);
  nor _49703_ (_42576_, _38225_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _49704_ (_42577_, _42576_, _42575_);
  or _49705_ (_42578_, _42577_, _42572_);
  and _49706_ (_39844_, _42578_, _42618_);
  or _49707_ (_42579_, _39844_, _42567_);
  and _49708_ (_42580_, _42579_, _42562_);
  and _49709_ (_02564_, _42580_, _42532_);
  not _49710_ (_42581_, _42476_);
  nor _49711_ (_42582_, _42487_, _42581_);
  nor _49712_ (_42583_, _42581_, _42480_);
  and _49713_ (_42584_, _42583_, _42582_);
  nor _49714_ (_42585_, _42495_, _42581_);
  nor _49715_ (_42586_, _42581_, _42501_);
  and _49716_ (_42587_, _42586_, _42585_);
  and _49717_ (_42588_, _42587_, _42584_);
  and _49718_ (_42589_, _42578_, _42476_);
  and _49719_ (_42590_, _42589_, _42588_);
  not _49720_ (_42591_, _42588_);
  and _49721_ (_42592_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _49722_ (_02574_, _42592_, _42590_);
  nor _49723_ (_42593_, _42586_, _42585_);
  nor _49724_ (_42594_, _42583_, _42582_);
  and _49725_ (_42595_, _42594_, _42476_);
  and _49726_ (_42596_, _42595_, _42593_);
  not _49727_ (_42597_, _42596_);
  and _49728_ (_42598_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _49729_ (_42599_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _29012_);
  and _49730_ (_42600_, _42599_, _28957_);
  not _49731_ (_42601_, _42600_);
  nor _49732_ (_42602_, _42601_, _31757_);
  not _49733_ (_42603_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _49734_ (_42604_, _38203_, _42603_);
  or _49735_ (_42606_, _19441_, _42603_);
  and _49736_ (_42608_, _42606_, _42601_);
  and _49737_ (_42610_, _42608_, _42604_);
  or _49738_ (_42612_, _42610_, _42602_);
  and _49739_ (_42614_, _42612_, _42596_);
  or _49740_ (_02798_, _42614_, _42598_);
  and _49741_ (_42617_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nand _49742_ (_42619_, _42599_, _28912_);
  nor _49743_ (_42620_, _42619_, _31757_);
  nor _49744_ (_42622_, _38191_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49745_ (_42624_, _42599_, _28847_);
  and _49746_ (_42625_, _42599_, _28935_);
  or _49747_ (_42626_, _42625_, _42569_);
  or _49748_ (_42627_, _42626_, _42624_);
  and _49749_ (_42628_, _42627_, _20427_);
  or _49750_ (_42629_, _42628_, _42622_);
  or _49751_ (_42630_, _42629_, _42620_);
  and _49752_ (_42631_, _42630_, _42596_);
  or _49753_ (_02803_, _42631_, _42617_);
  and _49754_ (_42632_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand _49755_ (_42633_, _42599_, _28858_);
  nor _49756_ (_42634_, _42633_, _31757_);
  nor _49757_ (_42635_, _38184_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49758_ (_42636_, _42599_, _28891_);
  or _49759_ (_42637_, _42636_, _42626_);
  and _49760_ (_42638_, _42637_, _19080_);
  or _49761_ (_42639_, _42638_, _42635_);
  or _49762_ (_42640_, _42639_, _42634_);
  and _49763_ (_42641_, _42640_, _42596_);
  or _49764_ (_02809_, _42641_, _42632_);
  and _49765_ (_42642_, _42625_, _32410_);
  nor _49766_ (_42643_, _38177_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _49767_ (_42644_, _42624_, _42569_);
  or _49768_ (_42645_, _42644_, _42636_);
  and _49769_ (_42646_, _42645_, _20112_);
  or _49770_ (_42647_, _42646_, _42643_);
  or _49771_ (_42648_, _42647_, _42642_);
  and _49772_ (_42649_, _42648_, _42596_);
  and _49773_ (_42650_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or _49774_ (_02814_, _42650_, _42649_);
  nand _49775_ (_42651_, _42569_, _28957_);
  nor _49776_ (_42652_, _42651_, _31757_);
  nor _49777_ (_42653_, _38169_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _49778_ (_42654_, _28957_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _49779_ (_42655_, _19277_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49780_ (_42656_, _42655_, _42654_);
  or _49781_ (_42657_, _42656_, _42653_);
  or _49782_ (_42658_, _42657_, _42652_);
  and _49783_ (_42659_, _42658_, _42596_);
  and _49784_ (_42660_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _49785_ (_02819_, _42660_, _42659_);
  nand _49786_ (_42661_, _42569_, _28912_);
  nor _49787_ (_42662_, _42661_, _31757_);
  nor _49788_ (_42663_, _38162_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _49789_ (_42664_, _28912_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _49790_ (_42665_, _20264_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49791_ (_42666_, _42665_, _42664_);
  or _49792_ (_42667_, _42666_, _42663_);
  or _49793_ (_42668_, _42667_, _42662_);
  and _49794_ (_42669_, _42668_, _42596_);
  and _49795_ (_42670_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _49796_ (_02824_, _42670_, _42669_);
  and _49797_ (_42671_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand _49798_ (_42672_, _42569_, _28858_);
  nor _49799_ (_42673_, _42672_, _31757_);
  nor _49800_ (_42674_, _38155_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _49801_ (_42675_, _28858_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _49802_ (_42676_, _19615_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49803_ (_42677_, _42676_, _42675_);
  or _49804_ (_42678_, _42677_, _42674_);
  or _49805_ (_42679_, _42678_, _42673_);
  and _49806_ (_42680_, _42679_, _42596_);
  or _49807_ (_02829_, _42680_, _42671_);
  and _49808_ (_42681_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and _49809_ (_42682_, _42596_, _42578_);
  or _49810_ (_02831_, _42682_, _42681_);
  and _49811_ (_42683_, _42612_, _42476_);
  and _49812_ (_42684_, _42582_, _42480_);
  and _49813_ (_42685_, _42684_, _42593_);
  and _49814_ (_42686_, _42685_, _42683_);
  not _49815_ (_42687_, _42685_);
  and _49816_ (_42688_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _49817_ (_02839_, _42688_, _42686_);
  and _49818_ (_42689_, _42630_, _42476_);
  and _49819_ (_42690_, _42685_, _42689_);
  and _49820_ (_42691_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _49821_ (_02842_, _42691_, _42690_);
  and _49822_ (_42692_, _42640_, _42476_);
  and _49823_ (_42693_, _42685_, _42692_);
  and _49824_ (_42694_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _49825_ (_02846_, _42694_, _42693_);
  and _49826_ (_42695_, _42648_, _42476_);
  and _49827_ (_42696_, _42685_, _42695_);
  and _49828_ (_42697_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _49829_ (_02850_, _42697_, _42696_);
  and _49830_ (_42698_, _42658_, _42476_);
  and _49831_ (_42699_, _42685_, _42698_);
  and _49832_ (_42700_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or _49833_ (_02853_, _42700_, _42699_);
  and _49834_ (_42701_, _42668_, _42476_);
  and _49835_ (_42702_, _42685_, _42701_);
  and _49836_ (_42703_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or _49837_ (_02856_, _42703_, _42702_);
  and _49838_ (_42704_, _42679_, _42476_);
  and _49839_ (_42705_, _42685_, _42704_);
  and _49840_ (_42706_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _49841_ (_02860_, _42706_, _42705_);
  and _49842_ (_42707_, _42685_, _42589_);
  and _49843_ (_42708_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _49844_ (_02862_, _42708_, _42707_);
  and _49845_ (_42709_, _42583_, _42487_);
  and _49846_ (_42710_, _42709_, _42593_);
  and _49847_ (_42711_, _42710_, _42683_);
  not _49848_ (_42712_, _42710_);
  and _49849_ (_42713_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _49850_ (_02868_, _42713_, _42711_);
  and _49851_ (_42714_, _42710_, _42689_);
  and _49852_ (_42715_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _49853_ (_02873_, _42715_, _42714_);
  and _49854_ (_42716_, _42710_, _42692_);
  and _49855_ (_42717_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _49856_ (_02876_, _42717_, _42716_);
  and _49857_ (_42718_, _42710_, _42695_);
  and _49858_ (_42719_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _49859_ (_02879_, _42719_, _42718_);
  and _49860_ (_42720_, _42710_, _42698_);
  and _49861_ (_42721_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _49862_ (_02884_, _42721_, _42720_);
  and _49863_ (_42722_, _42710_, _42701_);
  and _49864_ (_42723_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _49865_ (_02887_, _42723_, _42722_);
  and _49866_ (_42724_, _42710_, _42704_);
  and _49867_ (_42725_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _49868_ (_02890_, _42725_, _42724_);
  and _49869_ (_42726_, _42710_, _42589_);
  and _49870_ (_42727_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _49871_ (_02893_, _42727_, _42726_);
  and _49872_ (_42728_, _42593_, _42584_);
  and _49873_ (_42729_, _42728_, _42683_);
  not _49874_ (_42730_, _42728_);
  and _49875_ (_42731_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _49876_ (_02898_, _42731_, _42729_);
  and _49877_ (_42732_, _42728_, _42689_);
  and _49878_ (_42733_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _49879_ (_02902_, _42733_, _42732_);
  and _49880_ (_42734_, _42728_, _42692_);
  and _49881_ (_42735_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _49882_ (_02905_, _42735_, _42734_);
  and _49883_ (_42736_, _42728_, _42695_);
  and _49884_ (_42737_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _49885_ (_02908_, _42737_, _42736_);
  and _49886_ (_42738_, _42728_, _42698_);
  and _49887_ (_42739_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _49888_ (_02911_, _42739_, _42738_);
  and _49889_ (_42740_, _42728_, _42701_);
  and _49890_ (_42741_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _49891_ (_02915_, _42741_, _42740_);
  and _49892_ (_42742_, _42728_, _42704_);
  and _49893_ (_42743_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _49894_ (_02918_, _42743_, _42742_);
  and _49895_ (_42744_, _42728_, _42589_);
  and _49896_ (_42745_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _49897_ (_02921_, _42745_, _42744_);
  and _49898_ (_42746_, _42586_, _42495_);
  and _49899_ (_42747_, _42746_, _42594_);
  and _49900_ (_42748_, _42747_, _42683_);
  not _49901_ (_42749_, _42747_);
  and _49902_ (_42750_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _49903_ (_02929_, _42750_, _42748_);
  and _49904_ (_42751_, _42747_, _42689_);
  and _49905_ (_42752_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _49906_ (_02933_, _42752_, _42751_);
  and _49907_ (_42753_, _42747_, _42692_);
  and _49908_ (_42754_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _49909_ (_02937_, _42754_, _42753_);
  and _49910_ (_42755_, _42747_, _42695_);
  and _49911_ (_42756_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _49912_ (_02941_, _42756_, _42755_);
  and _49913_ (_42757_, _42747_, _42698_);
  and _49914_ (_42758_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _49915_ (_02945_, _42758_, _42757_);
  and _49916_ (_42759_, _42747_, _42701_);
  and _49917_ (_42760_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _49918_ (_02948_, _42760_, _42759_);
  and _49919_ (_42761_, _42747_, _42704_);
  and _49920_ (_42762_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _49921_ (_02952_, _42762_, _42761_);
  and _49922_ (_42763_, _42747_, _42589_);
  and _49923_ (_42764_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _49924_ (_02956_, _42764_, _42763_);
  and _49925_ (_42765_, _42746_, _42684_);
  and _49926_ (_42766_, _42765_, _42683_);
  not _49927_ (_42767_, _42765_);
  and _49928_ (_42768_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _49929_ (_02960_, _42768_, _42766_);
  and _49930_ (_42769_, _42765_, _42689_);
  and _49931_ (_42770_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _49932_ (_02964_, _42770_, _42769_);
  and _49933_ (_42771_, _42765_, _42692_);
  and _49934_ (_42772_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or _49935_ (_02969_, _42772_, _42771_);
  and _49936_ (_42773_, _42765_, _42695_);
  and _49937_ (_42774_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _49938_ (_02973_, _42774_, _42773_);
  and _49939_ (_42775_, _42765_, _42698_);
  and _49940_ (_42776_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or _49941_ (_02977_, _42776_, _42775_);
  and _49942_ (_42777_, _42765_, _42701_);
  and _49943_ (_42778_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or _49944_ (_02982_, _42778_, _42777_);
  and _49945_ (_42779_, _42765_, _42704_);
  and _49946_ (_42780_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or _49947_ (_02986_, _42780_, _42779_);
  and _49948_ (_42781_, _42765_, _42589_);
  and _49949_ (_42782_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _49950_ (_02988_, _42782_, _42781_);
  and _49951_ (_42783_, _42746_, _42709_);
  and _49952_ (_42784_, _42783_, _42683_);
  not _49953_ (_42785_, _42783_);
  and _49954_ (_42786_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _49955_ (_02993_, _42786_, _42784_);
  and _49956_ (_42787_, _42783_, _42689_);
  and _49957_ (_42788_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _49958_ (_02998_, _42788_, _42787_);
  and _49959_ (_42789_, _42783_, _42692_);
  and _49960_ (_42790_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _49961_ (_03002_, _42790_, _42789_);
  and _49962_ (_42791_, _42783_, _42695_);
  and _49963_ (_42792_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _49964_ (_03005_, _42792_, _42791_);
  and _49965_ (_42793_, _42783_, _42698_);
  and _49966_ (_42794_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _49967_ (_03010_, _42794_, _42793_);
  and _49968_ (_42795_, _42783_, _42701_);
  and _49969_ (_42796_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _49970_ (_03014_, _42796_, _42795_);
  and _49971_ (_42797_, _42783_, _42704_);
  and _49972_ (_42798_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _49973_ (_03017_, _42798_, _42797_);
  and _49974_ (_42799_, _42783_, _42589_);
  and _49975_ (_42800_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _49976_ (_03020_, _42800_, _42799_);
  and _49977_ (_42801_, _42746_, _42584_);
  and _49978_ (_42802_, _42801_, _42683_);
  not _49979_ (_42803_, _42801_);
  and _49980_ (_42804_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _49981_ (_03026_, _42804_, _42802_);
  and _49982_ (_42805_, _42801_, _42689_);
  and _49983_ (_42806_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _49984_ (_03030_, _42806_, _42805_);
  and _49985_ (_42807_, _42801_, _42692_);
  and _49986_ (_42808_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _49987_ (_03033_, _42808_, _42807_);
  and _49988_ (_42809_, _42801_, _42695_);
  and _49989_ (_42810_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _49990_ (_03037_, _42810_, _42809_);
  and _49991_ (_42811_, _42801_, _42698_);
  and _49992_ (_42812_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _49993_ (_03040_, _42812_, _42811_);
  and _49994_ (_42813_, _42801_, _42701_);
  and _49995_ (_42814_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _49996_ (_03043_, _42814_, _42813_);
  and _49997_ (_42815_, _42801_, _42704_);
  and _49998_ (_42816_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _49999_ (_03046_, _42816_, _42815_);
  and _50000_ (_42817_, _42801_, _42589_);
  and _50001_ (_42818_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _50002_ (_03049_, _42818_, _42817_);
  and _50003_ (_42819_, _42585_, _42501_);
  and _50004_ (_42820_, _42819_, _42594_);
  and _50005_ (_42821_, _42820_, _42683_);
  not _50006_ (_42822_, _42820_);
  and _50007_ (_42823_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or _50008_ (_03055_, _42823_, _42821_);
  and _50009_ (_42824_, _42820_, _42689_);
  and _50010_ (_42825_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _50011_ (_03058_, _42825_, _42824_);
  and _50012_ (_42826_, _42820_, _42692_);
  and _50013_ (_42827_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or _50014_ (_03062_, _42827_, _42826_);
  and _50015_ (_42828_, _42820_, _42695_);
  and _50016_ (_42829_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or _50017_ (_03065_, _42829_, _42828_);
  and _50018_ (_42830_, _42820_, _42698_);
  and _50019_ (_42831_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _50020_ (_03069_, _42831_, _42830_);
  and _50021_ (_42832_, _42820_, _42701_);
  and _50022_ (_42833_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _50023_ (_03072_, _42833_, _42832_);
  and _50024_ (_42834_, _42820_, _42704_);
  and _50025_ (_42835_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or _50026_ (_03076_, _42835_, _42834_);
  and _50027_ (_42836_, _42820_, _42589_);
  and _50028_ (_42837_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _50029_ (_03079_, _42837_, _42836_);
  and _50030_ (_42838_, _42819_, _42684_);
  and _50031_ (_42839_, _42838_, _42683_);
  not _50032_ (_42840_, _42838_);
  and _50033_ (_42841_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _50034_ (_03083_, _42841_, _42839_);
  and _50035_ (_42842_, _42838_, _42689_);
  and _50036_ (_42843_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _50037_ (_03087_, _42843_, _42842_);
  and _50038_ (_42844_, _42838_, _42692_);
  and _50039_ (_42845_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _50040_ (_03090_, _42845_, _42844_);
  and _50041_ (_42846_, _42838_, _42695_);
  and _50042_ (_42847_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _50043_ (_03094_, _42847_, _42846_);
  and _50044_ (_42848_, _42838_, _42698_);
  and _50045_ (_42849_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _50046_ (_03097_, _42849_, _42848_);
  and _50047_ (_42850_, _42838_, _42701_);
  and _50048_ (_42851_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _50049_ (_03101_, _42851_, _42850_);
  and _50050_ (_42852_, _42838_, _42704_);
  and _50051_ (_42853_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _50052_ (_03104_, _42853_, _42852_);
  and _50053_ (_42854_, _42838_, _42589_);
  and _50054_ (_42855_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _50055_ (_03107_, _42855_, _42854_);
  and _50056_ (_42856_, _42819_, _42709_);
  and _50057_ (_42857_, _42856_, _42683_);
  not _50058_ (_42858_, _42856_);
  and _50059_ (_42859_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _50060_ (_03112_, _42859_, _42857_);
  and _50061_ (_42860_, _42856_, _42689_);
  and _50062_ (_42861_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _50063_ (_03115_, _42861_, _42860_);
  and _50064_ (_42862_, _42856_, _42692_);
  and _50065_ (_42863_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _50066_ (_03119_, _42863_, _42862_);
  and _50067_ (_42864_, _42856_, _42695_);
  and _50068_ (_42865_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _50069_ (_03122_, _42865_, _42864_);
  and _50070_ (_42866_, _42856_, _42698_);
  and _50071_ (_42867_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _50072_ (_03126_, _42867_, _42866_);
  and _50073_ (_42868_, _42856_, _42701_);
  and _50074_ (_42869_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _50075_ (_03130_, _42869_, _42868_);
  and _50076_ (_42870_, _42856_, _42704_);
  and _50077_ (_42871_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _50078_ (_03133_, _42871_, _42870_);
  and _50079_ (_42872_, _42856_, _42589_);
  and _50080_ (_42873_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _50081_ (_03136_, _42873_, _42872_);
  and _50082_ (_42874_, _42819_, _42584_);
  and _50083_ (_42875_, _42874_, _42683_);
  not _50084_ (_42876_, _42874_);
  and _50085_ (_42877_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or _50086_ (_03140_, _42877_, _42875_);
  and _50087_ (_42878_, _42874_, _42689_);
  and _50088_ (_42879_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _50089_ (_03143_, _42879_, _42878_);
  and _50090_ (_42880_, _42874_, _42692_);
  and _50091_ (_42881_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or _50092_ (_03146_, _42881_, _42880_);
  and _50093_ (_42882_, _42874_, _42695_);
  and _50094_ (_42883_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _50095_ (_03149_, _42883_, _42882_);
  and _50096_ (_42884_, _42874_, _42698_);
  and _50097_ (_42885_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or _50098_ (_03153_, _42885_, _42884_);
  and _50099_ (_42886_, _42874_, _42701_);
  and _50100_ (_42887_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or _50101_ (_03156_, _42887_, _42886_);
  and _50102_ (_42888_, _42874_, _42704_);
  and _50103_ (_42889_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or _50104_ (_03159_, _42889_, _42888_);
  and _50105_ (_42890_, _42874_, _42589_);
  and _50106_ (_42891_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _50107_ (_03162_, _42891_, _42890_);
  and _50108_ (_42892_, _42594_, _42587_);
  and _50109_ (_42893_, _42892_, _42683_);
  not _50110_ (_42894_, _42892_);
  and _50111_ (_42895_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or _50112_ (_03166_, _42895_, _42893_);
  and _50113_ (_42896_, _42892_, _42689_);
  and _50114_ (_42897_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _50115_ (_03170_, _42897_, _42896_);
  and _50116_ (_42898_, _42892_, _42692_);
  and _50117_ (_42899_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or _50118_ (_03173_, _42899_, _42898_);
  and _50119_ (_42900_, _42892_, _42695_);
  and _50120_ (_42901_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or _50121_ (_03176_, _42901_, _42900_);
  and _50122_ (_42902_, _42892_, _42698_);
  and _50123_ (_42903_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or _50124_ (_03179_, _42903_, _42902_);
  and _50125_ (_42904_, _42892_, _42701_);
  and _50126_ (_42905_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or _50127_ (_03183_, _42905_, _42904_);
  and _50128_ (_42906_, _42892_, _42704_);
  and _50129_ (_42907_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or _50130_ (_03186_, _42907_, _42906_);
  and _50131_ (_42908_, _42892_, _42589_);
  and _50132_ (_42909_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _50133_ (_03188_, _42909_, _42908_);
  and _50134_ (_42910_, _42684_, _42587_);
  and _50135_ (_42911_, _42910_, _42683_);
  not _50136_ (_42912_, _42910_);
  and _50137_ (_42913_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _50138_ (_03193_, _42913_, _42911_);
  and _50139_ (_42914_, _42910_, _42689_);
  and _50140_ (_42915_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _50141_ (_03196_, _42915_, _42914_);
  and _50142_ (_42916_, _42910_, _42692_);
  and _50143_ (_42917_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _50144_ (_03200_, _42917_, _42916_);
  and _50145_ (_42918_, _42910_, _42695_);
  and _50146_ (_42919_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _50147_ (_03204_, _42919_, _42918_);
  and _50148_ (_42920_, _42910_, _42698_);
  and _50149_ (_42921_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _50150_ (_03207_, _42921_, _42920_);
  and _50151_ (_42922_, _42910_, _42701_);
  and _50152_ (_42923_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _50153_ (_03211_, _42923_, _42922_);
  and _50154_ (_42924_, _42910_, _42704_);
  and _50155_ (_42925_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _50156_ (_03214_, _42925_, _42924_);
  and _50157_ (_42926_, _42910_, _42589_);
  and _50158_ (_42927_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _50159_ (_03217_, _42927_, _42926_);
  and _50160_ (_42928_, _42709_, _42587_);
  and _50161_ (_42929_, _42928_, _42683_);
  not _50162_ (_42930_, _42928_);
  and _50163_ (_42931_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _50164_ (_03221_, _42931_, _42929_);
  and _50165_ (_42932_, _42928_, _42689_);
  and _50166_ (_42933_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _50167_ (_03225_, _42933_, _42932_);
  and _50168_ (_42934_, _42928_, _42692_);
  and _50169_ (_42935_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _50170_ (_03228_, _42935_, _42934_);
  and _50171_ (_42936_, _42928_, _42695_);
  and _50172_ (_42937_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _50173_ (_03232_, _42937_, _42936_);
  and _50174_ (_42938_, _42928_, _42698_);
  and _50175_ (_42939_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _50176_ (_03235_, _42939_, _42938_);
  and _50177_ (_42940_, _42928_, _42701_);
  and _50178_ (_42941_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _50179_ (_03238_, _42941_, _42940_);
  and _50180_ (_42942_, _42928_, _42704_);
  and _50181_ (_42943_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _50182_ (_03242_, _42943_, _42942_);
  and _50183_ (_42944_, _42928_, _42589_);
  and _50184_ (_42945_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _50185_ (_03244_, _42945_, _42944_);
  and _50186_ (_42946_, _42683_, _42588_);
  and _50187_ (_42947_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or _50188_ (_03248_, _42947_, _42946_);
  and _50189_ (_42948_, _42689_, _42588_);
  and _50190_ (_42949_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or _50191_ (_03251_, _42949_, _42948_);
  and _50192_ (_42950_, _42692_, _42588_);
  and _50193_ (_42951_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or _50194_ (_03255_, _42951_, _42950_);
  and _50195_ (_42952_, _42695_, _42588_);
  and _50196_ (_42953_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _50197_ (_03258_, _42953_, _42952_);
  and _50198_ (_42954_, _42698_, _42588_);
  and _50199_ (_42955_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or _50200_ (_03261_, _42955_, _42954_);
  and _50201_ (_42956_, _42701_, _42588_);
  and _50202_ (_42957_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or _50203_ (_03264_, _42957_, _42956_);
  and _50204_ (_42958_, _42704_, _42588_);
  and _50205_ (_42959_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or _50206_ (_03268_, _42959_, _42958_);
  and _50207_ (_42960_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and _50208_ (_42961_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _50209_ (_42962_, _42961_, _42309_);
  or _50210_ (_42963_, _42962_, _42960_);
  and _50211_ (_42964_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _50212_ (_42965_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _50213_ (_42966_, _42965_, _42455_);
  or _50214_ (_42967_, _42966_, _42964_);
  and _50215_ (_42968_, _42967_, _42963_);
  or _50216_ (_42969_, _42968_, _42215_);
  and _50217_ (_42970_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and _50218_ (_42971_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _50219_ (_42972_, _42971_, _42309_);
  or _50220_ (_42973_, _42972_, _42970_);
  and _50221_ (_42974_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and _50222_ (_42975_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _50223_ (_42976_, _42975_, _42455_);
  or _50224_ (_42977_, _42976_, _42974_);
  and _50225_ (_42978_, _42977_, _42973_);
  or _50226_ (_42979_, _42978_, _42214_);
  and _50227_ (_42980_, _42979_, _42466_);
  and _50228_ (_42981_, _42980_, _42969_);
  or _50229_ (_42982_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or _50230_ (_42983_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _50231_ (_42984_, _42983_, _42982_);
  or _50232_ (_42985_, _42984_, _42455_);
  or _50233_ (_42986_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or _50234_ (_42987_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and _50235_ (_42988_, _42987_, _42986_);
  or _50236_ (_42989_, _42988_, _42309_);
  and _50237_ (_42990_, _42989_, _42985_);
  or _50238_ (_42991_, _42990_, _42215_);
  or _50239_ (_42992_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or _50240_ (_42993_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _50241_ (_42994_, _42993_, _42992_);
  or _50242_ (_42995_, _42994_, _42455_);
  or _50243_ (_42996_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or _50244_ (_42997_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and _50245_ (_42998_, _42997_, _42996_);
  or _50246_ (_42999_, _42998_, _42309_);
  and _50247_ (_43000_, _42999_, _42995_);
  or _50248_ (_43001_, _43000_, _42214_);
  and _50249_ (_43002_, _43001_, _42454_);
  and _50250_ (_43003_, _43002_, _42991_);
  or _50251_ (_43004_, _43003_, _42981_);
  and _50252_ (_43005_, _43004_, _42560_);
  and _50253_ (_43006_, _42558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or _50254_ (_43007_, _43006_, _42565_);
  or _50255_ (_43008_, _43007_, _43005_);
  and _50256_ (_39864_, _42612_, _42618_);
  or _50257_ (_43009_, _39864_, _42567_);
  and _50258_ (_05053_, _43009_, _43008_);
  and _50259_ (_43010_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and _50260_ (_43011_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _50261_ (_43012_, _43011_, _42309_);
  or _50262_ (_43013_, _43012_, _43010_);
  and _50263_ (_43014_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and _50264_ (_43015_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _50265_ (_43016_, _43015_, _42455_);
  or _50266_ (_43017_, _43016_, _43014_);
  and _50267_ (_43018_, _43017_, _43013_);
  or _50268_ (_43019_, _43018_, _42215_);
  and _50269_ (_43020_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and _50270_ (_43021_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _50271_ (_43022_, _43021_, _42309_);
  or _50272_ (_43023_, _43022_, _43020_);
  and _50273_ (_43024_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and _50274_ (_43025_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _50275_ (_43026_, _43025_, _42455_);
  or _50276_ (_43027_, _43026_, _43024_);
  and _50277_ (_43028_, _43027_, _43023_);
  or _50278_ (_43029_, _43028_, _42214_);
  and _50279_ (_43030_, _43029_, _42466_);
  and _50280_ (_43031_, _43030_, _43019_);
  or _50281_ (_43032_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _50282_ (_43033_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _50283_ (_43034_, _43033_, _43032_);
  or _50284_ (_43035_, _43034_, _42455_);
  or _50285_ (_43036_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _50286_ (_43037_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and _50287_ (_43038_, _43037_, _43036_);
  or _50288_ (_43039_, _43038_, _42309_);
  and _50289_ (_43040_, _43039_, _43035_);
  or _50290_ (_43041_, _43040_, _42215_);
  or _50291_ (_43042_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _50292_ (_43043_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _50293_ (_43044_, _43043_, _43042_);
  or _50294_ (_43045_, _43044_, _42455_);
  or _50295_ (_43046_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or _50296_ (_43047_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and _50297_ (_43048_, _43047_, _43046_);
  or _50298_ (_43049_, _43048_, _42309_);
  and _50299_ (_43050_, _43049_, _43045_);
  or _50300_ (_43051_, _43050_, _42214_);
  and _50301_ (_43052_, _43051_, _42454_);
  and _50302_ (_43053_, _43052_, _43041_);
  or _50303_ (_43054_, _43053_, _43031_);
  or _50304_ (_43055_, _43054_, _42558_);
  or _50305_ (_43056_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _50306_ (_43057_, _43056_, _42567_);
  and _50307_ (_43058_, _43057_, _43055_);
  and _50308_ (_39865_, _42630_, _42618_);
  and _50309_ (_43059_, _39865_, _42565_);
  or _50310_ (_05055_, _43059_, _43058_);
  and _50311_ (_43060_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and _50312_ (_43061_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _50313_ (_43062_, _43061_, _42309_);
  or _50314_ (_43063_, _43062_, _43060_);
  and _50315_ (_43064_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _50316_ (_43065_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _50317_ (_43066_, _43065_, _42455_);
  or _50318_ (_43067_, _43066_, _43064_);
  and _50319_ (_43068_, _43067_, _43063_);
  or _50320_ (_43069_, _43068_, _42215_);
  and _50321_ (_43070_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and _50322_ (_43071_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _50323_ (_43072_, _43071_, _42309_);
  or _50324_ (_43073_, _43072_, _43070_);
  and _50325_ (_43074_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and _50326_ (_43075_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or _50327_ (_43076_, _43075_, _42455_);
  or _50328_ (_43077_, _43076_, _43074_);
  and _50329_ (_43078_, _43077_, _43073_);
  or _50330_ (_43079_, _43078_, _42214_);
  and _50331_ (_43080_, _43079_, _42466_);
  and _50332_ (_43081_, _43080_, _43069_);
  or _50333_ (_43082_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or _50334_ (_43083_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _50335_ (_43084_, _43083_, _43082_);
  or _50336_ (_43085_, _43084_, _42455_);
  or _50337_ (_43086_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or _50338_ (_43087_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and _50339_ (_43088_, _43087_, _43086_);
  or _50340_ (_43089_, _43088_, _42309_);
  and _50341_ (_43090_, _43089_, _43085_);
  or _50342_ (_43091_, _43090_, _42215_);
  or _50343_ (_43092_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or _50344_ (_43093_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _50345_ (_43094_, _43093_, _43092_);
  or _50346_ (_43095_, _43094_, _42455_);
  or _50347_ (_43096_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or _50348_ (_43097_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and _50349_ (_43098_, _43097_, _43096_);
  or _50350_ (_43099_, _43098_, _42309_);
  and _50351_ (_43100_, _43099_, _43095_);
  or _50352_ (_43101_, _43100_, _42214_);
  and _50353_ (_43102_, _43101_, _42454_);
  and _50354_ (_43103_, _43102_, _43091_);
  or _50355_ (_43104_, _43103_, _43081_);
  or _50356_ (_43105_, _43104_, _42558_);
  or _50357_ (_43106_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _50358_ (_43107_, _43106_, _42567_);
  and _50359_ (_43108_, _43107_, _43105_);
  and _50360_ (_39866_, _42640_, _42618_);
  and _50361_ (_43109_, _39866_, _42565_);
  or _50362_ (_05057_, _43109_, _43108_);
  and _50363_ (_43110_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _50364_ (_43111_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _50365_ (_43112_, _43111_, _42455_);
  or _50366_ (_43113_, _43112_, _43110_);
  and _50367_ (_43114_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and _50368_ (_43115_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _50369_ (_43116_, _43115_, _42309_);
  or _50370_ (_43117_, _43116_, _43114_);
  and _50371_ (_43118_, _43117_, _43113_);
  or _50372_ (_43119_, _43118_, _42215_);
  and _50373_ (_43120_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and _50374_ (_43121_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _50375_ (_43122_, _43121_, _42309_);
  or _50376_ (_43123_, _43122_, _43120_);
  and _50377_ (_43124_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and _50378_ (_43125_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _50379_ (_43126_, _43125_, _42455_);
  or _50380_ (_43127_, _43126_, _43124_);
  and _50381_ (_43128_, _43127_, _43123_);
  or _50382_ (_43129_, _43128_, _42214_);
  and _50383_ (_43130_, _43129_, _42466_);
  and _50384_ (_43131_, _43130_, _43119_);
  and _50385_ (_43132_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _50386_ (_43133_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _50387_ (_43134_, _43133_, _42309_);
  or _50388_ (_43135_, _43134_, _43132_);
  and _50389_ (_43136_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and _50390_ (_43137_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _50391_ (_43138_, _43137_, _42455_);
  or _50392_ (_43139_, _43138_, _43136_);
  and _50393_ (_43140_, _43139_, _43135_);
  or _50394_ (_43141_, _43140_, _42215_);
  and _50395_ (_43142_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _50396_ (_43143_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _50397_ (_43144_, _43143_, _42309_);
  or _50398_ (_43145_, _43144_, _43142_);
  and _50399_ (_43146_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _50400_ (_43147_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _50401_ (_43148_, _43147_, _42455_);
  or _50402_ (_43149_, _43148_, _43146_);
  and _50403_ (_43150_, _43149_, _43145_);
  or _50404_ (_43151_, _43150_, _42214_);
  and _50405_ (_43152_, _43151_, _42454_);
  and _50406_ (_43158_, _43152_, _43141_);
  or _50407_ (_43162_, _43158_, _43131_);
  and _50408_ (_43169_, _43162_, _42563_);
  and _50409_ (_43177_, _42648_, _42565_);
  and _50410_ (_43181_, _42558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or _50411_ (_43186_, _43181_, _43177_);
  or _50412_ (_43194_, _43186_, _43169_);
  and _50413_ (_05059_, _43194_, _42618_);
  and _50414_ (_43203_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and _50415_ (_43210_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or _50416_ (_43218_, _43210_, _42455_);
  or _50417_ (_43222_, _43218_, _43203_);
  and _50418_ (_43227_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and _50419_ (_43235_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _50420_ (_43241_, _43235_, _42309_);
  or _50421_ (_43244_, _43241_, _43227_);
  and _50422_ (_43248_, _43244_, _43222_);
  or _50423_ (_43259_, _43248_, _42215_);
  and _50424_ (_43263_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and _50425_ (_43270_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _50426_ (_43278_, _43270_, _42309_);
  or _50427_ (_43282_, _43278_, _43263_);
  and _50428_ (_43287_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and _50429_ (_43295_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or _50430_ (_43301_, _43295_, _42455_);
  or _50431_ (_43305_, _43301_, _43287_);
  and _50432_ (_43312_, _43305_, _43282_);
  or _50433_ (_43320_, _43312_, _42214_);
  and _50434_ (_43324_, _43320_, _42466_);
  and _50435_ (_43329_, _43324_, _43259_);
  and _50436_ (_43337_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _50437_ (_43343_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _50438_ (_43346_, _43343_, _42309_);
  or _50439_ (_43347_, _43346_, _43337_);
  and _50440_ (_43348_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _50441_ (_43349_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _50442_ (_43350_, _43349_, _42455_);
  or _50443_ (_43351_, _43350_, _43348_);
  and _50444_ (_43352_, _43351_, _43347_);
  or _50445_ (_43353_, _43352_, _42215_);
  and _50446_ (_43354_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _50447_ (_43355_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _50448_ (_43356_, _43355_, _42309_);
  or _50449_ (_43357_, _43356_, _43354_);
  and _50450_ (_43358_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _50451_ (_43359_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _50452_ (_43360_, _43359_, _42455_);
  or _50453_ (_43361_, _43360_, _43358_);
  and _50454_ (_43362_, _43361_, _43357_);
  or _50455_ (_43363_, _43362_, _42214_);
  and _50456_ (_43364_, _43363_, _42454_);
  and _50457_ (_43365_, _43364_, _43353_);
  or _50458_ (_43366_, _43365_, _43329_);
  and _50459_ (_43367_, _43366_, _42563_);
  and _50460_ (_43368_, _42658_, _42565_);
  and _50461_ (_43369_, _42558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or _50462_ (_43370_, _43369_, _43368_);
  or _50463_ (_43371_, _43370_, _43367_);
  and _50464_ (_05061_, _43371_, _42618_);
  and _50465_ (_43372_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and _50466_ (_43373_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _50467_ (_43374_, _43373_, _42309_);
  or _50468_ (_43375_, _43374_, _43372_);
  and _50469_ (_43376_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and _50470_ (_43377_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or _50471_ (_43378_, _43377_, _42455_);
  or _50472_ (_43379_, _43378_, _43376_);
  and _50473_ (_43380_, _43379_, _43375_);
  or _50474_ (_43381_, _43380_, _42215_);
  and _50475_ (_43382_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and _50476_ (_43383_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _50477_ (_43384_, _43383_, _42309_);
  or _50478_ (_43385_, _43384_, _43382_);
  and _50479_ (_43386_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and _50480_ (_43387_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or _50481_ (_43388_, _43387_, _42455_);
  or _50482_ (_43389_, _43388_, _43386_);
  and _50483_ (_43390_, _43389_, _43385_);
  or _50484_ (_43391_, _43390_, _42214_);
  and _50485_ (_43392_, _43391_, _42466_);
  and _50486_ (_43393_, _43392_, _43381_);
  or _50487_ (_43394_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _50488_ (_43395_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _50489_ (_43396_, _43395_, _43394_);
  or _50490_ (_43397_, _43396_, _42455_);
  or _50491_ (_43398_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or _50492_ (_43399_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and _50493_ (_43400_, _43399_, _43398_);
  or _50494_ (_43401_, _43400_, _42309_);
  and _50495_ (_43402_, _43401_, _43397_);
  or _50496_ (_43403_, _43402_, _42215_);
  or _50497_ (_43404_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or _50498_ (_43405_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _50499_ (_43406_, _43405_, _43404_);
  or _50500_ (_43407_, _43406_, _42455_);
  or _50501_ (_43408_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or _50502_ (_43409_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and _50503_ (_43410_, _43409_, _43408_);
  or _50504_ (_43411_, _43410_, _42309_);
  and _50505_ (_43412_, _43411_, _43407_);
  or _50506_ (_43413_, _43412_, _42214_);
  and _50507_ (_43414_, _43413_, _42454_);
  and _50508_ (_43415_, _43414_, _43403_);
  or _50509_ (_43416_, _43415_, _43393_);
  or _50510_ (_43417_, _43416_, _42558_);
  or _50511_ (_43418_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _50512_ (_43419_, _43418_, _42567_);
  and _50513_ (_43420_, _43419_, _43417_);
  and _50514_ (_39869_, _42668_, _42618_);
  and _50515_ (_43421_, _39869_, _42565_);
  or _50516_ (_05063_, _43421_, _43420_);
  and _50517_ (_43422_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and _50518_ (_43423_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _50519_ (_43424_, _43423_, _42309_);
  or _50520_ (_43425_, _43424_, _43422_);
  and _50521_ (_43426_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and _50522_ (_43427_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _50523_ (_43428_, _43427_, _42455_);
  or _50524_ (_43429_, _43428_, _43426_);
  and _50525_ (_43430_, _43429_, _43425_);
  or _50526_ (_43431_, _43430_, _42215_);
  and _50527_ (_43432_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and _50528_ (_43433_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _50529_ (_43434_, _43433_, _42309_);
  or _50530_ (_43435_, _43434_, _43432_);
  and _50531_ (_43436_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and _50532_ (_43437_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or _50533_ (_43438_, _43437_, _42455_);
  or _50534_ (_43439_, _43438_, _43436_);
  and _50535_ (_43440_, _43439_, _43435_);
  or _50536_ (_43441_, _43440_, _42214_);
  and _50537_ (_43442_, _43441_, _42466_);
  and _50538_ (_43443_, _43442_, _43431_);
  or _50539_ (_43444_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or _50540_ (_43445_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _50541_ (_43446_, _43445_, _43444_);
  or _50542_ (_43447_, _43446_, _42455_);
  or _50543_ (_43448_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or _50544_ (_43449_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and _50545_ (_43450_, _43449_, _43448_);
  or _50546_ (_43451_, _43450_, _42309_);
  and _50547_ (_43452_, _43451_, _43447_);
  or _50548_ (_43453_, _43452_, _42215_);
  or _50549_ (_43454_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or _50550_ (_43455_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _50551_ (_43456_, _43455_, _43454_);
  or _50552_ (_43457_, _43456_, _42455_);
  or _50553_ (_43458_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or _50554_ (_43459_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and _50555_ (_43460_, _43459_, _43458_);
  or _50556_ (_43461_, _43460_, _42309_);
  and _50557_ (_43462_, _43461_, _43457_);
  or _50558_ (_43463_, _43462_, _42214_);
  and _50559_ (_43464_, _43463_, _42454_);
  and _50560_ (_43465_, _43464_, _43453_);
  or _50561_ (_43466_, _43465_, _43443_);
  or _50562_ (_43467_, _43466_, _42558_);
  or _50563_ (_43468_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _50564_ (_43469_, _43468_, _42567_);
  and _50565_ (_43470_, _43469_, _43467_);
  and _50566_ (_39870_, _42679_, _42618_);
  and _50567_ (_43471_, _39870_, _42565_);
  or _50568_ (_05065_, _43471_, _43470_);
  or _50569_ (_43472_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not _50570_ (_43473_, \oc8051_gm_cxrom_1.cell0.valid );
  or _50571_ (_43474_, _43473_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand _50572_ (_43475_, _43474_, _43472_);
  nand _50573_ (_43476_, _43475_, _42618_);
  or _50574_ (_43477_, \oc8051_gm_cxrom_1.cell0.data [7], _42618_);
  and _50575_ (_05073_, _43477_, _43476_);
  or _50576_ (_43478_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or _50577_ (_43479_, \oc8051_gm_cxrom_1.cell0.data [0], _43473_);
  nand _50578_ (_43480_, _43479_, _43478_);
  nand _50579_ (_43481_, _43480_, _42618_);
  or _50580_ (_43482_, \oc8051_gm_cxrom_1.cell0.data [0], _42618_);
  and _50581_ (_05080_, _43482_, _43481_);
  or _50582_ (_43483_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or _50583_ (_43484_, \oc8051_gm_cxrom_1.cell0.data [1], _43473_);
  nand _50584_ (_43485_, _43484_, _43483_);
  nand _50585_ (_43486_, _43485_, _42618_);
  or _50586_ (_43487_, \oc8051_gm_cxrom_1.cell0.data [1], _42618_);
  and _50587_ (_05083_, _43487_, _43486_);
  or _50588_ (_43488_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or _50589_ (_43489_, \oc8051_gm_cxrom_1.cell0.data [2], _43473_);
  nand _50590_ (_43490_, _43489_, _43488_);
  nand _50591_ (_43491_, _43490_, _42618_);
  or _50592_ (_43492_, \oc8051_gm_cxrom_1.cell0.data [2], _42618_);
  and _50593_ (_05087_, _43492_, _43491_);
  or _50594_ (_43493_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or _50595_ (_43494_, \oc8051_gm_cxrom_1.cell0.data [3], _43473_);
  nand _50596_ (_43495_, _43494_, _43493_);
  nand _50597_ (_43496_, _43495_, _42618_);
  or _50598_ (_43497_, \oc8051_gm_cxrom_1.cell0.data [3], _42618_);
  and _50599_ (_05091_, _43497_, _43496_);
  or _50600_ (_43498_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or _50601_ (_43499_, \oc8051_gm_cxrom_1.cell0.data [4], _43473_);
  nand _50602_ (_43500_, _43499_, _43498_);
  nand _50603_ (_43501_, _43500_, _42618_);
  or _50604_ (_43502_, \oc8051_gm_cxrom_1.cell0.data [4], _42618_);
  and _50605_ (_05095_, _43502_, _43501_);
  or _50606_ (_43503_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or _50607_ (_43504_, \oc8051_gm_cxrom_1.cell0.data [5], _43473_);
  nand _50608_ (_43505_, _43504_, _43503_);
  nand _50609_ (_43506_, _43505_, _42618_);
  or _50610_ (_43507_, \oc8051_gm_cxrom_1.cell0.data [5], _42618_);
  and _50611_ (_05099_, _43507_, _43506_);
  or _50612_ (_43508_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or _50613_ (_43509_, \oc8051_gm_cxrom_1.cell0.data [6], _43473_);
  nand _50614_ (_43510_, _43509_, _43508_);
  nand _50615_ (_43511_, _43510_, _42618_);
  or _50616_ (_43512_, \oc8051_gm_cxrom_1.cell0.data [6], _42618_);
  and _50617_ (_05103_, _43512_, _43511_);
  or _50618_ (_43513_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not _50619_ (_43514_, \oc8051_gm_cxrom_1.cell1.valid );
  or _50620_ (_43515_, _43514_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand _50621_ (_43516_, _43515_, _43513_);
  nand _50622_ (_43517_, _43516_, _42618_);
  or _50623_ (_43518_, \oc8051_gm_cxrom_1.cell1.data [7], _42618_);
  and _50624_ (_05124_, _43518_, _43517_);
  or _50625_ (_43519_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or _50626_ (_43520_, \oc8051_gm_cxrom_1.cell1.data [0], _43514_);
  nand _50627_ (_43521_, _43520_, _43519_);
  nand _50628_ (_43522_, _43521_, _42618_);
  or _50629_ (_43523_, \oc8051_gm_cxrom_1.cell1.data [0], _42618_);
  and _50630_ (_05131_, _43523_, _43522_);
  or _50631_ (_43524_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or _50632_ (_43525_, \oc8051_gm_cxrom_1.cell1.data [1], _43514_);
  nand _50633_ (_43526_, _43525_, _43524_);
  nand _50634_ (_43527_, _43526_, _42618_);
  or _50635_ (_43528_, \oc8051_gm_cxrom_1.cell1.data [1], _42618_);
  and _50636_ (_05135_, _43528_, _43527_);
  or _50637_ (_43529_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or _50638_ (_43530_, \oc8051_gm_cxrom_1.cell1.data [2], _43514_);
  nand _50639_ (_43531_, _43530_, _43529_);
  nand _50640_ (_43532_, _43531_, _42618_);
  or _50641_ (_43533_, \oc8051_gm_cxrom_1.cell1.data [2], _42618_);
  and _50642_ (_05139_, _43533_, _43532_);
  or _50643_ (_00001_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or _50644_ (_00002_, \oc8051_gm_cxrom_1.cell1.data [3], _43514_);
  nand _50645_ (_00003_, _00002_, _00001_);
  nand _50646_ (_00004_, _00003_, _42618_);
  or _50647_ (_00005_, \oc8051_gm_cxrom_1.cell1.data [3], _42618_);
  and _50648_ (_05143_, _00005_, _00004_);
  or _50649_ (_00006_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or _50650_ (_00007_, \oc8051_gm_cxrom_1.cell1.data [4], _43514_);
  nand _50651_ (_00008_, _00007_, _00006_);
  nand _50652_ (_00009_, _00008_, _42618_);
  or _50653_ (_00010_, \oc8051_gm_cxrom_1.cell1.data [4], _42618_);
  and _50654_ (_05147_, _00010_, _00009_);
  or _50655_ (_00011_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or _50656_ (_00012_, \oc8051_gm_cxrom_1.cell1.data [5], _43514_);
  nand _50657_ (_00013_, _00012_, _00011_);
  nand _50658_ (_00014_, _00013_, _42618_);
  or _50659_ (_00015_, \oc8051_gm_cxrom_1.cell1.data [5], _42618_);
  and _50660_ (_05151_, _00015_, _00014_);
  or _50661_ (_00016_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or _50662_ (_00017_, \oc8051_gm_cxrom_1.cell1.data [6], _43514_);
  nand _50663_ (_00018_, _00017_, _00016_);
  nand _50664_ (_00019_, _00018_, _42618_);
  or _50665_ (_00020_, \oc8051_gm_cxrom_1.cell1.data [6], _42618_);
  and _50666_ (_05155_, _00020_, _00019_);
  or _50667_ (_00021_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not _50668_ (_00022_, \oc8051_gm_cxrom_1.cell2.valid );
  or _50669_ (_00023_, _00022_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand _50670_ (_00024_, _00023_, _00021_);
  nand _50671_ (_00025_, _00024_, _42618_);
  or _50672_ (_00026_, \oc8051_gm_cxrom_1.cell2.data [7], _42618_);
  and _50673_ (_05176_, _00026_, _00025_);
  or _50674_ (_00027_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or _50675_ (_00028_, \oc8051_gm_cxrom_1.cell2.data [0], _00022_);
  nand _50676_ (_00029_, _00028_, _00027_);
  nand _50677_ (_00030_, _00029_, _42618_);
  or _50678_ (_00031_, \oc8051_gm_cxrom_1.cell2.data [0], _42618_);
  and _50679_ (_05183_, _00031_, _00030_);
  or _50680_ (_00032_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or _50681_ (_00033_, \oc8051_gm_cxrom_1.cell2.data [1], _00022_);
  nand _50682_ (_00034_, _00033_, _00032_);
  nand _50683_ (_00035_, _00034_, _42618_);
  or _50684_ (_00036_, \oc8051_gm_cxrom_1.cell2.data [1], _42618_);
  and _50685_ (_05187_, _00036_, _00035_);
  or _50686_ (_00037_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or _50687_ (_00038_, \oc8051_gm_cxrom_1.cell2.data [2], _00022_);
  nand _50688_ (_00039_, _00038_, _00037_);
  nand _50689_ (_00040_, _00039_, _42618_);
  or _50690_ (_00041_, \oc8051_gm_cxrom_1.cell2.data [2], _42618_);
  and _50691_ (_05191_, _00041_, _00040_);
  or _50692_ (_00042_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or _50693_ (_00043_, \oc8051_gm_cxrom_1.cell2.data [3], _00022_);
  nand _50694_ (_00044_, _00043_, _00042_);
  nand _50695_ (_00045_, _00044_, _42618_);
  or _50696_ (_00046_, \oc8051_gm_cxrom_1.cell2.data [3], _42618_);
  and _50697_ (_05194_, _00046_, _00045_);
  or _50698_ (_00047_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or _50699_ (_00048_, \oc8051_gm_cxrom_1.cell2.data [4], _00022_);
  nand _50700_ (_00049_, _00048_, _00047_);
  nand _50701_ (_00050_, _00049_, _42618_);
  or _50702_ (_00051_, \oc8051_gm_cxrom_1.cell2.data [4], _42618_);
  and _50703_ (_05198_, _00051_, _00050_);
  or _50704_ (_00052_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or _50705_ (_00053_, \oc8051_gm_cxrom_1.cell2.data [5], _00022_);
  nand _50706_ (_00054_, _00053_, _00052_);
  nand _50707_ (_00055_, _00054_, _42618_);
  or _50708_ (_00056_, \oc8051_gm_cxrom_1.cell2.data [5], _42618_);
  and _50709_ (_05202_, _00056_, _00055_);
  or _50710_ (_00057_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or _50711_ (_00058_, \oc8051_gm_cxrom_1.cell2.data [6], _00022_);
  nand _50712_ (_00059_, _00058_, _00057_);
  nand _50713_ (_00060_, _00059_, _42618_);
  or _50714_ (_00061_, \oc8051_gm_cxrom_1.cell2.data [6], _42618_);
  and _50715_ (_05206_, _00061_, _00060_);
  or _50716_ (_00062_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not _50717_ (_00063_, \oc8051_gm_cxrom_1.cell3.valid );
  or _50718_ (_00064_, _00063_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand _50719_ (_00065_, _00064_, _00062_);
  nand _50720_ (_00066_, _00065_, _42618_);
  or _50721_ (_00067_, \oc8051_gm_cxrom_1.cell3.data [7], _42618_);
  and _50722_ (_05227_, _00067_, _00066_);
  or _50723_ (_00068_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or _50724_ (_00069_, \oc8051_gm_cxrom_1.cell3.data [0], _00063_);
  nand _50725_ (_00070_, _00069_, _00068_);
  nand _50726_ (_00071_, _00070_, _42618_);
  or _50727_ (_00072_, \oc8051_gm_cxrom_1.cell3.data [0], _42618_);
  and _50728_ (_05234_, _00072_, _00071_);
  or _50729_ (_00073_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or _50730_ (_00074_, \oc8051_gm_cxrom_1.cell3.data [1], _00063_);
  nand _50731_ (_00075_, _00074_, _00073_);
  nand _50732_ (_00076_, _00075_, _42618_);
  or _50733_ (_00077_, \oc8051_gm_cxrom_1.cell3.data [1], _42618_);
  and _50734_ (_05238_, _00077_, _00076_);
  or _50735_ (_00078_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or _50736_ (_00079_, \oc8051_gm_cxrom_1.cell3.data [2], _00063_);
  nand _50737_ (_00080_, _00079_, _00078_);
  nand _50738_ (_00081_, _00080_, _42618_);
  or _50739_ (_00082_, \oc8051_gm_cxrom_1.cell3.data [2], _42618_);
  and _50740_ (_05242_, _00082_, _00081_);
  or _50741_ (_00083_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or _50742_ (_00084_, \oc8051_gm_cxrom_1.cell3.data [3], _00063_);
  nand _50743_ (_00085_, _00084_, _00083_);
  nand _50744_ (_00086_, _00085_, _42618_);
  or _50745_ (_00087_, \oc8051_gm_cxrom_1.cell3.data [3], _42618_);
  and _50746_ (_05246_, _00087_, _00086_);
  or _50747_ (_00088_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or _50748_ (_00089_, \oc8051_gm_cxrom_1.cell3.data [4], _00063_);
  nand _50749_ (_00090_, _00089_, _00088_);
  nand _50750_ (_00091_, _00090_, _42618_);
  or _50751_ (_00092_, \oc8051_gm_cxrom_1.cell3.data [4], _42618_);
  and _50752_ (_05250_, _00092_, _00091_);
  or _50753_ (_00093_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or _50754_ (_00094_, \oc8051_gm_cxrom_1.cell3.data [5], _00063_);
  nand _50755_ (_00095_, _00094_, _00093_);
  nand _50756_ (_00096_, _00095_, _42618_);
  or _50757_ (_00097_, \oc8051_gm_cxrom_1.cell3.data [5], _42618_);
  and _50758_ (_05254_, _00097_, _00096_);
  or _50759_ (_00098_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or _50760_ (_00099_, \oc8051_gm_cxrom_1.cell3.data [6], _00063_);
  nand _50761_ (_00100_, _00099_, _00098_);
  nand _50762_ (_00101_, _00100_, _42618_);
  or _50763_ (_00102_, \oc8051_gm_cxrom_1.cell3.data [6], _42618_);
  and _50764_ (_05258_, _00102_, _00101_);
  or _50765_ (_00103_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not _50766_ (_00104_, \oc8051_gm_cxrom_1.cell4.valid );
  or _50767_ (_00105_, _00104_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand _50768_ (_00106_, _00105_, _00103_);
  nand _50769_ (_00107_, _00106_, _42618_);
  or _50770_ (_00108_, \oc8051_gm_cxrom_1.cell4.data [7], _42618_);
  and _50771_ (_05279_, _00108_, _00107_);
  or _50772_ (_00109_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or _50773_ (_00110_, \oc8051_gm_cxrom_1.cell4.data [0], _00104_);
  nand _50774_ (_00111_, _00110_, _00109_);
  nand _50775_ (_00112_, _00111_, _42618_);
  or _50776_ (_00113_, \oc8051_gm_cxrom_1.cell4.data [0], _42618_);
  and _50777_ (_05286_, _00113_, _00112_);
  or _50778_ (_00114_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or _50779_ (_00115_, \oc8051_gm_cxrom_1.cell4.data [1], _00104_);
  nand _50780_ (_00116_, _00115_, _00114_);
  nand _50781_ (_00117_, _00116_, _42618_);
  or _50782_ (_00118_, \oc8051_gm_cxrom_1.cell4.data [1], _42618_);
  and _50783_ (_05290_, _00118_, _00117_);
  or _50784_ (_00119_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or _50785_ (_00120_, \oc8051_gm_cxrom_1.cell4.data [2], _00104_);
  nand _50786_ (_00121_, _00120_, _00119_);
  nand _50787_ (_00122_, _00121_, _42618_);
  or _50788_ (_00123_, \oc8051_gm_cxrom_1.cell4.data [2], _42618_);
  and _50789_ (_05294_, _00123_, _00122_);
  or _50790_ (_00124_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or _50791_ (_00125_, \oc8051_gm_cxrom_1.cell4.data [3], _00104_);
  nand _50792_ (_00126_, _00125_, _00124_);
  nand _50793_ (_00127_, _00126_, _42618_);
  or _50794_ (_00128_, \oc8051_gm_cxrom_1.cell4.data [3], _42618_);
  and _50795_ (_05298_, _00128_, _00127_);
  or _50796_ (_00129_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or _50797_ (_00131_, \oc8051_gm_cxrom_1.cell4.data [4], _00104_);
  nand _50798_ (_00133_, _00131_, _00129_);
  nand _50799_ (_00135_, _00133_, _42618_);
  or _50800_ (_00137_, \oc8051_gm_cxrom_1.cell4.data [4], _42618_);
  and _50801_ (_05301_, _00137_, _00135_);
  or _50802_ (_00140_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or _50803_ (_00142_, \oc8051_gm_cxrom_1.cell4.data [5], _00104_);
  nand _50804_ (_00144_, _00142_, _00140_);
  nand _50805_ (_00146_, _00144_, _42618_);
  or _50806_ (_00148_, \oc8051_gm_cxrom_1.cell4.data [5], _42618_);
  and _50807_ (_05305_, _00148_, _00146_);
  or _50808_ (_00151_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or _50809_ (_00153_, \oc8051_gm_cxrom_1.cell4.data [6], _00104_);
  nand _50810_ (_00155_, _00153_, _00151_);
  nand _50811_ (_00157_, _00155_, _42618_);
  or _50812_ (_00159_, \oc8051_gm_cxrom_1.cell4.data [6], _42618_);
  and _50813_ (_05309_, _00159_, _00157_);
  or _50814_ (_00162_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not _50815_ (_00164_, \oc8051_gm_cxrom_1.cell5.valid );
  or _50816_ (_00166_, _00164_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand _50817_ (_00168_, _00166_, _00162_);
  nand _50818_ (_00170_, _00168_, _42618_);
  or _50819_ (_00172_, \oc8051_gm_cxrom_1.cell5.data [7], _42618_);
  and _50820_ (_05331_, _00172_, _00170_);
  or _50821_ (_00175_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or _50822_ (_00177_, \oc8051_gm_cxrom_1.cell5.data [0], _00164_);
  nand _50823_ (_00179_, _00177_, _00175_);
  nand _50824_ (_00181_, _00179_, _42618_);
  or _50825_ (_00183_, \oc8051_gm_cxrom_1.cell5.data [0], _42618_);
  and _50826_ (_05337_, _00183_, _00181_);
  or _50827_ (_00186_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or _50828_ (_00187_, \oc8051_gm_cxrom_1.cell5.data [1], _00164_);
  nand _50829_ (_00188_, _00187_, _00186_);
  nand _50830_ (_00189_, _00188_, _42618_);
  or _50831_ (_00190_, \oc8051_gm_cxrom_1.cell5.data [1], _42618_);
  and _50832_ (_05341_, _00190_, _00189_);
  or _50833_ (_00191_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or _50834_ (_00192_, \oc8051_gm_cxrom_1.cell5.data [2], _00164_);
  nand _50835_ (_00193_, _00192_, _00191_);
  nand _50836_ (_00194_, _00193_, _42618_);
  or _50837_ (_00195_, \oc8051_gm_cxrom_1.cell5.data [2], _42618_);
  and _50838_ (_05345_, _00195_, _00194_);
  or _50839_ (_00196_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or _50840_ (_00197_, \oc8051_gm_cxrom_1.cell5.data [3], _00164_);
  nand _50841_ (_00198_, _00197_, _00196_);
  nand _50842_ (_00199_, _00198_, _42618_);
  or _50843_ (_00200_, \oc8051_gm_cxrom_1.cell5.data [3], _42618_);
  and _50844_ (_05349_, _00200_, _00199_);
  or _50845_ (_00201_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or _50846_ (_00202_, \oc8051_gm_cxrom_1.cell5.data [4], _00164_);
  nand _50847_ (_00203_, _00202_, _00201_);
  nand _50848_ (_00204_, _00203_, _42618_);
  or _50849_ (_00205_, \oc8051_gm_cxrom_1.cell5.data [4], _42618_);
  and _50850_ (_05353_, _00205_, _00204_);
  or _50851_ (_00206_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or _50852_ (_00207_, \oc8051_gm_cxrom_1.cell5.data [5], _00164_);
  nand _50853_ (_00208_, _00207_, _00206_);
  nand _50854_ (_00209_, _00208_, _42618_);
  or _50855_ (_00210_, \oc8051_gm_cxrom_1.cell5.data [5], _42618_);
  and _50856_ (_05357_, _00210_, _00209_);
  or _50857_ (_00211_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or _50858_ (_00212_, \oc8051_gm_cxrom_1.cell5.data [6], _00164_);
  nand _50859_ (_00213_, _00212_, _00211_);
  nand _50860_ (_00214_, _00213_, _42618_);
  or _50861_ (_00215_, \oc8051_gm_cxrom_1.cell5.data [6], _42618_);
  and _50862_ (_05361_, _00215_, _00214_);
  or _50863_ (_00216_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not _50864_ (_00217_, \oc8051_gm_cxrom_1.cell6.valid );
  or _50865_ (_00218_, _00217_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand _50866_ (_00219_, _00218_, _00216_);
  nand _50867_ (_00220_, _00219_, _42618_);
  or _50868_ (_00221_, \oc8051_gm_cxrom_1.cell6.data [7], _42618_);
  and _50869_ (_05382_, _00221_, _00220_);
  or _50870_ (_00222_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or _50871_ (_00223_, \oc8051_gm_cxrom_1.cell6.data [0], _00217_);
  nand _50872_ (_00224_, _00223_, _00222_);
  nand _50873_ (_00225_, _00224_, _42618_);
  or _50874_ (_00226_, \oc8051_gm_cxrom_1.cell6.data [0], _42618_);
  and _50875_ (_05389_, _00226_, _00225_);
  or _50876_ (_00227_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or _50877_ (_00228_, \oc8051_gm_cxrom_1.cell6.data [1], _00217_);
  nand _50878_ (_00229_, _00228_, _00227_);
  nand _50879_ (_00230_, _00229_, _42618_);
  or _50880_ (_00231_, \oc8051_gm_cxrom_1.cell6.data [1], _42618_);
  and _50881_ (_05393_, _00231_, _00230_);
  or _50882_ (_00232_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or _50883_ (_00233_, \oc8051_gm_cxrom_1.cell6.data [2], _00217_);
  nand _50884_ (_00234_, _00233_, _00232_);
  nand _50885_ (_00235_, _00234_, _42618_);
  or _50886_ (_00236_, \oc8051_gm_cxrom_1.cell6.data [2], _42618_);
  and _50887_ (_05397_, _00236_, _00235_);
  or _50888_ (_00237_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or _50889_ (_00238_, \oc8051_gm_cxrom_1.cell6.data [3], _00217_);
  nand _50890_ (_00239_, _00238_, _00237_);
  nand _50891_ (_00240_, _00239_, _42618_);
  or _50892_ (_00241_, \oc8051_gm_cxrom_1.cell6.data [3], _42618_);
  and _50893_ (_05401_, _00241_, _00240_);
  or _50894_ (_00242_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or _50895_ (_00243_, \oc8051_gm_cxrom_1.cell6.data [4], _00217_);
  nand _50896_ (_00244_, _00243_, _00242_);
  nand _50897_ (_00245_, _00244_, _42618_);
  or _50898_ (_00246_, \oc8051_gm_cxrom_1.cell6.data [4], _42618_);
  and _50899_ (_05405_, _00246_, _00245_);
  or _50900_ (_00247_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or _50901_ (_00248_, \oc8051_gm_cxrom_1.cell6.data [5], _00217_);
  nand _50902_ (_00249_, _00248_, _00247_);
  nand _50903_ (_00250_, _00249_, _42618_);
  or _50904_ (_00251_, \oc8051_gm_cxrom_1.cell6.data [5], _42618_);
  and _50905_ (_05409_, _00251_, _00250_);
  or _50906_ (_00252_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or _50907_ (_00253_, \oc8051_gm_cxrom_1.cell6.data [6], _00217_);
  nand _50908_ (_00254_, _00253_, _00252_);
  nand _50909_ (_00255_, _00254_, _42618_);
  or _50910_ (_00256_, \oc8051_gm_cxrom_1.cell6.data [6], _42618_);
  and _50911_ (_05412_, _00256_, _00255_);
  or _50912_ (_00257_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not _50913_ (_00258_, \oc8051_gm_cxrom_1.cell7.valid );
  or _50914_ (_00259_, _00258_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand _50915_ (_00260_, _00259_, _00257_);
  nand _50916_ (_00261_, _00260_, _42618_);
  or _50917_ (_00262_, \oc8051_gm_cxrom_1.cell7.data [7], _42618_);
  and _50918_ (_05434_, _00262_, _00261_);
  or _50919_ (_00263_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or _50920_ (_00264_, \oc8051_gm_cxrom_1.cell7.data [0], _00258_);
  nand _50921_ (_00265_, _00264_, _00263_);
  nand _50922_ (_00266_, _00265_, _42618_);
  or _50923_ (_00267_, \oc8051_gm_cxrom_1.cell7.data [0], _42618_);
  and _50924_ (_05441_, _00267_, _00266_);
  or _50925_ (_00268_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or _50926_ (_00269_, \oc8051_gm_cxrom_1.cell7.data [1], _00258_);
  nand _50927_ (_00270_, _00269_, _00268_);
  nand _50928_ (_00271_, _00270_, _42618_);
  or _50929_ (_00272_, \oc8051_gm_cxrom_1.cell7.data [1], _42618_);
  and _50930_ (_05445_, _00272_, _00271_);
  or _50931_ (_00273_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or _50932_ (_00274_, \oc8051_gm_cxrom_1.cell7.data [2], _00258_);
  nand _50933_ (_00275_, _00274_, _00273_);
  nand _50934_ (_00276_, _00275_, _42618_);
  or _50935_ (_00277_, \oc8051_gm_cxrom_1.cell7.data [2], _42618_);
  and _50936_ (_05448_, _00277_, _00276_);
  or _50937_ (_00278_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or _50938_ (_00279_, \oc8051_gm_cxrom_1.cell7.data [3], _00258_);
  nand _50939_ (_00280_, _00279_, _00278_);
  nand _50940_ (_00281_, _00280_, _42618_);
  or _50941_ (_00282_, \oc8051_gm_cxrom_1.cell7.data [3], _42618_);
  and _50942_ (_05452_, _00282_, _00281_);
  or _50943_ (_00283_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or _50944_ (_00284_, \oc8051_gm_cxrom_1.cell7.data [4], _00258_);
  nand _50945_ (_00285_, _00284_, _00283_);
  nand _50946_ (_00286_, _00285_, _42618_);
  or _50947_ (_00287_, \oc8051_gm_cxrom_1.cell7.data [4], _42618_);
  and _50948_ (_05456_, _00287_, _00286_);
  or _50949_ (_00288_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or _50950_ (_00289_, \oc8051_gm_cxrom_1.cell7.data [5], _00258_);
  nand _50951_ (_00290_, _00289_, _00288_);
  nand _50952_ (_00291_, _00290_, _42618_);
  or _50953_ (_00292_, \oc8051_gm_cxrom_1.cell7.data [5], _42618_);
  and _50954_ (_05460_, _00292_, _00291_);
  or _50955_ (_00293_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or _50956_ (_00294_, \oc8051_gm_cxrom_1.cell7.data [6], _00258_);
  nand _50957_ (_00295_, _00294_, _00293_);
  nand _50958_ (_00296_, _00295_, _42618_);
  or _50959_ (_00297_, \oc8051_gm_cxrom_1.cell7.data [6], _42618_);
  and _50960_ (_05464_, _00297_, _00296_);
  or _50961_ (_00298_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not _50962_ (_00299_, \oc8051_gm_cxrom_1.cell8.valid );
  or _50963_ (_00300_, _00299_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand _50964_ (_00301_, _00300_, _00298_);
  nand _50965_ (_00302_, _00301_, _42618_);
  or _50966_ (_00303_, \oc8051_gm_cxrom_1.cell8.data [7], _42618_);
  and _50967_ (_05485_, _00303_, _00302_);
  or _50968_ (_00304_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or _50969_ (_00305_, \oc8051_gm_cxrom_1.cell8.data [0], _00299_);
  nand _50970_ (_00306_, _00305_, _00304_);
  nand _50971_ (_00307_, _00306_, _42618_);
  or _50972_ (_00308_, \oc8051_gm_cxrom_1.cell8.data [0], _42618_);
  and _50973_ (_05492_, _00308_, _00307_);
  or _50974_ (_00309_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or _50975_ (_00310_, \oc8051_gm_cxrom_1.cell8.data [1], _00299_);
  nand _50976_ (_00311_, _00310_, _00309_);
  nand _50977_ (_00312_, _00311_, _42618_);
  or _50978_ (_00313_, \oc8051_gm_cxrom_1.cell8.data [1], _42618_);
  and _50979_ (_05496_, _00313_, _00312_);
  or _50980_ (_00314_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or _50981_ (_00315_, \oc8051_gm_cxrom_1.cell8.data [2], _00299_);
  nand _50982_ (_00316_, _00315_, _00314_);
  nand _50983_ (_00317_, _00316_, _42618_);
  or _50984_ (_00318_, \oc8051_gm_cxrom_1.cell8.data [2], _42618_);
  and _50985_ (_05500_, _00318_, _00317_);
  or _50986_ (_00319_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or _50987_ (_00320_, \oc8051_gm_cxrom_1.cell8.data [3], _00299_);
  nand _50988_ (_00321_, _00320_, _00319_);
  nand _50989_ (_00322_, _00321_, _42618_);
  or _50990_ (_00323_, \oc8051_gm_cxrom_1.cell8.data [3], _42618_);
  and _50991_ (_05504_, _00323_, _00322_);
  or _50992_ (_00324_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or _50993_ (_00325_, \oc8051_gm_cxrom_1.cell8.data [4], _00299_);
  nand _50994_ (_00326_, _00325_, _00324_);
  nand _50995_ (_00327_, _00326_, _42618_);
  or _50996_ (_00328_, \oc8051_gm_cxrom_1.cell8.data [4], _42618_);
  and _50997_ (_05508_, _00328_, _00327_);
  or _50998_ (_00329_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or _50999_ (_00330_, \oc8051_gm_cxrom_1.cell8.data [5], _00299_);
  nand _51000_ (_00331_, _00330_, _00329_);
  nand _51001_ (_00332_, _00331_, _42618_);
  or _51002_ (_00333_, \oc8051_gm_cxrom_1.cell8.data [5], _42618_);
  and _51003_ (_05512_, _00333_, _00332_);
  or _51004_ (_00334_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or _51005_ (_00335_, \oc8051_gm_cxrom_1.cell8.data [6], _00299_);
  nand _51006_ (_00336_, _00335_, _00334_);
  nand _51007_ (_00337_, _00336_, _42618_);
  or _51008_ (_00338_, \oc8051_gm_cxrom_1.cell8.data [6], _42618_);
  and _51009_ (_05516_, _00338_, _00337_);
  or _51010_ (_00339_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not _51011_ (_00340_, \oc8051_gm_cxrom_1.cell9.valid );
  or _51012_ (_00341_, _00340_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand _51013_ (_00342_, _00341_, _00339_);
  nand _51014_ (_00343_, _00342_, _42618_);
  or _51015_ (_00344_, \oc8051_gm_cxrom_1.cell9.data [7], _42618_);
  and _51016_ (_05537_, _00344_, _00343_);
  or _51017_ (_00345_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or _51018_ (_00346_, \oc8051_gm_cxrom_1.cell9.data [0], _00340_);
  nand _51019_ (_00347_, _00346_, _00345_);
  nand _51020_ (_00348_, _00347_, _42618_);
  or _51021_ (_00349_, \oc8051_gm_cxrom_1.cell9.data [0], _42618_);
  and _51022_ (_05544_, _00349_, _00348_);
  or _51023_ (_00350_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or _51024_ (_00351_, \oc8051_gm_cxrom_1.cell9.data [1], _00340_);
  nand _51025_ (_00352_, _00351_, _00350_);
  nand _51026_ (_00353_, _00352_, _42618_);
  or _51027_ (_00354_, \oc8051_gm_cxrom_1.cell9.data [1], _42618_);
  and _51028_ (_05548_, _00354_, _00353_);
  or _51029_ (_00355_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or _51030_ (_00356_, \oc8051_gm_cxrom_1.cell9.data [2], _00340_);
  nand _51031_ (_00357_, _00356_, _00355_);
  nand _51032_ (_00358_, _00357_, _42618_);
  or _51033_ (_00359_, \oc8051_gm_cxrom_1.cell9.data [2], _42618_);
  and _51034_ (_05552_, _00359_, _00358_);
  or _51035_ (_00360_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or _51036_ (_00361_, \oc8051_gm_cxrom_1.cell9.data [3], _00340_);
  nand _51037_ (_00362_, _00361_, _00360_);
  nand _51038_ (_00363_, _00362_, _42618_);
  or _51039_ (_00364_, \oc8051_gm_cxrom_1.cell9.data [3], _42618_);
  and _51040_ (_05555_, _00364_, _00363_);
  or _51041_ (_00365_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or _51042_ (_00366_, \oc8051_gm_cxrom_1.cell9.data [4], _00340_);
  nand _51043_ (_00367_, _00366_, _00365_);
  nand _51044_ (_00368_, _00367_, _42618_);
  or _51045_ (_00369_, \oc8051_gm_cxrom_1.cell9.data [4], _42618_);
  and _51046_ (_05559_, _00369_, _00368_);
  or _51047_ (_00370_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or _51048_ (_00371_, \oc8051_gm_cxrom_1.cell9.data [5], _00340_);
  nand _51049_ (_00372_, _00371_, _00370_);
  nand _51050_ (_00373_, _00372_, _42618_);
  or _51051_ (_00374_, \oc8051_gm_cxrom_1.cell9.data [5], _42618_);
  and _51052_ (_05563_, _00374_, _00373_);
  or _51053_ (_00375_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or _51054_ (_00376_, \oc8051_gm_cxrom_1.cell9.data [6], _00340_);
  nand _51055_ (_00377_, _00376_, _00375_);
  nand _51056_ (_00378_, _00377_, _42618_);
  or _51057_ (_00379_, \oc8051_gm_cxrom_1.cell9.data [6], _42618_);
  and _51058_ (_05567_, _00379_, _00378_);
  or _51059_ (_00380_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not _51060_ (_00381_, \oc8051_gm_cxrom_1.cell10.valid );
  or _51061_ (_00382_, _00381_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand _51062_ (_00383_, _00382_, _00380_);
  nand _51063_ (_00384_, _00383_, _42618_);
  or _51064_ (_00385_, \oc8051_gm_cxrom_1.cell10.data [7], _42618_);
  and _51065_ (_05589_, _00385_, _00384_);
  or _51066_ (_00386_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or _51067_ (_00387_, \oc8051_gm_cxrom_1.cell10.data [0], _00381_);
  nand _51068_ (_00388_, _00387_, _00386_);
  nand _51069_ (_00389_, _00388_, _42618_);
  or _51070_ (_00390_, \oc8051_gm_cxrom_1.cell10.data [0], _42618_);
  and _51071_ (_05595_, _00390_, _00389_);
  or _51072_ (_00391_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or _51073_ (_00392_, \oc8051_gm_cxrom_1.cell10.data [1], _00381_);
  nand _51074_ (_00393_, _00392_, _00391_);
  nand _51075_ (_00394_, _00393_, _42618_);
  or _51076_ (_00395_, \oc8051_gm_cxrom_1.cell10.data [1], _42618_);
  and _51077_ (_05599_, _00395_, _00394_);
  or _51078_ (_00396_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or _51079_ (_00397_, \oc8051_gm_cxrom_1.cell10.data [2], _00381_);
  nand _51080_ (_00398_, _00397_, _00396_);
  nand _51081_ (_00399_, _00398_, _42618_);
  or _51082_ (_00400_, \oc8051_gm_cxrom_1.cell10.data [2], _42618_);
  and _51083_ (_05603_, _00400_, _00399_);
  or _51084_ (_00401_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or _51085_ (_00402_, \oc8051_gm_cxrom_1.cell10.data [3], _00381_);
  nand _51086_ (_00403_, _00402_, _00401_);
  nand _51087_ (_00404_, _00403_, _42618_);
  or _51088_ (_00405_, \oc8051_gm_cxrom_1.cell10.data [3], _42618_);
  and _51089_ (_05607_, _00405_, _00404_);
  or _51090_ (_00406_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or _51091_ (_00407_, \oc8051_gm_cxrom_1.cell10.data [4], _00381_);
  nand _51092_ (_00408_, _00407_, _00406_);
  nand _51093_ (_00409_, _00408_, _42618_);
  or _51094_ (_00410_, \oc8051_gm_cxrom_1.cell10.data [4], _42618_);
  and _51095_ (_05611_, _00410_, _00409_);
  or _51096_ (_00411_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or _51097_ (_00412_, \oc8051_gm_cxrom_1.cell10.data [5], _00381_);
  nand _51098_ (_00413_, _00412_, _00411_);
  nand _51099_ (_00414_, _00413_, _42618_);
  or _51100_ (_00415_, \oc8051_gm_cxrom_1.cell10.data [5], _42618_);
  and _51101_ (_05615_, _00415_, _00414_);
  or _51102_ (_00416_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or _51103_ (_00417_, \oc8051_gm_cxrom_1.cell10.data [6], _00381_);
  nand _51104_ (_00418_, _00417_, _00416_);
  nand _51105_ (_00419_, _00418_, _42618_);
  or _51106_ (_00420_, \oc8051_gm_cxrom_1.cell10.data [6], _42618_);
  and _51107_ (_05619_, _00420_, _00419_);
  or _51108_ (_00421_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not _51109_ (_00422_, \oc8051_gm_cxrom_1.cell11.valid );
  or _51110_ (_00423_, _00422_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand _51111_ (_00424_, _00423_, _00421_);
  nand _51112_ (_00425_, _00424_, _42618_);
  or _51113_ (_00426_, \oc8051_gm_cxrom_1.cell11.data [7], _42618_);
  and _51114_ (_05641_, _00426_, _00425_);
  or _51115_ (_00427_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or _51116_ (_00428_, \oc8051_gm_cxrom_1.cell11.data [0], _00422_);
  nand _51117_ (_00429_, _00428_, _00427_);
  nand _51118_ (_00430_, _00429_, _42618_);
  or _51119_ (_00431_, \oc8051_gm_cxrom_1.cell11.data [0], _42618_);
  and _51120_ (_05648_, _00431_, _00430_);
  or _51121_ (_00432_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or _51122_ (_00433_, \oc8051_gm_cxrom_1.cell11.data [1], _00422_);
  nand _51123_ (_00434_, _00433_, _00432_);
  nand _51124_ (_00435_, _00434_, _42618_);
  or _51125_ (_00436_, \oc8051_gm_cxrom_1.cell11.data [1], _42618_);
  and _51126_ (_05652_, _00436_, _00435_);
  or _51127_ (_00437_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or _51128_ (_00438_, \oc8051_gm_cxrom_1.cell11.data [2], _00422_);
  nand _51129_ (_00439_, _00438_, _00437_);
  nand _51130_ (_00440_, _00439_, _42618_);
  or _51131_ (_00441_, \oc8051_gm_cxrom_1.cell11.data [2], _42618_);
  and _51132_ (_05656_, _00441_, _00440_);
  or _51133_ (_00442_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or _51134_ (_00443_, \oc8051_gm_cxrom_1.cell11.data [3], _00422_);
  nand _51135_ (_00444_, _00443_, _00442_);
  nand _51136_ (_00445_, _00444_, _42618_);
  or _51137_ (_00446_, \oc8051_gm_cxrom_1.cell11.data [3], _42618_);
  and _51138_ (_05660_, _00446_, _00445_);
  or _51139_ (_00447_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or _51140_ (_00448_, \oc8051_gm_cxrom_1.cell11.data [4], _00422_);
  nand _51141_ (_00449_, _00448_, _00447_);
  nand _51142_ (_00450_, _00449_, _42618_);
  or _51143_ (_00451_, \oc8051_gm_cxrom_1.cell11.data [4], _42618_);
  and _51144_ (_05664_, _00451_, _00450_);
  or _51145_ (_00452_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or _51146_ (_00453_, \oc8051_gm_cxrom_1.cell11.data [5], _00422_);
  nand _51147_ (_00454_, _00453_, _00452_);
  nand _51148_ (_00455_, _00454_, _42618_);
  or _51149_ (_00456_, \oc8051_gm_cxrom_1.cell11.data [5], _42618_);
  and _51150_ (_05668_, _00456_, _00455_);
  or _51151_ (_00457_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or _51152_ (_00458_, \oc8051_gm_cxrom_1.cell11.data [6], _00422_);
  nand _51153_ (_00459_, _00458_, _00457_);
  nand _51154_ (_00460_, _00459_, _42618_);
  or _51155_ (_00461_, \oc8051_gm_cxrom_1.cell11.data [6], _42618_);
  and _51156_ (_05672_, _00461_, _00460_);
  or _51157_ (_00462_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not _51158_ (_00463_, \oc8051_gm_cxrom_1.cell12.valid );
  or _51159_ (_00464_, _00463_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand _51160_ (_00465_, _00464_, _00462_);
  nand _51161_ (_00466_, _00465_, _42618_);
  or _51162_ (_00467_, \oc8051_gm_cxrom_1.cell12.data [7], _42618_);
  and _51163_ (_05694_, _00467_, _00466_);
  or _51164_ (_00468_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or _51165_ (_00469_, \oc8051_gm_cxrom_1.cell12.data [0], _00463_);
  nand _51166_ (_00470_, _00469_, _00468_);
  nand _51167_ (_00471_, _00470_, _42618_);
  or _51168_ (_00472_, \oc8051_gm_cxrom_1.cell12.data [0], _42618_);
  and _51169_ (_05701_, _00472_, _00471_);
  or _51170_ (_00473_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or _51171_ (_00474_, \oc8051_gm_cxrom_1.cell12.data [1], _00463_);
  nand _51172_ (_00475_, _00474_, _00473_);
  nand _51173_ (_00476_, _00475_, _42618_);
  or _51174_ (_00477_, \oc8051_gm_cxrom_1.cell12.data [1], _42618_);
  and _51175_ (_05705_, _00477_, _00476_);
  or _51176_ (_00478_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or _51177_ (_00479_, \oc8051_gm_cxrom_1.cell12.data [2], _00463_);
  nand _51178_ (_00480_, _00479_, _00478_);
  nand _51179_ (_00481_, _00480_, _42618_);
  or _51180_ (_00482_, \oc8051_gm_cxrom_1.cell12.data [2], _42618_);
  and _51181_ (_05709_, _00482_, _00481_);
  or _51182_ (_00483_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or _51183_ (_00484_, \oc8051_gm_cxrom_1.cell12.data [3], _00463_);
  nand _51184_ (_00485_, _00484_, _00483_);
  nand _51185_ (_00486_, _00485_, _42618_);
  or _51186_ (_00487_, \oc8051_gm_cxrom_1.cell12.data [3], _42618_);
  and _51187_ (_05713_, _00487_, _00486_);
  or _51188_ (_00488_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or _51189_ (_00489_, \oc8051_gm_cxrom_1.cell12.data [4], _00463_);
  nand _51190_ (_00490_, _00489_, _00488_);
  nand _51191_ (_00491_, _00490_, _42618_);
  or _51192_ (_00492_, \oc8051_gm_cxrom_1.cell12.data [4], _42618_);
  and _51193_ (_05717_, _00492_, _00491_);
  or _51194_ (_00493_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or _51195_ (_00494_, \oc8051_gm_cxrom_1.cell12.data [5], _00463_);
  nand _51196_ (_00495_, _00494_, _00493_);
  nand _51197_ (_00496_, _00495_, _42618_);
  or _51198_ (_00497_, \oc8051_gm_cxrom_1.cell12.data [5], _42618_);
  and _51199_ (_05721_, _00497_, _00496_);
  or _51200_ (_00498_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or _51201_ (_00499_, \oc8051_gm_cxrom_1.cell12.data [6], _00463_);
  nand _51202_ (_00500_, _00499_, _00498_);
  nand _51203_ (_00501_, _00500_, _42618_);
  or _51204_ (_00502_, \oc8051_gm_cxrom_1.cell12.data [6], _42618_);
  and _51205_ (_05725_, _00502_, _00501_);
  or _51206_ (_00503_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not _51207_ (_00504_, \oc8051_gm_cxrom_1.cell13.valid );
  or _51208_ (_00505_, _00504_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand _51209_ (_00506_, _00505_, _00503_);
  nand _51210_ (_00507_, _00506_, _42618_);
  or _51211_ (_00508_, \oc8051_gm_cxrom_1.cell13.data [7], _42618_);
  and _51212_ (_05747_, _00508_, _00507_);
  or _51213_ (_00509_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or _51214_ (_00510_, \oc8051_gm_cxrom_1.cell13.data [0], _00504_);
  nand _51215_ (_00511_, _00510_, _00509_);
  nand _51216_ (_00512_, _00511_, _42618_);
  or _51217_ (_00513_, \oc8051_gm_cxrom_1.cell13.data [0], _42618_);
  and _51218_ (_05754_, _00513_, _00512_);
  or _51219_ (_00514_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or _51220_ (_00515_, \oc8051_gm_cxrom_1.cell13.data [1], _00504_);
  nand _51221_ (_00516_, _00515_, _00514_);
  nand _51222_ (_00517_, _00516_, _42618_);
  or _51223_ (_00518_, \oc8051_gm_cxrom_1.cell13.data [1], _42618_);
  and _51224_ (_05758_, _00518_, _00517_);
  or _51225_ (_00519_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or _51226_ (_00520_, \oc8051_gm_cxrom_1.cell13.data [2], _00504_);
  nand _51227_ (_00521_, _00520_, _00519_);
  nand _51228_ (_00522_, _00521_, _42618_);
  or _51229_ (_00523_, \oc8051_gm_cxrom_1.cell13.data [2], _42618_);
  and _51230_ (_05762_, _00523_, _00522_);
  or _51231_ (_00524_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or _51232_ (_00525_, \oc8051_gm_cxrom_1.cell13.data [3], _00504_);
  nand _51233_ (_00526_, _00525_, _00524_);
  nand _51234_ (_00527_, _00526_, _42618_);
  or _51235_ (_00528_, \oc8051_gm_cxrom_1.cell13.data [3], _42618_);
  and _51236_ (_05766_, _00528_, _00527_);
  or _51237_ (_00529_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or _51238_ (_00530_, \oc8051_gm_cxrom_1.cell13.data [4], _00504_);
  nand _51239_ (_00531_, _00530_, _00529_);
  nand _51240_ (_00532_, _00531_, _42618_);
  or _51241_ (_00533_, \oc8051_gm_cxrom_1.cell13.data [4], _42618_);
  and _51242_ (_05770_, _00533_, _00532_);
  or _51243_ (_00534_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or _51244_ (_00535_, \oc8051_gm_cxrom_1.cell13.data [5], _00504_);
  nand _51245_ (_00536_, _00535_, _00534_);
  nand _51246_ (_00537_, _00536_, _42618_);
  or _51247_ (_00538_, \oc8051_gm_cxrom_1.cell13.data [5], _42618_);
  and _51248_ (_05774_, _00538_, _00537_);
  or _51249_ (_00539_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or _51250_ (_00540_, \oc8051_gm_cxrom_1.cell13.data [6], _00504_);
  nand _51251_ (_00541_, _00540_, _00539_);
  nand _51252_ (_00542_, _00541_, _42618_);
  or _51253_ (_00544_, \oc8051_gm_cxrom_1.cell13.data [6], _42618_);
  and _51254_ (_05778_, _00544_, _00542_);
  or _51255_ (_00546_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not _51256_ (_00547_, \oc8051_gm_cxrom_1.cell14.valid );
  or _51257_ (_00549_, _00547_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand _51258_ (_00550_, _00549_, _00546_);
  nand _51259_ (_00552_, _00550_, _42618_);
  or _51260_ (_00553_, \oc8051_gm_cxrom_1.cell14.data [7], _42618_);
  and _51261_ (_05800_, _00553_, _00552_);
  or _51262_ (_00555_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or _51263_ (_00557_, \oc8051_gm_cxrom_1.cell14.data [0], _00547_);
  nand _51264_ (_00558_, _00557_, _00555_);
  nand _51265_ (_00560_, _00558_, _42618_);
  or _51266_ (_00561_, \oc8051_gm_cxrom_1.cell14.data [0], _42618_);
  and _51267_ (_05807_, _00561_, _00560_);
  or _51268_ (_00563_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or _51269_ (_00565_, \oc8051_gm_cxrom_1.cell14.data [1], _00547_);
  nand _51270_ (_00566_, _00565_, _00563_);
  nand _51271_ (_00568_, _00566_, _42618_);
  or _51272_ (_00569_, \oc8051_gm_cxrom_1.cell14.data [1], _42618_);
  and _51273_ (_05811_, _00569_, _00568_);
  or _51274_ (_00571_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or _51275_ (_00573_, \oc8051_gm_cxrom_1.cell14.data [2], _00547_);
  nand _51276_ (_00574_, _00573_, _00571_);
  nand _51277_ (_00576_, _00574_, _42618_);
  or _51278_ (_00577_, \oc8051_gm_cxrom_1.cell14.data [2], _42618_);
  and _51279_ (_05815_, _00577_, _00576_);
  or _51280_ (_00579_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or _51281_ (_00581_, \oc8051_gm_cxrom_1.cell14.data [3], _00547_);
  nand _51282_ (_00582_, _00581_, _00579_);
  nand _51283_ (_00584_, _00582_, _42618_);
  or _51284_ (_00585_, \oc8051_gm_cxrom_1.cell14.data [3], _42618_);
  and _51285_ (_05819_, _00585_, _00584_);
  or _51286_ (_00587_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or _51287_ (_00589_, \oc8051_gm_cxrom_1.cell14.data [4], _00547_);
  nand _51288_ (_00590_, _00589_, _00587_);
  nand _51289_ (_00592_, _00590_, _42618_);
  or _51290_ (_00593_, \oc8051_gm_cxrom_1.cell14.data [4], _42618_);
  and _51291_ (_05823_, _00593_, _00592_);
  or _51292_ (_00594_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or _51293_ (_00595_, \oc8051_gm_cxrom_1.cell14.data [5], _00547_);
  nand _51294_ (_00596_, _00595_, _00594_);
  nand _51295_ (_00597_, _00596_, _42618_);
  or _51296_ (_00598_, \oc8051_gm_cxrom_1.cell14.data [5], _42618_);
  and _51297_ (_05827_, _00598_, _00597_);
  or _51298_ (_00599_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or _51299_ (_00600_, \oc8051_gm_cxrom_1.cell14.data [6], _00547_);
  nand _51300_ (_00601_, _00600_, _00599_);
  nand _51301_ (_00602_, _00601_, _42618_);
  or _51302_ (_00603_, \oc8051_gm_cxrom_1.cell14.data [6], _42618_);
  and _51303_ (_05831_, _00603_, _00602_);
  or _51304_ (_00604_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not _51305_ (_00605_, \oc8051_gm_cxrom_1.cell15.valid );
  or _51306_ (_00606_, _00605_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand _51307_ (_00607_, _00606_, _00604_);
  nand _51308_ (_00608_, _00607_, _42618_);
  or _51309_ (_00609_, \oc8051_gm_cxrom_1.cell15.data [7], _42618_);
  and _51310_ (_05853_, _00609_, _00608_);
  or _51311_ (_00610_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or _51312_ (_00611_, \oc8051_gm_cxrom_1.cell15.data [0], _00605_);
  nand _51313_ (_00612_, _00611_, _00610_);
  nand _51314_ (_00613_, _00612_, _42618_);
  or _51315_ (_00614_, \oc8051_gm_cxrom_1.cell15.data [0], _42618_);
  and _51316_ (_05860_, _00614_, _00613_);
  or _51317_ (_00615_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or _51318_ (_00616_, \oc8051_gm_cxrom_1.cell15.data [1], _00605_);
  nand _51319_ (_00617_, _00616_, _00615_);
  nand _51320_ (_00618_, _00617_, _42618_);
  or _51321_ (_00619_, \oc8051_gm_cxrom_1.cell15.data [1], _42618_);
  and _51322_ (_05864_, _00619_, _00618_);
  or _51323_ (_00620_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or _51324_ (_00621_, \oc8051_gm_cxrom_1.cell15.data [2], _00605_);
  nand _51325_ (_00622_, _00621_, _00620_);
  nand _51326_ (_00623_, _00622_, _42618_);
  or _51327_ (_00624_, \oc8051_gm_cxrom_1.cell15.data [2], _42618_);
  and _51328_ (_05868_, _00624_, _00623_);
  or _51329_ (_00625_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or _51330_ (_00626_, \oc8051_gm_cxrom_1.cell15.data [3], _00605_);
  nand _51331_ (_00627_, _00626_, _00625_);
  nand _51332_ (_00628_, _00627_, _42618_);
  or _51333_ (_00629_, \oc8051_gm_cxrom_1.cell15.data [3], _42618_);
  and _51334_ (_05872_, _00629_, _00628_);
  or _51335_ (_00630_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or _51336_ (_00631_, \oc8051_gm_cxrom_1.cell15.data [4], _00605_);
  nand _51337_ (_00632_, _00631_, _00630_);
  nand _51338_ (_00633_, _00632_, _42618_);
  or _51339_ (_00634_, \oc8051_gm_cxrom_1.cell15.data [4], _42618_);
  and _51340_ (_05876_, _00634_, _00633_);
  or _51341_ (_00635_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or _51342_ (_00636_, \oc8051_gm_cxrom_1.cell15.data [5], _00605_);
  nand _51343_ (_00637_, _00636_, _00635_);
  nand _51344_ (_00638_, _00637_, _42618_);
  or _51345_ (_00639_, \oc8051_gm_cxrom_1.cell15.data [5], _42618_);
  and _51346_ (_05880_, _00639_, _00638_);
  or _51347_ (_00640_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or _51348_ (_00641_, \oc8051_gm_cxrom_1.cell15.data [6], _00605_);
  nand _51349_ (_00642_, _00641_, _00640_);
  nand _51350_ (_00643_, _00642_, _42618_);
  or _51351_ (_00644_, \oc8051_gm_cxrom_1.cell15.data [6], _42618_);
  and _51352_ (_05884_, _00644_, _00643_);
  nor _51353_ (_09659_, _37997_, rst);
  and _51354_ (_00645_, _38048_, _37987_);
  and _51355_ (_00646_, _00645_, _37890_);
  not _51356_ (_00647_, _00646_);
  and _51357_ (_00648_, _37970_, _37866_);
  and _51358_ (_00649_, _38049_, _38005_);
  nor _51359_ (_00650_, _00649_, _00648_);
  and _51360_ (_00651_, _00650_, _00647_);
  and _51361_ (_00652_, _38048_, _37889_);
  or _51362_ (_00653_, _37987_, _38005_);
  nand _51363_ (_00654_, _00653_, _00652_);
  and _51364_ (_00655_, _00654_, _00651_);
  and _51365_ (_00656_, _36958_, _42618_);
  not _51366_ (_00657_, _00656_);
  or _51367_ (_00658_, _00657_, _00648_);
  or _51368_ (_09662_, _00658_, _00655_);
  not _51369_ (_00659_, _37858_);
  and _51370_ (_00660_, _00659_, _37602_);
  and _51371_ (_00661_, _37832_, _37330_);
  and _51372_ (_00662_, _00661_, _00660_);
  not _51373_ (_00663_, _37954_);
  and _51374_ (_00664_, _00663_, _37931_);
  and _51375_ (_00665_, _00664_, _37884_);
  and _51376_ (_00666_, _00665_, _00662_);
  nor _51377_ (_00667_, _37858_, _37832_);
  and _51378_ (_00668_, _00667_, _37330_);
  and _51379_ (_00669_, _00668_, _37602_);
  not _51380_ (_00670_, _37884_);
  nor _51381_ (_00671_, _00663_, _37931_);
  and _51382_ (_00672_, _00671_, _00670_);
  and _51383_ (_00673_, _00672_, _00669_);
  and _51384_ (_00674_, _37908_, _37884_);
  nor _51385_ (_00675_, _37954_, _37931_);
  and _51386_ (_00676_, _00675_, _00674_);
  not _51387_ (_00677_, _37602_);
  and _51388_ (_00678_, _00668_, _00677_);
  and _51389_ (_00679_, _00678_, _00676_);
  or _51390_ (_00680_, _00679_, _00673_);
  or _51391_ (_00681_, _00680_, _00666_);
  nor _51392_ (_00682_, _37908_, _00670_);
  and _51393_ (_00683_, _00671_, _00682_);
  and _51394_ (_00684_, _00683_, _00668_);
  and _51395_ (_00685_, _37858_, _37832_);
  and _51396_ (_00686_, _37330_, _37602_);
  and _51397_ (_00687_, _00686_, _00685_);
  not _51398_ (_00688_, _00674_);
  and _51399_ (_00689_, _37954_, _37931_);
  and _51400_ (_00690_, _00689_, _00688_);
  and _51401_ (_00691_, _00690_, _00687_);
  or _51402_ (_00692_, _00691_, _00684_);
  and _51403_ (_00693_, _00671_, _37908_);
  and _51404_ (_00694_, _00685_, _37330_);
  and _51405_ (_00695_, _00694_, _00677_);
  and _51406_ (_00696_, _00695_, _00693_);
  not _51407_ (_00697_, _37330_);
  and _51408_ (_00698_, _00676_, _00697_);
  or _51409_ (_00699_, _00698_, _00696_);
  or _51410_ (_00700_, _00699_, _00692_);
  and _51411_ (_00701_, _00682_, _00664_);
  and _51412_ (_00702_, _00695_, _00701_);
  and _51413_ (_00703_, _37908_, _00670_);
  and _51414_ (_00704_, _00703_, _00671_);
  and _51415_ (_00705_, _00704_, _00662_);
  or _51416_ (_00706_, _00705_, _00702_);
  nor _51417_ (_00707_, _00659_, _37832_);
  nor _51418_ (_00708_, _00707_, _00697_);
  not _51419_ (_00709_, _00708_);
  and _51420_ (_00710_, _00709_, _00683_);
  not _51421_ (_00711_, _37908_);
  and _51422_ (_00712_, _00675_, _00711_);
  and _51423_ (_00713_, _00712_, _00662_);
  or _51424_ (_00714_, _00713_, _00710_);
  or _51425_ (_00715_, _00714_, _00706_);
  or _51426_ (_00716_, _00715_, _00700_);
  or _51427_ (_00717_, _00716_, _00681_);
  nor _51428_ (_00718_, _37908_, _37884_);
  and _51429_ (_00719_, _00718_, _00664_);
  nor _51430_ (_00720_, _00719_, _00677_);
  and _51431_ (_00721_, _00661_, _00659_);
  not _51432_ (_00722_, _00721_);
  nor _51433_ (_00723_, _00722_, _00720_);
  not _51434_ (_00724_, _00723_);
  and _51435_ (_00725_, _00703_, _00664_);
  and _51436_ (_00726_, _00725_, _00662_);
  and _51437_ (_00727_, _00689_, _00682_);
  and _51438_ (_00728_, _00727_, _00662_);
  nor _51439_ (_00729_, _00728_, _00726_);
  and _51440_ (_00730_, _00729_, _00724_);
  and _51441_ (_00731_, _00712_, _00694_);
  not _51442_ (_00732_, _00662_);
  and _51443_ (_00733_, _00689_, _00674_);
  and _51444_ (_00734_, _00689_, _00718_);
  nor _51445_ (_00735_, _00734_, _00733_);
  nor _51446_ (_00736_, _00735_, _00732_);
  and _51447_ (_00737_, _00733_, _00687_);
  or _51448_ (_00738_, _00737_, _00736_);
  nor _51449_ (_00739_, _00738_, _00731_);
  nand _51450_ (_00740_, _00739_, _00730_);
  or _51451_ (_00741_, _00740_, _00717_);
  and _51452_ (_00742_, _00741_, _36969_);
  not _51453_ (_00743_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _51454_ (_00744_, _36947_, _18772_);
  and _51455_ (_00745_, _00744_, _37988_);
  nor _51456_ (_00746_, _00745_, _00743_);
  or _51457_ (_00747_, _00746_, rst);
  or _51458_ (_09665_, _00747_, _00742_);
  nand _51459_ (_00748_, _37931_, _36893_);
  or _51460_ (_00749_, _36893_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _51461_ (_00750_, _00749_, _42618_);
  and _51462_ (_09668_, _00750_, _00748_);
  and _51463_ (_00751_, \oc8051_top_1.oc8051_sfr1.wait_data , _42618_);
  and _51464_ (_00752_, _00751_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or _51465_ (_00753_, _38034_, _38007_);
  and _51466_ (_00754_, _37866_, _38003_);
  or _51467_ (_00755_, _00754_, _00753_);
  and _51468_ (_00756_, _37978_, _38049_);
  and _51469_ (_00757_, _00648_, _37890_);
  or _51470_ (_00758_, _00757_, _00756_);
  and _51471_ (_00759_, _37985_, _37987_);
  and _51472_ (_00760_, _37975_, _37987_);
  or _51473_ (_00761_, _00760_, _00759_);
  or _51474_ (_00762_, _00761_, _00758_);
  nor _51475_ (_00763_, _00762_, _00755_);
  nand _51476_ (_00764_, _00763_, _38045_);
  and _51477_ (_00765_, _00764_, _00656_);
  or _51478_ (_09671_, _00765_, _00752_);
  and _51479_ (_00766_, _37971_, _37987_);
  or _51480_ (_00767_, _00766_, _37963_);
  and _51481_ (_00768_, _37395_, _37890_);
  and _51482_ (_00769_, _00768_, _38002_);
  or _51483_ (_00770_, _00769_, _38112_);
  and _51484_ (_00771_, _37977_, _38013_);
  and _51485_ (_00772_, _00771_, _38003_);
  or _51486_ (_00773_, _00772_, _00770_);
  or _51487_ (_00774_, _00773_, _00767_);
  and _51488_ (_00775_, _00774_, _36958_);
  and _51489_ (_00776_, _38092_, _00743_);
  not _51490_ (_00777_, _37981_);
  and _51491_ (_00778_, _00777_, _00776_);
  and _51492_ (_00779_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51493_ (_00780_, _00779_, _00778_);
  or _51494_ (_00781_, _00780_, _00775_);
  and _51495_ (_09674_, _00781_, _42618_);
  and _51496_ (_00782_, _00751_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _51497_ (_00783_, _37978_, _38046_);
  or _51498_ (_00784_, _38046_, _38020_);
  and _51499_ (_00785_, _00784_, _38015_);
  or _51500_ (_00786_, _00785_, _00783_);
  and _51501_ (_00787_, _00771_, _38024_);
  or _51502_ (_00788_, _00787_, _00786_);
  not _51503_ (_00789_, _38105_);
  and _51504_ (_00790_, _00784_, _37395_);
  and _51505_ (_00791_, _37395_, _37889_);
  and _51506_ (_00792_, _00791_, _38023_);
  or _51507_ (_00793_, _00792_, _00790_);
  or _51508_ (_00794_, _00793_, _00789_);
  not _51509_ (_00795_, _38084_);
  and _51510_ (_00796_, _37978_, _00795_);
  and _51511_ (_00797_, _38008_, _37395_);
  or _51512_ (_00798_, _00797_, _00767_);
  or _51513_ (_00799_, _00798_, _00796_);
  or _51514_ (_00800_, _00799_, _00794_);
  or _51515_ (_00801_, _00800_, _00788_);
  and _51516_ (_00802_, _00801_, _00656_);
  or _51517_ (_09677_, _00802_, _00782_);
  and _51518_ (_00803_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _51519_ (_00804_, _38081_, _36958_);
  or _51520_ (_00805_, _00804_, _00803_);
  or _51521_ (_00806_, _00805_, _00778_);
  and _51522_ (_09680_, _00806_, _42618_);
  and _51523_ (_00807_, _38024_, _38006_);
  and _51524_ (_00808_, _38014_, _37986_);
  and _51525_ (_00809_, _00808_, _37889_);
  or _51526_ (_00810_, _00809_, _00807_);
  or _51527_ (_00811_, _00810_, _00757_);
  and _51528_ (_00812_, _00810_, _37990_);
  or _51529_ (_00813_, _00812_, _36903_);
  and _51530_ (_00814_, _00813_, _00811_);
  not _51531_ (_00815_, _00651_);
  and _51532_ (_00816_, _00815_, _00776_);
  or _51533_ (_00817_, _00816_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51534_ (_00818_, _00817_, _00814_);
  or _51535_ (_00819_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18772_);
  and _51536_ (_00820_, _00819_, _42618_);
  and _51537_ (_09683_, _00820_, _00818_);
  and _51538_ (_00821_, _00751_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _51539_ (_00822_, _00769_, _38066_);
  and _51540_ (_00823_, _00791_, _38002_);
  or _51541_ (_00824_, _00792_, _00823_);
  or _51542_ (_00825_, _37963_, _38021_);
  or _51543_ (_00826_, _00825_, _00824_);
  or _51544_ (_00827_, _00826_, _00822_);
  and _51545_ (_00828_, _38052_, _38003_);
  and _51546_ (_00829_, _38102_, _38023_);
  or _51547_ (_00830_, _00787_, _00829_);
  or _51548_ (_00831_, _00830_, _00828_);
  or _51549_ (_00832_, _38034_, _38033_);
  or _51550_ (_00833_, _00832_, _38010_);
  or _51551_ (_00834_, _00833_, _00831_);
  or _51552_ (_00835_, _00834_, _00827_);
  and _51553_ (_00836_, _00835_, _00656_);
  or _51554_ (_09686_, _00836_, _00821_);
  and _51555_ (_00837_, _00751_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _51556_ (_00838_, _00771_, _38064_);
  and _51557_ (_00839_, _37866_, _38022_);
  or _51558_ (_00840_, _00839_, _00772_);
  or _51559_ (_00841_, _00840_, _00838_);
  or _51560_ (_00842_, _00841_, _00793_);
  not _51561_ (_00843_, _38029_);
  and _51562_ (_00844_, _37978_, _38017_);
  or _51563_ (_00845_, _00844_, _00843_);
  and _51564_ (_00846_, _38053_, _38001_);
  or _51565_ (_00847_, _00846_, _38118_);
  and _51566_ (_00848_, _38052_, _38020_);
  or _51567_ (_00849_, _00848_, _00847_);
  or _51568_ (_00850_, _00849_, _00845_);
  or _51569_ (_00851_, _00850_, _00842_);
  and _51570_ (_00852_, _00768_, _38001_);
  and _51571_ (_00853_, _00768_, _37966_);
  or _51572_ (_00854_, _00853_, _00852_);
  nor _51573_ (_00855_, _38104_, _38069_);
  nand _51574_ (_00856_, _00855_, _38019_);
  or _51575_ (_00857_, _00856_, _00854_);
  or _51576_ (_00858_, _00857_, _00788_);
  or _51577_ (_00859_, _00858_, _00851_);
  and _51578_ (_00860_, _00859_, _00656_);
  or _51579_ (_09689_, _00860_, _00837_);
  and _51580_ (_00861_, _37971_, _37395_);
  or _51581_ (_00862_, _00861_, _38110_);
  and _51582_ (_00863_, _37971_, _38052_);
  and _51583_ (_00864_, _38037_, _37395_);
  and _51584_ (_00865_, _00771_, _38037_);
  or _51585_ (_00866_, _00865_, _00864_);
  or _51586_ (_00867_, _00866_, _00863_);
  or _51587_ (_00868_, _00867_, _00862_);
  and _51588_ (_00869_, _00771_, _37971_);
  or _51589_ (_00870_, _00869_, _00868_);
  and _51590_ (_00871_, _00870_, _36958_);
  and _51591_ (_00872_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _51592_ (_00873_, _00872_, _37994_);
  or _51593_ (_00874_, _00873_, _00871_);
  and _51594_ (_09692_, _00874_, _42618_);
  nand _51595_ (_00875_, _38082_, _38070_);
  or _51596_ (_00876_, _00875_, _00785_);
  or _51597_ (_00877_, _38066_, _38035_);
  and _51598_ (_00878_, _37965_, _37889_);
  and _51599_ (_00879_, _00878_, _38015_);
  nor _51600_ (_00880_, _00879_, _38028_);
  nor _51601_ (_00881_, _00807_, _38025_);
  and _51602_ (_00882_, _00881_, _00880_);
  nand _51603_ (_00883_, _00882_, _38011_);
  or _51604_ (_00884_, _00883_, _00877_);
  or _51605_ (_00885_, _00884_, _00876_);
  and _51606_ (_00886_, _00791_, _37965_);
  or _51607_ (_00887_, _00886_, _38077_);
  and _51608_ (_00888_, _00768_, _37970_);
  or _51609_ (_00889_, _00888_, _00809_);
  or _51610_ (_00890_, _00889_, _00770_);
  or _51611_ (_00891_, _00890_, _00887_);
  and _51612_ (_00892_, _00878_, _38052_);
  or _51613_ (_00893_, _00892_, _38104_);
  or _51614_ (_00894_, _00893_, _38054_);
  or _51615_ (_00895_, _38106_, _38074_);
  or _51616_ (_00896_, _00895_, _00894_);
  or _51617_ (_00897_, _00896_, _00891_);
  or _51618_ (_00898_, _00897_, _00793_);
  or _51619_ (_00899_, _00898_, _00885_);
  and _51620_ (_00900_, _00899_, _36958_);
  and _51621_ (_00901_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51622_ (_00902_, _00812_, _00778_);
  and _51623_ (_00903_, _37990_, _38043_);
  or _51624_ (_00904_, _00903_, _00902_);
  or _51625_ (_00905_, _00904_, _00901_);
  or _51626_ (_00906_, _00905_, _00900_);
  and _51627_ (_09695_, _00906_, _42618_);
  nor _51628_ (_09754_, _38131_, rst);
  nor _51629_ (_09756_, _38097_, rst);
  or _51630_ (_09759_, _00657_, _00651_);
  nor _51631_ (_00907_, _00648_, _00645_);
  or _51632_ (_09762_, _00907_, _00657_);
  and _51633_ (_00908_, _00689_, _00711_);
  and _51634_ (_00909_, _00908_, _00687_);
  or _51635_ (_00910_, _00909_, _00673_);
  or _51636_ (_00911_, _00696_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _51637_ (_00912_, _00911_, _00910_);
  and _51638_ (_00913_, _00912_, _00745_);
  nor _51639_ (_00914_, _00744_, _37988_);
  or _51640_ (_00915_, _00914_, rst);
  or _51641_ (_09765_, _00915_, _00913_);
  nand _51642_ (_00916_, _37602_, _36893_);
  or _51643_ (_00917_, _36893_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _51644_ (_00918_, _00917_, _42618_);
  and _51645_ (_09768_, _00918_, _00916_);
  or _51646_ (_00919_, _37858_, _37993_);
  or _51647_ (_00920_, _36893_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _51648_ (_00921_, _00920_, _42618_);
  and _51649_ (_09771_, _00921_, _00919_);
  nand _51650_ (_00922_, _37832_, _36893_);
  or _51651_ (_00923_, _36893_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _51652_ (_00924_, _00923_, _42618_);
  and _51653_ (_09774_, _00924_, _00922_);
  nand _51654_ (_00926_, _37330_, _36893_);
  or _51655_ (_00927_, _36893_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _51656_ (_00928_, _00927_, _42618_);
  and _51657_ (_09777_, _00928_, _00926_);
  or _51658_ (_00929_, _37884_, _37993_);
  or _51659_ (_00930_, _36893_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _51660_ (_00931_, _00930_, _42618_);
  and _51661_ (_09780_, _00931_, _00929_);
  nand _51662_ (_00932_, _37908_, _36893_);
  or _51663_ (_00933_, _36893_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _51664_ (_00934_, _00933_, _42618_);
  and _51665_ (_09783_, _00934_, _00932_);
  nand _51666_ (_00935_, _37954_, _36893_);
  or _51667_ (_00936_, _36893_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _51668_ (_00937_, _00936_, _42618_);
  and _51669_ (_09786_, _00937_, _00935_);
  or _51670_ (_00938_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _18772_);
  and _51671_ (_00939_, _00938_, _42618_);
  and _51672_ (_00940_, _00939_, _00817_);
  not _51673_ (_00941_, _38061_);
  and _51674_ (_00942_, _00771_, _00941_);
  and _51675_ (_00943_, _00771_, _38017_);
  or _51676_ (_00944_, _00943_, _00766_);
  or _51677_ (_00945_, _00771_, _37395_);
  or _51678_ (_00946_, _38064_, _38049_);
  and _51679_ (_00947_, _00946_, _00945_);
  or _51680_ (_00948_, _00947_, _00944_);
  or _51681_ (_00949_, _00948_, _00942_);
  or _51682_ (_00950_, _38123_, _00863_);
  and _51683_ (_00952_, _38060_, _38052_);
  or _51684_ (_00953_, _00952_, _38118_);
  or _51685_ (_00954_, _00953_, _00950_);
  and _51686_ (_00955_, _00768_, _38016_);
  or _51687_ (_00956_, _00955_, _00839_);
  or _51688_ (_00957_, _00956_, _37963_);
  or _51689_ (_00958_, _00957_, _00862_);
  or _51690_ (_00959_, _00958_, _00954_);
  nor _51691_ (_00960_, _38061_, _37406_);
  or _51692_ (_00961_, _00960_, _00869_);
  or _51693_ (_00962_, _38023_, _38020_);
  or _51694_ (_00963_, _00962_, _00878_);
  and _51695_ (_00964_, _00963_, _37978_);
  or _51696_ (_00965_, _00964_, _00961_);
  or _51697_ (_00966_, _00965_, _00959_);
  or _51698_ (_00967_, _00966_, _00949_);
  and _51699_ (_00968_, _00967_, _00656_);
  or _51700_ (_09789_, _00968_, _00940_);
  and _51701_ (_00969_, _00751_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _51702_ (_00970_, _38064_, _38017_);
  and _51703_ (_00972_, _00970_, _38006_);
  and _51704_ (_00973_, _00791_, _37961_);
  nor _51705_ (_00974_, _00973_, _38103_);
  nand _51706_ (_00975_, _37978_, _00941_);
  nand _51707_ (_00976_, _00975_, _00974_);
  or _51708_ (_00977_, _00976_, _00972_);
  or _51709_ (_00978_, _00796_, _00758_);
  or _51710_ (_00979_, _00944_, _00854_);
  or _51711_ (_00980_, _00979_, _00978_);
  not _51712_ (_00981_, _38067_);
  and _51713_ (_00982_, _37978_, _38064_);
  or _51714_ (_00983_, _00982_, _00981_);
  or _51715_ (_00984_, _00983_, _00849_);
  or _51716_ (_00985_, _00984_, _00980_);
  or _51717_ (_00986_, _00985_, _00977_);
  and _51718_ (_00987_, _00986_, _00656_);
  or _51719_ (_34182_, _00987_, _00969_);
  or _51720_ (_00988_, _00895_, _00889_);
  or _51721_ (_00989_, _00988_, _00885_);
  and _51722_ (_00990_, _00989_, _36958_);
  and _51723_ (_00991_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51724_ (_00992_, _00991_, _00904_);
  or _51725_ (_00993_, _00992_, _00990_);
  and _51726_ (_34184_, _00993_, _42618_);
  and _51727_ (_00994_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51728_ (_00995_, _00994_, _00902_);
  and _51729_ (_00996_, _00995_, _42618_);
  and _51730_ (_00997_, _38068_, _37890_);
  or _51731_ (_00998_, _00997_, _38112_);
  or _51732_ (_00999_, _00998_, _00810_);
  or _51733_ (_01000_, _00999_, _00894_);
  and _51734_ (_01001_, _01000_, _00656_);
  or _51735_ (_34187_, _01001_, _00996_);
  or _51736_ (_01002_, _00648_, _37980_);
  and _51737_ (_01003_, _00771_, _38060_);
  and _51738_ (_01004_, _00865_, _37889_);
  or _51739_ (_01005_, _01004_, _01003_);
  or _51740_ (_01006_, _01005_, _01002_);
  or _51741_ (_01007_, _00861_, _38111_);
  and _51742_ (_01008_, _00652_, _38015_);
  and _51743_ (_01009_, _37978_, _37967_);
  and _51744_ (_01010_, _38060_, _38006_);
  or _51745_ (_01011_, _01010_, _01009_);
  or _51746_ (_01012_, _01011_, _01008_);
  or _51747_ (_01013_, _01012_, _01007_);
  or _51748_ (_01014_, _01013_, _01006_);
  and _51749_ (_01015_, _00771_, _38008_);
  or _51750_ (_01016_, _01015_, _00756_);
  and _51751_ (_01017_, _00652_, _37978_);
  or _51752_ (_01018_, _01017_, _37979_);
  or _51753_ (_01019_, _01018_, _01016_);
  and _51754_ (_01020_, _00962_, _37978_);
  or _51755_ (_01021_, _01020_, _01019_);
  and _51756_ (_01022_, _37978_, _38003_);
  or _51757_ (_01023_, _00839_, _01022_);
  or _51758_ (_01024_, _01023_, _00961_);
  or _51759_ (_01025_, _00844_, _00863_);
  and _51760_ (_01026_, _00865_, _37890_);
  or _51761_ (_01027_, _01026_, _00982_);
  or _51762_ (_01028_, _01027_, _01025_);
  or _51763_ (_01029_, _00892_, _00886_);
  or _51764_ (_01030_, _01029_, _37968_);
  or _51765_ (_01031_, _01030_, _00810_);
  or _51766_ (_01032_, _01031_, _01028_);
  or _51767_ (_01033_, _01032_, _01024_);
  or _51768_ (_01034_, _01033_, _01021_);
  or _51769_ (_01035_, _01034_, _01014_);
  and _51770_ (_01036_, _01035_, _36958_);
  and _51771_ (_01037_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51772_ (_01038_, _00816_, _37995_);
  or _51773_ (_01039_, _01038_, _01037_);
  or _51774_ (_01040_, _01039_, _01036_);
  and _51775_ (_34189_, _01040_, _42618_);
  and _51776_ (_01041_, _00791_, _38048_);
  or _51777_ (_01042_, _01041_, _00879_);
  nor _51778_ (_01043_, _01042_, _00863_);
  nand _51779_ (_01044_, _01043_, _37973_);
  and _51780_ (_01045_, _00970_, _37866_);
  or _51781_ (_01046_, _01045_, _38062_);
  or _51782_ (_01047_, _01046_, _01044_);
  or _51783_ (_01048_, _37980_, _38074_);
  and _51784_ (_01049_, _00652_, _38052_);
  or _51785_ (_01050_, _01049_, _00766_);
  or _51786_ (_01051_, _01050_, _01048_);
  or _51787_ (_01052_, _01051_, _01007_);
  or _51788_ (_01053_, _01052_, _01047_);
  or _51789_ (_01054_, _01024_, _01021_);
  or _51790_ (_01055_, _01054_, _01053_);
  and _51791_ (_01056_, _01055_, _36958_);
  and _51792_ (_01057_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51793_ (_01058_, _01057_, _01038_);
  or _51794_ (_01059_, _01058_, _01056_);
  and _51795_ (_34191_, _01059_, _42618_);
  and _51796_ (_01060_, _00751_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _51797_ (_01061_, _00828_, _00829_);
  or _51798_ (_01062_, _01061_, _01004_);
  nor _51799_ (_01063_, _00863_, _38080_);
  nand _51800_ (_01064_, _01063_, _42104_);
  or _51801_ (_01065_, _01064_, _01062_);
  not _51802_ (_01066_, _42102_);
  or _51803_ (_01067_, _00869_, _01066_);
  or _51804_ (_01068_, _01067_, _00877_);
  or _51805_ (_01069_, _01068_, _01065_);
  or _51806_ (_01070_, _00861_, _00769_);
  or _51807_ (_01071_, _38051_, _37395_);
  or _51808_ (_01072_, _01071_, _37866_);
  and _51809_ (_01073_, _01072_, _38038_);
  and _51810_ (_01074_, _38009_, _37657_);
  or _51811_ (_01075_, _01074_, _01073_);
  or _51812_ (_01076_, _01075_, _01070_);
  or _51813_ (_01077_, _38024_, _38020_);
  and _51814_ (_01078_, _01077_, _37866_);
  and _51815_ (_01079_, _37978_, _38020_);
  or _51816_ (_01080_, _01079_, _00787_);
  or _51817_ (_01081_, _01080_, _01078_);
  or _51818_ (_01082_, _01081_, _00826_);
  or _51819_ (_01083_, _01082_, _01076_);
  or _51820_ (_01084_, _01083_, _01069_);
  and _51821_ (_01085_, _01084_, _00656_);
  or _51822_ (_34193_, _01085_, _01060_);
  and _51823_ (_01086_, _00751_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _51824_ (_01087_, _37866_, _38024_);
  or _51825_ (_01088_, _01026_, _00848_);
  or _51826_ (_01089_, _01088_, _01087_);
  or _51827_ (_01090_, _01089_, _00845_);
  or _51828_ (_01091_, _01090_, _01006_);
  and _51829_ (_01092_, _38038_, _37866_);
  or _51830_ (_01093_, _01092_, _01079_);
  not _51831_ (_01094_, _38075_);
  or _51832_ (_01095_, _00960_, _01094_);
  or _51833_ (_01096_, _01095_, _01093_);
  or _51834_ (_01097_, _37968_, _38018_);
  or _51835_ (_01098_, _00846_, _00772_);
  or _51836_ (_01099_, _01098_, _01097_);
  or _51837_ (_01100_, _00852_, _36914_);
  or _51838_ (_01101_, _01100_, _37963_);
  or _51839_ (_01102_, _01101_, _38111_);
  or _51840_ (_01103_, _01102_, _01099_);
  or _51841_ (_01104_, _01103_, _01096_);
  or _51842_ (_01105_, _01104_, _01091_);
  or _51843_ (_01106_, _37980_, _36903_);
  nor _51844_ (_01107_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and _51845_ (_01108_, _01107_, _01106_);
  and _51846_ (_01109_, _01108_, _01105_);
  or _51847_ (_34195_, _01109_, _01086_);
  and _51848_ (_01110_, _00751_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not _51849_ (_01111_, _01003_);
  and _51850_ (_01112_, _01111_, _38075_);
  and _51851_ (_01113_, _38060_, _37395_);
  or _51852_ (_01114_, _01113_, _00869_);
  or _51853_ (_01115_, _01114_, _00952_);
  nor _51854_ (_01116_, _01115_, _00786_);
  nand _51855_ (_01117_, _01116_, _01112_);
  or _51856_ (_01118_, _01017_, _38009_);
  or _51857_ (_01119_, _01070_, _01016_);
  or _51858_ (_01120_, _01119_, _01118_);
  or _51859_ (_01121_, _00772_, _42103_);
  or _51860_ (_01122_, _00797_, _00787_);
  or _51861_ (_01123_, _01122_, _01121_);
  and _51862_ (_01124_, _38037_, _37866_);
  or _51863_ (_01125_, _01124_, _37980_);
  or _51864_ (_01126_, _01125_, _38115_);
  or _51865_ (_01127_, _01126_, _01123_);
  or _51866_ (_01128_, _01127_, _01120_);
  or _51867_ (_01129_, _01128_, _00794_);
  or _51868_ (_01130_, _01129_, _01117_);
  and _51869_ (_01131_, _01130_, _01108_);
  or _51870_ (_34197_, _01131_, _01110_);
  or _51871_ (_01132_, _01080_, _00822_);
  or _51872_ (_01133_, _01132_, _01118_);
  and _51873_ (_01134_, _01071_, _38060_);
  or _51874_ (_01135_, _01003_, _38074_);
  or _51875_ (_01136_, _01135_, _01134_);
  and _51876_ (_01137_, _37866_, _38023_);
  or _51877_ (_01138_, _38112_, _38104_);
  nor _51878_ (_01139_, _01138_, _01137_);
  nand _51879_ (_01140_, _01139_, _42102_);
  or _51880_ (_01141_, _01140_, _01136_);
  or _51881_ (_01142_, _00793_, _00786_);
  or _51882_ (_01143_, _01142_, _01141_);
  or _51883_ (_01144_, _01143_, _01133_);
  and _51884_ (_01145_, _01144_, _36958_);
  and _51885_ (_01146_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _51886_ (_01147_, _37979_, _18772_);
  or _51887_ (_01148_, _01147_, _01146_);
  or _51888_ (_01149_, _01148_, _01145_);
  and _51889_ (_34199_, _01149_, _42618_);
  and _51890_ (_01150_, _00751_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _51891_ (_01151_, _01078_, _42105_);
  or _51892_ (_01152_, _01093_, _01074_);
  or _51893_ (_01153_, _01152_, _01151_);
  or _51894_ (_01154_, _00754_, _38033_);
  not _51895_ (_01155_, _37986_);
  and _51896_ (_01156_, _38008_, _01155_);
  or _51897_ (_01157_, _01156_, _01154_);
  or _51898_ (_01158_, _01157_, _00868_);
  or _51899_ (_01159_, _01158_, _01067_);
  or _51900_ (_01160_, _01159_, _01153_);
  and _51901_ (_01161_, _01160_, _00656_);
  or _51902_ (_34201_, _01161_, _01150_);
  nor _51903_ (_38643_, _37931_, rst);
  nor _51904_ (_38644_, _42095_, rst);
  and _51905_ (_01162_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _51906_ (_01163_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _51907_ (_01164_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _51908_ (_01165_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _51909_ (_01166_, _01165_, _01164_);
  and _51910_ (_01167_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _51911_ (_01168_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _51912_ (_01169_, _01168_, _01167_);
  and _51913_ (_01170_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _51914_ (_01171_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _51915_ (_01172_, _01171_, _01170_);
  and _51916_ (_01173_, _01172_, _01169_);
  and _51917_ (_01174_, _01173_, _01166_);
  nor _51918_ (_01175_, _01174_, _37012_);
  nor _51919_ (_01176_, _01175_, _01163_);
  nor _51920_ (_01177_, _01176_, _42079_);
  nor _51921_ (_01178_, _01177_, _01162_);
  nor _51922_ (_38646_, _01178_, rst);
  nor _51923_ (_38656_, _37602_, rst);
  and _51924_ (_38658_, _37858_, _42618_);
  nor _51925_ (_38659_, _37832_, rst);
  nor _51926_ (_38660_, _37330_, rst);
  and _51927_ (_38661_, _37884_, _42618_);
  nor _51928_ (_38662_, _37908_, rst);
  nor _51929_ (_38663_, _37954_, rst);
  nor _51930_ (_38664_, _42391_, rst);
  nor _51931_ (_38665_, _42298_, rst);
  nor _51932_ (_38667_, _42207_, rst);
  nor _51933_ (_38668_, _42349_, rst);
  nor _51934_ (_38669_, _42253_, rst);
  nor _51935_ (_38670_, _42131_, rst);
  nor _51936_ (_38671_, _42446_, rst);
  and _51937_ (_01179_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _51938_ (_01180_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _51939_ (_01181_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _51940_ (_01182_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _51941_ (_01183_, _01182_, _01181_);
  and _51942_ (_01184_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _51943_ (_01185_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _51944_ (_01186_, _01185_, _01184_);
  and _51945_ (_01187_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _51946_ (_01188_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _51947_ (_01189_, _01188_, _01187_);
  and _51948_ (_01190_, _01189_, _01186_);
  and _51949_ (_01191_, _01190_, _01183_);
  nor _51950_ (_01192_, _01191_, _37012_);
  nor _51951_ (_01193_, _01192_, _01180_);
  nor _51952_ (_01194_, _01193_, _42079_);
  nor _51953_ (_01195_, _01194_, _01179_);
  nor _51954_ (_38673_, _01195_, rst);
  and _51955_ (_01196_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _51956_ (_01197_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _51957_ (_01198_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _51958_ (_01199_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _51959_ (_01200_, _01199_, _01198_);
  and _51960_ (_01201_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _51961_ (_01202_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _51962_ (_01203_, _01202_, _01201_);
  and _51963_ (_01204_, _01203_, _01200_);
  and _51964_ (_01205_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _51965_ (_01207_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _51966_ (_01209_, _01207_, _01205_);
  and _51967_ (_01211_, _01209_, _01204_);
  nor _51968_ (_01213_, _01211_, _37012_);
  nor _51969_ (_01215_, _01213_, _01197_);
  nor _51970_ (_01217_, _01215_, _42079_);
  nor _51971_ (_01219_, _01217_, _01196_);
  nor _51972_ (_38674_, _01219_, rst);
  and _51973_ (_01222_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _51974_ (_01224_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _51975_ (_01226_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _51976_ (_01228_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _51977_ (_01230_, _01228_, _01226_);
  and _51978_ (_01232_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _51979_ (_01234_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _51980_ (_01236_, _01234_, _01232_);
  and _51981_ (_01238_, _01236_, _01230_);
  and _51982_ (_01240_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _51983_ (_01242_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _51984_ (_01244_, _01242_, _01240_);
  and _51985_ (_01246_, _01244_, _01238_);
  nor _51986_ (_01248_, _01246_, _37012_);
  nor _51987_ (_01250_, _01248_, _01224_);
  nor _51988_ (_01252_, _01250_, _42079_);
  nor _51989_ (_01254_, _01252_, _01222_);
  nor _51990_ (_38675_, _01254_, rst);
  and _51991_ (_01257_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _51992_ (_01259_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _51993_ (_01261_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _51994_ (_01263_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _51995_ (_01265_, _01263_, _01261_);
  and _51996_ (_01267_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _51997_ (_01269_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _51998_ (_01271_, _01269_, _01267_);
  and _51999_ (_01273_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _52000_ (_01275_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _52001_ (_01277_, _01275_, _01273_);
  and _52002_ (_01279_, _01277_, _01271_);
  and _52003_ (_01281_, _01279_, _01265_);
  nor _52004_ (_01283_, _01281_, _37012_);
  nor _52005_ (_01285_, _01283_, _01259_);
  nor _52006_ (_01287_, _01285_, _42079_);
  nor _52007_ (_01289_, _01287_, _01257_);
  nor _52008_ (_38676_, _01289_, rst);
  and _52009_ (_01292_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _52010_ (_01294_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _52011_ (_01296_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _52012_ (_01298_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _52013_ (_01300_, _01298_, _01296_);
  and _52014_ (_01301_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _52015_ (_01302_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _52016_ (_01303_, _01302_, _01301_);
  and _52017_ (_01304_, _01303_, _01300_);
  and _52018_ (_01305_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _52019_ (_01306_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _52020_ (_01307_, _01306_, _01305_);
  and _52021_ (_01308_, _01307_, _01304_);
  nor _52022_ (_01309_, _01308_, _37012_);
  nor _52023_ (_01310_, _01309_, _01294_);
  nor _52024_ (_01311_, _01310_, _42079_);
  nor _52025_ (_01312_, _01311_, _01292_);
  nor _52026_ (_38677_, _01312_, rst);
  and _52027_ (_01313_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _52028_ (_01314_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _52029_ (_01315_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _52030_ (_01316_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _52031_ (_01317_, _01316_, _01315_);
  and _52032_ (_01318_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _52033_ (_01319_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _52034_ (_01320_, _01319_, _01318_);
  and _52035_ (_01321_, _01320_, _01317_);
  and _52036_ (_01322_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _52037_ (_01323_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _52038_ (_01324_, _01323_, _01322_);
  and _52039_ (_01325_, _01324_, _01321_);
  nor _52040_ (_01326_, _01325_, _37012_);
  nor _52041_ (_01327_, _01326_, _01314_);
  nor _52042_ (_01328_, _01327_, _42079_);
  nor _52043_ (_01329_, _01328_, _01313_);
  nor _52044_ (_38679_, _01329_, rst);
  and _52045_ (_01330_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _52046_ (_01331_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _52047_ (_01332_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _52048_ (_01333_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _52049_ (_01334_, _01333_, _01332_);
  and _52050_ (_01335_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _52051_ (_01336_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _52052_ (_01337_, _01336_, _01335_);
  and _52053_ (_01338_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _52054_ (_01339_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _52055_ (_01340_, _01339_, _01338_);
  and _52056_ (_01341_, _01340_, _01337_);
  and _52057_ (_01342_, _01341_, _01334_);
  nor _52058_ (_01343_, _01342_, _37012_);
  nor _52059_ (_01344_, _01343_, _01331_);
  nor _52060_ (_01345_, _01344_, _42079_);
  nor _52061_ (_01346_, _01345_, _01330_);
  nor _52062_ (_38680_, _01346_, rst);
  and _52063_ (_01347_, _36969_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _52064_ (_01348_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _52065_ (_01349_, _01347_, _38317_);
  and _52066_ (_01350_, _01349_, _42618_);
  and _52067_ (_38705_, _01350_, _01348_);
  not _52068_ (_01351_, _01347_);
  or _52069_ (_01352_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _52070_ (_01353_, _36969_, _42618_);
  and _52071_ (_01354_, _01353_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _52072_ (_01355_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _42618_);
  or _52073_ (_01356_, _01355_, _01354_);
  and _52074_ (_38706_, _01356_, _01352_);
  nor _52075_ (_38741_, _42100_, rst);
  nor _52076_ (_38744_, _42072_, rst);
  nor _52077_ (_01357_, _42354_, _27948_);
  and _52078_ (_01358_, _42354_, _27948_);
  nor _52079_ (_01359_, _01358_, _01357_);
  not _52080_ (_01360_, _01359_);
  nor _52081_ (_01361_, _42451_, _28376_);
  and _52082_ (_01362_, _42451_, _28376_);
  nor _52083_ (_01363_, _01362_, _01361_);
  not _52084_ (_01364_, _01363_);
  and _52085_ (_01365_, _01364_, _42548_);
  nor _52086_ (_01366_, _42259_, _27542_);
  and _52087_ (_01367_, _42259_, _27542_);
  nor _52088_ (_01368_, _01367_, _01366_);
  nor _52089_ (_01369_, _42164_, _27345_);
  and _52090_ (_01370_, _42164_, _27345_);
  nor _52091_ (_01371_, _01370_, _01369_);
  nor _52092_ (_01372_, _01371_, _01368_);
  and _52093_ (_01373_, _01372_, _01365_);
  and _52094_ (_01374_, _01373_, _01360_);
  nor _52095_ (_01375_, _42307_, _33107_);
  and _52096_ (_01376_, _42307_, _33107_);
  or _52097_ (_01377_, _01376_, _01375_);
  nor _52098_ (_01378_, _01377_, _38947_);
  nor _52099_ (_01379_, _42400_, _27795_);
  and _52100_ (_01380_, _42400_, _27795_);
  nor _52101_ (_01381_, _01380_, _01379_);
  nor _52102_ (_01382_, _42212_, _28069_);
  and _52103_ (_01383_, _42212_, _28069_);
  nor _52104_ (_01384_, _01383_, _01382_);
  nor _52105_ (_01385_, _01384_, _01381_);
  and _52106_ (_01386_, _01385_, _01378_);
  and _52107_ (_01387_, _01386_, _01374_);
  nor _52108_ (_01388_, _28244_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _52109_ (_01389_, _01388_, _01387_);
  not _52110_ (_01390_, _01389_);
  nor _52111_ (_01391_, _38045_, _38092_);
  nor _52112_ (_01392_, _31855_, _39551_);
  and _52113_ (_01393_, _01392_, _01374_);
  and _52114_ (_01394_, _01393_, _01391_);
  and _52115_ (_01395_, _38023_, _38006_);
  nor _52116_ (_01396_, _01395_, _00808_);
  nor _52117_ (_01397_, _01396_, _36914_);
  and _52118_ (_01398_, _33379_, _29987_);
  nand _52119_ (_01399_, _01398_, _34064_);
  nor _52120_ (_01400_, _01399_, _34760_);
  and _52121_ (_01401_, _01400_, _35577_);
  nand _52122_ (_01402_, _01401_, _36295_);
  nor _52123_ (_01403_, _01402_, _31996_);
  nor _52124_ (_01404_, _01391_, _37992_);
  and _52125_ (_01405_, _01404_, _01403_);
  and _52126_ (_01406_, _01405_, _30173_);
  not _52127_ (_01407_, _01406_);
  and _52128_ (_01408_, _01391_, _29143_);
  not _52129_ (_01409_, _01408_);
  not _52130_ (_01410_, _37992_);
  nor _52131_ (_01411_, _01391_, _38016_);
  nor _52132_ (_01412_, _01411_, _01410_);
  and _52133_ (_01413_, _01412_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _52134_ (_01414_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _52135_ (_01415_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _52136_ (_01416_, _01415_, _01414_);
  nor _52137_ (_01417_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _52138_ (_01418_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _52139_ (_01419_, _01418_, _01417_);
  and _52140_ (_01420_, _01419_, _01416_);
  and _52141_ (_01421_, _01420_, _38129_);
  nor _52142_ (_01422_, _01421_, _01413_);
  and _52143_ (_01423_, _01422_, _01409_);
  and _52144_ (_01424_, _01423_, _01407_);
  and _52145_ (_01425_, _00759_, _37890_);
  not _52146_ (_01426_, _01425_);
  and _52147_ (_01427_, _01426_, _38044_);
  nor _52148_ (_01428_, _01427_, _01424_);
  not _52149_ (_01429_, _01428_);
  not _52150_ (_01430_, _37987_);
  or _52151_ (_01431_, _38038_, _37967_);
  nor _52152_ (_01432_, _01431_, _38060_);
  nor _52153_ (_01433_, _01432_, _01430_);
  not _52154_ (_01434_, _01433_);
  nor _52155_ (_01435_, _01015_, _38021_);
  not _52156_ (_01436_, _01435_);
  nor _52157_ (_01437_, _01436_, _00823_);
  and _52158_ (_01438_, _01437_, _00974_);
  and _52159_ (_01439_, _01438_, _01434_);
  not _52160_ (_01440_, _01439_);
  and _52161_ (_01441_, _01440_, _01424_);
  or _52162_ (_01442_, _37968_, _38076_);
  or _52163_ (_01443_, _01442_, _00760_);
  nor _52164_ (_01444_, _01443_, _01441_);
  and _52165_ (_01445_, _01444_, _01429_);
  nor _52166_ (_01446_, _37990_, _38094_);
  nor _52167_ (_01447_, _01446_, _01445_);
  nor _52168_ (_01448_, _01447_, _01397_);
  not _52169_ (_01449_, _38889_);
  and _52170_ (_01450_, _01449_, _38129_);
  nor _52171_ (_01451_, _38624_, _38616_);
  and _52172_ (_01452_, _01451_, _38638_);
  not _52173_ (_01453_, _01452_);
  and _52174_ (_01454_, _01453_, _01412_);
  nor _52175_ (_01455_, _01454_, _01450_);
  not _52176_ (_01456_, _01455_);
  nor _52177_ (_01457_, _01456_, _01448_);
  not _52178_ (_01458_, _01457_);
  nor _52179_ (_01459_, _01458_, _01394_);
  and _52180_ (_01460_, _01459_, _01390_);
  nor _52181_ (_01461_, _38094_, rst);
  and _52182_ (_38748_, _01461_, _01460_);
  and _52183_ (_38749_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _42618_);
  and _52184_ (_38750_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _42618_);
  and _52185_ (_01462_, _38094_, _31147_);
  not _52186_ (_01463_, _38368_);
  and _52187_ (_01464_, _37968_, _37990_);
  and _52188_ (_01465_, _01464_, _01463_);
  nand _52189_ (_01466_, _00974_, _38045_);
  or _52190_ (_01467_, _01466_, _01436_);
  and _52191_ (_01468_, _01467_, _37990_);
  and _52192_ (_01469_, _01395_, _36903_);
  not _52193_ (_01470_, _01469_);
  and _52194_ (_01471_, _38037_, _36903_);
  and _52195_ (_01472_, _01471_, _37987_);
  nor _52196_ (_01473_, _01472_, _38094_);
  and _52197_ (_01474_, _01473_, _01470_);
  not _52198_ (_01475_, _01474_);
  nor _52199_ (_01476_, _01475_, _01468_);
  nor _52200_ (_01477_, _01464_, _01397_);
  nor _52201_ (_01478_, _00761_, _37968_);
  nand _52202_ (_01479_, _01478_, _01437_);
  or _52203_ (_01480_, _01479_, _01466_);
  and _52204_ (_01481_, _01480_, _37990_);
  nor _52205_ (_01482_, _01481_, _01472_);
  and _52206_ (_01483_, _01482_, _01477_);
  and _52207_ (_01484_, _01483_, _01476_);
  and _52208_ (_01485_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _52209_ (_01486_, _01469_, _42096_);
  or _52210_ (_01487_, _01486_, _01485_);
  or _52211_ (_01488_, _01487_, _01465_);
  or _52212_ (_01489_, _01488_, _01462_);
  and _52213_ (_01490_, _01476_, _42095_);
  not _52214_ (_01491_, _01178_);
  nor _52215_ (_01492_, _01476_, _01491_);
  nor _52216_ (_01493_, _01492_, _01490_);
  and _52217_ (_01494_, _01493_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _52218_ (_01495_, _01493_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _52219_ (_01496_, _01476_, _42446_);
  not _52220_ (_01497_, _01346_);
  nor _52221_ (_01498_, _01476_, _01497_);
  nor _52222_ (_01499_, _01498_, _01496_);
  nand _52223_ (_01500_, _01499_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _52224_ (_01501_, _01499_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _52225_ (_01502_, _01501_, _01500_);
  and _52226_ (_01503_, _01476_, _42131_);
  not _52227_ (_01504_, _01329_);
  nor _52228_ (_01505_, _01476_, _01504_);
  nor _52229_ (_01506_, _01505_, _01503_);
  and _52230_ (_01507_, _01506_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _52231_ (_01508_, _01506_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _52232_ (_01509_, _01476_, _42253_);
  not _52233_ (_01510_, _01312_);
  nor _52234_ (_01511_, _01476_, _01510_);
  nor _52235_ (_01512_, _01511_, _01509_);
  nand _52236_ (_01513_, _01512_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52237_ (_01514_, _01476_, _42349_);
  not _52238_ (_01515_, _01289_);
  nor _52239_ (_01516_, _01476_, _01515_);
  nor _52240_ (_01517_, _01516_, _01514_);
  and _52241_ (_01518_, _01517_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _52242_ (_01519_, _01517_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _52243_ (_01520_, _01476_, _42207_);
  not _52244_ (_01521_, _01254_);
  nor _52245_ (_01522_, _01476_, _01521_);
  nor _52246_ (_01523_, _01522_, _01520_);
  and _52247_ (_01524_, _01523_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _52248_ (_01525_, _01476_, _42298_);
  not _52249_ (_01526_, _01219_);
  nor _52250_ (_01527_, _01476_, _01526_);
  nor _52251_ (_01528_, _01527_, _01525_);
  and _52252_ (_01529_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _52253_ (_01530_, _01476_, _42391_);
  not _52254_ (_01531_, _01195_);
  nor _52255_ (_01532_, _01476_, _01531_);
  nor _52256_ (_01533_, _01532_, _01530_);
  and _52257_ (_01534_, _01533_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _52258_ (_01535_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _52259_ (_01536_, _01535_, _01529_);
  and _52260_ (_01537_, _01536_, _01534_);
  nor _52261_ (_01538_, _01537_, _01529_);
  not _52262_ (_01539_, _01538_);
  nor _52263_ (_01540_, _01523_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _52264_ (_01541_, _01540_, _01524_);
  and _52265_ (_01542_, _01541_, _01539_);
  nor _52266_ (_01543_, _01542_, _01524_);
  nor _52267_ (_01544_, _01543_, _01519_);
  or _52268_ (_01545_, _01544_, _01518_);
  or _52269_ (_01546_, _01512_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52270_ (_01547_, _01546_, _01513_);
  nand _52271_ (_01548_, _01547_, _01545_);
  and _52272_ (_01549_, _01548_, _01513_);
  nor _52273_ (_01550_, _01549_, _01508_);
  or _52274_ (_01551_, _01550_, _01507_);
  nand _52275_ (_01552_, _01551_, _01502_);
  and _52276_ (_01553_, _01552_, _01500_);
  nor _52277_ (_01554_, _01553_, _01495_);
  or _52278_ (_01555_, _01554_, _01494_);
  and _52279_ (_01556_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _52280_ (_01557_, _01556_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _52281_ (_01558_, _01557_, _01555_);
  and _52282_ (_01559_, _01558_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _52283_ (_01560_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52284_ (_01561_, _01560_, _01559_);
  nor _52285_ (_01562_, _01561_, _01493_);
  not _52286_ (_01563_, _01493_);
  nor _52287_ (_01564_, _01555_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _52288_ (_01565_, _01564_, _38291_);
  and _52289_ (_01566_, _01565_, _38296_);
  and _52290_ (_01567_, _01566_, _38281_);
  nor _52291_ (_01568_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52292_ (_01569_, _01568_, _01567_);
  nor _52293_ (_01570_, _01569_, _01563_);
  nor _52294_ (_01571_, _01570_, _01562_);
  or _52295_ (_01572_, _01493_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _52296_ (_01573_, _01493_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _52297_ (_01574_, _01573_, _01572_);
  and _52298_ (_01575_, _01574_, _01571_);
  or _52299_ (_01576_, _01575_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _52300_ (_01577_, _01575_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _52301_ (_01578_, _01477_);
  and _52302_ (_01579_, _01578_, _01476_);
  and _52303_ (_01580_, _37987_, _36903_);
  and _52304_ (_01581_, _01580_, _38037_);
  nor _52305_ (_01582_, _01481_, _01581_);
  nor _52306_ (_01583_, _01582_, _01579_);
  and _52307_ (_01584_, _01583_, _01577_);
  and _52308_ (_01585_, _01584_, _01576_);
  or _52309_ (_01586_, _01585_, _01489_);
  and _52310_ (_01587_, _01482_, _01579_);
  and _52311_ (_01588_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52312_ (_01589_, _01588_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _52313_ (_01590_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _52314_ (_01591_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _52315_ (_01592_, _01591_, _01590_);
  and _52316_ (_01593_, _01592_, _01589_);
  and _52317_ (_01594_, _01593_, _01557_);
  and _52318_ (_01595_, _01594_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _52319_ (_01596_, _01595_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52320_ (_01597_, _01596_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _52321_ (_01598_, _01597_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _52322_ (_01599_, _01598_, _38317_);
  or _52323_ (_01600_, _01598_, _38317_);
  and _52324_ (_01601_, _01600_, _01599_);
  nand _52325_ (_01602_, _01601_, _01587_);
  nand _52326_ (_01603_, _01602_, _01460_);
  or _52327_ (_01604_, _01603_, _01586_);
  and _52328_ (_01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _52329_ (_01606_, _37067_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _52330_ (_01607_, _01606_, _42079_);
  nor _52331_ (_01608_, _01607_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _52332_ (_01609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _52333_ (_01610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _52334_ (_01611_, _01610_, _01609_);
  not _52335_ (_01612_, _01611_);
  nor _52336_ (_01613_, _01612_, _01608_);
  and _52337_ (_01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _52338_ (_01615_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _52339_ (_01616_, _01615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _52340_ (_01617_, _01616_, _01613_);
  and _52341_ (_01618_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _52342_ (_01619_, _01618_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _52343_ (_01620_, _01619_, _01605_);
  and _52344_ (_01621_, _01620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _52345_ (_01622_, _01621_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _52346_ (_01623_, _01621_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _52347_ (_01624_, _01623_, _01622_);
  or _52348_ (_01625_, _01624_, _01460_);
  and _52349_ (_01627_, _01625_, _42618_);
  and _52350_ (_38751_, _01627_, _01604_);
  and _52351_ (_01629_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _42618_);
  and _52352_ (_01630_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _52353_ (_01632_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _52354_ (_01633_, _36958_, _01632_);
  not _52355_ (_01635_, _01633_);
  not _52356_ (_01636_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _52357_ (_01638_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _52358_ (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _52359_ (_01641_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _52360_ (_01642_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _52361_ (_01644_, _01642_, _01639_);
  and _52362_ (_01645_, _01644_, _01641_);
  nor _52363_ (_01647_, _01645_, _01639_);
  nor _52364_ (_01648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _52365_ (_01650_, _01648_, _01638_);
  not _52366_ (_01651_, _01650_);
  nor _52367_ (_01653_, _01651_, _01647_);
  nor _52368_ (_01654_, _01653_, _01638_);
  not _52369_ (_01656_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _52370_ (_01657_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _52371_ (_01658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _52372_ (_01659_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _52373_ (_01660_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _52374_ (_01661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _52375_ (_01662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _52376_ (_01663_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _52377_ (_01664_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _52378_ (_01665_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _52379_ (_01666_, _01665_, _01664_);
  and _52380_ (_01667_, _01666_, _01663_);
  and _52381_ (_01668_, _01667_, _01662_);
  and _52382_ (_01669_, _01668_, _01661_);
  and _52383_ (_01670_, _01669_, _01660_);
  and _52384_ (_01671_, _01670_, _01659_);
  and _52385_ (_01672_, _01671_, _01658_);
  and _52386_ (_01673_, _01672_, _01657_);
  and _52387_ (_01674_, _01673_, _01656_);
  and _52388_ (_01675_, _01674_, _01654_);
  and _52389_ (_01676_, _01675_, _01636_);
  nor _52390_ (_01677_, _01676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _52391_ (_01678_, _01676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _52392_ (_01679_, _01678_, _01677_);
  not _52393_ (_01680_, _01679_);
  nor _52394_ (_01681_, _01675_, _01636_);
  nor _52395_ (_01682_, _01681_, _01676_);
  not _52396_ (_01683_, _01682_);
  and _52397_ (_01684_, _01673_, _01654_);
  nor _52398_ (_01685_, _01684_, _01656_);
  or _52399_ (_01686_, _01685_, _01675_);
  and _52400_ (_01687_, _01672_, _01654_);
  nor _52401_ (_01688_, _01687_, _01657_);
  nor _52402_ (_01689_, _01688_, _01684_);
  not _52403_ (_01690_, _01689_);
  and _52404_ (_01691_, _01670_, _01654_);
  and _52405_ (_01692_, _01691_, _01659_);
  nor _52406_ (_01693_, _01692_, _01658_);
  nor _52407_ (_01694_, _01693_, _01687_);
  not _52408_ (_01695_, _01694_);
  nor _52409_ (_01696_, _01691_, _01659_);
  nor _52410_ (_01697_, _01696_, _01692_);
  not _52411_ (_01698_, _01697_);
  and _52412_ (_01699_, _01669_, _01654_);
  nor _52413_ (_01700_, _01699_, _01660_);
  nor _52414_ (_01701_, _01700_, _01691_);
  not _52415_ (_01702_, _01701_);
  and _52416_ (_01703_, _01667_, _01654_);
  nor _52417_ (_01704_, _01703_, _01662_);
  and _52418_ (_01705_, _01668_, _01654_);
  nor _52419_ (_01706_, _01705_, _01704_);
  not _52420_ (_01707_, _01706_);
  and _52421_ (_01708_, _01666_, _01654_);
  nor _52422_ (_01709_, _01708_, _01663_);
  nor _52423_ (_01710_, _01709_, _01703_);
  not _52424_ (_01711_, _01710_);
  and _52425_ (_01712_, _01665_, _01654_);
  nor _52426_ (_01713_, _01712_, _01664_);
  nor _52427_ (_01714_, _01713_, _01708_);
  not _52428_ (_01715_, _01714_);
  not _52429_ (_01716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _52430_ (_01717_, _01654_, _01716_);
  nor _52431_ (_01718_, _01654_, _01716_);
  nor _52432_ (_01719_, _01718_, _01717_);
  not _52433_ (_01720_, _01719_);
  not _52434_ (_01721_, _00730_);
  not _52435_ (_01722_, _00687_);
  and _52436_ (_01723_, _00675_, _00703_);
  not _52437_ (_01724_, _01723_);
  nor _52438_ (_01725_, _00683_, _00676_);
  and _52439_ (_01726_, _01725_, _01724_);
  and _52440_ (_01727_, _00718_, _00671_);
  and _52441_ (_01728_, _00671_, _00674_);
  or _52442_ (_01729_, _01728_, _01727_);
  nor _52443_ (_01730_, _00704_, _00701_);
  not _52444_ (_01731_, _01730_);
  nor _52445_ (_01732_, _01731_, _01729_);
  and _52446_ (_01733_, _01732_, _01726_);
  nor _52447_ (_01734_, _01733_, _01722_);
  nor _52448_ (_01735_, _01734_, _01721_);
  and _52449_ (_01736_, _00683_, _00669_);
  not _52450_ (_01737_, _01736_);
  nor _52451_ (_01738_, _00736_, _00679_);
  and _52452_ (_01739_, _01738_, _01737_);
  not _52453_ (_01740_, _01739_);
  or _52454_ (_01741_, _01728_, _00719_);
  nor _52455_ (_01742_, _01730_, _37602_);
  or _52456_ (_01743_, _01742_, _01741_);
  and _52457_ (_01744_, _01743_, _00668_);
  nor _52458_ (_01745_, _01744_, _01740_);
  and _52459_ (_01746_, _01745_, _01735_);
  nor _52460_ (_01747_, _00710_, _00698_);
  and _52461_ (_01748_, _00675_, _00718_);
  and _52462_ (_01749_, _01748_, _00678_);
  nor _52463_ (_01750_, _01749_, _00666_);
  and _52464_ (_01751_, _01750_, _01747_);
  and _52465_ (_01752_, _00683_, _00678_);
  and _52466_ (_01753_, _00674_, _00664_);
  and _52467_ (_01754_, _00695_, _01753_);
  nor _52468_ (_01755_, _01754_, _01752_);
  and _52469_ (_01756_, _00689_, _37908_);
  and _52470_ (_01757_, _01756_, _00687_);
  nor _52471_ (_01758_, _01757_, _00705_);
  and _52472_ (_01759_, _01758_, _01755_);
  and _52473_ (_01760_, _01759_, _01751_);
  not _52474_ (_01761_, _00678_);
  and _52475_ (_01762_, _00675_, _00682_);
  not _52476_ (_01763_, _01762_);
  nor _52477_ (_01764_, _01723_, _00725_);
  and _52478_ (_01765_, _01764_, _01763_);
  nor _52479_ (_01766_, _01765_, _01761_);
  not _52480_ (_01767_, _01766_);
  and _52481_ (_01768_, _00719_, _00694_);
  and _52482_ (_01769_, _00725_, _00695_);
  nor _52483_ (_01770_, _01769_, _01768_);
  and _52484_ (_01771_, _00704_, _00697_);
  and _52485_ (_01772_, _00689_, _00678_);
  nor _52486_ (_01773_, _01772_, _01771_);
  and _52487_ (_01774_, _01773_, _01770_);
  and _52488_ (_01775_, _01774_, _01767_);
  and _52489_ (_01776_, _01775_, _01760_);
  nor _52490_ (_01777_, _00672_, _00701_);
  and _52491_ (_01778_, _00707_, _37330_);
  not _52492_ (_01779_, _01778_);
  nor _52493_ (_01780_, _01779_, _01777_);
  not _52494_ (_01781_, _01780_);
  not _52495_ (_01782_, _01753_);
  nor _52496_ (_01783_, _00687_, _00668_);
  nor _52497_ (_01784_, _01783_, _01782_);
  and _52498_ (_01785_, _00671_, _00662_);
  and _52499_ (_01786_, _01785_, _37884_);
  nor _52500_ (_01787_, _01786_, _01784_);
  and _52501_ (_01788_, _01787_, _01781_);
  not _52502_ (_01789_, _00725_);
  nor _52503_ (_01790_, _00687_, _00669_);
  nor _52504_ (_01791_, _01790_, _01789_);
  not _52505_ (_01792_, _00669_);
  nor _52506_ (_01793_, _00908_, _00701_);
  nor _52507_ (_01794_, _01793_, _01792_);
  nor _52508_ (_01795_, _01794_, _01791_);
  nor _52509_ (_01796_, _01727_, _00701_);
  nor _52510_ (_01797_, _01796_, _37330_);
  and _52511_ (_01798_, _00675_, _37908_);
  nor _52512_ (_01799_, _01798_, _01727_);
  nor _52513_ (_01800_, _01799_, _00732_);
  nor _52514_ (_01801_, _01800_, _01797_);
  and _52515_ (_01802_, _01801_, _01795_);
  and _52516_ (_01803_, _01802_, _01788_);
  and _52517_ (_01804_, _01803_, _01776_);
  and _52518_ (_01805_, _01804_, _01746_);
  nor _52519_ (_01806_, _01644_, _01641_);
  nor _52520_ (_01807_, _01806_, _01645_);
  not _52521_ (_01808_, _01807_);
  nor _52522_ (_01809_, _01808_, _01805_);
  and _52523_ (_01810_, _01755_, _01739_);
  nor _52524_ (_01811_, _01730_, _01761_);
  not _52525_ (_01812_, _01811_);
  nor _52526_ (_01813_, _01757_, _00710_);
  and _52527_ (_01814_, _01813_, _01812_);
  nor _52528_ (_01815_, _01769_, _00728_);
  and _52529_ (_01816_, _01728_, _00662_);
  and _52530_ (_01817_, _00719_, _00695_);
  nor _52531_ (_01818_, _01817_, _01816_);
  and _52532_ (_01819_, _01818_, _01815_);
  and _52533_ (_01820_, _01819_, _01814_);
  and _52534_ (_01821_, _01820_, _01810_);
  not _52535_ (_01822_, _01821_);
  nor _52536_ (_01823_, _01822_, _01805_);
  not _52537_ (_01824_, _01823_);
  nor _52538_ (_01825_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _52539_ (_01826_, _01825_, _01641_);
  and _52540_ (_01827_, _01826_, _01824_);
  and _52541_ (_01828_, _01808_, _01805_);
  nor _52542_ (_01829_, _01828_, _01809_);
  and _52543_ (_01830_, _01829_, _01827_);
  nor _52544_ (_01831_, _01830_, _01809_);
  not _52545_ (_01832_, _01831_);
  and _52546_ (_01833_, _01651_, _01647_);
  nor _52547_ (_01834_, _01833_, _01653_);
  and _52548_ (_01835_, _01834_, _01832_);
  and _52549_ (_01836_, _01835_, _01720_);
  not _52550_ (_01837_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _52551_ (_01838_, _01717_, _01837_);
  or _52552_ (_01839_, _01838_, _01712_);
  and _52553_ (_01840_, _01839_, _01836_);
  and _52554_ (_01841_, _01840_, _01715_);
  and _52555_ (_01842_, _01841_, _01711_);
  and _52556_ (_01843_, _01842_, _01707_);
  nor _52557_ (_01844_, _01705_, _01661_);
  or _52558_ (_01845_, _01844_, _01699_);
  and _52559_ (_01846_, _01845_, _01843_);
  and _52560_ (_01847_, _01846_, _01702_);
  and _52561_ (_01848_, _01847_, _01698_);
  and _52562_ (_01849_, _01848_, _01695_);
  and _52563_ (_01850_, _01849_, _01690_);
  and _52564_ (_01851_, _01850_, _01686_);
  nand _52565_ (_01852_, _01851_, _01683_);
  nand _52566_ (_01853_, _01852_, _01680_);
  or _52567_ (_01854_, _01852_, _01680_);
  and _52568_ (_01855_, _01854_, _01853_);
  or _52569_ (_01856_, _01855_, _01635_);
  or _52570_ (_01857_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _52571_ (_01858_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _52572_ (_01859_, _01858_, _01857_);
  and _52573_ (_01860_, _01859_, _01856_);
  or _52574_ (_38753_, _01860_, _01630_);
  nor _52575_ (_01861_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _52576_ (_38754_, _01861_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _52577_ (_38755_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _42618_);
  nor _52578_ (_01862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _52579_ (_01863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _52580_ (_01864_, _01863_, _01862_);
  nor _52581_ (_01865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _52582_ (_01866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _52583_ (_01867_, _01866_, _01865_);
  and _52584_ (_01868_, _01867_, _01864_);
  nor _52585_ (_01869_, _01868_, rst);
  and _52586_ (_01870_, \oc8051_top_1.oc8051_rom1.ea_int , _36925_);
  nand _52587_ (_01871_, _01870_, _36958_);
  and _52588_ (_01872_, _01871_, _38755_);
  or _52589_ (_38756_, _01872_, _01869_);
  and _52590_ (_01873_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _52591_ (_01874_, _01873_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _52592_ (_38758_, _01874_, _42618_);
  nor _52593_ (_01875_, _01608_, _42079_);
  nor _52594_ (_01876_, _01805_, _37155_);
  nor _52595_ (_01877_, _01823_, _37111_);
  and _52596_ (_01878_, _01805_, _37155_);
  nor _52597_ (_01879_, _01878_, _01876_);
  and _52598_ (_01880_, _01879_, _01877_);
  nor _52599_ (_01881_, _01880_, _01876_);
  nor _52600_ (_01882_, _01881_, _42079_);
  and _52601_ (_01883_, _01882_, _37023_);
  nor _52602_ (_01884_, _01882_, _37023_);
  nor _52603_ (_01885_, _01884_, _01883_);
  nor _52604_ (_01886_, _01885_, _01875_);
  and _52605_ (_01887_, _37166_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _52606_ (_01888_, _01887_, _01875_);
  nor _52607_ (_01889_, _01888_, _01821_);
  or _52608_ (_01890_, _01889_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _52609_ (_01891_, _01890_, _01886_);
  and _52610_ (_38759_, _01891_, _42618_);
  or _52611_ (_01892_, _37559_, _37927_);
  nor _52612_ (_01893_, _01892_, _37286_);
  not _52613_ (_01894_, _37852_);
  and _52614_ (_01895_, _01894_, _37950_);
  and _52615_ (_01896_, _01895_, _37820_);
  not _52616_ (_01897_, _01353_);
  nor _52617_ (_01898_, _01897_, _37878_);
  and _52618_ (_01899_, _01898_, _37904_);
  and _52619_ (_01900_, _01899_, _01896_);
  and _52620_ (_38762_, _01900_, _01893_);
  nor _52621_ (_01901_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _52622_ (_01902_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _52623_ (_01903_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _52624_ (_38765_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _42618_);
  and _52625_ (_01904_, _38765_, _01903_);
  or _52626_ (_38763_, _01904_, _01902_);
  not _52627_ (_01905_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _52628_ (_01906_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _52629_ (_01907_, _01906_, _01905_);
  and _52630_ (_01908_, _01906_, _01905_);
  nor _52631_ (_01909_, _01908_, _01907_);
  not _52632_ (_01910_, _01909_);
  and _52633_ (_01911_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _52634_ (_01912_, _01911_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _52635_ (_01913_, _01911_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _52636_ (_01914_, _01913_, _01912_);
  or _52637_ (_01915_, _01914_, _01906_);
  and _52638_ (_01916_, _01915_, _01910_);
  nor _52639_ (_01917_, _01907_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _52640_ (_01918_, _01907_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _52641_ (_01919_, _01918_, _01917_);
  or _52642_ (_01920_, _01912_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _52643_ (_38767_, _01920_, _42618_);
  and _52644_ (_01921_, _38767_, _01919_);
  and _52645_ (_38766_, _01921_, _01916_);
  not _52646_ (_01922_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _52647_ (_01923_, _01608_, _01922_);
  and _52648_ (_01924_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _52649_ (_01925_, _01923_);
  and _52650_ (_01926_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _52651_ (_01927_, _01926_, _01924_);
  and _52652_ (_38768_, _01927_, _42618_);
  and _52653_ (_01928_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _52654_ (_01929_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _52655_ (_01930_, _01929_, _01928_);
  and _52656_ (_38769_, _01930_, _42618_);
  and _52657_ (_01931_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _52658_ (_01932_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52659_ (_01933_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _01932_);
  and _52660_ (_01934_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _52661_ (_01935_, _01934_, _01931_);
  and _52662_ (_38770_, _01935_, _42618_);
  and _52663_ (_01936_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52664_ (_01937_, _01936_, _01933_);
  and _52665_ (_38771_, _01937_, _42618_);
  or _52666_ (_01938_, _01932_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _52667_ (_38773_, _01938_, _42618_);
  not _52668_ (_01939_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _52669_ (_01940_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _52670_ (_01941_, _01940_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52671_ (_01942_, _01932_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _52672_ (_01943_, _01942_, _42618_);
  and _52673_ (_38774_, _01943_, _01941_);
  or _52674_ (_01944_, _01932_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _52675_ (_38775_, _01944_, _42618_);
  nor _52676_ (_01945_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _52677_ (_01946_, _01945_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52678_ (_01947_, _01946_, _42618_);
  and _52679_ (_01948_, _38765_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _52680_ (_38776_, _01948_, _01947_);
  and _52681_ (_01949_, _01922_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _52682_ (_01950_, _01949_, _01946_);
  and _52683_ (_38777_, _01950_, _42618_);
  nand _52684_ (_01951_, _01946_, _38368_);
  or _52685_ (_01952_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _52686_ (_01953_, _01952_, _42618_);
  and _52687_ (_38778_, _01953_, _01951_);
  nand _52688_ (_01954_, _37999_, _42618_);
  nor _52689_ (_38779_, _01954_, _38133_);
  or _52690_ (_01955_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _52691_ (_01956_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand _52692_ (_01957_, _01347_, _01956_);
  and _52693_ (_01958_, _01957_, _42618_);
  and _52694_ (_38816_, _01958_, _01955_);
  or _52695_ (_01959_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _52696_ (_01960_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _52697_ (_01961_, _01347_, _01960_);
  and _52698_ (_01962_, _01961_, _42618_);
  and _52699_ (_38817_, _01962_, _01959_);
  or _52700_ (_01963_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _52701_ (_01964_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _52702_ (_01965_, _01347_, _01964_);
  and _52703_ (_01966_, _01965_, _42618_);
  and _52704_ (_38818_, _01966_, _01963_);
  or _52705_ (_01967_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _52706_ (_01968_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _52707_ (_01969_, _01347_, _01968_);
  and _52708_ (_01970_, _01969_, _42618_);
  and _52709_ (_38819_, _01970_, _01967_);
  or _52710_ (_01971_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _52711_ (_01972_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52712_ (_01973_, _01972_, _42618_);
  and _52713_ (_38820_, _01973_, _01971_);
  or _52714_ (_01974_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not _52715_ (_01975_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand _52716_ (_01976_, _01347_, _01975_);
  and _52717_ (_01977_, _01976_, _42618_);
  and _52718_ (_38822_, _01977_, _01974_);
  or _52719_ (_01978_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not _52720_ (_01979_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand _52721_ (_01980_, _01347_, _01979_);
  and _52722_ (_01981_, _01980_, _42618_);
  and _52723_ (_38823_, _01981_, _01978_);
  or _52724_ (_01982_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _52725_ (_01983_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand _52726_ (_01984_, _01347_, _01983_);
  and _52727_ (_01985_, _01984_, _42618_);
  and _52728_ (_38824_, _01985_, _01982_);
  or _52729_ (_01986_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _52730_ (_01987_, _01347_, _38285_);
  and _52731_ (_01988_, _01987_, _42618_);
  and _52732_ (_38825_, _01988_, _01986_);
  or _52733_ (_01989_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _52734_ (_01990_, _01347_, _38291_);
  and _52735_ (_01991_, _01990_, _42618_);
  and _52736_ (_38826_, _01991_, _01989_);
  or _52737_ (_01992_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _52738_ (_01993_, _01347_, _38296_);
  and _52739_ (_01994_, _01993_, _42618_);
  and _52740_ (_38827_, _01994_, _01992_);
  or _52741_ (_01995_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _52742_ (_01996_, _01347_, _38281_);
  and _52743_ (_01997_, _01996_, _42618_);
  and _52744_ (_38828_, _01997_, _01995_);
  or _52745_ (_01998_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _52746_ (_01999_, _01347_, _38302_);
  and _52747_ (_02000_, _01999_, _42618_);
  and _52748_ (_38829_, _02000_, _01998_);
  or _52749_ (_02001_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _52750_ (_02002_, _01347_, _38307_);
  and _52751_ (_02003_, _02002_, _42618_);
  and _52752_ (_38830_, _02003_, _02001_);
  or _52753_ (_02004_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _52754_ (_02005_, _01347_, _38312_);
  and _52755_ (_02006_, _02005_, _42618_);
  and _52756_ (_38831_, _02006_, _02004_);
  and _52757_ (_02007_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _52758_ (_02008_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _52759_ (_02009_, _02008_, _02007_);
  and _52760_ (_38836_, _02009_, _42618_);
  and _52761_ (_02010_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _52762_ (_02011_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _52763_ (_02012_, _02011_, _02010_);
  and _52764_ (_38837_, _02012_, _42618_);
  and _52765_ (_02013_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _52766_ (_02014_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _52767_ (_02015_, _02014_, _02013_);
  and _52768_ (_38838_, _02015_, _42618_);
  and _52769_ (_02016_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _52770_ (_02017_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _52771_ (_02018_, _02017_, _02016_);
  and _52772_ (_38839_, _02018_, _42618_);
  and _52773_ (_02019_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _52774_ (_02020_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or _52775_ (_02021_, _02020_, _02019_);
  and _52776_ (_38840_, _02021_, _42618_);
  and _52777_ (_02022_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _52778_ (_02023_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or _52779_ (_02024_, _02023_, _02022_);
  and _52780_ (_38841_, _02024_, _42618_);
  and _52781_ (_02025_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _52782_ (_02026_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or _52783_ (_02027_, _02026_, _02025_);
  and _52784_ (_38842_, _02027_, _42618_);
  and _52785_ (_02028_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _52786_ (_02029_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or _52787_ (_02030_, _02029_, _02028_);
  and _52788_ (_38843_, _02030_, _42618_);
  and _52789_ (_02031_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _52790_ (_02032_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or _52791_ (_02033_, _02032_, _02031_);
  and _52792_ (_38844_, _02033_, _42618_);
  and _52793_ (_02034_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _52794_ (_02035_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or _52795_ (_02036_, _02035_, _02034_);
  and _52796_ (_38845_, _02036_, _42618_);
  and _52797_ (_02037_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _52798_ (_02038_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or _52799_ (_02039_, _02038_, _02037_);
  and _52800_ (_38847_, _02039_, _42618_);
  and _52801_ (_02040_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _52802_ (_02041_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or _52803_ (_02042_, _02041_, _02040_);
  and _52804_ (_38848_, _02042_, _42618_);
  and _52805_ (_02043_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _52806_ (_02044_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or _52807_ (_02045_, _02044_, _02043_);
  and _52808_ (_38849_, _02045_, _42618_);
  and _52809_ (_02046_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _52810_ (_02047_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or _52811_ (_02048_, _02047_, _02046_);
  and _52812_ (_38850_, _02048_, _42618_);
  and _52813_ (_02049_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _52814_ (_02050_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or _52815_ (_02051_, _02050_, _02049_);
  and _52816_ (_38851_, _02051_, _42618_);
  and _52817_ (_39027_, _37657_, _42618_);
  and _52818_ (_39028_, _37863_, _42618_);
  and _52819_ (_39029_, _37837_, _42618_);
  nor _52820_ (_39030_, _42022_, rst);
  and _52821_ (_02052_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _52822_ (_02053_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or _52823_ (_02054_, _02053_, _02052_);
  and _52824_ (_39031_, _02054_, _42618_);
  and _52825_ (_02055_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _52826_ (_02056_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _52827_ (_02057_, _02056_, _01923_);
  or _52828_ (_02058_, _02057_, _02055_);
  and _52829_ (_39032_, _02058_, _42618_);
  and _52830_ (_02059_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _52831_ (_02060_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _52832_ (_02061_, _02060_, _02059_);
  and _52833_ (_39033_, _02061_, _42618_);
  and _52834_ (_02062_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _52835_ (_02063_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or _52836_ (_02064_, _02063_, _02062_);
  and _52837_ (_39034_, _02064_, _42618_);
  and _52838_ (_02065_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _52839_ (_02066_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _52840_ (_02067_, _02066_, _02065_);
  and _52841_ (_39036_, _02067_, _42618_);
  and _52842_ (_02068_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _52843_ (_02069_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _52844_ (_02070_, _02069_, _01923_);
  or _52845_ (_02071_, _02070_, _02068_);
  and _52846_ (_39037_, _02071_, _42618_);
  and _52847_ (_02072_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _52848_ (_02073_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or _52849_ (_02074_, _02073_, _02072_);
  and _52850_ (_39038_, _02074_, _42618_);
  and _52851_ (_02075_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _52852_ (_02076_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or _52853_ (_02077_, _02076_, _02075_);
  and _52854_ (_39039_, _02077_, _42618_);
  and _52855_ (_02078_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and _52856_ (_02079_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _52857_ (_02080_, _02079_, _02078_);
  and _52858_ (_39040_, _02080_, _42618_);
  and _52859_ (_02081_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and _52860_ (_02082_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _52861_ (_02083_, _02082_, _02081_);
  and _52862_ (_39041_, _02083_, _42618_);
  and _52863_ (_02084_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and _52864_ (_02085_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _52865_ (_02086_, _02085_, _02084_);
  and _52866_ (_39042_, _02086_, _42618_);
  and _52867_ (_02087_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and _52868_ (_02088_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _52869_ (_02089_, _02088_, _02087_);
  and _52870_ (_39043_, _02089_, _42618_);
  and _52871_ (_02090_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and _52872_ (_02091_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _52873_ (_02092_, _02091_, _02090_);
  and _52874_ (_39044_, _02092_, _42618_);
  and _52875_ (_02093_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and _52876_ (_02094_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _52877_ (_02095_, _02094_, _02093_);
  and _52878_ (_39045_, _02095_, _42618_);
  and _52879_ (_02096_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and _52880_ (_02097_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _52881_ (_02098_, _02097_, _02096_);
  and _52882_ (_39047_, _02098_, _42618_);
  and _52883_ (_02099_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and _52884_ (_02100_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _52885_ (_02101_, _02100_, _02099_);
  and _52886_ (_39048_, _02101_, _42618_);
  and _52887_ (_02102_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _52888_ (_02103_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _52889_ (_02104_, _02103_, _02102_);
  and _52890_ (_39049_, _02104_, _42618_);
  and _52891_ (_02105_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _52892_ (_02106_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _52893_ (_02107_, _02106_, _02105_);
  and _52894_ (_39050_, _02107_, _42618_);
  and _52895_ (_02108_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _52896_ (_02109_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _52897_ (_02110_, _02109_, _02108_);
  and _52898_ (_39051_, _02110_, _42618_);
  and _52899_ (_02112_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _52900_ (_02114_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _52901_ (_02116_, _02114_, _02112_);
  and _52902_ (_39052_, _02116_, _42618_);
  and _52903_ (_02119_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _52904_ (_02121_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _52905_ (_02123_, _02121_, _02119_);
  and _52906_ (_39053_, _02123_, _42618_);
  and _52907_ (_02126_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _52908_ (_02128_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _52909_ (_02130_, _02128_, _02126_);
  and _52910_ (_39054_, _02130_, _42618_);
  and _52911_ (_02133_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _52912_ (_02135_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _52913_ (_02137_, _02135_, _02133_);
  and _52914_ (_39055_, _02137_, _42618_);
  and _52915_ (_02140_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _52916_ (_02142_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _52917_ (_02144_, _02142_, _02140_);
  and _52918_ (_39056_, _02144_, _42618_);
  and _52919_ (_02147_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _52920_ (_02149_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _52921_ (_02151_, _02149_, _02147_);
  and _52922_ (_39058_, _02151_, _42618_);
  and _52923_ (_02154_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _52924_ (_02156_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _52925_ (_02158_, _02156_, _02154_);
  and _52926_ (_39059_, _02158_, _42618_);
  and _52927_ (_02161_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _52928_ (_02163_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _52929_ (_02165_, _02163_, _02161_);
  and _52930_ (_39060_, _02165_, _42618_);
  and _52931_ (_02168_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _52932_ (_02170_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _52933_ (_02172_, _02170_, _02168_);
  and _52934_ (_39061_, _02172_, _42618_);
  and _52935_ (_02173_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _52936_ (_02174_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _52937_ (_02175_, _02174_, _02173_);
  and _52938_ (_39062_, _02175_, _42618_);
  and _52939_ (_02176_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _52940_ (_02177_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _52941_ (_02178_, _02177_, _02176_);
  and _52942_ (_39063_, _02178_, _42618_);
  and _52943_ (_02179_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _52944_ (_02180_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _52945_ (_02181_, _02180_, _02179_);
  and _52946_ (_39064_, _02181_, _42618_);
  nor _52947_ (_39065_, _42374_, rst);
  nor _52948_ (_39067_, _42280_, rst);
  nor _52949_ (_39068_, _42184_, rst);
  nor _52950_ (_39069_, _42327_, rst);
  nor _52951_ (_39070_, _42233_, rst);
  nor _52952_ (_39071_, _42160_, rst);
  nor _52953_ (_39073_, _42428_, rst);
  and _52954_ (_39089_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _42618_);
  and _52955_ (_39090_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _42618_);
  and _52956_ (_39091_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _42618_);
  and _52957_ (_39092_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _42618_);
  and _52958_ (_39093_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _42618_);
  and _52959_ (_39095_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _42618_);
  and _52960_ (_39096_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _42618_);
  or _52961_ (_02182_, _01484_, _01464_);
  and _52962_ (_02183_, _02182_, _32334_);
  and _52963_ (_02184_, _01587_, _42392_);
  and _52964_ (_02185_, _01469_, _01531_);
  and _52965_ (_02186_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _52966_ (_02187_, _02186_, _02185_);
  or _52967_ (_02188_, _02187_, _02184_);
  nor _52968_ (_02189_, _01533_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _52969_ (_02190_, _02189_, _01534_);
  and _52970_ (_02191_, _02190_, _01583_);
  nor _52971_ (_02192_, _02191_, _02188_);
  nand _52972_ (_02193_, _02192_, _01460_);
  or _52973_ (_02194_, _02193_, _02183_);
  or _52974_ (_02195_, _01460_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _52975_ (_02196_, _02195_, _42618_);
  and _52976_ (_39097_, _02196_, _02194_);
  and _52977_ (_02197_, _02182_, _33031_);
  and _52978_ (_02198_, _01587_, _42299_);
  and _52979_ (_02199_, _01469_, _01526_);
  and _52980_ (_02200_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _52981_ (_02201_, _02200_, _02199_);
  or _52982_ (_02202_, _02201_, _02198_);
  or _52983_ (_02203_, _02202_, _02197_);
  nor _52984_ (_02204_, _01536_, _01534_);
  nor _52985_ (_02205_, _02204_, _01537_);
  nand _52986_ (_02206_, _02205_, _01583_);
  nand _52987_ (_02207_, _02206_, _01460_);
  or _52988_ (_02208_, _02207_, _02203_);
  or _52989_ (_02209_, _01460_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _52990_ (_02210_, _02209_, _42618_);
  and _52991_ (_39098_, _02210_, _02208_);
  and _52992_ (_02211_, _02182_, _33728_);
  and _52993_ (_02212_, _01587_, _42208_);
  and _52994_ (_02213_, _01469_, _01521_);
  or _52995_ (_02214_, _02213_, _02212_);
  or _52996_ (_02215_, _01541_, _01539_);
  not _52997_ (_02216_, _01542_);
  and _52998_ (_02217_, _01583_, _02216_);
  and _52999_ (_02218_, _02217_, _02215_);
  or _53000_ (_02219_, _02218_, _02214_);
  or _53001_ (_02220_, _02219_, _02211_);
  nand _53002_ (_02221_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nand _53003_ (_02222_, _02221_, _01460_);
  or _53004_ (_02223_, _02222_, _02220_);
  not _53005_ (_02224_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _53006_ (_02225_, _01608_, _02224_);
  and _53007_ (_02226_, _01608_, _02224_);
  nor _53008_ (_02227_, _02226_, _02225_);
  or _53009_ (_02228_, _02227_, _01460_);
  and _53010_ (_02229_, _02228_, _42618_);
  and _53011_ (_39099_, _02229_, _02223_);
  and _53012_ (_02230_, _02182_, _34489_);
  and _53013_ (_02231_, _01587_, _42350_);
  and _53014_ (_02232_, _01469_, _01515_);
  or _53015_ (_02233_, _02232_, _02231_);
  or _53016_ (_02234_, _01519_, _01518_);
  or _53017_ (_02235_, _02234_, _01543_);
  nand _53018_ (_02236_, _02234_, _01543_);
  and _53019_ (_02237_, _02236_, _01583_);
  and _53020_ (_02238_, _02237_, _02235_);
  or _53021_ (_02239_, _02238_, _02233_);
  or _53022_ (_02240_, _02239_, _02230_);
  nand _53023_ (_02241_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand _53024_ (_02242_, _02241_, _01460_);
  or _53025_ (_02243_, _02242_, _02240_);
  and _53026_ (_02244_, _02225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53027_ (_02245_, _02225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53028_ (_02246_, _02245_, _02244_);
  or _53029_ (_02247_, _02246_, _01460_);
  and _53030_ (_02248_, _02247_, _42618_);
  and _53031_ (_39100_, _02248_, _02243_);
  and _53032_ (_02249_, _02182_, _35251_);
  and _53033_ (_02250_, _01469_, _01510_);
  and _53034_ (_02251_, _01587_, _42254_);
  or _53035_ (_02252_, _02251_, _02250_);
  or _53036_ (_02253_, _01547_, _01545_);
  and _53037_ (_02254_, _01583_, _01548_);
  and _53038_ (_02255_, _02254_, _02253_);
  or _53039_ (_02256_, _02255_, _02252_);
  or _53040_ (_02257_, _02256_, _02249_);
  nand _53041_ (_02258_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nand _53042_ (_02259_, _02258_, _01460_);
  or _53043_ (_02260_, _02259_, _02257_);
  and _53044_ (_02261_, _02244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53045_ (_02262_, _02244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53046_ (_02263_, _02262_, _02261_);
  or _53047_ (_02264_, _02263_, _01460_);
  and _53048_ (_02265_, _02264_, _42618_);
  and _53049_ (_39101_, _02265_, _02260_);
  and _53050_ (_02266_, _02182_, _36057_);
  and _53051_ (_02267_, _01587_, _42132_);
  and _53052_ (_02268_, _01469_, _01504_);
  and _53053_ (_02269_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _53054_ (_02270_, _02269_, _02268_);
  or _53055_ (_02271_, _02270_, _02267_);
  or _53056_ (_02272_, _02271_, _02266_);
  or _53057_ (_02273_, _01508_, _01507_);
  or _53058_ (_02274_, _02273_, _01549_);
  nand _53059_ (_02275_, _02273_, _01549_);
  and _53060_ (_02276_, _02275_, _02274_);
  nand _53061_ (_02277_, _02276_, _01583_);
  nand _53062_ (_02278_, _02277_, _01460_);
  or _53063_ (_02279_, _02278_, _02272_);
  nor _53064_ (_02280_, _02261_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _53065_ (_02281_, _02280_, _01613_);
  or _53066_ (_02282_, _02281_, _01460_);
  and _53067_ (_02283_, _02282_, _42618_);
  and _53068_ (_39102_, _02283_, _02279_);
  nor _53069_ (_02284_, _01613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _53070_ (_02285_, _01613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _53071_ (_02286_, _02285_, _02284_);
  or _53072_ (_02287_, _02286_, _01460_);
  and _53073_ (_02288_, _02287_, _42618_);
  not _53074_ (_02289_, _01460_);
  and _53075_ (_02290_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _53076_ (_02291_, _02182_, _36698_);
  and _53077_ (_02292_, _01469_, _01497_);
  and _53078_ (_02293_, _01587_, _42447_);
  or _53079_ (_02294_, _02293_, _02292_);
  or _53080_ (_02295_, _01551_, _01502_);
  and _53081_ (_02296_, _01583_, _01552_);
  and _53082_ (_02297_, _02296_, _02295_);
  or _53083_ (_02298_, _02297_, _02294_);
  or _53084_ (_02299_, _02298_, _02291_);
  or _53085_ (_02300_, _02299_, _02290_);
  or _53086_ (_02301_, _02300_, _02289_);
  and _53087_ (_39103_, _02301_, _02288_);
  or _53088_ (_02302_, _01494_, _01495_);
  or _53089_ (_02303_, _02302_, _01553_);
  nand _53090_ (_02304_, _02302_, _01553_);
  and _53091_ (_02305_, _02304_, _02303_);
  and _53092_ (_02306_, _02305_, _01583_);
  and _53093_ (_02307_, _02182_, _31147_);
  and _53094_ (_02308_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _53095_ (_02309_, _01469_, _01491_);
  and _53096_ (_02310_, _01587_, _42096_);
  or _53097_ (_02311_, _02310_, _02309_);
  or _53098_ (_02312_, _02311_, _02308_);
  or _53099_ (_02313_, _02312_, _02307_);
  or _53100_ (_02314_, _02313_, _02306_);
  or _53101_ (_02315_, _02314_, _02289_);
  nor _53102_ (_02316_, _02285_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _53103_ (_02317_, _02285_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _53104_ (_02318_, _02317_, _02316_);
  or _53105_ (_02319_, _02318_, _01460_);
  and _53106_ (_02320_, _02319_, _42618_);
  and _53107_ (_39104_, _02320_, _02315_);
  and _53108_ (_02321_, _38094_, _32334_);
  and _53109_ (_02322_, _01555_, _38285_);
  nor _53110_ (_02323_, _01555_, _38285_);
  nor _53111_ (_02324_, _02323_, _02322_);
  nor _53112_ (_02325_, _02324_, _01493_);
  and _53113_ (_02326_, _02324_, _01493_);
  or _53114_ (_02327_, _02326_, _02325_);
  and _53115_ (_02328_, _02327_, _01583_);
  not _53116_ (_02329_, _38405_);
  and _53117_ (_02330_, _01464_, _02329_);
  and _53118_ (_02331_, _01587_, _00711_);
  and _53119_ (_02332_, _01469_, _42392_);
  or _53120_ (_02333_, _02332_, _02331_);
  and _53121_ (_02334_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _53122_ (_02335_, _02334_, _02333_);
  or _53123_ (_02336_, _02335_, _02330_);
  or _53124_ (_02337_, _02336_, _02328_);
  or _53125_ (_02338_, _02337_, _02321_);
  or _53126_ (_02339_, _02338_, _02289_);
  or _53127_ (_02340_, _02317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand _53128_ (_02341_, _01615_, _01613_);
  and _53129_ (_02342_, _02341_, _02340_);
  or _53130_ (_02343_, _02342_, _01460_);
  and _53131_ (_02344_, _02343_, _42618_);
  and _53132_ (_39106_, _02344_, _02339_);
  and _53133_ (_02345_, _38094_, _33031_);
  not _53134_ (_02346_, _38436_);
  and _53135_ (_02347_, _01464_, _02346_);
  and _53136_ (_02348_, _01587_, _00663_);
  and _53137_ (_02349_, _01469_, _42299_);
  or _53138_ (_02350_, _02349_, _02348_);
  and _53139_ (_02351_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _53140_ (_02352_, _02351_, _02350_);
  or _53141_ (_02353_, _02352_, _02347_);
  and _53142_ (_02355_, _01555_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _53143_ (_02356_, _02355_, _01563_);
  and _53144_ (_02357_, _01564_, _01493_);
  nor _53145_ (_02358_, _02357_, _02356_);
  nand _53146_ (_02359_, _02358_, _38291_);
  or _53147_ (_02360_, _02358_, _38291_);
  and _53148_ (_02361_, _02360_, _02359_);
  and _53149_ (_02362_, _02361_, _01583_);
  or _53150_ (_02363_, _02362_, _02353_);
  or _53151_ (_02364_, _02363_, _02289_);
  or _53152_ (_02365_, _02364_, _02345_);
  nand _53153_ (_02366_, _02341_, _01660_);
  or _53154_ (_02367_, _02341_, _01660_);
  and _53155_ (_02368_, _02367_, _02366_);
  or _53156_ (_02369_, _02368_, _01460_);
  and _53157_ (_02370_, _02369_, _42618_);
  and _53158_ (_39107_, _02370_, _02365_);
  and _53159_ (_02371_, _38094_, _33728_);
  not _53160_ (_02372_, _38466_);
  and _53161_ (_02373_, _01464_, _02372_);
  and _53162_ (_02374_, _01469_, _42208_);
  not _53163_ (_02375_, _37931_);
  and _53164_ (_02376_, _01587_, _02375_);
  and _53165_ (_02377_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _53166_ (_02378_, _02377_, _02376_);
  or _53167_ (_02379_, _02378_, _02374_);
  or _53168_ (_02380_, _02379_, _02373_);
  and _53169_ (_02381_, _01565_, _01493_);
  and _53170_ (_02382_, _02356_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _53171_ (_02383_, _02382_, _02381_);
  nand _53172_ (_02384_, _02383_, _38296_);
  or _53173_ (_02385_, _02383_, _38296_);
  and _53174_ (_02386_, _02385_, _02384_);
  and _53175_ (_02387_, _02386_, _01583_);
  or _53176_ (_02388_, _02387_, _02380_);
  or _53177_ (_02389_, _02388_, _02371_);
  or _53178_ (_02390_, _02389_, _02289_);
  nor _53179_ (_02391_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _53180_ (_02392_, _02391_, _01618_);
  or _53181_ (_02393_, _02392_, _01460_);
  and _53182_ (_02394_, _02393_, _42618_);
  and _53183_ (_39108_, _02394_, _02390_);
  and _53184_ (_02395_, _01558_, _01563_);
  and _53185_ (_02396_, _01566_, _01493_);
  nor _53186_ (_02397_, _02396_, _02395_);
  nand _53187_ (_02398_, _02397_, _38281_);
  or _53188_ (_02399_, _02397_, _38281_);
  and _53189_ (_02400_, _02399_, _02398_);
  and _53190_ (_02401_, _02400_, _01583_);
  and _53191_ (_02402_, _38094_, _34489_);
  not _53192_ (_02403_, _38497_);
  and _53193_ (_02404_, _01464_, _02403_);
  and _53194_ (_02405_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _53195_ (_02406_, _01594_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _53196_ (_02407_, _02406_, _01595_);
  and _53197_ (_02408_, _02407_, _01587_);
  and _53198_ (_02409_, _01469_, _42350_);
  or _53199_ (_02410_, _02409_, _02408_);
  or _53200_ (_02411_, _02410_, _02405_);
  or _53201_ (_02412_, _02411_, _02404_);
  or _53202_ (_02413_, _02412_, _02402_);
  or _53203_ (_02414_, _02413_, _02401_);
  or _53204_ (_02415_, _02414_, _02289_);
  nor _53205_ (_02416_, _01618_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _53206_ (_02417_, _02416_, _01619_);
  or _53207_ (_02418_, _02417_, _01460_);
  and _53208_ (_02419_, _02418_, _42618_);
  and _53209_ (_39109_, _02419_, _02415_);
  nor _53210_ (_02420_, _01595_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _53211_ (_02421_, _02420_, _01596_);
  and _53212_ (_02422_, _02421_, _01587_);
  and _53213_ (_02423_, _01559_, _01563_);
  and _53214_ (_02424_, _01567_, _01493_);
  nor _53215_ (_02425_, _02424_, _02423_);
  or _53216_ (_02426_, _02425_, _38302_);
  nand _53217_ (_02427_, _02425_, _38302_);
  and _53218_ (_02428_, _02427_, _01583_);
  and _53219_ (_02429_, _02428_, _02426_);
  and _53220_ (_02430_, _38094_, _35251_);
  not _53221_ (_02431_, _38528_);
  and _53222_ (_02432_, _01464_, _02431_);
  and _53223_ (_02433_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _53224_ (_02434_, _01469_, _42254_);
  or _53225_ (_02435_, _02434_, _02433_);
  or _53226_ (_02436_, _02435_, _02432_);
  or _53227_ (_02437_, _02436_, _02430_);
  or _53228_ (_02438_, _02437_, _02429_);
  or _53229_ (_02439_, _02438_, _02422_);
  or _53230_ (_02440_, _02439_, _02289_);
  nor _53231_ (_02441_, _01619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _53232_ (_02442_, _01619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _53233_ (_02443_, _02442_, _02441_);
  or _53234_ (_02444_, _02443_, _01460_);
  and _53235_ (_02445_, _02444_, _42618_);
  and _53236_ (_39110_, _02445_, _02440_);
  nor _53237_ (_02446_, _01596_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _53238_ (_02447_, _02446_, _01597_);
  and _53239_ (_02448_, _02447_, _01587_);
  and _53240_ (_02449_, _38094_, _36057_);
  not _53241_ (_02450_, _38561_);
  and _53242_ (_02451_, _01464_, _02450_);
  and _53243_ (_02452_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _53244_ (_02453_, _01469_, _42132_);
  or _53245_ (_02454_, _02453_, _02452_);
  or _53246_ (_02455_, _02454_, _02451_);
  or _53247_ (_02456_, _02455_, _02449_);
  or _53248_ (_02457_, _02456_, _02448_);
  and _53249_ (_02458_, _02423_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _53250_ (_02459_, _02424_, _38302_);
  nor _53251_ (_02460_, _02459_, _02458_);
  or _53252_ (_02461_, _02460_, _38307_);
  nand _53253_ (_02462_, _02460_, _38307_);
  and _53254_ (_02463_, _02462_, _01583_);
  and _53255_ (_02464_, _02463_, _02461_);
  or _53256_ (_02465_, _02464_, _02289_);
  or _53257_ (_02466_, _02465_, _02457_);
  or _53258_ (_02467_, _02442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand _53259_ (_02468_, _02442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _53260_ (_02469_, _02468_, _02467_);
  or _53261_ (_02470_, _02469_, _01460_);
  and _53262_ (_02471_, _02470_, _42618_);
  and _53263_ (_39111_, _02471_, _02466_);
  or _53264_ (_02472_, _01597_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _53265_ (_02473_, _02472_, _01598_);
  and _53266_ (_02474_, _02473_, _01587_);
  and _53267_ (_02475_, _38094_, _36698_);
  and _53268_ (_02476_, _01464_, _38589_);
  and _53269_ (_02477_, _01469_, _42447_);
  and _53270_ (_02478_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _53271_ (_02479_, _02478_, _02477_);
  or _53272_ (_02480_, _02479_, _02476_);
  or _53273_ (_02481_, _02480_, _02475_);
  or _53274_ (_02482_, _01571_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _53275_ (_02483_, _01571_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _53276_ (_02484_, _02483_, _01583_);
  and _53277_ (_02485_, _02484_, _02482_);
  or _53278_ (_02486_, _02485_, _02481_);
  or _53279_ (_02487_, _02486_, _02474_);
  or _53280_ (_02488_, _02487_, _02289_);
  nor _53281_ (_02489_, _01620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _53282_ (_02490_, _02489_, _01621_);
  or _53283_ (_02491_, _02490_, _01460_);
  and _53284_ (_02492_, _02491_, _42618_);
  and _53285_ (_39112_, _02492_, _02488_);
  and _53286_ (_02493_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _53287_ (_02494_, _01826_, _01824_);
  nor _53288_ (_02495_, _02494_, _01827_);
  or _53289_ (_02496_, _02495_, _01635_);
  or _53290_ (_02497_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _53291_ (_02498_, _02497_, _01858_);
  and _53292_ (_02499_, _02498_, _02496_);
  or _53293_ (_39113_, _02499_, _02493_);
  nor _53294_ (_02500_, _01829_, _01827_);
  nor _53295_ (_02501_, _02500_, _01830_);
  or _53296_ (_02502_, _02501_, _01635_);
  or _53297_ (_02503_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _53298_ (_02504_, _02503_, _01858_);
  and _53299_ (_02505_, _02504_, _02502_);
  and _53300_ (_02506_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _53301_ (_39114_, _02506_, _02505_);
  and _53302_ (_02507_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _53303_ (_02508_, _01834_, _01832_);
  nor _53304_ (_02509_, _02508_, _01835_);
  or _53305_ (_02510_, _02509_, _01635_);
  or _53306_ (_02511_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _53307_ (_02512_, _02511_, _01858_);
  and _53308_ (_02513_, _02512_, _02510_);
  or _53309_ (_39115_, _02513_, _02507_);
  and _53310_ (_02514_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53311_ (_02515_, _01835_, _01720_);
  nor _53312_ (_02516_, _02515_, _01836_);
  or _53313_ (_02517_, _02516_, _01635_);
  or _53314_ (_02518_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _53315_ (_02519_, _02518_, _01858_);
  and _53316_ (_02520_, _02519_, _02517_);
  or _53317_ (_39117_, _02520_, _02514_);
  and _53318_ (_02521_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53319_ (_02522_, _01839_, _01836_);
  nor _53320_ (_02523_, _02522_, _01840_);
  or _53321_ (_02524_, _02523_, _01635_);
  or _53322_ (_02525_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _53323_ (_02526_, _02525_, _01858_);
  and _53324_ (_02527_, _02526_, _02524_);
  or _53325_ (_39118_, _02527_, _02521_);
  and _53326_ (_02528_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _53327_ (_02529_, _01840_, _01715_);
  nor _53328_ (_02530_, _02529_, _01841_);
  or _53329_ (_02531_, _02530_, _01635_);
  or _53330_ (_02532_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _53331_ (_02533_, _02532_, _01858_);
  and _53332_ (_02534_, _02533_, _02531_);
  or _53333_ (_39119_, _02534_, _02528_);
  nor _53334_ (_02535_, _01841_, _01711_);
  nor _53335_ (_02536_, _02535_, _01842_);
  or _53336_ (_02537_, _02536_, _01635_);
  or _53337_ (_02538_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _53338_ (_02539_, _02538_, _01858_);
  and _53339_ (_02540_, _02539_, _02537_);
  and _53340_ (_02541_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _53341_ (_39120_, _02541_, _02540_);
  nor _53342_ (_02543_, _01842_, _01707_);
  nor _53343_ (_02544_, _02543_, _01843_);
  or _53344_ (_02545_, _02544_, _01635_);
  or _53345_ (_02546_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _53346_ (_02547_, _02546_, _01858_);
  and _53347_ (_02548_, _02547_, _02545_);
  and _53348_ (_02549_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _53349_ (_39121_, _02549_, _02548_);
  and _53350_ (_02550_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _53351_ (_02551_, _01845_, _01843_);
  nor _53352_ (_02552_, _02551_, _01846_);
  or _53353_ (_02553_, _02552_, _01635_);
  or _53354_ (_02554_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _53355_ (_02555_, _02554_, _01858_);
  and _53356_ (_02556_, _02555_, _02553_);
  or _53357_ (_39122_, _02556_, _02550_);
  nor _53358_ (_02557_, _01846_, _01702_);
  nor _53359_ (_02558_, _02557_, _01847_);
  or _53360_ (_02559_, _02558_, _01635_);
  or _53361_ (_02560_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _53362_ (_02561_, _02560_, _01858_);
  and _53363_ (_02562_, _02561_, _02559_);
  and _53364_ (_02563_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _53365_ (_39123_, _02563_, _02562_);
  nor _53366_ (_02565_, _01847_, _01698_);
  nor _53367_ (_02566_, _02565_, _01848_);
  or _53368_ (_02567_, _02566_, _01635_);
  or _53369_ (_02568_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _53370_ (_02569_, _02568_, _01858_);
  and _53371_ (_02570_, _02569_, _02567_);
  and _53372_ (_02571_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _53373_ (_39124_, _02571_, _02570_);
  nor _53374_ (_02572_, _01848_, _01695_);
  nor _53375_ (_02573_, _02572_, _01849_);
  or _53376_ (_02575_, _02573_, _01635_);
  or _53377_ (_02576_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _53378_ (_02577_, _02576_, _01858_);
  and _53379_ (_02578_, _02577_, _02575_);
  and _53380_ (_02579_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _53381_ (_39125_, _02579_, _02578_);
  or _53382_ (_02580_, _01849_, _01690_);
  nor _53383_ (_02581_, _01850_, _01635_);
  and _53384_ (_02582_, _02581_, _02580_);
  nor _53385_ (_02583_, _01633_, _38302_);
  or _53386_ (_02584_, _02583_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _53387_ (_02585_, _02584_, _02582_);
  or _53388_ (_02586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _36925_);
  and _53389_ (_02587_, _02586_, _42618_);
  and _53390_ (_39126_, _02587_, _02585_);
  nor _53391_ (_02588_, _01850_, _01686_);
  nor _53392_ (_02589_, _02588_, _01851_);
  or _53393_ (_02590_, _02589_, _01635_);
  or _53394_ (_02591_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _53395_ (_02592_, _02591_, _01858_);
  and _53396_ (_02593_, _02592_, _02590_);
  and _53397_ (_02594_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _53398_ (_39128_, _02594_, _02593_);
  or _53399_ (_02595_, _01851_, _01683_);
  and _53400_ (_02596_, _02595_, _01852_);
  or _53401_ (_02597_, _02596_, _01635_);
  or _53402_ (_02598_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _53403_ (_02599_, _02598_, _01858_);
  and _53404_ (_02600_, _02599_, _02597_);
  and _53405_ (_02601_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _53406_ (_39129_, _02601_, _02600_);
  and _53407_ (_02602_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _53408_ (_02603_, _02602_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _53409_ (_39130_, _02603_, _42618_);
  and _53410_ (_02604_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _53411_ (_02605_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _53412_ (_39131_, _02605_, _42618_);
  and _53413_ (_02606_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _53414_ (_02607_, _02606_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _53415_ (_39132_, _02607_, _42618_);
  and _53416_ (_02608_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _53417_ (_02609_, _02608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _53418_ (_39133_, _02609_, _42618_);
  and _53419_ (_02610_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _53420_ (_02611_, _02610_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _53421_ (_39134_, _02611_, _42618_);
  and _53422_ (_02612_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _53423_ (_02613_, _02612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _53424_ (_39135_, _02613_, _42618_);
  and _53425_ (_02614_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _53426_ (_02615_, _02614_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _53427_ (_39136_, _02615_, _42618_);
  nor _53428_ (_02616_, _01823_, _42079_);
  nand _53429_ (_02617_, _02616_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _53430_ (_02618_, _02616_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _53431_ (_02619_, _02618_, _01858_);
  and _53432_ (_39137_, _02619_, _02617_);
  nor _53433_ (_02620_, _01879_, _01877_);
  nor _53434_ (_02621_, _02620_, _01880_);
  or _53435_ (_02622_, _02621_, _42079_);
  or _53436_ (_02623_, _36958_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _53437_ (_02624_, _02623_, _01858_);
  and _53438_ (_39139_, _02624_, _02622_);
  and _53439_ (_02625_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _53440_ (_02626_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _53441_ (_02627_, _02626_, _38765_);
  or _53442_ (_39155_, _02627_, _02625_);
  and _53443_ (_02628_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _53444_ (_02629_, _02056_, _38765_);
  or _53445_ (_39156_, _02629_, _02628_);
  and _53446_ (_02630_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _53447_ (_02631_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _53448_ (_02632_, _02631_, _38765_);
  or _53449_ (_39157_, _02632_, _02630_);
  and _53450_ (_02633_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _53451_ (_02634_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _53452_ (_02635_, _02634_, _38765_);
  or _53453_ (_39158_, _02635_, _02633_);
  and _53454_ (_02636_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _53455_ (_02637_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _53456_ (_02638_, _02637_, _38765_);
  or _53457_ (_39159_, _02638_, _02636_);
  and _53458_ (_02639_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _53459_ (_02640_, _02069_, _38765_);
  or _53460_ (_39161_, _02640_, _02639_);
  and _53461_ (_02641_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _53462_ (_02642_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _53463_ (_02643_, _02642_, _38765_);
  or _53464_ (_39162_, _02643_, _02641_);
  and _53465_ (_39163_, _01909_, _42618_);
  nor _53466_ (_39164_, _01919_, rst);
  and _53467_ (_39165_, _01915_, _42618_);
  and _53468_ (_02644_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _53469_ (_02645_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or _53470_ (_02646_, _02645_, _02644_);
  and _53471_ (_39166_, _02646_, _42618_);
  and _53472_ (_02647_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _53473_ (_02648_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or _53474_ (_02649_, _02648_, _02647_);
  and _53475_ (_39167_, _02649_, _42618_);
  and _53476_ (_02650_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _53477_ (_02651_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or _53478_ (_02652_, _02651_, _02650_);
  and _53479_ (_39168_, _02652_, _42618_);
  and _53480_ (_02653_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _53481_ (_02654_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or _53482_ (_02655_, _02654_, _02653_);
  and _53483_ (_39169_, _02655_, _42618_);
  and _53484_ (_02656_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _53485_ (_02657_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or _53486_ (_02658_, _02657_, _02656_);
  and _53487_ (_39170_, _02658_, _42618_);
  and _53488_ (_02659_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _53489_ (_02660_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or _53490_ (_02661_, _02660_, _02659_);
  and _53491_ (_39171_, _02661_, _42618_);
  and _53492_ (_02662_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _53493_ (_02663_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or _53494_ (_02664_, _02663_, _02662_);
  and _53495_ (_39172_, _02664_, _42618_);
  and _53496_ (_02665_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _53497_ (_02666_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or _53498_ (_02667_, _02666_, _02665_);
  and _53499_ (_39173_, _02667_, _42618_);
  and _53500_ (_02668_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _53501_ (_02669_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or _53502_ (_02670_, _02669_, _02668_);
  and _53503_ (_39174_, _02670_, _42618_);
  and _53504_ (_02671_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _53505_ (_02672_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _53506_ (_02673_, _02672_, _02671_);
  and _53507_ (_39175_, _02673_, _42618_);
  and _53508_ (_02674_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _53509_ (_02675_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _53510_ (_02676_, _02675_, _02674_);
  and _53511_ (_39176_, _02676_, _42618_);
  and _53512_ (_02677_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _53513_ (_02678_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _53514_ (_02679_, _02678_, _02677_);
  and _53515_ (_39177_, _02679_, _42618_);
  and _53516_ (_02680_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _53517_ (_02681_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _53518_ (_02682_, _02681_, _02680_);
  and _53519_ (_39178_, _02682_, _42618_);
  and _53520_ (_02683_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _53521_ (_02684_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _53522_ (_02685_, _02684_, _02683_);
  and _53523_ (_39179_, _02685_, _42618_);
  and _53524_ (_02686_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _53525_ (_02687_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _53526_ (_02688_, _02687_, _02686_);
  and _53527_ (_39180_, _02688_, _42618_);
  and _53528_ (_02689_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _53529_ (_02690_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _53530_ (_02691_, _02690_, _02689_);
  and _53531_ (_39182_, _02691_, _42618_);
  and _53532_ (_02692_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _53533_ (_02693_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _53534_ (_02694_, _02693_, _02692_);
  and _53535_ (_39183_, _02694_, _42618_);
  and _53536_ (_02695_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _53537_ (_02696_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _53538_ (_02697_, _02696_, _02695_);
  and _53539_ (_39184_, _02697_, _42618_);
  and _53540_ (_02698_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _53541_ (_02699_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _53542_ (_02701_, _02699_, _02698_);
  and _53543_ (_39185_, _02701_, _42618_);
  and _53544_ (_02702_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _53545_ (_02703_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _53546_ (_02704_, _02703_, _02702_);
  and _53547_ (_39186_, _02704_, _42618_);
  and _53548_ (_02705_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _53549_ (_02706_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _53550_ (_02707_, _02706_, _02705_);
  and _53551_ (_39187_, _02707_, _42618_);
  and _53552_ (_02708_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _53553_ (_02709_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _53554_ (_02710_, _02709_, _02708_);
  and _53555_ (_39188_, _02710_, _42618_);
  and _53556_ (_02711_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _53557_ (_02712_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _53558_ (_02713_, _02712_, _02711_);
  and _53559_ (_39189_, _02713_, _42618_);
  and _53560_ (_02714_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _53561_ (_02715_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _53562_ (_02716_, _02715_, _02714_);
  and _53563_ (_39190_, _02716_, _42618_);
  and _53564_ (_02717_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _53565_ (_02718_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _53566_ (_02719_, _02718_, _02717_);
  and _53567_ (_39191_, _02719_, _42618_);
  and _53568_ (_02720_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _53569_ (_02721_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _53570_ (_02722_, _02721_, _02720_);
  and _53571_ (_39193_, _02722_, _42618_);
  and _53572_ (_02723_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _53573_ (_02724_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _53574_ (_02725_, _02724_, _02723_);
  and _53575_ (_39194_, _02725_, _42618_);
  and _53576_ (_02726_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _53577_ (_02727_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _53578_ (_02728_, _02727_, _02726_);
  and _53579_ (_39195_, _02728_, _42618_);
  and _53580_ (_02729_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _53581_ (_02730_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _53582_ (_02731_, _02730_, _02729_);
  and _53583_ (_39196_, _02731_, _42618_);
  and _53584_ (_02732_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _53585_ (_02733_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _53586_ (_02734_, _02733_, _02732_);
  and _53587_ (_39197_, _02734_, _42618_);
  and _53588_ (_02735_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _53589_ (_02736_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _53590_ (_02737_, _02736_, _02735_);
  and _53591_ (_39198_, _02737_, _42618_);
  and _53592_ (_02738_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53593_ (_02739_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _53594_ (_02740_, _02739_, _02738_);
  and _53595_ (_39199_, _02740_, _42618_);
  and _53596_ (_02741_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53597_ (_02742_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _53598_ (_02743_, _02742_, _02741_);
  and _53599_ (_39200_, _02743_, _42618_);
  and _53600_ (_02744_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53601_ (_02745_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _53602_ (_02746_, _02745_, _02744_);
  and _53603_ (_39201_, _02746_, _42618_);
  and _53604_ (_02747_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53605_ (_02748_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _53606_ (_02749_, _02748_, _02747_);
  and _53607_ (_39202_, _02749_, _42618_);
  and _53608_ (_02750_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53609_ (_02751_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _53610_ (_02752_, _02751_, _02750_);
  and _53611_ (_39204_, _02752_, _42618_);
  and _53612_ (_02753_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53613_ (_02754_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _53614_ (_02755_, _02754_, _02753_);
  and _53615_ (_39205_, _02755_, _42618_);
  and _53616_ (_02756_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53617_ (_02757_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _53618_ (_02758_, _02757_, _02756_);
  and _53619_ (_39206_, _02758_, _42618_);
  and _53620_ (_02759_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53621_ (_02760_, _42374_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53622_ (_02761_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _53623_ (_02762_, _02761_, _01932_);
  and _53624_ (_02763_, _02762_, _02760_);
  or _53625_ (_02764_, _02763_, _02759_);
  and _53626_ (_39207_, _02764_, _42618_);
  and _53627_ (_02765_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53628_ (_02766_, _42280_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53629_ (_02767_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _53630_ (_02768_, _02767_, _01932_);
  and _53631_ (_02769_, _02768_, _02766_);
  or _53632_ (_02770_, _02769_, _02765_);
  and _53633_ (_39208_, _02770_, _42618_);
  and _53634_ (_02771_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53635_ (_02772_, _42184_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53636_ (_02773_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _53637_ (_02774_, _02773_, _01932_);
  and _53638_ (_02775_, _02774_, _02772_);
  or _53639_ (_02776_, _02775_, _02771_);
  and _53640_ (_39209_, _02776_, _42618_);
  and _53641_ (_02777_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53642_ (_02778_, _42327_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53643_ (_02779_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _53644_ (_02780_, _02779_, _01932_);
  and _53645_ (_02781_, _02780_, _02778_);
  or _53646_ (_02782_, _02781_, _02777_);
  and _53647_ (_39210_, _02782_, _42618_);
  and _53648_ (_02783_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53649_ (_02784_, _42233_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53650_ (_02785_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _53651_ (_02786_, _02785_, _01932_);
  and _53652_ (_02787_, _02786_, _02784_);
  or _53653_ (_02788_, _02787_, _02783_);
  and _53654_ (_39211_, _02788_, _42618_);
  and _53655_ (_02789_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53656_ (_02790_, _42160_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53657_ (_02791_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _53658_ (_02792_, _02791_, _01932_);
  and _53659_ (_02793_, _02792_, _02790_);
  or _53660_ (_02794_, _02793_, _02789_);
  and _53661_ (_39212_, _02794_, _42618_);
  and _53662_ (_02795_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53663_ (_02796_, _42428_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53664_ (_02797_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _53665_ (_02799_, _02797_, _01932_);
  and _53666_ (_02800_, _02799_, _02796_);
  or _53667_ (_02801_, _02800_, _02795_);
  and _53668_ (_39213_, _02801_, _42618_);
  and _53669_ (_02802_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53670_ (_02804_, _42072_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53671_ (_02805_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _53672_ (_02806_, _02805_, _01932_);
  and _53673_ (_02807_, _02806_, _02804_);
  or _53674_ (_02808_, _02807_, _02802_);
  and _53675_ (_39215_, _02808_, _42618_);
  and _53676_ (_02810_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _53677_ (_02811_, _02810_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53678_ (_02812_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _01932_);
  and _53679_ (_02813_, _02812_, _42618_);
  and _53680_ (_39216_, _02813_, _02811_);
  and _53681_ (_02815_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _53682_ (_02816_, _02815_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53683_ (_02817_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _01932_);
  and _53684_ (_02818_, _02817_, _42618_);
  and _53685_ (_39217_, _02818_, _02816_);
  and _53686_ (_02820_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _53687_ (_02821_, _02820_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53688_ (_02822_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _01932_);
  and _53689_ (_02823_, _02822_, _42618_);
  and _53690_ (_39218_, _02823_, _02821_);
  and _53691_ (_02825_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _53692_ (_02826_, _02825_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53693_ (_02827_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _01932_);
  and _53694_ (_02828_, _02827_, _42618_);
  and _53695_ (_39219_, _02828_, _02826_);
  and _53696_ (_02830_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _53697_ (_02832_, _02830_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53698_ (_02833_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _01932_);
  and _53699_ (_02834_, _02833_, _42618_);
  and _53700_ (_39220_, _02834_, _02832_);
  and _53701_ (_02835_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _53702_ (_02837_, _02835_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53703_ (_02838_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _01932_);
  and _53704_ (_02840_, _02838_, _42618_);
  and _53705_ (_39221_, _02840_, _02837_);
  and _53706_ (_02841_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _53707_ (_02843_, _02841_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53708_ (_02844_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _01932_);
  and _53709_ (_02845_, _02844_, _42618_);
  and _53710_ (_39222_, _02845_, _02843_);
  nand _53711_ (_02847_, _01946_, _32323_);
  or _53712_ (_02849_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _53713_ (_02851_, _02849_, _42618_);
  and _53714_ (_39223_, _02851_, _02847_);
  nand _53715_ (_02852_, _01946_, _33020_);
  or _53716_ (_02854_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _53717_ (_02855_, _02854_, _42618_);
  and _53718_ (_39224_, _02855_, _02852_);
  nand _53719_ (_02857_, _01946_, _33717_);
  or _53720_ (_02858_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _53721_ (_02859_, _02858_, _42618_);
  and _53722_ (_39226_, _02859_, _02857_);
  nand _53723_ (_02861_, _01946_, _34478_);
  or _53724_ (_02863_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _53725_ (_02864_, _02863_, _42618_);
  and _53726_ (_39227_, _02864_, _02861_);
  nand _53727_ (_02865_, _01946_, _35240_);
  or _53728_ (_02866_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _53729_ (_02867_, _02866_, _42618_);
  and _53730_ (_39228_, _02867_, _02865_);
  nand _53731_ (_02869_, _01946_, _36046_);
  or _53732_ (_02871_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _53733_ (_02872_, _02871_, _42618_);
  and _53734_ (_39229_, _02872_, _02869_);
  not _53735_ (_02874_, _01946_);
  or _53736_ (_02875_, _02874_, _36698_);
  or _53737_ (_02877_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _53738_ (_02878_, _02877_, _42618_);
  and _53739_ (_39230_, _02878_, _02875_);
  nand _53740_ (_02880_, _01946_, _31136_);
  or _53741_ (_02881_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _53742_ (_02883_, _02881_, _42618_);
  and _53743_ (_39231_, _02883_, _02880_);
  nand _53744_ (_02885_, _01946_, _38405_);
  or _53745_ (_02886_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _53746_ (_02888_, _02886_, _42618_);
  and _53747_ (_39232_, _02888_, _02885_);
  nand _53748_ (_02889_, _01946_, _38436_);
  or _53749_ (_02891_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _53750_ (_02892_, _02891_, _42618_);
  and _53751_ (_39233_, _02892_, _02889_);
  nand _53752_ (_02895_, _01946_, _38466_);
  or _53753_ (_02896_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _53754_ (_02897_, _02896_, _42618_);
  and _53755_ (_39234_, _02897_, _02895_);
  nand _53756_ (_02899_, _01946_, _38497_);
  or _53757_ (_02900_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _53758_ (_02901_, _02900_, _42618_);
  and _53759_ (_39235_, _02901_, _02899_);
  nand _53760_ (_02903_, _01946_, _38528_);
  or _53761_ (_02904_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _53762_ (_02906_, _02904_, _42618_);
  and _53763_ (_39237_, _02906_, _02903_);
  nand _53764_ (_02907_, _01946_, _38561_);
  or _53765_ (_02909_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _53766_ (_02910_, _02909_, _42618_);
  and _53767_ (_39238_, _02910_, _02907_);
  or _53768_ (_02912_, _02874_, _38589_);
  or _53769_ (_02913_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _53770_ (_02914_, _02913_, _42618_);
  and _53771_ (_39239_, _02914_, _02912_);
  nor _53772_ (_39457_, _42115_, rst);
  and _53773_ (_02917_, _42030_, _38137_);
  and _53774_ (_02919_, _02917_, _28091_);
  and _53775_ (_02920_, _02919_, _42032_);
  nand _53776_ (_02922_, _02920_, _38225_);
  or _53777_ (_02923_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _53778_ (_02924_, _02923_, _42618_);
  and _53779_ (_39458_, _02924_, _02922_);
  and _53780_ (_02925_, _02917_, _39011_);
  not _53781_ (_02926_, _02925_);
  nor _53782_ (_02928_, _02926_, _38225_);
  not _53783_ (_02930_, _42032_);
  and _53784_ (_02931_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _53785_ (_02932_, _02931_, _02930_);
  or _53786_ (_02934_, _02932_, _02928_);
  or _53787_ (_02935_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _53788_ (_02936_, _02935_, _42618_);
  and _53789_ (_39459_, _02936_, _02934_);
  and _53790_ (_02938_, _38813_, _31790_);
  and _53791_ (_02939_, _02917_, _02938_);
  and _53792_ (_02942_, _02939_, _42032_);
  nand _53793_ (_02943_, _02942_, _38225_);
  or _53794_ (_02944_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _53795_ (_02946_, _02944_, _42618_);
  and _53796_ (_39460_, _02946_, _02943_);
  and _53797_ (_02947_, _02917_, _41127_);
  and _53798_ (_02949_, _02947_, _42032_);
  not _53799_ (_02950_, _02949_);
  nor _53800_ (_02951_, _02950_, _38225_);
  and _53801_ (_02953_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _53802_ (_02955_, _02953_, _02951_);
  and _53803_ (_39462_, _02955_, _42618_);
  and _53804_ (_02957_, _42030_, _38629_);
  and _53805_ (_02958_, _02957_, _28091_);
  and _53806_ (_02959_, _02958_, _42032_);
  not _53807_ (_02961_, _02959_);
  nor _53808_ (_02962_, _02961_, _38225_);
  nor _53809_ (_02963_, _02925_, _02919_);
  not _53810_ (_02965_, _02939_);
  and _53811_ (_02966_, _02965_, _02963_);
  not _53812_ (_02968_, _02947_);
  and _53813_ (_02970_, _02968_, _02966_);
  not _53814_ (_02971_, _02958_);
  and _53815_ (_02972_, _02971_, _02970_);
  or _53816_ (_02974_, _02972_, _02930_);
  or _53817_ (_02975_, _02974_, _02919_);
  and _53818_ (_02976_, _02975_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or _53819_ (_02978_, _02947_, _02939_);
  or _53820_ (_02979_, _02978_, _02925_);
  and _53821_ (_02980_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _53822_ (_02983_, _02980_, _02979_);
  or _53823_ (_02984_, _02983_, _02976_);
  or _53824_ (_02985_, _02984_, _02962_);
  and _53825_ (_39463_, _02985_, _42618_);
  and _53826_ (_02987_, _02957_, _39011_);
  nor _53827_ (_02989_, _02987_, _02958_);
  and _53828_ (_02990_, _02989_, _02968_);
  and _53829_ (_02991_, _02990_, _02966_);
  or _53830_ (_02992_, _02958_, _02978_);
  and _53831_ (_02994_, _02992_, _42032_);
  nand _53832_ (_02996_, _02963_, _42032_);
  or _53833_ (_02997_, _02996_, _02994_);
  or _53834_ (_02999_, _02997_, _02991_);
  and _53835_ (_03000_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _53836_ (_03001_, _02987_, _42032_);
  and _53837_ (_03003_, _03001_, _41608_);
  or _53838_ (_03004_, _03003_, _03000_);
  and _53839_ (_39464_, _03004_, _42618_);
  and _53840_ (_03006_, _02957_, _02938_);
  and _53841_ (_03007_, _03006_, _42032_);
  not _53842_ (_03009_, _03007_);
  and _53843_ (_03011_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor _53844_ (_03012_, _03009_, _38225_);
  or _53845_ (_03013_, _03012_, _03011_);
  and _53846_ (_39465_, _03013_, _42618_);
  and _53847_ (_03015_, _02957_, _41127_);
  and _53848_ (_03016_, _03015_, _42032_);
  not _53849_ (_03018_, _03016_);
  nor _53850_ (_03019_, _03018_, _38225_);
  not _53851_ (_03021_, _03006_);
  and _53852_ (_03023_, _03021_, _02989_);
  nor _53853_ (_03024_, _03015_, _03006_);
  and _53854_ (_03025_, _03024_, _02991_);
  nand _53855_ (_03027_, _02970_, _42032_);
  nor _53856_ (_03028_, _03027_, _03025_);
  nand _53857_ (_03029_, _03028_, _03023_);
  and _53858_ (_03031_, _03029_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or _53859_ (_03032_, _03031_, _03019_);
  and _53860_ (_39466_, _03032_, _42618_);
  nand _53861_ (_03034_, _02920_, _38203_);
  or _53862_ (_03035_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _53863_ (_03036_, _03035_, _42618_);
  and _53864_ (_39555_, _03036_, _03034_);
  nand _53865_ (_03038_, _02920_, _38191_);
  or _53866_ (_03039_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _53867_ (_03041_, _03039_, _42618_);
  and _53868_ (_39556_, _03041_, _03038_);
  nand _53869_ (_03042_, _02920_, _38184_);
  or _53870_ (_03044_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _53871_ (_03045_, _03044_, _42618_);
  and _53872_ (_39557_, _03045_, _03042_);
  nand _53873_ (_03047_, _02920_, _38177_);
  or _53874_ (_03048_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _53875_ (_03050_, _03048_, _42618_);
  and _53876_ (_39558_, _03050_, _03047_);
  nand _53877_ (_03051_, _02920_, _38169_);
  or _53878_ (_03052_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _53879_ (_03053_, _03052_, _42618_);
  and _53880_ (_39559_, _03053_, _03051_);
  nand _53881_ (_03054_, _02920_, _38162_);
  or _53882_ (_03056_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _53883_ (_03057_, _03056_, _42618_);
  and _53884_ (_39560_, _03057_, _03054_);
  nand _53885_ (_03059_, _02920_, _38155_);
  or _53886_ (_03060_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _53887_ (_03061_, _03060_, _42618_);
  and _53888_ (_39561_, _03061_, _03059_);
  and _53889_ (_03063_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _53890_ (_03064_, _02926_, _38203_);
  or _53891_ (_03066_, _03064_, _02930_);
  or _53892_ (_03067_, _03066_, _03063_);
  or _53893_ (_03068_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _53894_ (_03070_, _03068_, _42618_);
  and _53895_ (_39562_, _03070_, _03067_);
  nor _53896_ (_03071_, _02926_, _38191_);
  and _53897_ (_03073_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _53898_ (_03074_, _03073_, _02930_);
  or _53899_ (_03075_, _03074_, _03071_);
  or _53900_ (_03077_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _53901_ (_03078_, _03077_, _42618_);
  and _53902_ (_39563_, _03078_, _03075_);
  nor _53903_ (_03080_, _02926_, _38184_);
  and _53904_ (_03081_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _53905_ (_03082_, _03081_, _02930_);
  or _53906_ (_03084_, _03082_, _03080_);
  or _53907_ (_03085_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _53908_ (_03086_, _03085_, _42618_);
  and _53909_ (_39564_, _03086_, _03084_);
  nor _53910_ (_03088_, _02926_, _38177_);
  and _53911_ (_03089_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _53912_ (_03091_, _03089_, _02930_);
  or _53913_ (_03092_, _03091_, _03088_);
  or _53914_ (_03093_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _53915_ (_03095_, _03093_, _42618_);
  and _53916_ (_39566_, _03095_, _03092_);
  nor _53917_ (_03096_, _02926_, _38169_);
  and _53918_ (_03098_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _53919_ (_03099_, _03098_, _02930_);
  or _53920_ (_03100_, _03099_, _03096_);
  or _53921_ (_03102_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _53922_ (_03103_, _03102_, _42618_);
  and _53923_ (_39567_, _03103_, _03100_);
  nor _53924_ (_03105_, _02926_, _38162_);
  and _53925_ (_03106_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _53926_ (_03108_, _03106_, _02930_);
  or _53927_ (_03109_, _03108_, _03105_);
  or _53928_ (_03110_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _53929_ (_03111_, _03110_, _42618_);
  and _53930_ (_39568_, _03111_, _03109_);
  nor _53931_ (_03113_, _02926_, _38155_);
  and _53932_ (_03114_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _53933_ (_03116_, _03114_, _02930_);
  or _53934_ (_03117_, _03116_, _03113_);
  or _53935_ (_03118_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _53936_ (_03120_, _03118_, _42618_);
  and _53937_ (_39569_, _03120_, _03117_);
  nand _53938_ (_03121_, _02942_, _38203_);
  or _53939_ (_03123_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _53940_ (_03124_, _03123_, _03121_);
  and _53941_ (_39570_, _03124_, _42618_);
  not _53942_ (_03127_, _02942_);
  nor _53943_ (_03128_, _03127_, _38191_);
  and _53944_ (_03129_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or _53945_ (_03131_, _03129_, _03128_);
  and _53946_ (_39571_, _03131_, _42618_);
  nor _53947_ (_03132_, _03127_, _38184_);
  and _53948_ (_03134_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or _53949_ (_03135_, _03134_, _03132_);
  and _53950_ (_39572_, _03135_, _42618_);
  nor _53951_ (_03137_, _03127_, _38177_);
  and _53952_ (_03138_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or _53953_ (_03139_, _03138_, _03137_);
  and _53954_ (_39573_, _03139_, _42618_);
  nand _53955_ (_03141_, _02942_, _38169_);
  or _53956_ (_03142_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _53957_ (_03144_, _03142_, _42618_);
  and _53958_ (_39574_, _03144_, _03141_);
  nor _53959_ (_03145_, _03127_, _38162_);
  and _53960_ (_03147_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _53961_ (_03148_, _03147_, _03145_);
  and _53962_ (_39575_, _03148_, _42618_);
  nor _53963_ (_03150_, _03127_, _38155_);
  and _53964_ (_03151_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _53965_ (_03152_, _03151_, _03150_);
  and _53966_ (_39577_, _03152_, _42618_);
  and _53967_ (_03154_, _02949_, _38204_);
  and _53968_ (_03155_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _53969_ (_03157_, _03155_, _03154_);
  and _53970_ (_39578_, _03157_, _42618_);
  nor _53971_ (_03158_, _02950_, _38191_);
  and _53972_ (_03160_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _53973_ (_03161_, _03160_, _03158_);
  and _53974_ (_39579_, _03161_, _42618_);
  and _53975_ (_03163_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _53976_ (_03164_, _02950_, _38184_);
  or _53977_ (_03165_, _03164_, _03163_);
  and _53978_ (_39580_, _03165_, _42618_);
  nor _53979_ (_03167_, _02950_, _38177_);
  and _53980_ (_03168_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _53981_ (_03169_, _03168_, _03167_);
  and _53982_ (_39581_, _03169_, _42618_);
  nor _53983_ (_03171_, _02950_, _38169_);
  and _53984_ (_03172_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or _53985_ (_03174_, _03172_, _03171_);
  and _53986_ (_39582_, _03174_, _42618_);
  nor _53987_ (_03175_, _02950_, _38162_);
  and _53988_ (_03177_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or _53989_ (_03178_, _03177_, _03175_);
  and _53990_ (_39583_, _03178_, _42618_);
  nor _53991_ (_03180_, _02950_, _38155_);
  and _53992_ (_03181_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _53993_ (_03182_, _03181_, _03180_);
  and _53994_ (_39584_, _03182_, _42618_);
  and _53995_ (_03184_, _02959_, _38204_);
  and _53996_ (_03185_, _02961_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or _53997_ (_03187_, _03185_, _03184_);
  and _53998_ (_39585_, _03187_, _42618_);
  and _53999_ (_03189_, _02971_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _54000_ (_03190_, _02971_, _38191_);
  or _54001_ (_03191_, _03190_, _03189_);
  or _54002_ (_03192_, _03191_, _02930_);
  or _54003_ (_03194_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _54004_ (_03195_, _03194_, _42618_);
  and _54005_ (_39586_, _03195_, _03192_);
  nor _54006_ (_03197_, _02971_, _38184_);
  and _54007_ (_03198_, _02971_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or _54008_ (_03199_, _03198_, _02930_);
  or _54009_ (_03201_, _03199_, _03197_);
  or _54010_ (_03202_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _54011_ (_03203_, _03202_, _42618_);
  and _54012_ (_39588_, _03203_, _03201_);
  and _54013_ (_03205_, _02975_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _54014_ (_03206_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _54015_ (_03208_, _03206_, _02979_);
  nor _54016_ (_03209_, _02961_, _38177_);
  or _54017_ (_03210_, _03209_, _03208_);
  or _54018_ (_03212_, _03210_, _03205_);
  and _54019_ (_39589_, _03212_, _42618_);
  and _54020_ (_03213_, _02975_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _54021_ (_03215_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _54022_ (_03216_, _03215_, _02979_);
  nor _54023_ (_03218_, _02961_, _38169_);
  or _54024_ (_03219_, _03218_, _03216_);
  or _54025_ (_03220_, _03219_, _03213_);
  and _54026_ (_39590_, _03220_, _42618_);
  nor _54027_ (_03222_, _02961_, _38162_);
  and _54028_ (_03223_, _02961_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or _54029_ (_03224_, _03223_, _03222_);
  and _54030_ (_39591_, _03224_, _42618_);
  nor _54031_ (_03226_, _02961_, _38155_);
  and _54032_ (_03227_, _02975_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _54033_ (_03229_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _54034_ (_03230_, _03229_, _02979_);
  or _54035_ (_03231_, _03230_, _03227_);
  or _54036_ (_03233_, _03231_, _03226_);
  and _54037_ (_39592_, _03233_, _42618_);
  and _54038_ (_03234_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _54039_ (_03236_, _03001_, _38204_);
  or _54040_ (_03237_, _03236_, _03234_);
  and _54041_ (_39593_, _03237_, _42618_);
  and _54042_ (_03239_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _54043_ (_03240_, _03001_, _42278_);
  or _54044_ (_03241_, _03240_, _03239_);
  and _54045_ (_39594_, _03241_, _42618_);
  and _54046_ (_03243_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _54047_ (_03245_, _03001_, _39884_);
  or _54048_ (_03246_, _03245_, _03243_);
  and _54049_ (_39595_, _03246_, _42618_);
  and _54050_ (_03247_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _54051_ (_03249_, _03001_, _39896_);
  or _54052_ (_03250_, _03249_, _03247_);
  and _54053_ (_39596_, _03250_, _42618_);
  and _54054_ (_03252_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _54055_ (_03253_, _03001_, _39907_);
  or _54056_ (_03254_, _03253_, _03252_);
  and _54057_ (_39597_, _03254_, _42618_);
  and _54058_ (_03256_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _54059_ (_03257_, _03001_, _39920_);
  or _54060_ (_03259_, _03257_, _03256_);
  and _54061_ (_39599_, _03259_, _42618_);
  and _54062_ (_03260_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _54063_ (_03262_, _03001_, _39933_);
  or _54064_ (_03263_, _03262_, _03260_);
  and _54065_ (_39600_, _03263_, _42618_);
  and _54066_ (_03265_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _54067_ (_03266_, _03007_, _38204_);
  or _54068_ (_03267_, _03266_, _03265_);
  and _54069_ (_39601_, _03267_, _42618_);
  and _54070_ (_03269_, _03023_, _02970_);
  nor _54071_ (_03270_, _03269_, _02930_);
  nand _54072_ (_03271_, _03270_, _02966_);
  and _54073_ (_03272_, _03271_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _54074_ (_03273_, _03009_, _38191_);
  nand _54075_ (_03274_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _54076_ (_03275_, _03274_, _02990_);
  or _54077_ (_03276_, _03275_, _03273_);
  or _54078_ (_03277_, _03276_, _03272_);
  and _54079_ (_39602_, _03277_, _42618_);
  nor _54080_ (_03278_, _03009_, _38184_);
  and _54081_ (_03279_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or _54082_ (_03280_, _03279_, _03278_);
  and _54083_ (_39603_, _03280_, _42618_);
  nor _54084_ (_03281_, _03009_, _38177_);
  and _54085_ (_03282_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or _54086_ (_03283_, _03282_, _03281_);
  and _54087_ (_39604_, _03283_, _42618_);
  nor _54088_ (_03284_, _03009_, _38169_);
  and _54089_ (_03285_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or _54090_ (_03286_, _03285_, _03284_);
  and _54091_ (_39605_, _03286_, _42618_);
  nor _54092_ (_03287_, _03009_, _38162_);
  and _54093_ (_03288_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _54094_ (_03289_, _03288_, _03287_);
  and _54095_ (_39606_, _03289_, _42618_);
  nor _54096_ (_03290_, _03009_, _38155_);
  and _54097_ (_03291_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _54098_ (_03292_, _03291_, _03290_);
  and _54099_ (_39607_, _03292_, _42618_);
  and _54100_ (_03293_, _03024_, _02989_);
  or _54101_ (_03294_, _03293_, _02930_);
  and _54102_ (_03295_, _03294_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _54103_ (_03296_, _03016_, _38204_);
  nand _54104_ (_03297_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _54105_ (_03298_, _03297_, _03023_);
  or _54106_ (_03299_, _03298_, _03296_);
  or _54107_ (_03300_, _03299_, _03295_);
  and _54108_ (_39608_, _03300_, _42618_);
  and _54109_ (_03301_, _03029_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor _54110_ (_03302_, _03018_, _38191_);
  or _54111_ (_03303_, _03302_, _03301_);
  and _54112_ (_39610_, _03303_, _42618_);
  and _54113_ (_03304_, _03294_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _54114_ (_03305_, _03018_, _38184_);
  nand _54115_ (_03306_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _54116_ (_03307_, _03306_, _03023_);
  or _54117_ (_03308_, _03307_, _03305_);
  or _54118_ (_03309_, _03308_, _03304_);
  and _54119_ (_39611_, _03309_, _42618_);
  and _54120_ (_03310_, _03294_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _54121_ (_03311_, _03018_, _38177_);
  nand _54122_ (_03312_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _54123_ (_03313_, _03312_, _03023_);
  or _54124_ (_03314_, _03313_, _03311_);
  or _54125_ (_03315_, _03314_, _03310_);
  and _54126_ (_39612_, _03315_, _42618_);
  nor _54127_ (_03316_, _03018_, _38169_);
  and _54128_ (_03317_, _03018_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or _54129_ (_03318_, _03317_, _03316_);
  and _54130_ (_39613_, _03318_, _42618_);
  and _54131_ (_03319_, _03018_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _54132_ (_03320_, _03018_, _38162_);
  or _54133_ (_03321_, _03320_, _03319_);
  and _54134_ (_39614_, _03321_, _42618_);
  and _54135_ (_03322_, _03294_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _54136_ (_03323_, _03018_, _38155_);
  nand _54137_ (_03324_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _54138_ (_03325_, _03324_, _03023_);
  or _54139_ (_03326_, _03325_, _03323_);
  or _54140_ (_03327_, _03326_, _03322_);
  and _54141_ (_39615_, _03327_, _42618_);
  not _54142_ (_03329_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _54143_ (_03330_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _54144_ (_03331_, _03330_, _03329_);
  and _54145_ (_03332_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _42618_);
  and _54146_ (_39679_, _03332_, _03331_);
  nor _54147_ (_03333_, _03331_, rst);
  nand _54148_ (_03334_, _03330_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _54149_ (_03335_, _03330_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _54150_ (_03336_, _03335_, _03334_);
  and _54151_ (_39681_, _03336_, _03333_);
  nor _54152_ (_03337_, _42451_, _42164_);
  not _54153_ (_03338_, _42100_);
  and _54154_ (_03339_, _42259_, _03338_);
  and _54155_ (_03340_, _03339_, _42354_);
  and _54156_ (_03341_, _03340_, _03337_);
  and _54157_ (_03342_, _03341_, _38785_);
  nor _54158_ (_03343_, _03342_, _01393_);
  nor _54159_ (_03344_, _42212_, _38162_);
  and _54160_ (_03345_, _42212_, _42278_);
  or _54161_ (_03346_, _03345_, _03344_);
  not _54162_ (_03347_, _42400_);
  and _54163_ (_03348_, _03347_, _42307_);
  and _54164_ (_03349_, _03348_, _03346_);
  or _54165_ (_03350_, _42212_, _39933_);
  nor _54166_ (_03351_, _03347_, _42307_);
  nand _54167_ (_03352_, _42212_, _38184_);
  and _54168_ (_03353_, _03352_, _03351_);
  and _54169_ (_03354_, _03353_, _03350_);
  nor _54170_ (_03355_, _42212_, _38225_);
  and _54171_ (_03356_, _42212_, _39896_);
  or _54172_ (_03357_, _03356_, _03355_);
  nor _54173_ (_03358_, _42400_, _42307_);
  and _54174_ (_03359_, _03358_, _03357_);
  nand _54175_ (_03360_, _42212_, _38203_);
  and _54176_ (_03361_, _42400_, _42307_);
  or _54177_ (_03362_, _42212_, _39907_);
  and _54178_ (_03363_, _03362_, _03361_);
  and _54179_ (_03364_, _03363_, _03360_);
  or _54180_ (_03365_, _03364_, _03359_);
  or _54181_ (_03366_, _03365_, _03354_);
  nor _54182_ (_03367_, _03366_, _03349_);
  nor _54183_ (_03368_, _03367_, _03343_);
  nor _54184_ (_03369_, _42451_, _42165_);
  nor _54185_ (_03370_, _42259_, _42100_);
  and _54186_ (_03371_, _03370_, _42354_);
  and _54187_ (_03372_, _03371_, _03369_);
  nor _54188_ (_03373_, _38899_, _38887_);
  and _54189_ (_03374_, _38899_, _38887_);
  nor _54190_ (_03375_, _03374_, _03373_);
  and _54191_ (_03376_, _38872_, _38857_);
  nor _54192_ (_03377_, _38872_, _38857_);
  or _54193_ (_03378_, _03377_, _03376_);
  nor _54194_ (_03379_, _03378_, _03375_);
  and _54195_ (_03380_, _03378_, _03375_);
  nor _54196_ (_03381_, _03380_, _03379_);
  nor _54197_ (_03382_, _38923_, _38911_);
  and _54198_ (_03383_, _38923_, _38911_);
  nor _54199_ (_03384_, _03383_, _03382_);
  not _54200_ (_03385_, _38809_);
  nor _54201_ (_03386_, _38933_, _03385_);
  and _54202_ (_03387_, _38933_, _03385_);
  nor _54203_ (_03388_, _03387_, _03386_);
  nor _54204_ (_03389_, _03388_, _03384_);
  and _54205_ (_03390_, _03388_, _03384_);
  or _54206_ (_03391_, _03390_, _03389_);
  nor _54207_ (_03392_, _03391_, _03381_);
  and _54208_ (_03393_, _03391_, _03381_);
  nor _54209_ (_03394_, _03393_, _03392_);
  nand _54210_ (_03395_, _03394_, _42212_);
  or _54211_ (_03396_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _54212_ (_03397_, _03396_, _03361_);
  and _54213_ (_03398_, _03397_, _03395_);
  not _54214_ (_03399_, _42212_);
  and _54215_ (_03400_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _54216_ (_03401_, _03358_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _54217_ (_03402_, _03401_, _03400_);
  and _54218_ (_03403_, _03402_, _03399_);
  nor _54219_ (_03404_, _42212_, _34086_);
  and _54220_ (_03405_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _54221_ (_03406_, _03405_, _03404_);
  and _54222_ (_03407_, _03406_, _03351_);
  and _54223_ (_03408_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _54224_ (_03409_, _03358_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _54225_ (_03410_, _03409_, _03408_);
  and _54226_ (_03411_, _03410_, _42212_);
  or _54227_ (_03412_, _03411_, _03407_);
  or _54228_ (_03413_, _03412_, _03403_);
  or _54229_ (_03414_, _03413_, _03398_);
  and _54230_ (_03415_, _03414_, _03372_);
  and _54231_ (_03416_, _01387_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _54232_ (_03417_, _03358_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _54233_ (_03418_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _54234_ (_03419_, _03418_, _03417_);
  and _54235_ (_03420_, _03419_, _03399_);
  or _54236_ (_03421_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _54237_ (_03422_, _42212_, _38815_);
  and _54238_ (_03423_, _03422_, _03361_);
  and _54239_ (_03424_, _03423_, _03421_);
  and _54240_ (_03425_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _54241_ (_03426_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _54242_ (_03427_, _03426_, _03425_);
  and _54243_ (_03428_, _03427_, _03351_);
  or _54244_ (_03429_, _03428_, _03424_);
  and _54245_ (_03430_, _03358_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _54246_ (_03431_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _54247_ (_03432_, _03431_, _03430_);
  and _54248_ (_03433_, _03432_, _42212_);
  or _54249_ (_03434_, _03433_, _03429_);
  or _54250_ (_03435_, _03434_, _03420_);
  and _54251_ (_03436_, _03435_, _03341_);
  or _54252_ (_03437_, _03436_, _03416_);
  and _54253_ (_03438_, _03369_, _03339_);
  and _54254_ (_03439_, _03438_, _42355_);
  and _54255_ (_03440_, _03361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _54256_ (_03441_, _03351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _54257_ (_03442_, _03441_, _03440_);
  and _54258_ (_03443_, _03442_, _03399_);
  and _54259_ (_03444_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _54260_ (_03445_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _54261_ (_03446_, _03445_, _03444_);
  and _54262_ (_03447_, _03446_, _03358_);
  and _54263_ (_03448_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nor _54264_ (_03449_, _42212_, _41014_);
  or _54265_ (_03450_, _03449_, _03448_);
  and _54266_ (_03451_, _03450_, _03348_);
  or _54267_ (_03452_, _03451_, _03447_);
  and _54268_ (_03453_, _03361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _54269_ (_03454_, _03351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _54270_ (_03455_, _03454_, _03453_);
  and _54271_ (_03456_, _03455_, _42212_);
  or _54272_ (_03457_, _03456_, _03452_);
  or _54273_ (_03458_, _03457_, _03443_);
  and _54274_ (_03459_, _03458_, _03439_);
  and _54275_ (_03460_, _42451_, _42164_);
  and _54276_ (_03461_, _03460_, _03340_);
  nor _54277_ (_03462_, _00790_, _38035_);
  and _54278_ (_03463_, _03462_, _00855_);
  nor _54279_ (_03464_, _00853_, _38109_);
  and _54280_ (_03465_, _38053_, _37985_);
  not _54281_ (_03466_, _03465_);
  and _54282_ (_03467_, _03466_, _03464_);
  and _54283_ (_03468_, _38016_, _37395_);
  nor _54284_ (_03469_, _03468_, _38065_);
  nor _54285_ (_03470_, _00792_, _38047_);
  and _54286_ (_03471_, _03470_, _03469_);
  and _54287_ (_03472_, _03471_, _03467_);
  and _54288_ (_03473_, _03472_, _01112_);
  and _54289_ (_03474_, _03473_, _03463_);
  and _54290_ (_03475_, _03474_, _38032_);
  nor _54291_ (_03476_, _03475_, _36914_);
  nor _54292_ (_03477_, _03476_, p0_in[0]);
  and _54293_ (_03478_, _03476_, _39007_);
  nor _54294_ (_03479_, _03478_, _03477_);
  or _54295_ (_03480_, _03479_, _03399_);
  nor _54296_ (_03481_, _03476_, p0_in[4]);
  and _54297_ (_03482_, _03476_, _39258_);
  nor _54298_ (_03483_, _03482_, _03481_);
  or _54299_ (_03484_, _03483_, _42212_);
  and _54300_ (_03485_, _03484_, _03361_);
  and _54301_ (_03486_, _03485_, _03480_);
  or _54302_ (_03487_, _03476_, p0_in[3]);
  not _54303_ (_03488_, _03476_);
  or _54304_ (_03489_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _54305_ (_03490_, _03489_, _03487_);
  or _54306_ (_03491_, _03490_, _03399_);
  or _54307_ (_03492_, _03476_, p0_in[7]);
  or _54308_ (_03493_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _54309_ (_03494_, _03493_, _03492_);
  or _54310_ (_03495_, _03494_, _42212_);
  and _54311_ (_03496_, _03495_, _03358_);
  and _54312_ (_03497_, _03496_, _03491_);
  or _54313_ (_03498_, _03497_, _03486_);
  or _54314_ (_03499_, _03476_, p0_in[5]);
  or _54315_ (_03500_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _54316_ (_03501_, _03500_, _03499_);
  and _54317_ (_03502_, _03501_, _03399_);
  or _54318_ (_03503_, _03476_, p0_in[1]);
  or _54319_ (_03504_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _54320_ (_03505_, _03504_, _03503_);
  and _54321_ (_03506_, _03505_, _42212_);
  or _54322_ (_03507_, _03506_, _03502_);
  and _54323_ (_03508_, _03507_, _03348_);
  or _54324_ (_03509_, _03476_, p0_in[2]);
  nand _54325_ (_03510_, _03476_, _39024_);
  and _54326_ (_03511_, _03510_, _03509_);
  or _54327_ (_03512_, _03511_, _03399_);
  or _54328_ (_03513_, _03476_, p0_in[6]);
  or _54329_ (_03514_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _54330_ (_03515_, _03514_, _03513_);
  or _54331_ (_03516_, _03515_, _42212_);
  and _54332_ (_03517_, _03516_, _03351_);
  and _54333_ (_03518_, _03517_, _03512_);
  or _54334_ (_03519_, _03518_, _03508_);
  or _54335_ (_03520_, _03519_, _03498_);
  and _54336_ (_03521_, _03520_, _03461_);
  or _54337_ (_03522_, _03521_, _03459_);
  or _54338_ (_03523_, _03522_, _03437_);
  and _54339_ (_03524_, _42451_, _42165_);
  and _54340_ (_03525_, _03370_, _42355_);
  or _54341_ (_03526_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand _54342_ (_03528_, _42212_, _40470_);
  and _54343_ (_03529_, _03528_, _03358_);
  and _54344_ (_03530_, _03529_, _03526_);
  and _54345_ (_03531_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _54346_ (_03532_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _54347_ (_03533_, _03532_, _03531_);
  and _54348_ (_03534_, _03533_, _03351_);
  or _54349_ (_03535_, _03534_, _03530_);
  and _54350_ (_03536_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor _54351_ (_03537_, _42212_, _40465_);
  or _54352_ (_03538_, _03537_, _03536_);
  and _54353_ (_03539_, _03538_, _03361_);
  and _54354_ (_03540_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _54355_ (_03541_, _42212_, _40467_);
  or _54356_ (_03542_, _03541_, _03540_);
  and _54357_ (_03543_, _03542_, _03348_);
  or _54358_ (_03544_, _03543_, _03539_);
  or _54359_ (_03545_, _03544_, _03535_);
  and _54360_ (_03546_, _03545_, _03525_);
  or _54361_ (_03547_, _03476_, p2_in[3]);
  or _54362_ (_03548_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _54363_ (_03549_, _03548_, _03547_);
  or _54364_ (_03550_, _03549_, _03399_);
  or _54365_ (_03551_, _03476_, p2_in[7]);
  or _54366_ (_03552_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _54367_ (_03553_, _03552_, _03551_);
  or _54368_ (_03554_, _03553_, _42212_);
  and _54369_ (_03555_, _03554_, _03358_);
  and _54370_ (_03556_, _03555_, _03550_);
  or _54371_ (_03557_, _03476_, p2_in[6]);
  or _54372_ (_03558_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _54373_ (_03559_, _03558_, _03557_);
  and _54374_ (_03560_, _03559_, _03399_);
  or _54375_ (_03561_, _03476_, p2_in[2]);
  or _54376_ (_03562_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _54377_ (_03563_, _03562_, _03561_);
  and _54378_ (_03564_, _03563_, _42212_);
  or _54379_ (_03565_, _03564_, _03560_);
  and _54380_ (_03566_, _03565_, _03351_);
  or _54381_ (_03567_, _03566_, _03556_);
  nor _54382_ (_03568_, _03476_, p2_in[0]);
  and _54383_ (_03569_, _03476_, _39376_);
  nor _54384_ (_03570_, _03569_, _03568_);
  or _54385_ (_03571_, _03570_, _03399_);
  nor _54386_ (_03572_, _03476_, p2_in[4]);
  and _54387_ (_03573_, _03476_, _39425_);
  nor _54388_ (_03574_, _03573_, _03572_);
  or _54389_ (_03575_, _03574_, _42212_);
  and _54390_ (_03576_, _03575_, _03361_);
  and _54391_ (_03577_, _03576_, _03571_);
  or _54392_ (_03578_, _03476_, p2_in[5]);
  or _54393_ (_03579_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _54394_ (_03580_, _03579_, _03578_);
  and _54395_ (_03581_, _03580_, _03399_);
  or _54396_ (_03582_, _03476_, p2_in[1]);
  or _54397_ (_03583_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _54398_ (_03584_, _03583_, _03582_);
  and _54399_ (_03585_, _03584_, _42212_);
  or _54400_ (_03586_, _03585_, _03581_);
  and _54401_ (_03587_, _03586_, _03348_);
  or _54402_ (_03588_, _03587_, _03577_);
  or _54403_ (_03589_, _03588_, _03567_);
  and _54404_ (_03590_, _03589_, _03340_);
  or _54405_ (_03591_, _03590_, _03546_);
  and _54406_ (_03592_, _03591_, _03524_);
  and _54407_ (_03593_, _03525_, _03460_);
  and _54408_ (_03594_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor _54409_ (_03595_, _42212_, _41017_);
  or _54410_ (_03596_, _03595_, _03594_);
  and _54411_ (_03597_, _03596_, _03358_);
  and _54412_ (_03598_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor _54413_ (_03599_, _42212_, _41443_);
  or _54414_ (_03600_, _03599_, _03598_);
  and _54415_ (_03601_, _03600_, _03348_);
  or _54416_ (_03602_, _03601_, _03597_);
  and _54417_ (_03603_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _54418_ (_03604_, _42212_, _41042_);
  or _54419_ (_03605_, _03604_, _03603_);
  and _54420_ (_03606_, _03605_, _03361_);
  and _54421_ (_03607_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _54422_ (_03608_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _54423_ (_03609_, _03608_, _03607_);
  and _54424_ (_03610_, _03609_, _03351_);
  or _54425_ (_03611_, _03610_, _03606_);
  or _54426_ (_03612_, _03611_, _03602_);
  and _54427_ (_03613_, _03612_, _03593_);
  nor _54428_ (_03614_, _03439_, _03371_);
  not _54429_ (_03615_, _03369_);
  nand _54430_ (_03616_, _03615_, _03340_);
  and _54431_ (_03617_, _42451_, _03338_);
  nand _54432_ (_03618_, _03617_, _42355_);
  and _54433_ (_03619_, _03618_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _54434_ (_03620_, _03619_, _03616_);
  and _54435_ (_03621_, _03620_, _03614_);
  and _54436_ (_03622_, _03524_, _03371_);
  or _54437_ (_03623_, _03476_, p3_in[3]);
  or _54438_ (_03624_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _54439_ (_03625_, _03624_, _03623_);
  or _54440_ (_03626_, _03625_, _03399_);
  or _54441_ (_03627_, _03476_, p3_in[7]);
  or _54442_ (_03628_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _54443_ (_03629_, _03628_, _03627_);
  or _54444_ (_03630_, _03629_, _42212_);
  and _54445_ (_03631_, _03630_, _03358_);
  and _54446_ (_03632_, _03631_, _03626_);
  or _54447_ (_03633_, _03476_, p3_in[5]);
  or _54448_ (_03634_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _54449_ (_03635_, _03634_, _03633_);
  and _54450_ (_03636_, _03635_, _03399_);
  or _54451_ (_03637_, _03476_, p3_in[1]);
  or _54452_ (_03638_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _54453_ (_03639_, _03638_, _03637_);
  and _54454_ (_03640_, _03639_, _42212_);
  or _54455_ (_03641_, _03640_, _03636_);
  and _54456_ (_03642_, _03641_, _03348_);
  or _54457_ (_03643_, _03642_, _03632_);
  nor _54458_ (_03644_, _03476_, p3_in[0]);
  and _54459_ (_03645_, _03476_, _39471_);
  nor _54460_ (_03646_, _03645_, _03644_);
  or _54461_ (_03647_, _03646_, _03399_);
  nor _54462_ (_03648_, _03476_, p3_in[4]);
  and _54463_ (_03649_, _03476_, _39520_);
  nor _54464_ (_03650_, _03649_, _03648_);
  or _54465_ (_03651_, _03650_, _42212_);
  and _54466_ (_03652_, _03651_, _03361_);
  and _54467_ (_03653_, _03652_, _03647_);
  or _54468_ (_03654_, _03476_, p3_in[6]);
  or _54469_ (_03655_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _54470_ (_03656_, _03655_, _03654_);
  and _54471_ (_03657_, _03656_, _03399_);
  or _54472_ (_03658_, _03476_, p3_in[2]);
  or _54473_ (_03659_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _54474_ (_03660_, _03659_, _03658_);
  and _54475_ (_03661_, _03660_, _42212_);
  or _54476_ (_03662_, _03661_, _03657_);
  and _54477_ (_03663_, _03662_, _03351_);
  or _54478_ (_03664_, _03663_, _03653_);
  or _54479_ (_03665_, _03664_, _03643_);
  and _54480_ (_03666_, _03665_, _03622_);
  or _54481_ (_03667_, _03666_, _03621_);
  or _54482_ (_03668_, _03667_, _03613_);
  or _54483_ (_03669_, _03668_, _03592_);
  or _54484_ (_03670_, _03669_, _03523_);
  and _54485_ (_03671_, _03339_, _42355_);
  and _54486_ (_03672_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nor _54487_ (_03673_, _42212_, _39713_);
  or _54488_ (_03674_, _03673_, _03672_);
  and _54489_ (_03675_, _03674_, _03361_);
  or _54490_ (_03676_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _54491_ (_03677_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _54492_ (_03678_, _03677_, _03358_);
  and _54493_ (_03679_, _03678_, _03676_);
  or _54494_ (_03680_, _03679_, _03675_);
  and _54495_ (_03681_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _54496_ (_03682_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _54497_ (_03683_, _03682_, _03681_);
  and _54498_ (_03684_, _03683_, _03348_);
  nand _54499_ (_03685_, _42212_, _40896_);
  or _54500_ (_03686_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _54501_ (_03687_, _03686_, _03351_);
  and _54502_ (_03688_, _03687_, _03685_);
  or _54503_ (_03689_, _03688_, _03684_);
  or _54504_ (_03690_, _03689_, _03680_);
  and _54505_ (_03691_, _03690_, _03460_);
  and _54506_ (_03692_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nor _54507_ (_03693_, _42212_, _40446_);
  or _54508_ (_03694_, _03693_, _03692_);
  and _54509_ (_03695_, _03694_, _03361_);
  or _54510_ (_03696_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _54511_ (_03697_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _54512_ (_03698_, _03697_, _03358_);
  and _54513_ (_03699_, _03698_, _03696_);
  or _54514_ (_03700_, _03699_, _03695_);
  and _54515_ (_03701_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nor _54516_ (_03702_, _42212_, _40450_);
  or _54517_ (_03703_, _03702_, _03701_);
  and _54518_ (_03704_, _03703_, _03348_);
  or _54519_ (_03705_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _54520_ (_03706_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _54521_ (_03707_, _03706_, _03351_);
  and _54522_ (_03708_, _03707_, _03705_);
  or _54523_ (_03709_, _03708_, _03704_);
  or _54524_ (_03710_, _03709_, _03700_);
  and _54525_ (_03711_, _03710_, _03524_);
  or _54526_ (_03712_, _03711_, _03691_);
  and _54527_ (_03713_, _03712_, _03671_);
  and _54528_ (_03714_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor _54529_ (_03715_, _42212_, _35273_);
  or _54530_ (_03716_, _03715_, _03714_);
  and _54531_ (_03717_, _03716_, _03361_);
  and _54532_ (_03718_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor _54533_ (_03719_, _42212_, _36078_);
  or _54534_ (_03720_, _03719_, _03718_);
  and _54535_ (_03721_, _03720_, _03348_);
  or _54536_ (_03722_, _03721_, _03717_);
  and _54537_ (_03723_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor _54538_ (_03724_, _42212_, _31233_);
  or _54539_ (_03725_, _03724_, _03723_);
  and _54540_ (_03726_, _03725_, _03358_);
  nor _54541_ (_03727_, _42212_, _36719_);
  and _54542_ (_03729_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _54543_ (_03730_, _03729_, _03727_);
  and _54544_ (_03731_, _03730_, _03351_);
  or _54545_ (_03732_, _03731_, _03726_);
  or _54546_ (_03733_, _03732_, _03722_);
  and _54547_ (_03734_, _03733_, _03337_);
  or _54548_ (_03735_, _03476_, p1_in[5]);
  or _54549_ (_03736_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _54550_ (_03737_, _03736_, _03735_);
  and _54551_ (_03738_, _03737_, _03399_);
  or _54552_ (_03739_, _03476_, p1_in[1]);
  or _54553_ (_03740_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _54554_ (_03741_, _03740_, _03739_);
  and _54555_ (_03742_, _03741_, _42212_);
  or _54556_ (_03743_, _03742_, _03738_);
  and _54557_ (_03744_, _03743_, _03348_);
  or _54558_ (_03745_, _03476_, p1_in[2]);
  or _54559_ (_03746_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _54560_ (_03747_, _03746_, _03745_);
  or _54561_ (_03748_, _03747_, _03399_);
  or _54562_ (_03749_, _03476_, p1_in[6]);
  or _54563_ (_03750_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _54564_ (_03751_, _03750_, _03749_);
  or _54565_ (_03752_, _03751_, _42212_);
  and _54566_ (_03753_, _03752_, _03351_);
  and _54567_ (_03754_, _03753_, _03748_);
  or _54568_ (_03755_, _03476_, p1_in[3]);
  or _54569_ (_03756_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _54570_ (_03757_, _03756_, _03755_);
  or _54571_ (_03758_, _03757_, _03399_);
  or _54572_ (_03759_, _03476_, p1_in[7]);
  or _54573_ (_03760_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _54574_ (_03761_, _03760_, _03759_);
  or _54575_ (_03762_, _03761_, _42212_);
  and _54576_ (_03763_, _03762_, _03358_);
  and _54577_ (_03764_, _03763_, _03758_);
  nor _54578_ (_03765_, _03476_, p1_in[0]);
  and _54579_ (_03766_, _03476_, _39294_);
  nor _54580_ (_03767_, _03766_, _03765_);
  or _54581_ (_03768_, _03767_, _03399_);
  nor _54582_ (_03769_, _03476_, p1_in[4]);
  and _54583_ (_03770_, _03476_, _39343_);
  nor _54584_ (_03771_, _03770_, _03769_);
  or _54585_ (_03772_, _03771_, _42212_);
  and _54586_ (_03773_, _03772_, _03361_);
  and _54587_ (_03774_, _03773_, _03768_);
  or _54588_ (_03775_, _03774_, _03764_);
  or _54589_ (_03776_, _03775_, _03754_);
  or _54590_ (_03777_, _03776_, _03744_);
  and _54591_ (_03778_, _03777_, _03460_);
  or _54592_ (_03779_, _03778_, _03734_);
  and _54593_ (_03780_, _03779_, _03371_);
  or _54594_ (_03781_, _03780_, _03713_);
  or _54595_ (_03782_, _03781_, _03670_);
  or _54596_ (_03783_, _03782_, _03415_);
  nand _54597_ (_03784_, _03416_, _31757_);
  and _54598_ (_03785_, _03784_, _03343_);
  and _54599_ (_03786_, _03785_, _03783_);
  or _54600_ (_03787_, _03786_, _03368_);
  and _54601_ (_39682_, _03787_, _42618_);
  and _54602_ (_03788_, _42354_, _42212_);
  and _54603_ (_03789_, _03788_, _03361_);
  and _54604_ (_03790_, _03339_, _03337_);
  and _54605_ (_03791_, _03790_, _03789_);
  and _54606_ (_03792_, _03791_, _38785_);
  and _54607_ (_03793_, _03358_, _03399_);
  not _54608_ (_03794_, _03793_);
  and _54609_ (_03795_, _03794_, _38795_);
  and _54610_ (_03796_, _03795_, _01374_);
  nor _54611_ (_03797_, _03796_, _03792_);
  and _54612_ (_03798_, _03797_, _01390_);
  and _54613_ (_03799_, _03460_, _03339_);
  and _54614_ (_03800_, _03788_, _03358_);
  and _54615_ (_03801_, _03800_, _03799_);
  and _54616_ (_03802_, _03801_, _38276_);
  not _54617_ (_03803_, _03802_);
  and _54618_ (_03804_, _03791_, _38782_);
  nor _54619_ (_03805_, _42451_, _42100_);
  and _54620_ (_03806_, _42260_, _42164_);
  and _54621_ (_03807_, _03806_, _03805_);
  and _54622_ (_03808_, _03807_, _03789_);
  and _54623_ (_03809_, _03808_, _38624_);
  nor _54624_ (_03810_, _03809_, _03804_);
  and _54625_ (_03811_, _03810_, _03803_);
  nor _54626_ (_03812_, _03811_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _54627_ (_03813_, _03812_);
  and _54628_ (_03814_, _03813_, _03798_);
  and _54629_ (_03815_, _03788_, _03351_);
  and _54630_ (_03816_, _03815_, _03799_);
  and _54631_ (_03817_, _03816_, _38276_);
  or _54632_ (_03818_, _03817_, rst);
  nor _54633_ (_39683_, _03818_, _03814_);
  nand _54634_ (_03819_, _03817_, _31136_);
  and _54635_ (_03820_, _42355_, _42212_);
  and _54636_ (_03821_, _03820_, _03358_);
  and _54637_ (_03822_, _03821_, _03438_);
  and _54638_ (_03823_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _54639_ (_03824_, _03820_, _03361_);
  and _54640_ (_03825_, _03824_, _03799_);
  and _54641_ (_03826_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _54642_ (_03827_, _03826_, _03823_);
  and _54643_ (_03828_, _03524_, _03339_);
  and _54644_ (_03829_, _03828_, _03824_);
  and _54645_ (_03830_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _54646_ (_03831_, _03793_, _42354_);
  nor _54647_ (_03832_, _42259_, _42164_);
  and _54648_ (_03833_, _03832_, _03617_);
  and _54649_ (_03834_, _03833_, _03831_);
  and _54650_ (_03835_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _54651_ (_03836_, _03835_, _03830_);
  or _54652_ (_03837_, _03836_, _03827_);
  nor _54653_ (_03838_, _42354_, _42212_);
  and _54654_ (_03839_, _03838_, _03361_);
  and _54655_ (_03840_, _03839_, _03438_);
  and _54656_ (_03841_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _54657_ (_03842_, _03824_, _03438_);
  and _54658_ (_03843_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _54659_ (_03844_, _03843_, _03841_);
  and _54660_ (_03845_, _03838_, _03348_);
  and _54661_ (_03846_, _03845_, _03438_);
  and _54662_ (_03847_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _54663_ (_03848_, _03820_, _03351_);
  and _54664_ (_03849_, _03848_, _03438_);
  and _54665_ (_03850_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _54666_ (_03851_, _03850_, _03847_);
  or _54667_ (_03852_, _03851_, _03844_);
  or _54668_ (_03853_, _03852_, _03837_);
  and _54669_ (_03854_, _03460_, _03370_);
  and _54670_ (_03855_, _03820_, _03348_);
  and _54671_ (_03856_, _03855_, _03854_);
  and _54672_ (_03857_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _54673_ (_03858_, _03854_, _03824_);
  and _54674_ (_03859_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _54675_ (_03860_, _03859_, _03857_);
  and _54676_ (_03861_, _03839_, _03799_);
  and _54677_ (_03862_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _54678_ (_03863_, _03831_, _03799_);
  and _54679_ (_03864_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _54680_ (_03865_, _03864_, _03862_);
  or _54681_ (_03866_, _03865_, _03860_);
  and _54682_ (_03867_, _03821_, _03799_);
  and _54683_ (_03868_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _54684_ (_03869_, _03855_, _03799_);
  and _54685_ (_03870_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _54686_ (_03871_, _03870_, _03868_);
  and _54687_ (_03872_, _03845_, _03799_);
  and _54688_ (_03873_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _54689_ (_03874_, _03848_, _03799_);
  and _54690_ (_03875_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _54691_ (_03876_, _03875_, _03873_);
  or _54692_ (_03877_, _03876_, _03871_);
  or _54693_ (_03878_, _03877_, _03866_);
  or _54694_ (_03879_, _03878_, _03853_);
  and _54695_ (_03880_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _54696_ (_03881_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or _54697_ (_03882_, _03881_, _03880_);
  and _54698_ (_03883_, _03832_, _03805_);
  and _54699_ (_03884_, _03883_, _03789_);
  and _54700_ (_03885_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _54701_ (_03886_, _03788_, _03348_);
  and _54702_ (_03887_, _03886_, _03799_);
  and _54703_ (_03888_, _03887_, _38227_);
  or _54704_ (_03889_, _03888_, _03885_);
  or _54705_ (_03890_, _03889_, _03882_);
  and _54706_ (_03891_, _03828_, _03789_);
  and _54707_ (_03892_, _03891_, _03553_);
  and _54708_ (_03893_, _03833_, _03789_);
  and _54709_ (_03894_, _03893_, _03629_);
  or _54710_ (_03895_, _03894_, _03892_);
  and _54711_ (_03896_, _03799_, _03789_);
  and _54712_ (_03897_, _03896_, _03494_);
  and _54713_ (_03898_, _03854_, _03789_);
  and _54714_ (_03899_, _03898_, _03761_);
  or _54715_ (_03900_, _03899_, _03897_);
  or _54716_ (_03901_, _03900_, _03895_);
  or _54717_ (_03902_, _03901_, _03890_);
  and _54718_ (_03903_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _54719_ (_03904_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _54720_ (_03905_, _03904_, _03903_);
  or _54721_ (_03906_, _03905_, _03902_);
  or _54722_ (_03907_, _03906_, _03879_);
  and _54723_ (_03908_, _03907_, _03814_);
  not _54724_ (_03909_, _03814_);
  nor _54725_ (_03910_, _03842_, _03840_);
  nor _54726_ (_03911_, _03849_, _03846_);
  and _54727_ (_03912_, _03911_, _03910_);
  nor _54728_ (_03913_, _03825_, _03822_);
  nor _54729_ (_03914_, _03834_, _03829_);
  and _54730_ (_03915_, _03914_, _03913_);
  and _54731_ (_03916_, _03915_, _03912_);
  nor _54732_ (_03917_, _03869_, _03867_);
  nor _54733_ (_03918_, _03874_, _03872_);
  and _54734_ (_03919_, _03918_, _03917_);
  nor _54735_ (_03920_, _03863_, _03861_);
  nor _54736_ (_03921_, _03858_, _03856_);
  and _54737_ (_03922_, _03921_, _03920_);
  and _54738_ (_03923_, _03922_, _03919_);
  and _54739_ (_03924_, _03923_, _03916_);
  nor _54740_ (_03925_, _03816_, _03801_);
  nor _54741_ (_03926_, _03887_, _03884_);
  and _54742_ (_03928_, _03926_, _03925_);
  nor _54743_ (_03929_, _03893_, _03891_);
  nor _54744_ (_03930_, _03898_, _03896_);
  and _54745_ (_03931_, _03930_, _03929_);
  and _54746_ (_03932_, _03931_, _03928_);
  nor _54747_ (_03933_, _03808_, _03791_);
  and _54748_ (_03934_, _03933_, _03932_);
  and _54749_ (_03935_, _03934_, _03924_);
  or _54750_ (_03936_, _03935_, _03909_);
  and _54751_ (_03937_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _54752_ (_03938_, _03937_, _03908_);
  or _54753_ (_03939_, _03938_, _03817_);
  and _54754_ (_03940_, _03939_, _42618_);
  and _54755_ (_39684_, _03940_, _03819_);
  nor _54756_ (_39764_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _54757_ (_03941_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _54758_ (_03942_, _03330_, rst);
  and _54759_ (_39765_, _03942_, _03941_);
  nor _54760_ (_03943_, _03330_, _03329_);
  or _54761_ (_03944_, _03943_, _03331_);
  and _54762_ (_03945_, _03334_, _42618_);
  and _54763_ (_39766_, _03945_, _03944_);
  nand _54764_ (_03946_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _54765_ (_03947_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _54766_ (_03948_, _03947_, _03946_);
  nand _54767_ (_03949_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _54768_ (_03950_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _54769_ (_03951_, _03950_, _03949_);
  and _54770_ (_03952_, _03951_, _03948_);
  nand _54771_ (_03953_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _54772_ (_03954_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _54773_ (_03955_, _03954_, _03953_);
  nand _54774_ (_03956_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _54775_ (_03957_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _54776_ (_03958_, _03957_, _03956_);
  and _54777_ (_03959_, _03958_, _03955_);
  and _54778_ (_03960_, _03959_, _03952_);
  nand _54779_ (_03961_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand _54780_ (_03962_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _54781_ (_03963_, _03962_, _03961_);
  nand _54782_ (_03964_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _54783_ (_03965_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _54784_ (_03966_, _03965_, _03964_);
  and _54785_ (_03967_, _03966_, _03963_);
  nand _54786_ (_03968_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _54787_ (_03969_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _54788_ (_03970_, _03969_, _03968_);
  nand _54789_ (_03971_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand _54790_ (_03972_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _54791_ (_03973_, _03972_, _03971_);
  and _54792_ (_03974_, _03973_, _03970_);
  and _54793_ (_03975_, _03974_, _03967_);
  and _54794_ (_03976_, _03975_, _03960_);
  nand _54795_ (_03977_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _54796_ (_03978_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _54797_ (_03979_, _03978_, _03977_);
  nand _54798_ (_03980_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _54799_ (_03981_, _03887_, _42395_);
  and _54800_ (_03982_, _03981_, _03980_);
  and _54801_ (_03983_, _03982_, _03979_);
  nand _54802_ (_03984_, _03891_, _03570_);
  nand _54803_ (_03985_, _03893_, _03646_);
  and _54804_ (_03986_, _03985_, _03984_);
  nand _54805_ (_03987_, _03898_, _03767_);
  nand _54806_ (_03988_, _03896_, _03479_);
  and _54807_ (_03989_, _03988_, _03987_);
  and _54808_ (_03990_, _03989_, _03986_);
  and _54809_ (_03991_, _03990_, _03983_);
  not _54810_ (_03992_, _03808_);
  or _54811_ (_03993_, _03992_, _03394_);
  nand _54812_ (_03994_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _54813_ (_03995_, _03994_, _03993_);
  and _54814_ (_03996_, _03995_, _03991_);
  and _54815_ (_03997_, _03996_, _03976_);
  nor _54816_ (_03998_, _03997_, _03909_);
  not _54817_ (_03999_, _03817_);
  nand _54818_ (_04000_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _54819_ (_04001_, _04000_, _03999_);
  or _54820_ (_04002_, _04001_, _03998_);
  nand _54821_ (_04003_, _03817_, _32323_);
  and _54822_ (_04004_, _04003_, _42618_);
  and _54823_ (_39768_, _04004_, _04002_);
  nand _54824_ (_04005_, _03817_, _33020_);
  or _54825_ (_04006_, _03798_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _54826_ (_04007_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _54827_ (_04008_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _54828_ (_04009_, _04008_, _04007_);
  and _54829_ (_04010_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _54830_ (_04011_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _54831_ (_04012_, _04011_, _04010_);
  or _54832_ (_04013_, _04012_, _04009_);
  and _54833_ (_04014_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _54834_ (_04015_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _54835_ (_04016_, _04015_, _04014_);
  and _54836_ (_04017_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _54837_ (_04018_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _54838_ (_04019_, _04018_, _04017_);
  or _54839_ (_04020_, _04019_, _04016_);
  or _54840_ (_04021_, _04020_, _04013_);
  and _54841_ (_04022_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _54842_ (_04024_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _54843_ (_04025_, _04024_, _04022_);
  and _54844_ (_04026_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _54845_ (_04027_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _54846_ (_04028_, _04027_, _04026_);
  or _54847_ (_04029_, _04028_, _04025_);
  and _54848_ (_04030_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _54849_ (_04031_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _54850_ (_04032_, _04031_, _04030_);
  and _54851_ (_04033_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _54852_ (_04034_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _54853_ (_04035_, _04034_, _04033_);
  or _54854_ (_04036_, _04035_, _04032_);
  or _54855_ (_04037_, _04036_, _04029_);
  or _54856_ (_04038_, _04037_, _04021_);
  and _54857_ (_04039_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _54858_ (_04040_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or _54859_ (_04041_, _04040_, _04039_);
  and _54860_ (_04042_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _54861_ (_04043_, _03887_, _42302_);
  or _54862_ (_04044_, _04043_, _04042_);
  or _54863_ (_04045_, _04044_, _04041_);
  and _54864_ (_04046_, _03891_, _03584_);
  and _54865_ (_04047_, _03893_, _03639_);
  or _54866_ (_04048_, _04047_, _04046_);
  and _54867_ (_04049_, _03896_, _03505_);
  and _54868_ (_04050_, _03898_, _03741_);
  or _54869_ (_04051_, _04050_, _04049_);
  or _54870_ (_04052_, _04051_, _04048_);
  or _54871_ (_04053_, _04052_, _04045_);
  and _54872_ (_04054_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _54873_ (_04055_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _54874_ (_04056_, _04055_, _04054_);
  or _54875_ (_04057_, _04056_, _04053_);
  or _54876_ (_04058_, _04057_, _04038_);
  and _54877_ (_04059_, _04058_, _03813_);
  and _54878_ (_04060_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or _54879_ (_04061_, _04060_, _04059_);
  and _54880_ (_04062_, _04061_, _04006_);
  or _54881_ (_04063_, _04062_, _03817_);
  and _54882_ (_04064_, _04063_, _42618_);
  and _54883_ (_39769_, _04064_, _04005_);
  nand _54884_ (_04065_, _03817_, _33717_);
  or _54885_ (_04066_, _03798_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _54886_ (_04067_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _54887_ (_04068_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _54888_ (_04069_, _04068_, _04067_);
  and _54889_ (_04070_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _54890_ (_04071_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _54891_ (_04072_, _04071_, _04070_);
  or _54892_ (_04073_, _04072_, _04069_);
  and _54893_ (_04074_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _54894_ (_04075_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or _54895_ (_04076_, _04075_, _04074_);
  and _54896_ (_04077_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _54897_ (_04078_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _54898_ (_04079_, _04078_, _04077_);
  or _54899_ (_04080_, _04079_, _04076_);
  or _54900_ (_04081_, _04080_, _04073_);
  and _54901_ (_04082_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _54902_ (_04083_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _54903_ (_04084_, _04083_, _04082_);
  and _54904_ (_04085_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _54905_ (_04086_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _54906_ (_04087_, _04086_, _04085_);
  or _54907_ (_04088_, _04087_, _04084_);
  and _54908_ (_04089_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _54909_ (_04090_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _54910_ (_04091_, _04090_, _04089_);
  and _54911_ (_04092_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _54912_ (_04093_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _54913_ (_04094_, _04093_, _04092_);
  or _54914_ (_04095_, _04094_, _04091_);
  or _54915_ (_04096_, _04095_, _04088_);
  or _54916_ (_04097_, _04096_, _04081_);
  and _54917_ (_04098_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _54918_ (_04099_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or _54919_ (_04100_, _04099_, _04098_);
  and _54920_ (_04101_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _54921_ (_04102_, _03887_, _42192_);
  or _54922_ (_04103_, _04102_, _04101_);
  or _54923_ (_04104_, _04103_, _04100_);
  and _54924_ (_04105_, _03891_, _03563_);
  and _54925_ (_04106_, _03893_, _03660_);
  or _54926_ (_04107_, _04106_, _04105_);
  and _54927_ (_04108_, _03898_, _03747_);
  and _54928_ (_04109_, _03896_, _03511_);
  or _54929_ (_04110_, _04109_, _04108_);
  or _54930_ (_04111_, _04110_, _04107_);
  or _54931_ (_04112_, _04111_, _04104_);
  and _54932_ (_04113_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _54933_ (_04114_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _54934_ (_04115_, _04114_, _04113_);
  or _54935_ (_04116_, _04115_, _04112_);
  or _54936_ (_04117_, _04116_, _04097_);
  and _54937_ (_04118_, _04117_, _03813_);
  and _54938_ (_04119_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or _54939_ (_04120_, _04119_, _04118_);
  and _54940_ (_04121_, _04120_, _04066_);
  or _54941_ (_04122_, _04121_, _03817_);
  and _54942_ (_04124_, _04122_, _42618_);
  and _54943_ (_39770_, _04124_, _04065_);
  nand _54944_ (_04125_, _03817_, _34478_);
  and _54945_ (_04126_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _54946_ (_04127_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _54947_ (_04128_, _04127_, _04126_);
  and _54948_ (_04129_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _54949_ (_04130_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _54950_ (_04131_, _04130_, _04129_);
  or _54951_ (_04132_, _04131_, _04128_);
  and _54952_ (_04133_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _54953_ (_04134_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _54954_ (_04135_, _04134_, _04133_);
  and _54955_ (_04136_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _54956_ (_04137_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _54957_ (_04138_, _04137_, _04136_);
  or _54958_ (_04139_, _04138_, _04135_);
  or _54959_ (_04140_, _04139_, _04132_);
  and _54960_ (_04141_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _54961_ (_04142_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or _54962_ (_04143_, _04142_, _04141_);
  and _54963_ (_04144_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _54964_ (_04145_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _54965_ (_04146_, _04145_, _04144_);
  or _54966_ (_04147_, _04146_, _04143_);
  and _54967_ (_04148_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _54968_ (_04149_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _54969_ (_04150_, _04149_, _04148_);
  and _54970_ (_04151_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _54971_ (_04152_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or _54972_ (_04153_, _04152_, _04151_);
  or _54973_ (_04154_, _04153_, _04150_);
  or _54974_ (_04155_, _04154_, _04147_);
  or _54975_ (_04156_, _04155_, _04140_);
  and _54976_ (_04157_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _54977_ (_04158_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _54978_ (_04159_, _04158_, _04157_);
  and _54979_ (_04160_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _54980_ (_04161_, _03887_, _42331_);
  or _54981_ (_04162_, _04161_, _04160_);
  or _54982_ (_04163_, _04162_, _04159_);
  and _54983_ (_04164_, _03891_, _03549_);
  and _54984_ (_04165_, _03893_, _03625_);
  or _54985_ (_04166_, _04165_, _04164_);
  and _54986_ (_04167_, _03896_, _03490_);
  and _54987_ (_04168_, _03898_, _03757_);
  or _54988_ (_04169_, _04168_, _04167_);
  or _54989_ (_04170_, _04169_, _04166_);
  or _54990_ (_04171_, _04170_, _04163_);
  and _54991_ (_04172_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _54992_ (_04173_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _54993_ (_04174_, _04173_, _04172_);
  or _54994_ (_04175_, _04174_, _04171_);
  or _54995_ (_04176_, _04175_, _04156_);
  and _54996_ (_04177_, _04176_, _03814_);
  and _54997_ (_04178_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or _54998_ (_04179_, _04178_, _04177_);
  or _54999_ (_04180_, _04179_, _03817_);
  and _55000_ (_04181_, _04180_, _42618_);
  and _55001_ (_39771_, _04181_, _04125_);
  nand _55002_ (_04182_, _03817_, _35240_);
  nand _55003_ (_04183_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand _55004_ (_04184_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _55005_ (_04185_, _04184_, _04183_);
  nand _55006_ (_04186_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand _55007_ (_04187_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _55008_ (_04188_, _04187_, _04186_);
  and _55009_ (_04189_, _04188_, _04185_);
  nand _55010_ (_04190_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nand _55011_ (_04191_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _55012_ (_04192_, _04191_, _04190_);
  nand _55013_ (_04193_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _55014_ (_04194_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _55015_ (_04195_, _04194_, _04193_);
  and _55016_ (_04196_, _04195_, _04192_);
  and _55017_ (_04197_, _04196_, _04189_);
  nand _55018_ (_04198_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand _55019_ (_04199_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _55020_ (_04200_, _04199_, _04198_);
  nand _55021_ (_04201_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _55022_ (_04202_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _55023_ (_04203_, _04202_, _04201_);
  and _55024_ (_04204_, _04203_, _04200_);
  nand _55025_ (_04205_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand _55026_ (_04206_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and _55027_ (_04207_, _04206_, _04205_);
  nand _55028_ (_04208_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _55029_ (_04209_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _55030_ (_04210_, _04209_, _04208_);
  and _55031_ (_04211_, _04210_, _04207_);
  and _55032_ (_04212_, _04211_, _04204_);
  and _55033_ (_04213_, _04212_, _04197_);
  nand _55034_ (_04214_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand _55035_ (_04215_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _55036_ (_04216_, _04215_, _04214_);
  nand _55037_ (_04217_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _55038_ (_04218_, _03887_, _42237_);
  and _55039_ (_04219_, _04218_, _04217_);
  and _55040_ (_04220_, _04219_, _04216_);
  nand _55041_ (_04221_, _03891_, _03574_);
  nand _55042_ (_04223_, _03893_, _03650_);
  and _55043_ (_04224_, _04223_, _04221_);
  nand _55044_ (_04225_, _03896_, _03483_);
  nand _55045_ (_04226_, _03898_, _03771_);
  and _55046_ (_04227_, _04226_, _04225_);
  and _55047_ (_04228_, _04227_, _04224_);
  and _55048_ (_04229_, _04228_, _04220_);
  nand _55049_ (_04230_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _55050_ (_04231_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _55051_ (_04232_, _04231_, _04230_);
  and _55052_ (_04233_, _04232_, _04229_);
  nand _55053_ (_04234_, _04233_, _04213_);
  and _55054_ (_04235_, _04234_, _03814_);
  and _55055_ (_04236_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or _55056_ (_04237_, _04236_, _03817_);
  or _55057_ (_04238_, _04237_, _04235_);
  and _55058_ (_04239_, _04238_, _42618_);
  and _55059_ (_39772_, _04239_, _04182_);
  nand _55060_ (_04240_, _03817_, _36046_);
  and _55061_ (_04241_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _55062_ (_04242_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _55063_ (_04243_, _04242_, _04241_);
  and _55064_ (_04244_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _55065_ (_04245_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _55066_ (_04246_, _04245_, _04244_);
  or _55067_ (_04247_, _04246_, _04243_);
  and _55068_ (_04248_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _55069_ (_04249_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _55070_ (_04250_, _04249_, _04248_);
  and _55071_ (_04251_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _55072_ (_04252_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _55073_ (_04253_, _04252_, _04251_);
  or _55074_ (_04254_, _04253_, _04250_);
  or _55075_ (_04255_, _04254_, _04247_);
  and _55076_ (_04256_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _55077_ (_04257_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or _55078_ (_04258_, _04257_, _04256_);
  and _55079_ (_04259_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _55080_ (_04260_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _55081_ (_04261_, _04260_, _04259_);
  or _55082_ (_04262_, _04261_, _04258_);
  and _55083_ (_04263_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _55084_ (_04264_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _55085_ (_04265_, _04264_, _04263_);
  and _55086_ (_04266_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _55087_ (_04267_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _55088_ (_04268_, _04267_, _04266_);
  or _55089_ (_04269_, _04268_, _04265_);
  or _55090_ (_04270_, _04269_, _04262_);
  or _55091_ (_04271_, _04270_, _04255_);
  and _55092_ (_04272_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _55093_ (_04273_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or _55094_ (_04274_, _04273_, _04272_);
  and _55095_ (_04275_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _55096_ (_04276_, _03887_, _42137_);
  or _55097_ (_04277_, _04276_, _04275_);
  or _55098_ (_04278_, _04277_, _04274_);
  and _55099_ (_04279_, _03891_, _03580_);
  and _55100_ (_04280_, _03893_, _03635_);
  or _55101_ (_04281_, _04280_, _04279_);
  and _55102_ (_04282_, _03898_, _03737_);
  and _55103_ (_04283_, _03896_, _03501_);
  or _55104_ (_04284_, _04283_, _04282_);
  or _55105_ (_04285_, _04284_, _04281_);
  or _55106_ (_04286_, _04285_, _04278_);
  and _55107_ (_04287_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _55108_ (_04288_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _55109_ (_04289_, _04288_, _04287_);
  or _55110_ (_04290_, _04289_, _04286_);
  or _55111_ (_04291_, _04290_, _04271_);
  and _55112_ (_04292_, _04291_, _03814_);
  and _55113_ (_04293_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or _55114_ (_04294_, _04293_, _04292_);
  or _55115_ (_04295_, _04294_, _03817_);
  and _55116_ (_04296_, _04295_, _42618_);
  and _55117_ (_39773_, _04296_, _04240_);
  and _55118_ (_04297_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _55119_ (_04298_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _55120_ (_04299_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _55121_ (_04300_, _04299_, _04298_);
  and _55122_ (_04301_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _55123_ (_04302_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _55124_ (_04303_, _04302_, _04301_);
  or _55125_ (_04304_, _04303_, _04300_);
  and _55126_ (_04305_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _55127_ (_04306_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or _55128_ (_04307_, _04306_, _04305_);
  and _55129_ (_04308_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _55130_ (_04309_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _55131_ (_04310_, _04309_, _04308_);
  or _55132_ (_04311_, _04310_, _04307_);
  or _55133_ (_04312_, _04311_, _04304_);
  and _55134_ (_04313_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _55135_ (_04314_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _55136_ (_04315_, _04314_, _04313_);
  and _55137_ (_04316_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _55138_ (_04317_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _55139_ (_04318_, _04317_, _04316_);
  or _55140_ (_04319_, _04318_, _04315_);
  and _55141_ (_04320_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _55142_ (_04322_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _55143_ (_04323_, _04322_, _04320_);
  and _55144_ (_04324_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _55145_ (_04325_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _55146_ (_04326_, _04325_, _04324_);
  or _55147_ (_04327_, _04326_, _04323_);
  or _55148_ (_04328_, _04327_, _04319_);
  or _55149_ (_04329_, _04328_, _04312_);
  and _55150_ (_04330_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _55151_ (_04331_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or _55152_ (_04332_, _04331_, _04330_);
  and _55153_ (_04333_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _55154_ (_04334_, _03887_, _42408_);
  or _55155_ (_04335_, _04334_, _04333_);
  or _55156_ (_04336_, _04335_, _04332_);
  and _55157_ (_04337_, _03891_, _03559_);
  and _55158_ (_04338_, _03893_, _03656_);
  or _55159_ (_04339_, _04338_, _04337_);
  and _55160_ (_04340_, _03896_, _03515_);
  and _55161_ (_04341_, _03898_, _03751_);
  or _55162_ (_04342_, _04341_, _04340_);
  or _55163_ (_04343_, _04342_, _04339_);
  or _55164_ (_04344_, _04343_, _04336_);
  and _55165_ (_04345_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _55166_ (_04346_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _55167_ (_04347_, _04346_, _04345_);
  or _55168_ (_04348_, _04347_, _04344_);
  or _55169_ (_04349_, _04348_, _04329_);
  and _55170_ (_04350_, _04349_, _03814_);
  or _55171_ (_04351_, _04350_, _04297_);
  and _55172_ (_04352_, _04351_, _03999_);
  and _55173_ (_04353_, _03817_, _36698_);
  or _55174_ (_04354_, _04353_, _04352_);
  and _55175_ (_39774_, _04354_, _42618_);
  and _55176_ (_39843_, _42558_, _42618_);
  nor _55177_ (_39846_, _42212_, rst);
  and _55178_ (_39867_, _42648_, _42618_);
  and _55179_ (_39868_, _42658_, _42618_);
  nor _55180_ (_39871_, _42400_, rst);
  nor _55181_ (_39872_, _42307_, rst);
  not _55182_ (_04355_, _00342_);
  nor _55183_ (_04356_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _55184_ (_04357_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55185_ (_04358_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04357_);
  nor _55186_ (_04359_, _04358_, _04356_);
  nor _55187_ (_04360_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55188_ (_04361_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04357_);
  nor _55189_ (_04362_, _04361_, _04360_);
  nor _55190_ (_04363_, _04362_, _04359_);
  and _55191_ (_04364_, _04362_, _04359_);
  nor _55192_ (_04365_, _02227_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55193_ (_04366_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04357_);
  nor _55194_ (_04367_, _04366_, _04365_);
  and _55195_ (_04368_, _04367_, _04364_);
  nor _55196_ (_04369_, _04367_, _04364_);
  nor _55197_ (_04370_, _04369_, _04368_);
  nor _55198_ (_04371_, _02246_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55199_ (_04372_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04357_);
  nor _55200_ (_04373_, _04372_, _04371_);
  not _55201_ (_04374_, _04373_);
  and _55202_ (_04375_, _04374_, _04368_);
  nor _55203_ (_04376_, _04374_, _04368_);
  nor _55204_ (_04377_, _04376_, _04375_);
  nor _55205_ (_04378_, _04377_, _04370_);
  and _55206_ (_04379_, _04378_, _04363_);
  and _55207_ (_04380_, _04379_, _04355_);
  not _55208_ (_04381_, _43516_);
  not _55209_ (_04382_, _04370_);
  and _55210_ (_04383_, _04377_, _04382_);
  and _55211_ (_04384_, _04383_, _04363_);
  and _55212_ (_04385_, _04384_, _04381_);
  or _55213_ (_04386_, _04385_, _04380_);
  not _55214_ (_04387_, _00424_);
  not _55215_ (_04388_, _04359_);
  and _55216_ (_04389_, _04362_, _04388_);
  and _55217_ (_04390_, _04378_, _04389_);
  and _55218_ (_04391_, _04390_, _04387_);
  not _55219_ (_04392_, _00065_);
  and _55220_ (_04393_, _04383_, _04389_);
  and _55221_ (_04394_, _04393_, _04392_);
  or _55222_ (_04395_, _04394_, _04391_);
  or _55223_ (_04396_, _04395_, _04386_);
  not _55224_ (_04397_, _00168_);
  and _55225_ (_04398_, _04374_, _04370_);
  and _55226_ (_04399_, _04398_, _04363_);
  and _55227_ (_04400_, _04399_, _04397_);
  not _55228_ (_04401_, _00550_);
  nor _55229_ (_04402_, _04362_, _04388_);
  and _55230_ (_04403_, _04373_, _04370_);
  and _55231_ (_04404_, _04403_, _04402_);
  and _55232_ (_04405_, _04404_, _04401_);
  not _55233_ (_04406_, _00106_);
  and _55234_ (_04407_, _04398_, _04364_);
  and _55235_ (_04408_, _04407_, _04406_);
  or _55236_ (_04409_, _04408_, _04405_);
  or _55237_ (_04410_, _04409_, _04400_);
  not _55238_ (_04411_, _00465_);
  and _55239_ (_04412_, _04376_, _04364_);
  and _55240_ (_04413_, _04412_, _04411_);
  not _55241_ (_04415_, _00260_);
  and _55242_ (_04416_, _04367_, _04389_);
  and _55243_ (_04417_, _04416_, _04374_);
  and _55244_ (_04418_, _04417_, _04415_);
  not _55245_ (_04419_, _43475_);
  and _55246_ (_04420_, _04373_, _04368_);
  and _55247_ (_04421_, _04420_, _04419_);
  or _55248_ (_04422_, _04421_, _04418_);
  not _55249_ (_04423_, _00607_);
  and _55250_ (_04424_, _04416_, _04373_);
  and _55251_ (_04425_, _04424_, _04423_);
  not _55252_ (_04426_, _00301_);
  and _55253_ (_04427_, _04375_, _04426_);
  or _55254_ (_04428_, _04427_, _04425_);
  or _55255_ (_04429_, _04428_, _04422_);
  or _55256_ (_04430_, _04429_, _04413_);
  not _55257_ (_04431_, _00506_);
  and _55258_ (_04432_, _04403_, _04363_);
  and _55259_ (_04433_, _04432_, _04431_);
  not _55260_ (_04434_, _00219_);
  and _55261_ (_04435_, _04398_, _04402_);
  and _55262_ (_04436_, _04435_, _04434_);
  or _55263_ (_04437_, _04436_, _04433_);
  or _55264_ (_04438_, _04437_, _04430_);
  not _55265_ (_04439_, _00383_);
  and _55266_ (_04440_, _04378_, _04402_);
  and _55267_ (_04441_, _04440_, _04439_);
  not _55268_ (_04442_, _00024_);
  and _55269_ (_04443_, _04383_, _04402_);
  and _55270_ (_04444_, _04443_, _04442_);
  or _55271_ (_04445_, _04444_, _04441_);
  or _55272_ (_04446_, _04445_, _04438_);
  or _55273_ (_04447_, _04446_, _04410_);
  or _55274_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04447_, _04396_);
  and _55275_ (_04448_, _04393_, _04406_);
  and _55276_ (_04449_, _04384_, _04442_);
  or _55277_ (_04450_, _04449_, _04448_);
  and _55278_ (_04451_, _04440_, _04387_);
  and _55279_ (_04452_, _04443_, _04392_);
  or _55280_ (_04453_, _04452_, _04451_);
  or _55281_ (_04454_, _04453_, _04450_);
  and _55282_ (_04455_, _04404_, _04423_);
  and _55283_ (_04456_, _04432_, _04401_);
  and _55284_ (_04457_, _04435_, _04415_);
  or _55285_ (_04458_, _04457_, _04456_);
  or _55286_ (_04459_, _04458_, _04455_);
  and _55287_ (_04460_, _04407_, _04397_);
  and _55288_ (_04461_, _04399_, _04434_);
  or _55289_ (_04462_, _04461_, _04460_);
  and _55290_ (_04463_, _04412_, _04431_);
  and _55291_ (_04464_, _04375_, _04355_);
  and _55292_ (_04465_, _04424_, _04419_);
  or _55293_ (_04466_, _04465_, _04464_);
  and _55294_ (_04467_, _04417_, _04426_);
  and _55295_ (_04468_, _04420_, _04381_);
  or _55296_ (_04469_, _04468_, _04467_);
  or _55297_ (_04470_, _04469_, _04466_);
  or _55298_ (_04471_, _04470_, _04463_);
  or _55299_ (_04472_, _04471_, _04462_);
  and _55300_ (_04473_, _04390_, _04411_);
  and _55301_ (_04474_, _04379_, _04439_);
  or _55302_ (_04475_, _04474_, _04473_);
  or _55303_ (_04476_, _04475_, _04472_);
  or _55304_ (_04477_, _04476_, _04459_);
  or _55305_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04477_, _04454_);
  and _55306_ (_04478_, _04379_, _04387_);
  and _55307_ (_04479_, _04384_, _04392_);
  or _55308_ (_04480_, _04479_, _04478_);
  and _55309_ (_04481_, _04393_, _04397_);
  and _55310_ (_04482_, _04443_, _04406_);
  or _55311_ (_04483_, _04482_, _04481_);
  or _55312_ (_04484_, _04483_, _04480_);
  and _55313_ (_04485_, _04435_, _04426_);
  and _55314_ (_04486_, _04407_, _04434_);
  and _55315_ (_04487_, _04404_, _04419_);
  or _55316_ (_04488_, _04487_, _04486_);
  or _55317_ (_04489_, _04488_, _04485_);
  and _55318_ (_04490_, _04412_, _04401_);
  and _55319_ (_04491_, _04417_, _04355_);
  and _55320_ (_04492_, _04420_, _04442_);
  or _55321_ (_04493_, _04492_, _04491_);
  and _55322_ (_04494_, _04375_, _04439_);
  and _55323_ (_04495_, _04424_, _04381_);
  or _55324_ (_04496_, _04495_, _04494_);
  or _55325_ (_04497_, _04496_, _04493_);
  or _55326_ (_04498_, _04497_, _04490_);
  and _55327_ (_04499_, _04432_, _04423_);
  and _55328_ (_04500_, _04399_, _04415_);
  or _55329_ (_04501_, _04500_, _04499_);
  or _55330_ (_04502_, _04501_, _04498_);
  and _55331_ (_04503_, _04440_, _04411_);
  and _55332_ (_04504_, _04390_, _04431_);
  or _55333_ (_04505_, _04504_, _04503_);
  or _55334_ (_04506_, _04505_, _04502_);
  or _55335_ (_04507_, _04506_, _04489_);
  or _55336_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04507_, _04484_);
  and _55337_ (_04508_, _04440_, _04355_);
  and _55338_ (_04509_, _04384_, _04419_);
  or _55339_ (_04510_, _04509_, _04508_);
  and _55340_ (_04511_, _04379_, _04426_);
  and _55341_ (_04513_, _04443_, _04381_);
  or _55342_ (_04514_, _04513_, _04511_);
  or _55343_ (_04515_, _04514_, _04510_);
  and _55344_ (_04516_, _04407_, _04392_);
  and _55345_ (_04517_, _04399_, _04406_);
  or _55346_ (_04518_, _04517_, _04516_);
  and _55347_ (_04519_, _04435_, _04397_);
  or _55348_ (_04520_, _04519_, _04518_);
  and _55349_ (_04521_, _04412_, _04387_);
  and _55350_ (_04522_, _04424_, _04401_);
  and _55351_ (_04523_, _04375_, _04415_);
  or _55352_ (_04524_, _04523_, _04522_);
  and _55353_ (_04525_, _04420_, _04423_);
  and _55354_ (_04526_, _04417_, _04434_);
  or _55355_ (_04527_, _04526_, _04525_);
  or _55356_ (_04528_, _04527_, _04524_);
  or _55357_ (_04529_, _04528_, _04521_);
  and _55358_ (_04530_, _04404_, _04431_);
  and _55359_ (_04531_, _04432_, _04411_);
  or _55360_ (_04532_, _04531_, _04530_);
  or _55361_ (_04533_, _04532_, _04529_);
  and _55362_ (_04534_, _04390_, _04439_);
  and _55363_ (_04535_, _04393_, _04442_);
  or _55364_ (_04536_, _04535_, _04534_);
  or _55365_ (_04537_, _04536_, _04533_);
  or _55366_ (_04538_, _04537_, _04520_);
  or _55367_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04538_, _04515_);
  not _55368_ (_04539_, _00029_);
  and _55369_ (_04540_, _04393_, _04539_);
  not _55370_ (_04541_, _00388_);
  and _55371_ (_04542_, _04390_, _04541_);
  or _55372_ (_04543_, _04542_, _04540_);
  not _55373_ (_04544_, _43480_);
  and _55374_ (_04545_, _04384_, _04544_);
  not _55375_ (_04546_, _00306_);
  and _55376_ (_04547_, _04379_, _04546_);
  or _55377_ (_04548_, _04547_, _04545_);
  or _55378_ (_04549_, _04548_, _04543_);
  not _55379_ (_04550_, _00470_);
  and _55380_ (_04551_, _04432_, _04550_);
  not _55381_ (_04552_, _00179_);
  and _55382_ (_04553_, _04435_, _04552_);
  not _55383_ (_04554_, _00511_);
  and _55384_ (_04555_, _04404_, _04554_);
  or _55385_ (_04556_, _04555_, _04553_);
  or _55386_ (_04557_, _04556_, _04551_);
  not _55387_ (_04558_, _00070_);
  and _55388_ (_04559_, _04407_, _04558_);
  not _55389_ (_04560_, _00111_);
  and _55390_ (_04561_, _04399_, _04560_);
  or _55391_ (_04562_, _04561_, _04559_);
  not _55392_ (_04563_, _00429_);
  and _55393_ (_04564_, _04412_, _04563_);
  not _55394_ (_04565_, _00612_);
  and _55395_ (_04566_, _04420_, _04565_);
  not _55396_ (_04567_, _00265_);
  and _55397_ (_04568_, _04375_, _04567_);
  or _55398_ (_04569_, _04568_, _04566_);
  not _55399_ (_04570_, _00224_);
  and _55400_ (_04571_, _04417_, _04570_);
  not _55401_ (_04572_, _00558_);
  and _55402_ (_04573_, _04424_, _04572_);
  or _55403_ (_04574_, _04573_, _04571_);
  or _55404_ (_04575_, _04574_, _04569_);
  or _55405_ (_04576_, _04575_, _04564_);
  or _55406_ (_04577_, _04576_, _04562_);
  not _55407_ (_04578_, _43521_);
  and _55408_ (_04579_, _04443_, _04578_);
  not _55409_ (_04580_, _00347_);
  and _55410_ (_04581_, _04440_, _04580_);
  or _55411_ (_04582_, _04581_, _04579_);
  or _55412_ (_04583_, _04582_, _04577_);
  or _55413_ (_04584_, _04583_, _04557_);
  or _55414_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _04584_, _04549_);
  not _55415_ (_04585_, _00352_);
  and _55416_ (_04586_, _04440_, _04585_);
  not _55417_ (_04587_, _00311_);
  and _55418_ (_04588_, _04379_, _04587_);
  or _55419_ (_04589_, _04588_, _04586_);
  not _55420_ (_04590_, _43485_);
  and _55421_ (_04591_, _04384_, _04590_);
  not _55422_ (_04592_, _00393_);
  and _55423_ (_04593_, _04390_, _04592_);
  or _55424_ (_04594_, _04593_, _04591_);
  or _55425_ (_04595_, _04594_, _04589_);
  not _55426_ (_04596_, _00516_);
  and _55427_ (_04597_, _04404_, _04596_);
  not _55428_ (_04598_, _00075_);
  and _55429_ (_04599_, _04407_, _04598_);
  not _55430_ (_04600_, _00475_);
  and _55431_ (_04601_, _04432_, _04600_);
  or _55432_ (_04602_, _04601_, _04599_);
  or _55433_ (_04603_, _04602_, _04597_);
  not _55434_ (_04604_, _43526_);
  and _55435_ (_04605_, _04443_, _04604_);
  not _55436_ (_04606_, _00034_);
  and _55437_ (_04607_, _04393_, _04606_);
  or _55438_ (_04608_, _04607_, _04605_);
  not _55439_ (_04609_, _00434_);
  and _55440_ (_04610_, _04412_, _04609_);
  not _55441_ (_04612_, _00617_);
  and _55442_ (_04613_, _04420_, _04612_);
  not _55443_ (_04614_, _00270_);
  and _55444_ (_04615_, _04375_, _04614_);
  or _55445_ (_04616_, _04615_, _04613_);
  not _55446_ (_04617_, _00229_);
  and _55447_ (_04618_, _04417_, _04617_);
  not _55448_ (_04619_, _00566_);
  and _55449_ (_04620_, _04424_, _04619_);
  or _55450_ (_04621_, _04620_, _04618_);
  or _55451_ (_04622_, _04621_, _04616_);
  or _55452_ (_04623_, _04622_, _04610_);
  not _55453_ (_04624_, _00188_);
  and _55454_ (_04625_, _04435_, _04624_);
  not _55455_ (_04626_, _00116_);
  and _55456_ (_04627_, _04399_, _04626_);
  or _55457_ (_04628_, _04627_, _04625_);
  or _55458_ (_04629_, _04628_, _04623_);
  or _55459_ (_04630_, _04629_, _04608_);
  or _55460_ (_04631_, _04630_, _04603_);
  or _55461_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _04631_, _04595_);
  not _55462_ (_04632_, _00316_);
  and _55463_ (_04633_, _04379_, _04632_);
  not _55464_ (_04634_, _43531_);
  and _55465_ (_04635_, _04443_, _04634_);
  or _55466_ (_04636_, _04635_, _04633_);
  not _55467_ (_04637_, _00357_);
  and _55468_ (_04638_, _04440_, _04637_);
  not _55469_ (_04639_, _43490_);
  and _55470_ (_04640_, _04384_, _04639_);
  or _55471_ (_04641_, _04640_, _04638_);
  or _55472_ (_04642_, _04641_, _04636_);
  not _55473_ (_04643_, _00121_);
  and _55474_ (_04644_, _04399_, _04643_);
  not _55475_ (_04645_, _00521_);
  and _55476_ (_04646_, _04404_, _04645_);
  not _55477_ (_04647_, _00080_);
  and _55478_ (_04648_, _04407_, _04647_);
  or _55479_ (_04649_, _04648_, _04646_);
  or _55480_ (_04650_, _04649_, _04644_);
  not _55481_ (_04651_, _00439_);
  and _55482_ (_04652_, _04412_, _04651_);
  not _55483_ (_04653_, _00574_);
  and _55484_ (_04654_, _04424_, _04653_);
  not _55485_ (_04655_, _00275_);
  and _55486_ (_04656_, _04375_, _04655_);
  or _55487_ (_04657_, _04656_, _04654_);
  not _55488_ (_04658_, _00622_);
  and _55489_ (_04659_, _04420_, _04658_);
  not _55490_ (_04660_, _00234_);
  and _55491_ (_04661_, _04417_, _04660_);
  or _55492_ (_04662_, _04661_, _04659_);
  or _55493_ (_04663_, _04662_, _04657_);
  or _55494_ (_04664_, _04663_, _04652_);
  not _55495_ (_04665_, _00480_);
  and _55496_ (_04666_, _04432_, _04665_);
  not _55497_ (_04667_, _00193_);
  and _55498_ (_04668_, _04435_, _04667_);
  or _55499_ (_04669_, _04668_, _04666_);
  or _55500_ (_04670_, _04669_, _04664_);
  not _55501_ (_04671_, _00398_);
  and _55502_ (_04672_, _04390_, _04671_);
  not _55503_ (_04673_, _00039_);
  and _55504_ (_04674_, _04393_, _04673_);
  or _55505_ (_04675_, _04674_, _04672_);
  or _55506_ (_04676_, _04675_, _04670_);
  or _55507_ (_04677_, _04676_, _04650_);
  or _55508_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _04677_, _04642_);
  not _55509_ (_04678_, _00403_);
  and _55510_ (_04679_, _04390_, _04678_);
  not _55511_ (_04680_, _00003_);
  and _55512_ (_04681_, _04443_, _04680_);
  or _55513_ (_04682_, _04681_, _04679_);
  not _55514_ (_04683_, _00321_);
  and _55515_ (_04684_, _04379_, _04683_);
  not _55516_ (_04685_, _43495_);
  and _55517_ (_04686_, _04384_, _04685_);
  or _55518_ (_04687_, _04686_, _04684_);
  or _55519_ (_04688_, _04687_, _04682_);
  not _55520_ (_04689_, _00526_);
  and _55521_ (_04690_, _04404_, _04689_);
  not _55522_ (_04691_, _00485_);
  and _55523_ (_04692_, _04432_, _04691_);
  not _55524_ (_04693_, _00085_);
  and _55525_ (_04694_, _04407_, _04693_);
  or _55526_ (_04695_, _04694_, _04692_);
  or _55527_ (_04696_, _04695_, _04690_);
  not _55528_ (_04697_, _00444_);
  and _55529_ (_04698_, _04412_, _04697_);
  not _55530_ (_04699_, _00627_);
  and _55531_ (_04700_, _04420_, _04699_);
  not _55532_ (_04701_, _00239_);
  and _55533_ (_04702_, _04417_, _04701_);
  or _55534_ (_04703_, _04702_, _04700_);
  not _55535_ (_04704_, _00582_);
  and _55536_ (_04705_, _04424_, _04704_);
  not _55537_ (_04706_, _00280_);
  and _55538_ (_04707_, _04375_, _04706_);
  or _55539_ (_04708_, _04707_, _04705_);
  or _55540_ (_04709_, _04708_, _04703_);
  or _55541_ (_04710_, _04709_, _04698_);
  not _55542_ (_04711_, _00198_);
  and _55543_ (_04712_, _04435_, _04711_);
  not _55544_ (_04713_, _00126_);
  and _55545_ (_04714_, _04399_, _04713_);
  or _55546_ (_04715_, _04714_, _04712_);
  or _55547_ (_04716_, _04715_, _04710_);
  not _55548_ (_04717_, _00362_);
  and _55549_ (_04718_, _04440_, _04717_);
  not _55550_ (_04719_, _00044_);
  and _55551_ (_04720_, _04393_, _04719_);
  or _55552_ (_04721_, _04720_, _04718_);
  or _55553_ (_04722_, _04721_, _04716_);
  or _55554_ (_04723_, _04722_, _04696_);
  or _55555_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _04723_, _04688_);
  not _55556_ (_04724_, _00326_);
  and _55557_ (_04725_, _04379_, _04724_);
  not _55558_ (_04726_, _00008_);
  and _55559_ (_04727_, _04443_, _04726_);
  or _55560_ (_04728_, _04727_, _04725_);
  not _55561_ (_04729_, _00367_);
  and _55562_ (_04730_, _04440_, _04729_);
  not _55563_ (_04731_, _43500_);
  and _55564_ (_04732_, _04384_, _04731_);
  or _55565_ (_04733_, _04732_, _04730_);
  or _55566_ (_04734_, _04733_, _04728_);
  not _55567_ (_04735_, _00133_);
  and _55568_ (_04736_, _04399_, _04735_);
  not _55569_ (_04737_, _00531_);
  and _55570_ (_04738_, _04404_, _04737_);
  not _55571_ (_04739_, _00090_);
  and _55572_ (_04740_, _04407_, _04739_);
  or _55573_ (_04741_, _04740_, _04738_);
  or _55574_ (_04742_, _04741_, _04736_);
  not _55575_ (_04743_, _00449_);
  and _55576_ (_04744_, _04412_, _04743_);
  not _55577_ (_04745_, _00590_);
  and _55578_ (_04746_, _04424_, _04745_);
  not _55579_ (_04747_, _00285_);
  and _55580_ (_04748_, _04375_, _04747_);
  or _55581_ (_04749_, _04748_, _04746_);
  not _55582_ (_04750_, _00632_);
  and _55583_ (_04751_, _04420_, _04750_);
  not _55584_ (_04752_, _00244_);
  and _55585_ (_04753_, _04417_, _04752_);
  or _55586_ (_04754_, _04753_, _04751_);
  or _55587_ (_04755_, _04754_, _04749_);
  or _55588_ (_04756_, _04755_, _04744_);
  not _55589_ (_04757_, _00490_);
  and _55590_ (_04758_, _04432_, _04757_);
  not _55591_ (_04759_, _00203_);
  and _55592_ (_04760_, _04435_, _04759_);
  or _55593_ (_04761_, _04760_, _04758_);
  or _55594_ (_04762_, _04761_, _04756_);
  not _55595_ (_04763_, _00408_);
  and _55596_ (_04764_, _04390_, _04763_);
  not _55597_ (_04765_, _00049_);
  and _55598_ (_04766_, _04393_, _04765_);
  or _55599_ (_04767_, _04766_, _04764_);
  or _55600_ (_04768_, _04767_, _04762_);
  or _55601_ (_04769_, _04768_, _04742_);
  or _55602_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _04769_, _04734_);
  not _55603_ (_04770_, _00331_);
  and _55604_ (_04771_, _04379_, _04770_);
  not _55605_ (_04772_, _00013_);
  and _55606_ (_04773_, _04443_, _04772_);
  or _55607_ (_04774_, _04773_, _04771_);
  not _55608_ (_04775_, _00372_);
  and _55609_ (_04776_, _04440_, _04775_);
  not _55610_ (_04777_, _43505_);
  and _55611_ (_04778_, _04384_, _04777_);
  or _55612_ (_04779_, _04778_, _04776_);
  or _55613_ (_04780_, _04779_, _04774_);
  not _55614_ (_04781_, _00095_);
  and _55615_ (_04782_, _04407_, _04781_);
  not _55616_ (_04783_, _00536_);
  and _55617_ (_04784_, _04404_, _04783_);
  not _55618_ (_04785_, _00495_);
  and _55619_ (_04786_, _04432_, _04785_);
  or _55620_ (_04787_, _04786_, _04784_);
  or _55621_ (_04788_, _04787_, _04782_);
  not _55622_ (_04789_, _00454_);
  and _55623_ (_04790_, _04412_, _04789_);
  not _55624_ (_04791_, _00596_);
  and _55625_ (_04792_, _04424_, _04791_);
  not _55626_ (_04793_, _00290_);
  and _55627_ (_04794_, _04375_, _04793_);
  or _55628_ (_04795_, _04794_, _04792_);
  not _55629_ (_04796_, _00637_);
  and _55630_ (_04797_, _04420_, _04796_);
  not _55631_ (_04798_, _00249_);
  and _55632_ (_04799_, _04417_, _04798_);
  or _55633_ (_04800_, _04799_, _04797_);
  or _55634_ (_04801_, _04800_, _04795_);
  or _55635_ (_04802_, _04801_, _04790_);
  not _55636_ (_04803_, _00208_);
  and _55637_ (_04804_, _04435_, _04803_);
  not _55638_ (_04805_, _00144_);
  and _55639_ (_04806_, _04399_, _04805_);
  or _55640_ (_04807_, _04806_, _04804_);
  or _55641_ (_04808_, _04807_, _04802_);
  not _55642_ (_04809_, _00413_);
  and _55643_ (_04810_, _04390_, _04809_);
  not _55644_ (_04811_, _00054_);
  and _55645_ (_04812_, _04393_, _04811_);
  or _55646_ (_04813_, _04812_, _04810_);
  or _55647_ (_04814_, _04813_, _04808_);
  or _55648_ (_04815_, _04814_, _04788_);
  or _55649_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _04815_, _04780_);
  not _55650_ (_04816_, _00336_);
  and _55651_ (_04817_, _04379_, _04816_);
  not _55652_ (_04818_, _00018_);
  and _55653_ (_04819_, _04443_, _04818_);
  or _55654_ (_04820_, _04819_, _04817_);
  not _55655_ (_04821_, _00377_);
  and _55656_ (_04822_, _04440_, _04821_);
  not _55657_ (_04823_, _43510_);
  and _55658_ (_04824_, _04384_, _04823_);
  or _55659_ (_04825_, _04824_, _04822_);
  or _55660_ (_04826_, _04825_, _04820_);
  not _55661_ (_04827_, _00155_);
  and _55662_ (_04828_, _04399_, _04827_);
  not _55663_ (_04829_, _00541_);
  and _55664_ (_04830_, _04404_, _04829_);
  not _55665_ (_04831_, _00100_);
  and _55666_ (_04832_, _04407_, _04831_);
  or _55667_ (_04833_, _04832_, _04830_);
  or _55668_ (_04834_, _04833_, _04828_);
  not _55669_ (_04835_, _00459_);
  and _55670_ (_04836_, _04412_, _04835_);
  not _55671_ (_04837_, _00601_);
  and _55672_ (_04838_, _04424_, _04837_);
  not _55673_ (_04839_, _00295_);
  and _55674_ (_04840_, _04375_, _04839_);
  or _55675_ (_04841_, _04840_, _04838_);
  not _55676_ (_04842_, _00642_);
  and _55677_ (_04843_, _04420_, _04842_);
  not _55678_ (_04844_, _00254_);
  and _55679_ (_04845_, _04417_, _04844_);
  or _55680_ (_04846_, _04845_, _04843_);
  or _55681_ (_04847_, _04846_, _04841_);
  or _55682_ (_04848_, _04847_, _04836_);
  not _55683_ (_04849_, _00500_);
  and _55684_ (_04850_, _04432_, _04849_);
  not _55685_ (_04851_, _00213_);
  and _55686_ (_04852_, _04435_, _04851_);
  or _55687_ (_04853_, _04852_, _04850_);
  or _55688_ (_04854_, _04853_, _04848_);
  not _55689_ (_04855_, _00418_);
  and _55690_ (_04856_, _04390_, _04855_);
  not _55691_ (_04857_, _00059_);
  and _55692_ (_04858_, _04393_, _04857_);
  or _55693_ (_04859_, _04858_, _04856_);
  or _55694_ (_04860_, _04859_, _04854_);
  or _55695_ (_04861_, _04860_, _04834_);
  or _55696_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _04861_, _04826_);
  and _55697_ (_04862_, _04393_, _04552_);
  and _55698_ (_04863_, _04384_, _04558_);
  or _55699_ (_04864_, _04863_, _04862_);
  and _55700_ (_04865_, _04390_, _04554_);
  and _55701_ (_04866_, _04379_, _04563_);
  or _55702_ (_04867_, _04866_, _04865_);
  or _55703_ (_04868_, _04867_, _04864_);
  and _55704_ (_04869_, _04404_, _04544_);
  and _55705_ (_04870_, _04432_, _04565_);
  and _55706_ (_04871_, _04435_, _04546_);
  or _55707_ (_04872_, _04871_, _04870_);
  or _55708_ (_04873_, _04872_, _04869_);
  and _55709_ (_04874_, _04399_, _04567_);
  and _55710_ (_04875_, _04407_, _04570_);
  or _55711_ (_04876_, _04875_, _04874_);
  and _55712_ (_04877_, _04412_, _04572_);
  and _55713_ (_04878_, _04417_, _04580_);
  and _55714_ (_04879_, _04420_, _04539_);
  or _55715_ (_04880_, _04879_, _04878_);
  and _55716_ (_04881_, _04375_, _04541_);
  and _55717_ (_04882_, _04424_, _04578_);
  or _55718_ (_04883_, _04882_, _04881_);
  or _55719_ (_04884_, _04883_, _04880_);
  or _55720_ (_04885_, _04884_, _04877_);
  or _55721_ (_04886_, _04885_, _04876_);
  and _55722_ (_04887_, _04440_, _04550_);
  and _55723_ (_04888_, _04443_, _04560_);
  or _55724_ (_04889_, _04888_, _04887_);
  or _55725_ (_04890_, _04889_, _04886_);
  or _55726_ (_04891_, _04890_, _04873_);
  or _55727_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04891_, _04868_);
  and _55728_ (_04892_, _04384_, _04598_);
  and _55729_ (_04893_, _04443_, _04626_);
  or _55730_ (_04894_, _04893_, _04892_);
  and _55731_ (_04895_, _04390_, _04596_);
  and _55732_ (_04896_, _04393_, _04624_);
  or _55733_ (_04897_, _04896_, _04895_);
  or _55734_ (_04898_, _04897_, _04894_);
  and _55735_ (_04899_, _04404_, _04590_);
  and _55736_ (_04900_, _04432_, _04612_);
  and _55737_ (_04901_, _04435_, _04587_);
  or _55738_ (_04902_, _04901_, _04900_);
  or _55739_ (_04903_, _04902_, _04899_);
  and _55740_ (_04904_, _04440_, _04600_);
  and _55741_ (_04905_, _04379_, _04609_);
  or _55742_ (_04906_, _04905_, _04904_);
  and _55743_ (_04907_, _04399_, _04614_);
  and _55744_ (_04908_, _04407_, _04617_);
  or _55745_ (_04909_, _04908_, _04907_);
  and _55746_ (_04910_, _04412_, _04619_);
  and _55747_ (_04911_, _04417_, _04585_);
  and _55748_ (_04912_, _04375_, _04592_);
  or _55749_ (_04913_, _04912_, _04911_);
  and _55750_ (_04914_, _04424_, _04604_);
  and _55751_ (_04915_, _04420_, _04606_);
  or _55752_ (_04916_, _04915_, _04914_);
  or _55753_ (_04917_, _04916_, _04913_);
  or _55754_ (_04918_, _04917_, _04910_);
  or _55755_ (_04919_, _04918_, _04909_);
  or _55756_ (_04920_, _04919_, _04906_);
  or _55757_ (_04921_, _04920_, _04903_);
  or _55758_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04921_, _04898_);
  and _55759_ (_04922_, _04443_, _04643_);
  and _55760_ (_04923_, _04384_, _04647_);
  or _55761_ (_04924_, _04923_, _04922_);
  and _55762_ (_04925_, _04390_, _04645_);
  and _55763_ (_04926_, _04379_, _04651_);
  or _55764_ (_04927_, _04926_, _04925_);
  or _55765_ (_04928_, _04927_, _04924_);
  and _55766_ (_04929_, _04435_, _04632_);
  and _55767_ (_04930_, _04399_, _04655_);
  and _55768_ (_04931_, _04404_, _04639_);
  or _55769_ (_04932_, _04931_, _04930_);
  or _55770_ (_04933_, _04932_, _04929_);
  and _55771_ (_04934_, _04412_, _04653_);
  and _55772_ (_04935_, _04375_, _04671_);
  and _55773_ (_04936_, _04424_, _04634_);
  or _55774_ (_04937_, _04936_, _04935_);
  and _55775_ (_04938_, _04417_, _04637_);
  and _55776_ (_04939_, _04420_, _04673_);
  or _55777_ (_04940_, _04939_, _04938_);
  or _55778_ (_04941_, _04940_, _04937_);
  or _55779_ (_04942_, _04941_, _04934_);
  and _55780_ (_04943_, _04432_, _04658_);
  and _55781_ (_04944_, _04407_, _04660_);
  or _55782_ (_04945_, _04944_, _04943_);
  or _55783_ (_04946_, _04945_, _04942_);
  and _55784_ (_04947_, _04440_, _04665_);
  and _55785_ (_04948_, _04393_, _04667_);
  or _55786_ (_04949_, _04948_, _04947_);
  or _55787_ (_04950_, _04949_, _04946_);
  or _55788_ (_04951_, _04950_, _04933_);
  or _55789_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04951_, _04928_);
  and _55790_ (_04952_, _04440_, _04691_);
  and _55791_ (_04953_, _04384_, _04693_);
  or _55792_ (_04954_, _04953_, _04952_);
  and _55793_ (_04955_, _04379_, _04697_);
  and _55794_ (_04956_, _04443_, _04713_);
  or _55795_ (_04957_, _04956_, _04955_);
  or _55796_ (_04958_, _04957_, _04954_);
  and _55797_ (_04959_, _04432_, _04699_);
  and _55798_ (_04960_, _04435_, _04683_);
  and _55799_ (_04961_, _04404_, _04685_);
  or _55800_ (_04962_, _04961_, _04960_);
  or _55801_ (_04963_, _04962_, _04959_);
  and _55802_ (_04964_, _04399_, _04706_);
  and _55803_ (_04965_, _04407_, _04701_);
  or _55804_ (_04966_, _04965_, _04964_);
  and _55805_ (_04967_, _04412_, _04704_);
  and _55806_ (_04968_, _04417_, _04717_);
  and _55807_ (_04969_, _04420_, _04719_);
  or _55808_ (_04970_, _04969_, _04968_);
  and _55809_ (_04971_, _04375_, _04678_);
  and _55810_ (_04972_, _04424_, _04680_);
  or _55811_ (_04973_, _04972_, _04971_);
  or _55812_ (_04974_, _04973_, _04970_);
  or _55813_ (_04975_, _04974_, _04967_);
  or _55814_ (_04976_, _04975_, _04966_);
  and _55815_ (_04977_, _04390_, _04689_);
  and _55816_ (_04978_, _04393_, _04711_);
  or _55817_ (_04979_, _04978_, _04977_);
  or _55818_ (_04980_, _04979_, _04976_);
  or _55819_ (_04981_, _04980_, _04963_);
  or _55820_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04981_, _04958_);
  and _55821_ (_04982_, _04379_, _04743_);
  and _55822_ (_04983_, _04384_, _04739_);
  or _55823_ (_04984_, _04983_, _04982_);
  and _55824_ (_04985_, _04393_, _04759_);
  and _55825_ (_04986_, _04443_, _04735_);
  or _55826_ (_04987_, _04986_, _04985_);
  or _55827_ (_04988_, _04987_, _04984_);
  and _55828_ (_04989_, _04435_, _04724_);
  and _55829_ (_04990_, _04407_, _04752_);
  and _55830_ (_04991_, _04404_, _04731_);
  or _55831_ (_04992_, _04991_, _04990_);
  or _55832_ (_04993_, _04992_, _04989_);
  and _55833_ (_04994_, _04412_, _04745_);
  and _55834_ (_04995_, _04417_, _04729_);
  and _55835_ (_04996_, _04420_, _04765_);
  or _55836_ (_04997_, _04996_, _04995_);
  and _55837_ (_04998_, _04375_, _04763_);
  and _55838_ (_04999_, _04424_, _04726_);
  or _55839_ (_05000_, _04999_, _04998_);
  or _55840_ (_05001_, _05000_, _04997_);
  or _55841_ (_05002_, _05001_, _04994_);
  and _55842_ (_05003_, _04432_, _04750_);
  and _55843_ (_05004_, _04399_, _04747_);
  or _55844_ (_05005_, _05004_, _05003_);
  or _55845_ (_05006_, _05005_, _05002_);
  and _55846_ (_05007_, _04440_, _04757_);
  and _55847_ (_05008_, _04390_, _04737_);
  or _55848_ (_05009_, _05008_, _05007_);
  or _55849_ (_05010_, _05009_, _05006_);
  or _55850_ (_05011_, _05010_, _04993_);
  or _55851_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _05011_, _04988_);
  and _55852_ (_05012_, _04443_, _04805_);
  and _55853_ (_05013_, _04384_, _04781_);
  or _55854_ (_05014_, _05013_, _05012_);
  and _55855_ (_05015_, _04440_, _04785_);
  and _55856_ (_05016_, _04393_, _04803_);
  or _55857_ (_05017_, _05016_, _05015_);
  or _55858_ (_05018_, _05017_, _05014_);
  and _55859_ (_05019_, _04407_, _04798_);
  and _55860_ (_05020_, _04435_, _04770_);
  and _55861_ (_05021_, _04404_, _04777_);
  or _55862_ (_05022_, _05021_, _05020_);
  or _55863_ (_05023_, _05022_, _05019_);
  and _55864_ (_05024_, _04412_, _04791_);
  and _55865_ (_05025_, _04375_, _04809_);
  and _55866_ (_05026_, _04424_, _04772_);
  or _55867_ (_05027_, _05026_, _05025_);
  and _55868_ (_05028_, _04417_, _04775_);
  and _55869_ (_05029_, _04420_, _04811_);
  or _55870_ (_05030_, _05029_, _05028_);
  or _55871_ (_05031_, _05030_, _05027_);
  or _55872_ (_05032_, _05031_, _05024_);
  and _55873_ (_05033_, _04432_, _04796_);
  and _55874_ (_05034_, _04399_, _04793_);
  or _55875_ (_05035_, _05034_, _05033_);
  or _55876_ (_05036_, _05035_, _05032_);
  and _55877_ (_05037_, _04379_, _04789_);
  and _55878_ (_05038_, _04390_, _04783_);
  or _55879_ (_05039_, _05038_, _05037_);
  or _55880_ (_05040_, _05039_, _05036_);
  or _55881_ (_05041_, _05040_, _05023_);
  or _55882_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _05041_, _05018_);
  and _55883_ (_05042_, _04443_, _04827_);
  and _55884_ (_05043_, _04384_, _04831_);
  or _55885_ (_05044_, _05043_, _05042_);
  and _55886_ (_05045_, _04390_, _04829_);
  and _55887_ (_05046_, _04379_, _04835_);
  or _55888_ (_05047_, _05046_, _05045_);
  or _55889_ (_05048_, _05047_, _05044_);
  and _55890_ (_05049_, _04407_, _04844_);
  and _55891_ (_05050_, _04432_, _04842_);
  and _55892_ (_05051_, _04404_, _04823_);
  or _55893_ (_05052_, _05051_, _05050_);
  or _55894_ (_05054_, _05052_, _05049_);
  and _55895_ (_05056_, _04399_, _04839_);
  and _55896_ (_05058_, _04435_, _04816_);
  or _55897_ (_05060_, _05058_, _05056_);
  and _55898_ (_05062_, _04412_, _04837_);
  and _55899_ (_05064_, _04417_, _04821_);
  and _55900_ (_05066_, _04420_, _04857_);
  or _55901_ (_05067_, _05066_, _05064_);
  and _55902_ (_05068_, _04375_, _04855_);
  and _55903_ (_05069_, _04424_, _04818_);
  or _55904_ (_05070_, _05069_, _05068_);
  or _55905_ (_05071_, _05070_, _05067_);
  or _55906_ (_05072_, _05071_, _05062_);
  or _55907_ (_05074_, _05072_, _05060_);
  and _55908_ (_05075_, _04440_, _04849_);
  and _55909_ (_05077_, _04393_, _04851_);
  or _55910_ (_05078_, _05077_, _05075_);
  or _55911_ (_05079_, _05078_, _05074_);
  or _55912_ (_05081_, _05079_, _05054_);
  or _55913_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _05081_, _05048_);
  and _55914_ (_05082_, _04390_, _04563_);
  and _55915_ (_05084_, _04393_, _04558_);
  or _55916_ (_05085_, _05084_, _05082_);
  and _55917_ (_05086_, _04379_, _04580_);
  and _55918_ (_05088_, _04384_, _04578_);
  or _55919_ (_05089_, _05088_, _05086_);
  or _55920_ (_05090_, _05089_, _05085_);
  and _55921_ (_05092_, _04407_, _04560_);
  and _55922_ (_05093_, _04404_, _04572_);
  and _55923_ (_05094_, _04435_, _04570_);
  or _55924_ (_05096_, _05094_, _05093_);
  or _55925_ (_05097_, _05096_, _05092_);
  and _55926_ (_05098_, _04412_, _04550_);
  and _55927_ (_05100_, _04375_, _04546_);
  and _55928_ (_05101_, _04417_, _04567_);
  or _55929_ (_05102_, _05101_, _05100_);
  and _55930_ (_05104_, _04424_, _04565_);
  and _55931_ (_05105_, _04420_, _04544_);
  or _55932_ (_05106_, _05105_, _05104_);
  or _55933_ (_05107_, _05106_, _05102_);
  or _55934_ (_05108_, _05107_, _05098_);
  and _55935_ (_05109_, _04432_, _04554_);
  and _55936_ (_05110_, _04399_, _04552_);
  or _55937_ (_05111_, _05110_, _05109_);
  or _55938_ (_05112_, _05111_, _05108_);
  and _55939_ (_05113_, _04440_, _04541_);
  and _55940_ (_05114_, _04443_, _04539_);
  or _55941_ (_05115_, _05114_, _05113_);
  or _55942_ (_05116_, _05115_, _05112_);
  or _55943_ (_05117_, _05116_, _05097_);
  or _55944_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _05117_, _05090_);
  and _55945_ (_05118_, _04390_, _04609_);
  and _55946_ (_05119_, _04393_, _04598_);
  or _55947_ (_05120_, _05119_, _05118_);
  and _55948_ (_05121_, _04379_, _04585_);
  and _55949_ (_05122_, _04384_, _04604_);
  or _55950_ (_05123_, _05122_, _05121_);
  or _55951_ (_05125_, _05123_, _05120_);
  and _55952_ (_05126_, _04435_, _04617_);
  and _55953_ (_05128_, _04404_, _04619_);
  and _55954_ (_05129_, _04407_, _04626_);
  or _55955_ (_05130_, _05129_, _05128_);
  or _55956_ (_05132_, _05130_, _05126_);
  and _55957_ (_05133_, _04412_, _04600_);
  and _55958_ (_05134_, _04375_, _04587_);
  and _55959_ (_05136_, _04417_, _04614_);
  or _55960_ (_05137_, _05136_, _05134_);
  and _55961_ (_05138_, _04424_, _04612_);
  and _55962_ (_05140_, _04420_, _04590_);
  or _55963_ (_05141_, _05140_, _05138_);
  or _55964_ (_05142_, _05141_, _05137_);
  or _55965_ (_05144_, _05142_, _05133_);
  and _55966_ (_05145_, _04432_, _04596_);
  and _55967_ (_05146_, _04399_, _04624_);
  or _55968_ (_05148_, _05146_, _05145_);
  or _55969_ (_05149_, _05148_, _05144_);
  and _55970_ (_05150_, _04440_, _04592_);
  and _55971_ (_05152_, _04443_, _04606_);
  or _55972_ (_05153_, _05152_, _05150_);
  or _55973_ (_05154_, _05153_, _05149_);
  or _55974_ (_05156_, _05154_, _05132_);
  or _55975_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _05156_, _05125_);
  and _55976_ (_05157_, _04379_, _04637_);
  and _55977_ (_05158_, _04384_, _04634_);
  or _55978_ (_05159_, _05158_, _05157_);
  and _55979_ (_05160_, _04390_, _04651_);
  and _55980_ (_05161_, _04393_, _04647_);
  or _55981_ (_05162_, _05161_, _05160_);
  or _55982_ (_05163_, _05162_, _05159_);
  and _55983_ (_05164_, _04432_, _04645_);
  and _55984_ (_05165_, _04399_, _04667_);
  and _55985_ (_05166_, _04435_, _04660_);
  or _55986_ (_05167_, _05166_, _05165_);
  or _55987_ (_05168_, _05167_, _05164_);
  and _55988_ (_05169_, _04412_, _04665_);
  and _55989_ (_05170_, _04417_, _04655_);
  and _55990_ (_05171_, _04420_, _04639_);
  or _55991_ (_05172_, _05171_, _05170_);
  and _55992_ (_05173_, _04424_, _04658_);
  and _55993_ (_05174_, _04375_, _04632_);
  or _55994_ (_05175_, _05174_, _05173_);
  or _55995_ (_05177_, _05175_, _05172_);
  or _55996_ (_05178_, _05177_, _05169_);
  and _55997_ (_05180_, _04404_, _04653_);
  and _55998_ (_05181_, _04407_, _04643_);
  or _55999_ (_05182_, _05181_, _05180_);
  or _56000_ (_05184_, _05182_, _05178_);
  and _56001_ (_05185_, _04440_, _04671_);
  and _56002_ (_05186_, _04443_, _04673_);
  or _56003_ (_05188_, _05186_, _05185_);
  or _56004_ (_05189_, _05188_, _05184_);
  or _56005_ (_05190_, _05189_, _05168_);
  or _56006_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05190_, _05163_);
  and _56007_ (_05192_, _04443_, _04719_);
  and _56008_ (_05193_, _04384_, _04680_);
  or _56009_ (_05195_, _05193_, _05192_);
  and _56010_ (_05196_, _04390_, _04697_);
  and _56011_ (_05197_, _04393_, _04693_);
  or _56012_ (_05199_, _05197_, _05196_);
  or _56013_ (_05200_, _05199_, _05195_);
  and _56014_ (_05201_, _04407_, _04713_);
  and _56015_ (_05203_, _04399_, _04711_);
  and _56016_ (_05204_, _04435_, _04701_);
  or _56017_ (_05205_, _05204_, _05203_);
  or _56018_ (_05207_, _05205_, _05201_);
  and _56019_ (_05208_, _04440_, _04678_);
  and _56020_ (_05209_, _04379_, _04717_);
  or _56021_ (_05210_, _05209_, _05208_);
  and _56022_ (_05211_, _04404_, _04704_);
  and _56023_ (_05212_, _04432_, _04689_);
  or _56024_ (_05213_, _05212_, _05211_);
  and _56025_ (_05214_, _04412_, _04691_);
  and _56026_ (_05215_, _04424_, _04699_);
  and _56027_ (_05216_, _04417_, _04706_);
  or _56028_ (_05217_, _05216_, _05215_);
  and _56029_ (_05218_, _04375_, _04683_);
  and _56030_ (_05219_, _04420_, _04685_);
  or _56031_ (_05220_, _05219_, _05218_);
  or _56032_ (_05221_, _05220_, _05217_);
  or _56033_ (_05222_, _05221_, _05214_);
  or _56034_ (_05223_, _05222_, _05213_);
  or _56035_ (_05224_, _05223_, _05210_);
  or _56036_ (_05225_, _05224_, _05207_);
  or _56037_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05225_, _05200_);
  and _56038_ (_05226_, _04379_, _04729_);
  and _56039_ (_05228_, _04384_, _04726_);
  or _56040_ (_05229_, _05228_, _05226_);
  and _56041_ (_05231_, _04390_, _04743_);
  and _56042_ (_05232_, _04443_, _04765_);
  or _56043_ (_05233_, _05232_, _05231_);
  or _56044_ (_05235_, _05233_, _05229_);
  and _56045_ (_05236_, _04404_, _04745_);
  and _56046_ (_05237_, _04432_, _04737_);
  and _56047_ (_05239_, _04399_, _04759_);
  or _56048_ (_05240_, _05239_, _05237_);
  or _56049_ (_05241_, _05240_, _05236_);
  and _56050_ (_05243_, _04412_, _04757_);
  and _56051_ (_05244_, _04417_, _04747_);
  and _56052_ (_05245_, _04420_, _04731_);
  or _56053_ (_05247_, _05245_, _05244_);
  and _56054_ (_05248_, _04424_, _04750_);
  and _56055_ (_05249_, _04375_, _04724_);
  or _56056_ (_05251_, _05249_, _05248_);
  or _56057_ (_05252_, _05251_, _05247_);
  or _56058_ (_05253_, _05252_, _05243_);
  and _56059_ (_05255_, _04435_, _04752_);
  and _56060_ (_05256_, _04407_, _04735_);
  or _56061_ (_05257_, _05256_, _05255_);
  or _56062_ (_05259_, _05257_, _05253_);
  and _56063_ (_05260_, _04440_, _04763_);
  and _56064_ (_05261_, _04393_, _04739_);
  or _56065_ (_05262_, _05261_, _05260_);
  or _56066_ (_05263_, _05262_, _05259_);
  or _56067_ (_05264_, _05263_, _05241_);
  or _56068_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05264_, _05235_);
  and _56069_ (_05265_, _04390_, _04789_);
  and _56070_ (_05266_, _04440_, _04809_);
  or _56071_ (_05267_, _05266_, _05265_);
  and _56072_ (_05268_, _04393_, _04781_);
  and _56073_ (_05269_, _04384_, _04772_);
  or _56074_ (_05270_, _05269_, _05268_);
  or _56075_ (_05271_, _05270_, _05267_);
  and _56076_ (_05272_, _04407_, _04805_);
  and _56077_ (_05273_, _04404_, _04791_);
  and _56078_ (_05274_, _04435_, _04798_);
  or _56079_ (_05275_, _05274_, _05273_);
  or _56080_ (_05276_, _05275_, _05272_);
  and _56081_ (_05277_, _04412_, _04785_);
  and _56082_ (_05278_, _04424_, _04796_);
  and _56083_ (_05280_, _04375_, _04770_);
  or _56084_ (_05281_, _05280_, _05278_);
  and _56085_ (_05283_, _04417_, _04793_);
  and _56086_ (_05284_, _04420_, _04777_);
  or _56087_ (_05285_, _05284_, _05283_);
  or _56088_ (_05287_, _05285_, _05281_);
  or _56089_ (_05288_, _05287_, _05277_);
  and _56090_ (_05289_, _04432_, _04783_);
  and _56091_ (_05291_, _04399_, _04803_);
  or _56092_ (_05292_, _05291_, _05289_);
  or _56093_ (_05293_, _05292_, _05288_);
  and _56094_ (_05295_, _04379_, _04775_);
  and _56095_ (_05296_, _04443_, _04811_);
  or _56096_ (_05297_, _05296_, _05295_);
  or _56097_ (_05299_, _05297_, _05293_);
  or _56098_ (_05300_, _05299_, _05276_);
  or _56099_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05300_, _05271_);
  and _56100_ (_05302_, _04379_, _04821_);
  and _56101_ (_05303_, _04384_, _04818_);
  or _56102_ (_05304_, _05303_, _05302_);
  and _56103_ (_05306_, _04390_, _04835_);
  and _56104_ (_05307_, _04393_, _04831_);
  or _56105_ (_05308_, _05307_, _05306_);
  or _56106_ (_05310_, _05308_, _05304_);
  and _56107_ (_05311_, _04404_, _04837_);
  and _56108_ (_05312_, _04432_, _04829_);
  and _56109_ (_05313_, _04407_, _04827_);
  or _56110_ (_05314_, _05313_, _05312_);
  or _56111_ (_05315_, _05314_, _05311_);
  and _56112_ (_05316_, _04435_, _04844_);
  and _56113_ (_05317_, _04399_, _04851_);
  or _56114_ (_05318_, _05317_, _05316_);
  and _56115_ (_05319_, _04412_, _04849_);
  and _56116_ (_05320_, _04375_, _04816_);
  and _56117_ (_05321_, _04417_, _04839_);
  or _56118_ (_05322_, _05321_, _05320_);
  and _56119_ (_05323_, _04424_, _04842_);
  and _56120_ (_05324_, _04420_, _04823_);
  or _56121_ (_05325_, _05324_, _05323_);
  or _56122_ (_05326_, _05325_, _05322_);
  or _56123_ (_05327_, _05326_, _05319_);
  or _56124_ (_05328_, _05327_, _05318_);
  and _56125_ (_05329_, _04440_, _04855_);
  and _56126_ (_05330_, _04443_, _04857_);
  or _56127_ (_05332_, _05330_, _05329_);
  or _56128_ (_05333_, _05332_, _05328_);
  or _56129_ (_05335_, _05333_, _05315_);
  or _56130_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05335_, _05310_);
  and _56131_ (_05336_, _04379_, _04541_);
  and _56132_ (_05338_, _04384_, _04539_);
  or _56133_ (_05339_, _05338_, _05336_);
  and _56134_ (_05340_, _04390_, _04550_);
  and _56135_ (_05342_, _04393_, _04560_);
  or _56136_ (_05343_, _05342_, _05340_);
  or _56137_ (_05344_, _05343_, _05339_);
  and _56138_ (_05346_, _04432_, _04572_);
  and _56139_ (_05347_, _04435_, _04567_);
  and _56140_ (_05348_, _04399_, _04570_);
  or _56141_ (_05350_, _05348_, _05347_);
  or _56142_ (_05351_, _05350_, _05346_);
  and _56143_ (_05352_, _04412_, _04554_);
  and _56144_ (_05354_, _04417_, _04546_);
  and _56145_ (_05355_, _04420_, _04578_);
  or _56146_ (_05356_, _05355_, _05354_);
  and _56147_ (_05358_, _04375_, _04580_);
  and _56148_ (_05359_, _04424_, _04544_);
  or _56149_ (_05360_, _05359_, _05358_);
  or _56150_ (_05362_, _05360_, _05356_);
  or _56151_ (_05363_, _05362_, _05352_);
  and _56152_ (_05364_, _04404_, _04565_);
  and _56153_ (_05365_, _04407_, _04552_);
  or _56154_ (_05366_, _05365_, _05364_);
  or _56155_ (_05367_, _05366_, _05363_);
  and _56156_ (_05368_, _04440_, _04563_);
  and _56157_ (_05369_, _04443_, _04558_);
  or _56158_ (_05370_, _05369_, _05368_);
  or _56159_ (_05371_, _05370_, _05367_);
  or _56160_ (_05372_, _05371_, _05351_);
  or _56161_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _05372_, _05344_);
  and _56162_ (_05373_, _04440_, _04609_);
  and _56163_ (_05374_, _04393_, _04626_);
  or _56164_ (_05375_, _05374_, _05373_);
  and _56165_ (_05376_, _04390_, _04600_);
  and _56166_ (_05377_, _04384_, _04606_);
  or _56167_ (_05378_, _05377_, _05376_);
  or _56168_ (_05379_, _05378_, _05375_);
  and _56169_ (_05380_, _04407_, _04624_);
  and _56170_ (_05381_, _04432_, _04619_);
  and _56171_ (_05383_, _04399_, _04617_);
  or _56172_ (_05384_, _05383_, _05381_);
  or _56173_ (_05386_, _05384_, _05380_);
  and _56174_ (_05387_, _04412_, _04596_);
  and _56175_ (_05388_, _04417_, _04587_);
  and _56176_ (_05390_, _04420_, _04604_);
  or _56177_ (_05391_, _05390_, _05388_);
  and _56178_ (_05392_, _04375_, _04585_);
  and _56179_ (_05394_, _04424_, _04590_);
  or _56180_ (_05395_, _05394_, _05392_);
  or _56181_ (_05396_, _05395_, _05391_);
  or _56182_ (_05398_, _05396_, _05387_);
  and _56183_ (_05399_, _04404_, _04612_);
  and _56184_ (_05400_, _04435_, _04614_);
  or _56185_ (_05402_, _05400_, _05399_);
  or _56186_ (_05403_, _05402_, _05398_);
  and _56187_ (_05404_, _04379_, _04592_);
  and _56188_ (_05406_, _04443_, _04598_);
  or _56189_ (_05407_, _05406_, _05404_);
  or _56190_ (_05408_, _05407_, _05403_);
  or _56191_ (_05410_, _05408_, _05386_);
  or _56192_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _05410_, _05379_);
  and _56193_ (_05411_, _04393_, _04643_);
  and _56194_ (_05413_, _04384_, _04673_);
  or _56195_ (_05414_, _05413_, _05411_);
  and _56196_ (_05415_, _04390_, _04665_);
  and _56197_ (_05416_, _04379_, _04671_);
  or _56198_ (_05417_, _05416_, _05415_);
  or _56199_ (_05418_, _05417_, _05414_);
  and _56200_ (_05419_, _04399_, _04660_);
  and _56201_ (_05420_, _04435_, _04655_);
  and _56202_ (_05421_, _04407_, _04667_);
  or _56203_ (_05422_, _05421_, _05420_);
  or _56204_ (_05423_, _05422_, _05419_);
  and _56205_ (_05424_, _04412_, _04645_);
  and _56206_ (_05425_, _04417_, _04632_);
  and _56207_ (_05426_, _04420_, _04634_);
  or _56208_ (_05427_, _05426_, _05425_);
  and _56209_ (_05428_, _04375_, _04637_);
  and _56210_ (_05429_, _04424_, _04639_);
  or _56211_ (_05430_, _05429_, _05428_);
  or _56212_ (_05431_, _05430_, _05427_);
  or _56213_ (_05432_, _05431_, _05424_);
  and _56214_ (_05433_, _04404_, _04658_);
  and _56215_ (_05435_, _04432_, _04653_);
  or _56216_ (_05436_, _05435_, _05433_);
  or _56217_ (_05438_, _05436_, _05432_);
  and _56218_ (_05439_, _04440_, _04651_);
  and _56219_ (_05440_, _04443_, _04647_);
  or _56220_ (_05442_, _05440_, _05439_);
  or _56221_ (_05443_, _05442_, _05438_);
  or _56222_ (_05444_, _05443_, _05423_);
  or _56223_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _05444_, _05418_);
  and _56224_ (_05446_, _04379_, _04678_);
  and _56225_ (_05447_, _04384_, _04719_);
  or _56226_ (_05449_, _05447_, _05446_);
  and _56227_ (_05450_, _04390_, _04691_);
  and _56228_ (_05451_, _04393_, _04713_);
  or _56229_ (_05453_, _05451_, _05450_);
  or _56230_ (_05454_, _05453_, _05449_);
  and _56231_ (_05455_, _04435_, _04706_);
  and _56232_ (_05457_, _04404_, _04699_);
  and _56233_ (_05458_, _04399_, _04701_);
  or _56234_ (_05459_, _05458_, _05457_);
  or _56235_ (_05461_, _05459_, _05455_);
  and _56236_ (_05462_, _04412_, _04689_);
  and _56237_ (_05463_, _04417_, _04683_);
  and _56238_ (_05465_, _04420_, _04680_);
  or _56239_ (_05466_, _05465_, _05463_);
  and _56240_ (_05467_, _04375_, _04717_);
  and _56241_ (_05468_, _04424_, _04685_);
  or _56242_ (_05469_, _05468_, _05467_);
  or _56243_ (_05470_, _05469_, _05466_);
  or _56244_ (_05471_, _05470_, _05462_);
  and _56245_ (_05472_, _04432_, _04704_);
  and _56246_ (_05473_, _04407_, _04711_);
  or _56247_ (_05474_, _05473_, _05472_);
  or _56248_ (_05475_, _05474_, _05471_);
  and _56249_ (_05476_, _04440_, _04697_);
  and _56250_ (_05477_, _04443_, _04693_);
  or _56251_ (_05478_, _05477_, _05476_);
  or _56252_ (_05479_, _05478_, _05475_);
  or _56253_ (_05480_, _05479_, _05461_);
  or _56254_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _05480_, _05454_);
  and _56255_ (_05481_, _04379_, _04763_);
  and _56256_ (_05482_, _04384_, _04765_);
  or _56257_ (_05483_, _05482_, _05481_);
  and _56258_ (_05484_, _04390_, _04757_);
  and _56259_ (_05486_, _04393_, _04735_);
  or _56260_ (_05487_, _05486_, _05484_);
  or _56261_ (_05489_, _05487_, _05483_);
  and _56262_ (_05490_, _04435_, _04747_);
  and _56263_ (_05491_, _04404_, _04750_);
  and _56264_ (_05493_, _04399_, _04752_);
  or _56265_ (_05494_, _05493_, _05491_);
  or _56266_ (_05495_, _05494_, _05490_);
  and _56267_ (_05497_, _04412_, _04737_);
  and _56268_ (_05498_, _04417_, _04724_);
  and _56269_ (_05499_, _04420_, _04726_);
  or _56270_ (_05501_, _05499_, _05498_);
  and _56271_ (_05502_, _04375_, _04729_);
  and _56272_ (_05503_, _04424_, _04731_);
  or _56273_ (_05505_, _05503_, _05502_);
  or _56274_ (_05506_, _05505_, _05501_);
  or _56275_ (_05507_, _05506_, _05497_);
  and _56276_ (_05509_, _04432_, _04745_);
  and _56277_ (_05510_, _04407_, _04759_);
  or _56278_ (_05511_, _05510_, _05509_);
  or _56279_ (_05513_, _05511_, _05507_);
  and _56280_ (_05514_, _04440_, _04743_);
  and _56281_ (_05515_, _04443_, _04739_);
  or _56282_ (_05517_, _05515_, _05514_);
  or _56283_ (_05518_, _05517_, _05513_);
  or _56284_ (_05519_, _05518_, _05495_);
  or _56285_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _05519_, _05489_);
  and _56286_ (_05520_, _04390_, _04785_);
  and _56287_ (_05521_, _04393_, _04805_);
  or _56288_ (_05522_, _05521_, _05520_);
  and _56289_ (_05523_, _04379_, _04809_);
  and _56290_ (_05524_, _04384_, _04811_);
  or _56291_ (_05525_, _05524_, _05523_);
  or _56292_ (_05526_, _05525_, _05522_);
  and _56293_ (_05527_, _04435_, _04793_);
  and _56294_ (_05528_, _04404_, _04796_);
  and _56295_ (_05529_, _04407_, _04803_);
  or _56296_ (_05530_, _05529_, _05528_);
  or _56297_ (_05531_, _05530_, _05527_);
  and _56298_ (_05532_, _04412_, _04783_);
  and _56299_ (_05533_, _04375_, _04775_);
  and _56300_ (_05534_, _04417_, _04770_);
  or _56301_ (_05535_, _05534_, _05533_);
  and _56302_ (_05536_, _04424_, _04777_);
  and _56303_ (_05538_, _04420_, _04772_);
  or _56304_ (_05539_, _05538_, _05536_);
  or _56305_ (_05541_, _05539_, _05535_);
  or _56306_ (_05542_, _05541_, _05532_);
  and _56307_ (_05543_, _04432_, _04791_);
  and _56308_ (_05545_, _04399_, _04798_);
  or _56309_ (_05546_, _05545_, _05543_);
  or _56310_ (_05547_, _05546_, _05542_);
  and _56311_ (_05549_, _04440_, _04789_);
  and _56312_ (_05550_, _04443_, _04781_);
  or _56313_ (_05551_, _05550_, _05549_);
  or _56314_ (_05553_, _05551_, _05547_);
  or _56315_ (_05554_, _05553_, _05531_);
  or _56316_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _05554_, _05526_);
  and _56317_ (_05556_, _04393_, _04827_);
  and _56318_ (_05557_, _04384_, _04857_);
  or _56319_ (_05558_, _05557_, _05556_);
  and _56320_ (_05560_, _04390_, _04849_);
  and _56321_ (_05561_, _04379_, _04855_);
  or _56322_ (_05562_, _05561_, _05560_);
  or _56323_ (_05564_, _05562_, _05558_);
  and _56324_ (_05565_, _04435_, _04839_);
  and _56325_ (_05566_, _04404_, _04842_);
  and _56326_ (_05568_, _04399_, _04844_);
  or _56327_ (_05569_, _05568_, _05566_);
  or _56328_ (_05570_, _05569_, _05565_);
  and _56329_ (_05571_, _04412_, _04829_);
  and _56330_ (_05572_, _04375_, _04821_);
  and _56331_ (_05573_, _04420_, _04818_);
  or _56332_ (_05574_, _05573_, _05572_);
  and _56333_ (_05575_, _04417_, _04816_);
  and _56334_ (_05576_, _04424_, _04823_);
  or _56335_ (_05577_, _05576_, _05575_);
  or _56336_ (_05578_, _05577_, _05574_);
  or _56337_ (_05579_, _05578_, _05571_);
  and _56338_ (_05580_, _04432_, _04837_);
  and _56339_ (_05581_, _04407_, _04851_);
  or _56340_ (_05582_, _05581_, _05580_);
  or _56341_ (_05583_, _05582_, _05579_);
  and _56342_ (_05584_, _04440_, _04835_);
  and _56343_ (_05585_, _04443_, _04831_);
  or _56344_ (_05586_, _05585_, _05584_);
  or _56345_ (_05587_, _05586_, _05583_);
  or _56346_ (_05588_, _05587_, _05570_);
  or _56347_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _05588_, _05564_);
  nand _56348_ (_05590_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not _56349_ (_05592_, \oc8051_golden_model_1.PC [3]);
  or _56350_ (_05593_, \oc8051_golden_model_1.PC [2], _05592_);
  or _56351_ (_05594_, _05593_, _05590_);
  or _56352_ (_05596_, _05594_, _00459_);
  not _56353_ (_05597_, \oc8051_golden_model_1.PC [1]);
  or _56354_ (_05598_, _05597_, \oc8051_golden_model_1.PC [0]);
  or _56355_ (_05600_, _05598_, _05593_);
  or _56356_ (_05601_, _05600_, _00418_);
  and _56357_ (_05602_, _05601_, _05596_);
  not _56358_ (_05604_, \oc8051_golden_model_1.PC [2]);
  or _56359_ (_05605_, _05604_, \oc8051_golden_model_1.PC [3]);
  or _56360_ (_05606_, _05605_, _05590_);
  or _56361_ (_05608_, _05606_, _00295_);
  or _56362_ (_05609_, _05605_, _05598_);
  or _56363_ (_05610_, _05609_, _00254_);
  and _56364_ (_05612_, _05610_, _05608_);
  and _56365_ (_05613_, _05612_, _05602_);
  nand _56366_ (_05614_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _56367_ (_05616_, _05614_, _05590_);
  or _56368_ (_05617_, _05616_, _00642_);
  or _56369_ (_05618_, _05614_, _05598_);
  or _56370_ (_05620_, _05618_, _00601_);
  and _56371_ (_05621_, _05620_, _05617_);
  or _56372_ (_05622_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _56373_ (_05623_, _05622_, _05590_);
  or _56374_ (_05624_, _05623_, _00100_);
  or _56375_ (_05625_, _05622_, _05598_);
  or _56376_ (_05626_, _05625_, _00059_);
  and _56377_ (_05627_, _05626_, _05624_);
  and _56378_ (_05628_, _05627_, _05621_);
  and _56379_ (_05629_, _05628_, _05613_);
  not _56380_ (_05630_, \oc8051_golden_model_1.PC [0]);
  or _56381_ (_05631_, \oc8051_golden_model_1.PC [1], _05630_);
  or _56382_ (_05632_, _05631_, _05614_);
  or _56383_ (_05633_, _05632_, _00541_);
  or _56384_ (_05634_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or _56385_ (_05635_, _05634_, _05614_);
  or _56386_ (_05636_, _05635_, _00500_);
  and _56387_ (_05637_, _05636_, _05633_);
  or _56388_ (_05638_, _05622_, _05634_);
  or _56389_ (_05639_, _05638_, _43510_);
  or _56390_ (_05640_, _05622_, _05631_);
  or _56391_ (_05642_, _05640_, _00018_);
  and _56392_ (_05643_, _05642_, _05639_);
  and _56393_ (_05645_, _05643_, _05637_);
  or _56394_ (_05646_, _05631_, _05593_);
  or _56395_ (_05647_, _05646_, _00377_);
  or _56396_ (_05649_, _05634_, _05593_);
  or _56397_ (_05650_, _05649_, _00336_);
  and _56398_ (_05651_, _05650_, _05647_);
  or _56399_ (_05653_, _05631_, _05605_);
  or _56400_ (_05654_, _05653_, _00213_);
  or _56401_ (_05655_, _05634_, _05605_);
  or _56402_ (_05657_, _05655_, _00155_);
  and _56403_ (_05658_, _05657_, _05654_);
  and _56404_ (_05659_, _05658_, _05651_);
  and _56405_ (_05661_, _05659_, _05645_);
  nand _56406_ (_05662_, _05661_, _05629_);
  or _56407_ (_05663_, _05594_, _00424_);
  or _56408_ (_05665_, _05600_, _00383_);
  and _56409_ (_05666_, _05665_, _05663_);
  or _56410_ (_05667_, _05606_, _00260_);
  or _56411_ (_05669_, _05609_, _00219_);
  and _56412_ (_05670_, _05669_, _05667_);
  and _56413_ (_05671_, _05670_, _05666_);
  or _56414_ (_05673_, _05616_, _00607_);
  or _56415_ (_05674_, _05618_, _00550_);
  and _56416_ (_05675_, _05674_, _05673_);
  or _56417_ (_05676_, _05623_, _00065_);
  or _56418_ (_05677_, _05625_, _00024_);
  and _56419_ (_05678_, _05677_, _05676_);
  and _56420_ (_05679_, _05678_, _05675_);
  and _56421_ (_05680_, _05679_, _05671_);
  or _56422_ (_05681_, _05632_, _00506_);
  or _56423_ (_05682_, _05635_, _00465_);
  and _56424_ (_05683_, _05682_, _05681_);
  or _56425_ (_05684_, _05638_, _43475_);
  or _56426_ (_05685_, _05640_, _43516_);
  and _56427_ (_05686_, _05685_, _05684_);
  and _56428_ (_05687_, _05686_, _05683_);
  or _56429_ (_05688_, _05646_, _00342_);
  or _56430_ (_05689_, _05649_, _00301_);
  and _56431_ (_05690_, _05689_, _05688_);
  or _56432_ (_05691_, _05653_, _00168_);
  or _56433_ (_05692_, _05655_, _00106_);
  and _56434_ (_05693_, _05692_, _05691_);
  and _56435_ (_05695_, _05693_, _05690_);
  and _56436_ (_05696_, _05695_, _05687_);
  nand _56437_ (_05698_, _05696_, _05680_);
  or _56438_ (_05699_, _05698_, _05662_);
  or _56439_ (_05700_, _05594_, _00449_);
  or _56440_ (_05702_, _05600_, _00408_);
  and _56441_ (_05703_, _05702_, _05700_);
  or _56442_ (_05704_, _05606_, _00285_);
  or _56443_ (_05706_, _05609_, _00244_);
  and _56444_ (_05707_, _05706_, _05704_);
  and _56445_ (_05708_, _05707_, _05703_);
  or _56446_ (_05710_, _05616_, _00632_);
  or _56447_ (_05711_, _05618_, _00590_);
  and _56448_ (_05712_, _05711_, _05710_);
  or _56449_ (_05714_, _05623_, _00090_);
  or _56450_ (_05715_, _05625_, _00049_);
  and _56451_ (_05716_, _05715_, _05714_);
  and _56452_ (_05718_, _05716_, _05712_);
  and _56453_ (_05719_, _05718_, _05708_);
  or _56454_ (_05720_, _05632_, _00531_);
  or _56455_ (_05722_, _05635_, _00490_);
  and _56456_ (_05723_, _05722_, _05720_);
  or _56457_ (_05724_, _05638_, _43500_);
  or _56458_ (_05726_, _05640_, _00008_);
  and _56459_ (_05727_, _05726_, _05724_);
  and _56460_ (_05728_, _05727_, _05723_);
  or _56461_ (_05729_, _05646_, _00367_);
  or _56462_ (_05730_, _05649_, _00326_);
  and _56463_ (_05731_, _05730_, _05729_);
  or _56464_ (_05732_, _05653_, _00203_);
  or _56465_ (_05733_, _05655_, _00133_);
  and _56466_ (_05734_, _05733_, _05732_);
  and _56467_ (_05735_, _05734_, _05731_);
  and _56468_ (_05736_, _05735_, _05728_);
  and _56469_ (_05737_, _05736_, _05719_);
  or _56470_ (_05738_, _05594_, _00454_);
  or _56471_ (_05739_, _05600_, _00413_);
  and _56472_ (_05740_, _05739_, _05738_);
  or _56473_ (_05741_, _05606_, _00290_);
  or _56474_ (_05742_, _05609_, _00249_);
  and _56475_ (_05743_, _05742_, _05741_);
  and _56476_ (_05744_, _05743_, _05740_);
  or _56477_ (_05745_, _05616_, _00637_);
  or _56478_ (_05746_, _05618_, _00596_);
  and _56479_ (_05748_, _05746_, _05745_);
  or _56480_ (_05749_, _05623_, _00095_);
  or _56481_ (_05751_, _05625_, _00054_);
  and _56482_ (_05752_, _05751_, _05749_);
  and _56483_ (_05753_, _05752_, _05748_);
  and _56484_ (_05755_, _05753_, _05744_);
  or _56485_ (_05756_, _05632_, _00536_);
  or _56486_ (_05757_, _05635_, _00495_);
  and _56487_ (_05759_, _05757_, _05756_);
  or _56488_ (_05760_, _05638_, _43505_);
  or _56489_ (_05761_, _05640_, _00013_);
  and _56490_ (_05763_, _05761_, _05760_);
  and _56491_ (_05764_, _05763_, _05759_);
  or _56492_ (_05765_, _05646_, _00372_);
  or _56493_ (_05767_, _05649_, _00331_);
  and _56494_ (_05768_, _05767_, _05765_);
  or _56495_ (_05769_, _05653_, _00208_);
  or _56496_ (_05771_, _05655_, _00144_);
  and _56497_ (_05772_, _05771_, _05769_);
  and _56498_ (_05773_, _05772_, _05768_);
  and _56499_ (_05775_, _05773_, _05764_);
  nand _56500_ (_05776_, _05775_, _05755_);
  or _56501_ (_05777_, _05776_, _05737_);
  nor _56502_ (_05779_, _05777_, _05699_);
  or _56503_ (_05780_, _05594_, _00429_);
  or _56504_ (_05781_, _05600_, _00388_);
  and _56505_ (_05782_, _05781_, _05780_);
  or _56506_ (_05783_, _05606_, _00265_);
  or _56507_ (_05784_, _05609_, _00224_);
  and _56508_ (_05785_, _05784_, _05783_);
  and _56509_ (_05786_, _05785_, _05782_);
  or _56510_ (_05787_, _05616_, _00612_);
  or _56511_ (_05788_, _05618_, _00558_);
  and _56512_ (_05789_, _05788_, _05787_);
  or _56513_ (_05790_, _05623_, _00070_);
  or _56514_ (_05791_, _05625_, _00029_);
  and _56515_ (_05792_, _05791_, _05790_);
  and _56516_ (_05793_, _05792_, _05789_);
  and _56517_ (_05794_, _05793_, _05786_);
  or _56518_ (_05795_, _05632_, _00511_);
  or _56519_ (_05796_, _05635_, _00470_);
  and _56520_ (_05797_, _05796_, _05795_);
  or _56521_ (_05798_, _05638_, _43480_);
  or _56522_ (_05799_, _05640_, _43521_);
  and _56523_ (_05801_, _05799_, _05798_);
  and _56524_ (_05802_, _05801_, _05797_);
  or _56525_ (_05804_, _05646_, _00347_);
  or _56526_ (_05805_, _05649_, _00306_);
  and _56527_ (_05806_, _05805_, _05804_);
  or _56528_ (_05808_, _05653_, _00179_);
  or _56529_ (_05809_, _05655_, _00111_);
  and _56530_ (_05810_, _05809_, _05808_);
  and _56531_ (_05812_, _05810_, _05806_);
  and _56532_ (_05813_, _05812_, _05802_);
  and _56533_ (_05814_, _05813_, _05794_);
  or _56534_ (_05816_, _05594_, _00434_);
  or _56535_ (_05817_, _05600_, _00393_);
  and _56536_ (_05818_, _05817_, _05816_);
  or _56537_ (_05820_, _05606_, _00270_);
  or _56538_ (_05821_, _05609_, _00229_);
  and _56539_ (_05822_, _05821_, _05820_);
  and _56540_ (_05824_, _05822_, _05818_);
  or _56541_ (_05825_, _05616_, _00617_);
  or _56542_ (_05826_, _05618_, _00566_);
  and _56543_ (_05828_, _05826_, _05825_);
  or _56544_ (_05829_, _05623_, _00075_);
  or _56545_ (_05830_, _05625_, _00034_);
  and _56546_ (_05832_, _05830_, _05829_);
  and _56547_ (_05833_, _05832_, _05828_);
  and _56548_ (_05834_, _05833_, _05824_);
  or _56549_ (_05835_, _05632_, _00516_);
  or _56550_ (_05836_, _05635_, _00475_);
  and _56551_ (_05837_, _05836_, _05835_);
  or _56552_ (_05838_, _05638_, _43485_);
  or _56553_ (_05839_, _05640_, _43526_);
  and _56554_ (_05840_, _05839_, _05838_);
  and _56555_ (_05841_, _05840_, _05837_);
  or _56556_ (_05842_, _05646_, _00352_);
  or _56557_ (_05843_, _05649_, _00311_);
  and _56558_ (_05844_, _05843_, _05842_);
  or _56559_ (_05845_, _05653_, _00188_);
  or _56560_ (_05846_, _05655_, _00116_);
  and _56561_ (_05847_, _05846_, _05845_);
  and _56562_ (_05848_, _05847_, _05844_);
  and _56563_ (_05849_, _05848_, _05841_);
  nand _56564_ (_05850_, _05849_, _05834_);
  not _56565_ (_05851_, _05850_);
  and _56566_ (_05852_, _05851_, _05814_);
  or _56567_ (_05854_, _05594_, _00439_);
  or _56568_ (_05855_, _05600_, _00398_);
  and _56569_ (_05857_, _05855_, _05854_);
  or _56570_ (_05858_, _05606_, _00275_);
  or _56571_ (_05859_, _05609_, _00234_);
  and _56572_ (_05861_, _05859_, _05858_);
  and _56573_ (_05862_, _05861_, _05857_);
  or _56574_ (_05863_, _05616_, _00622_);
  or _56575_ (_05865_, _05618_, _00574_);
  and _56576_ (_05866_, _05865_, _05863_);
  or _56577_ (_05867_, _05623_, _00080_);
  or _56578_ (_05869_, _05625_, _00039_);
  and _56579_ (_05870_, _05869_, _05867_);
  and _56580_ (_05871_, _05870_, _05866_);
  and _56581_ (_05873_, _05871_, _05862_);
  or _56582_ (_05874_, _05632_, _00521_);
  or _56583_ (_05875_, _05635_, _00480_);
  and _56584_ (_05877_, _05875_, _05874_);
  or _56585_ (_05878_, _05638_, _43490_);
  or _56586_ (_05879_, _05640_, _43531_);
  and _56587_ (_05881_, _05879_, _05878_);
  and _56588_ (_05882_, _05881_, _05877_);
  or _56589_ (_05883_, _05646_, _00357_);
  or _56590_ (_05885_, _05649_, _00316_);
  and _56591_ (_05886_, _05885_, _05883_);
  or _56592_ (_05887_, _05653_, _00193_);
  or _56593_ (_05888_, _05655_, _00121_);
  and _56594_ (_05889_, _05888_, _05887_);
  and _56595_ (_05890_, _05889_, _05886_);
  and _56596_ (_05891_, _05890_, _05882_);
  nand _56597_ (_05892_, _05891_, _05873_);
  or _56598_ (_05893_, _05594_, _00444_);
  or _56599_ (_05894_, _05600_, _00403_);
  and _56600_ (_05895_, _05894_, _05893_);
  or _56601_ (_05896_, _05606_, _00280_);
  or _56602_ (_05897_, _05609_, _00239_);
  and _56603_ (_05898_, _05897_, _05896_);
  and _56604_ (_05899_, _05898_, _05895_);
  or _56605_ (_05900_, _05616_, _00627_);
  or _56606_ (_05901_, _05618_, _00582_);
  and _56607_ (_05902_, _05901_, _05900_);
  or _56608_ (_05903_, _05623_, _00085_);
  or _56609_ (_05904_, _05625_, _00044_);
  and _56610_ (_05905_, _05904_, _05903_);
  and _56611_ (_05906_, _05905_, _05902_);
  and _56612_ (_05907_, _05906_, _05899_);
  or _56613_ (_05908_, _05632_, _00526_);
  or _56614_ (_05909_, _05635_, _00485_);
  and _56615_ (_05910_, _05909_, _05908_);
  or _56616_ (_05911_, _05638_, _43495_);
  or _56617_ (_05912_, _05640_, _00003_);
  and _56618_ (_05913_, _05912_, _05911_);
  and _56619_ (_05914_, _05913_, _05910_);
  or _56620_ (_05915_, _05646_, _00362_);
  or _56621_ (_05916_, _05649_, _00321_);
  and _56622_ (_05917_, _05916_, _05915_);
  or _56623_ (_05918_, _05653_, _00198_);
  or _56624_ (_05919_, _05655_, _00126_);
  and _56625_ (_05920_, _05919_, _05918_);
  and _56626_ (_05921_, _05920_, _05917_);
  and _56627_ (_05922_, _05921_, _05914_);
  nand _56628_ (_05923_, _05922_, _05907_);
  or _56629_ (_05924_, _05923_, _05892_);
  not _56630_ (_05925_, _05924_);
  and _56631_ (_05926_, _05925_, _05852_);
  and _56632_ (_05927_, _05926_, _05779_);
  not _56633_ (_05928_, _05927_);
  nor _56634_ (_05929_, _05614_, _05597_);
  and _56635_ (_05930_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _56636_ (_05931_, _05930_, \oc8051_golden_model_1.PC [3]);
  nor _56637_ (_05932_, _05931_, _05929_);
  or _56638_ (_05933_, _05850_, _05814_);
  or _56639_ (_05934_, _05933_, _05924_);
  not _56640_ (_05935_, _05934_);
  nand _56641_ (_05936_, _05736_, _05719_);
  or _56642_ (_05937_, _05776_, _05936_);
  nor _56643_ (_05938_, _05937_, _05699_);
  and _56644_ (_05939_, _05938_, _05935_);
  and _56645_ (_05940_, _05935_, _05779_);
  nor _56646_ (_05941_, _05940_, _05939_);
  and _56647_ (_05942_, _05696_, _05680_);
  or _56648_ (_05943_, _05942_, _05662_);
  nor _56649_ (_05944_, _05943_, _05937_);
  not _56650_ (_05945_, _05944_);
  or _56651_ (_05946_, _05945_, _05934_);
  and _56652_ (_05947_, _05661_, _05629_);
  or _56653_ (_05948_, _05698_, _05947_);
  and _56654_ (_05949_, _05775_, _05755_);
  or _56655_ (_05950_, _05949_, _05737_);
  or _56656_ (_05951_, _05950_, _05948_);
  or _56657_ (_05952_, _05951_, _05934_);
  or _56658_ (_05953_, _05949_, _05936_);
  or _56659_ (_05954_, _05948_, _05953_);
  or _56660_ (_05955_, _05954_, _05934_);
  and _56661_ (_05956_, _05955_, _05952_);
  and _56662_ (_05957_, _05956_, _05946_);
  or _56663_ (_05958_, _05950_, _05699_);
  or _56664_ (_05959_, _05958_, _05934_);
  or _56665_ (_05960_, _05948_, _05777_);
  or _56666_ (_05961_, _05960_, _05934_);
  and _56667_ (_05962_, _05961_, _05959_);
  or _56668_ (_05963_, _05953_, _05699_);
  or _56669_ (_05964_, _05963_, _05934_);
  or _56670_ (_05965_, _05948_, _05937_);
  or _56671_ (_05966_, _05965_, _05934_);
  and _56672_ (_05967_, _05966_, _05964_);
  and _56673_ (_05968_, _05967_, _05962_);
  and _56674_ (_05969_, _05968_, _05957_);
  and _56675_ (_05970_, _05969_, _05941_);
  or _56676_ (_05971_, _05970_, _05932_);
  or _56677_ (_05972_, _05851_, _05814_);
  or _56678_ (_05973_, _05972_, _05924_);
  nor _56679_ (_05974_, _05973_, _05945_);
  not _56680_ (_05975_, _05974_);
  nor _56681_ (_05976_, _05943_, _05777_);
  not _56682_ (_05977_, _05976_);
  or _56683_ (_05978_, _05977_, _05934_);
  not _56684_ (_05979_, _05892_);
  or _56685_ (_05980_, _05923_, _05979_);
  or _56686_ (_05981_, _05980_, _05933_);
  or _56687_ (_05982_, _05981_, _05945_);
  and _56688_ (_05983_, _05982_, _05978_);
  or _56689_ (_05984_, _05977_, _05973_);
  and _56690_ (_05985_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  and _56691_ (_05986_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and _56692_ (_05987_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _56693_ (_05988_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _56694_ (_05989_, _05988_, _05986_);
  and _56695_ (_05990_, _05989_, _05987_);
  nor _56696_ (_05991_, _05990_, _05986_);
  nor _56697_ (_05992_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _56698_ (_05993_, _05992_, _05985_);
  not _56699_ (_05994_, _05993_);
  nor _56700_ (_05995_, _05994_, _05991_);
  nor _56701_ (_05996_, _05995_, _05985_);
  and _56702_ (_05997_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _56703_ (_05998_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _56704_ (_05999_, _05998_, _05997_);
  not _56705_ (_06000_, _05999_);
  nor _56706_ (_06001_, _06000_, _05996_);
  and _56707_ (_06002_, _06000_, _05996_);
  nor _56708_ (_06003_, _06002_, _06001_);
  not _56709_ (_06004_, _06003_);
  or _56710_ (_06005_, _06004_, _05984_);
  or _56711_ (_06006_, _05943_, _05950_);
  or _56712_ (_06007_, _06006_, _05934_);
  or _56713_ (_06008_, _05942_, _05947_);
  or _56714_ (_06009_, _06008_, _05777_);
  or _56715_ (_06010_, _06009_, _05934_);
  and _56716_ (_06011_, _06010_, _06007_);
  or _56717_ (_06012_, _06008_, _05937_);
  or _56718_ (_06013_, _06012_, _05934_);
  or _56719_ (_06014_, _06008_, _05953_);
  or _56720_ (_06015_, _06014_, _05934_);
  and _56721_ (_06016_, _06015_, _06013_);
  or _56722_ (_06017_, _06008_, _05950_);
  or _56723_ (_06018_, _06017_, _05934_);
  or _56724_ (_06019_, _05943_, _05953_);
  or _56725_ (_06020_, _06019_, _05934_);
  and _56726_ (_06021_, _06020_, _06018_);
  and _56727_ (_06022_, _06021_, _06016_);
  and _56728_ (_06023_, _06022_, _06011_);
  not _56729_ (_06024_, _05606_);
  nor _56730_ (_06025_, _05590_, _05604_);
  nor _56731_ (_06026_, _06025_, _05592_);
  nor _56732_ (_06027_, _06026_, _06024_);
  not _56733_ (_06028_, _06027_);
  and _56734_ (_06029_, _05984_, _06028_);
  nand _56735_ (_06030_, _06029_, _06023_);
  nand _56736_ (_06031_, _06030_, _06005_);
  nand _56737_ (_06032_, _06031_, _05983_);
  not _56738_ (_06033_, _05932_);
  and _56739_ (_06034_, _06023_, _05983_);
  or _56740_ (_06035_, _06034_, _06033_);
  nand _56741_ (_06036_, _06035_, _06032_);
  nand _56742_ (_06037_, _06036_, _05975_);
  not _56743_ (_06038_, _05970_);
  and _56744_ (_06039_, _05590_, _05604_);
  nor _56745_ (_06040_, _06039_, _06025_);
  and _56746_ (_06041_, _06040_, \oc8051_golden_model_1.ACC [2]);
  not _56747_ (_06042_, \oc8051_golden_model_1.ACC [1]);
  and _56748_ (_06043_, _05631_, _05598_);
  nor _56749_ (_06044_, _06043_, _06042_);
  and _56750_ (_06045_, \oc8051_golden_model_1.ACC [0], _05630_);
  and _56751_ (_06046_, _06043_, _06042_);
  nor _56752_ (_06047_, _06046_, _06044_);
  and _56753_ (_06048_, _06047_, _06045_);
  nor _56754_ (_06049_, _06048_, _06044_);
  nor _56755_ (_06050_, _06040_, \oc8051_golden_model_1.ACC [2]);
  nor _56756_ (_06051_, _06050_, _06041_);
  not _56757_ (_06052_, _06051_);
  nor _56758_ (_06053_, _06052_, _06049_);
  nor _56759_ (_06054_, _06053_, _06041_);
  not _56760_ (_06055_, \oc8051_golden_model_1.ACC [3]);
  nor _56761_ (_06056_, _06027_, _06055_);
  and _56762_ (_06057_, _06027_, _06055_);
  nor _56763_ (_06058_, _06057_, _06056_);
  and _56764_ (_06059_, _06058_, _06054_);
  nor _56765_ (_06060_, _06058_, _06054_);
  nor _56766_ (_06061_, _06060_, _06059_);
  nor _56767_ (_06062_, _06061_, _05975_);
  nor _56768_ (_06063_, _06062_, _06038_);
  nand _56769_ (_06064_, _06063_, _06037_);
  nand _56770_ (_06065_, _06064_, _05971_);
  and _56771_ (_06066_, _06052_, _06049_);
  nor _56772_ (_06067_, _06066_, _06053_);
  and _56773_ (_06068_, _06067_, _05974_);
  and _56774_ (_06069_, _05994_, _05991_);
  nor _56775_ (_06070_, _06069_, _05995_);
  not _56776_ (_06071_, _06070_);
  or _56777_ (_06072_, _06071_, _05984_);
  and _56778_ (_06073_, _06072_, _05983_);
  not _56779_ (_06074_, _06040_);
  nand _56780_ (_06075_, _06074_, _06023_);
  nand _56781_ (_06076_, _06075_, _05984_);
  nand _56782_ (_06077_, _06076_, _06073_);
  nor _56783_ (_06078_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _56784_ (_06079_, _06078_, _05930_);
  or _56785_ (_06080_, _06079_, _06034_);
  and _56786_ (_06081_, _06080_, _05975_);
  and _56787_ (_06082_, _06081_, _06077_);
  or _56788_ (_06083_, _06082_, _06068_);
  nand _56789_ (_06084_, _06083_, _05970_);
  not _56790_ (_06085_, _06079_);
  or _56791_ (_06086_, _06085_, _05970_);
  and _56792_ (_06087_, _06086_, _06084_);
  or _56793_ (_06088_, _06087_, _06065_);
  nor _56794_ (_06089_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _56795_ (_06090_, _06089_, _05987_);
  or _56796_ (_06091_, _06090_, _05984_);
  and _56797_ (_06092_, _05984_, \oc8051_golden_model_1.PC [0]);
  nand _56798_ (_06093_, _06092_, _06023_);
  nand _56799_ (_06094_, _06093_, _06091_);
  and _56800_ (_06095_, _05983_, _05975_);
  and _56801_ (_06096_, _06095_, _06094_);
  not _56802_ (_06097_, \oc8051_golden_model_1.ACC [0]);
  and _56803_ (_06098_, _06097_, \oc8051_golden_model_1.PC [0]);
  nor _56804_ (_06099_, _06098_, _06045_);
  nor _56805_ (_06100_, _06099_, _05975_);
  or _56806_ (_06101_, _06100_, _06096_);
  nand _56807_ (_06102_, _06101_, _05970_);
  nand _56808_ (_06103_, _06034_, _05970_);
  nand _56809_ (_06104_, _06103_, _05630_);
  nand _56810_ (_06105_, _06104_, _06102_);
  or _56811_ (_06106_, _06034_, \oc8051_golden_model_1.PC [1]);
  nor _56812_ (_06107_, _05989_, _05987_);
  nor _56813_ (_06108_, _06107_, _05990_);
  not _56814_ (_06109_, _06108_);
  or _56815_ (_06110_, _06109_, _05984_);
  not _56816_ (_06111_, _06043_);
  and _56817_ (_06112_, _06111_, _05984_);
  nand _56818_ (_06113_, _06112_, _06023_);
  nand _56819_ (_06114_, _06113_, _06110_);
  and _56820_ (_06115_, _05983_, _05970_);
  nand _56821_ (_06116_, _06115_, _06114_);
  nand _56822_ (_06117_, _06116_, _06106_);
  nand _56823_ (_06118_, _06117_, _05975_);
  nor _56824_ (_06119_, _06047_, _06045_);
  nor _56825_ (_06120_, _06119_, _06048_);
  and _56826_ (_06121_, _06120_, _05974_);
  nor _56827_ (_06122_, _05970_, \oc8051_golden_model_1.PC [1]);
  nor _56828_ (_06123_, _06122_, _06121_);
  and _56829_ (_06124_, _06123_, _06118_);
  or _56830_ (_06125_, _06124_, _06105_);
  or _56831_ (_06126_, _06125_, _06088_);
  or _56832_ (_06127_, _06126_, _00607_);
  nand _56833_ (_06128_, _06123_, _06118_);
  or _56834_ (_06129_, _06128_, _06105_);
  and _56835_ (_06130_, _06064_, _05971_);
  nand _56836_ (_06131_, _06086_, _06084_);
  or _56837_ (_06132_, _06131_, _06130_);
  or _56838_ (_06133_, _06132_, _06129_);
  or _56839_ (_06134_, _06133_, _43516_);
  and _56840_ (_06135_, _06134_, _06127_);
  or _56841_ (_06136_, _06131_, _06065_);
  or _56842_ (_06137_, _06136_, _06125_);
  or _56843_ (_06138_, _06137_, _00424_);
  or _56844_ (_06139_, _06132_, _06125_);
  or _56845_ (_06140_, _06139_, _00065_);
  and _56846_ (_06141_, _06140_, _06138_);
  and _56847_ (_06142_, _06141_, _06135_);
  or _56848_ (_06143_, _06136_, _06129_);
  or _56849_ (_06144_, _06143_, _00342_);
  and _56850_ (_06145_, _06104_, _06102_);
  or _56851_ (_06146_, _06124_, _06145_);
  or _56852_ (_06147_, _06132_, _06146_);
  or _56853_ (_06148_, _06147_, _00024_);
  and _56854_ (_06149_, _06148_, _06144_);
  or _56855_ (_06150_, _06087_, _06130_);
  or _56856_ (_06151_, _06150_, _06125_);
  or _56857_ (_06152_, _06151_, _00260_);
  or _56858_ (_06153_, _06150_, _06129_);
  or _56859_ (_06154_, _06153_, _00168_);
  and _56860_ (_06155_, _06154_, _06152_);
  and _56861_ (_06156_, _06155_, _06149_);
  and _56862_ (_06157_, _06156_, _06142_);
  or _56863_ (_06158_, _06128_, _06145_);
  or _56864_ (_06159_, _06150_, _06158_);
  or _56865_ (_06160_, _06159_, _00106_);
  or _56866_ (_06161_, _06132_, _06158_);
  or _56867_ (_06162_, _06161_, _43475_);
  and _56868_ (_06163_, _06162_, _06160_);
  or _56869_ (_06164_, _06146_, _06088_);
  or _56870_ (_06165_, _06164_, _00550_);
  or _56871_ (_06166_, _06136_, _06146_);
  or _56872_ (_06167_, _06166_, _00383_);
  and _56873_ (_06168_, _06167_, _06165_);
  and _56874_ (_06169_, _06168_, _06163_);
  or _56875_ (_06170_, _06129_, _06088_);
  or _56876_ (_06171_, _06170_, _00506_);
  or _56877_ (_06172_, _06158_, _06136_);
  or _56878_ (_06173_, _06172_, _00301_);
  and _56879_ (_06174_, _06173_, _06171_);
  or _56880_ (_06175_, _06158_, _06088_);
  or _56881_ (_06176_, _06175_, _00465_);
  or _56882_ (_06177_, _06150_, _06146_);
  or _56883_ (_06178_, _06177_, _00219_);
  and _56884_ (_06179_, _06178_, _06176_);
  and _56885_ (_06180_, _06179_, _06174_);
  and _56886_ (_06181_, _06180_, _06169_);
  nand _56887_ (_06182_, _06181_, _06157_);
  or _56888_ (_06183_, _06151_, _00280_);
  or _56889_ (_06184_, _06139_, _00085_);
  and _56890_ (_06185_, _06184_, _06183_);
  or _56891_ (_06186_, _06170_, _00526_);
  or _56892_ (_06187_, _06175_, _00485_);
  and _56893_ (_06188_, _06187_, _06186_);
  and _56894_ (_06189_, _06188_, _06185_);
  or _56895_ (_06190_, _06147_, _00044_);
  or _56896_ (_06191_, _06133_, _00003_);
  and _56897_ (_06192_, _06191_, _06190_);
  or _56898_ (_06193_, _06153_, _00198_);
  or _56899_ (_06194_, _06159_, _00126_);
  and _56900_ (_06195_, _06194_, _06193_);
  and _56901_ (_06196_, _06195_, _06192_);
  and _56902_ (_06197_, _06196_, _06189_);
  or _56903_ (_06198_, _06137_, _00444_);
  or _56904_ (_06199_, _06166_, _00403_);
  and _56905_ (_06200_, _06199_, _06198_);
  or _56906_ (_06201_, _06126_, _00627_);
  or _56907_ (_06202_, _06143_, _00362_);
  and _56908_ (_06203_, _06202_, _06201_);
  and _56909_ (_06204_, _06203_, _06200_);
  or _56910_ (_06205_, _06177_, _00239_);
  or _56911_ (_06206_, _06161_, _43495_);
  and _56912_ (_06207_, _06206_, _06205_);
  or _56913_ (_06208_, _06164_, _00582_);
  or _56914_ (_06209_, _06172_, _00321_);
  and _56915_ (_06210_, _06209_, _06208_);
  and _56916_ (_06211_, _06210_, _06207_);
  and _56917_ (_06212_, _06211_, _06204_);
  and _56918_ (_06213_, _06212_, _06197_);
  or _56919_ (_06214_, _06213_, _06182_);
  nor _56920_ (_06215_, _06214_, _05928_);
  nor _56921_ (_06216_, _05959_, \oc8051_golden_model_1.SP [0]);
  not _56922_ (_06217_, _05952_);
  nor _56923_ (_06218_, _05981_, _05951_);
  not _56924_ (_06219_, _06218_);
  nor _56925_ (_06220_, _06219_, _06182_);
  or _56926_ (_06221_, _06177_, _00224_);
  or _56927_ (_06222_, _06153_, _00179_);
  and _56928_ (_06223_, _06222_, _06221_);
  or _56929_ (_06224_, _06139_, _00070_);
  or _56930_ (_06225_, _06147_, _00029_);
  and _56931_ (_06226_, _06225_, _06224_);
  and _56932_ (_06227_, _06226_, _06223_);
  or _56933_ (_06228_, _06143_, _00347_);
  or _56934_ (_06229_, _06172_, _00306_);
  and _56935_ (_06230_, _06229_, _06228_);
  or _56936_ (_06231_, _06170_, _00511_);
  or _56937_ (_06232_, _06175_, _00470_);
  and _56938_ (_06233_, _06232_, _06231_);
  and _56939_ (_06234_, _06233_, _06230_);
  and _56940_ (_06235_, _06234_, _06227_);
  or _56941_ (_06236_, _06161_, _43480_);
  or _56942_ (_06237_, _06133_, _43521_);
  and _56943_ (_06238_, _06237_, _06236_);
  or _56944_ (_06239_, _06151_, _00265_);
  or _56945_ (_06240_, _06159_, _00111_);
  and _56946_ (_06241_, _06240_, _06239_);
  and _56947_ (_06242_, _06241_, _06238_);
  or _56948_ (_06243_, _06126_, _00612_);
  or _56949_ (_06244_, _06164_, _00558_);
  and _56950_ (_06245_, _06244_, _06243_);
  or _56951_ (_06246_, _06137_, _00429_);
  or _56952_ (_06247_, _06166_, _00388_);
  and _56953_ (_06248_, _06247_, _06246_);
  and _56954_ (_06249_, _06248_, _06245_);
  and _56955_ (_06250_, _06249_, _06242_);
  and _56956_ (_06251_, _06250_, _06235_);
  not _56957_ (_06252_, _06251_);
  and _56958_ (_06253_, _06252_, _06220_);
  not _56959_ (_06254_, _05978_);
  and _56960_ (_06255_, _05850_, _05814_);
  and _56961_ (_06256_, _06255_, _05925_);
  and _56962_ (_06257_, _06256_, _05976_);
  not _56963_ (_06258_, _06257_);
  nor _56964_ (_06259_, _06258_, _06214_);
  not _56965_ (_06260_, _06006_);
  and _56966_ (_06261_, _06256_, _06260_);
  not _56967_ (_06262_, _06261_);
  nor _56968_ (_06263_, _06262_, _06214_);
  nor _56969_ (_06264_, _06262_, _06182_);
  not _56970_ (_06265_, _06264_);
  not _56971_ (_06266_, _06012_);
  and _56972_ (_06267_, _06266_, _05926_);
  and _56973_ (_06268_, _06256_, _06266_);
  not _56974_ (_06269_, _06268_);
  nor _56975_ (_06270_, _06269_, _06214_);
  not _56976_ (_06271_, _06009_);
  and _56977_ (_06272_, _06256_, _06271_);
  not _56978_ (_06273_, _06272_);
  or _56979_ (_06274_, _06273_, _06214_);
  nor _56980_ (_06275_, _06273_, _06182_);
  not _56981_ (_06276_, _06018_);
  not _56982_ (_06277_, _05938_);
  nor _56983_ (_06278_, _05981_, _06277_);
  not _56984_ (_06279_, _06278_);
  not _56985_ (_06280_, _05963_);
  and _56986_ (_06281_, _06256_, _06280_);
  not _56987_ (_06282_, _06281_);
  nor _56988_ (_06283_, _05981_, _05963_);
  and _56989_ (_06284_, _06283_, _06213_);
  not _56990_ (_06285_, _06283_);
  not _56991_ (_06286_, _06182_);
  nor _56992_ (_06287_, _06151_, _00295_);
  nor _56993_ (_06288_, _06139_, _00100_);
  nor _56994_ (_06289_, _06288_, _06287_);
  nor _56995_ (_06290_, _06170_, _00541_);
  nor _56996_ (_06291_, _06175_, _00500_);
  nor _56997_ (_06292_, _06291_, _06290_);
  and _56998_ (_06293_, _06292_, _06289_);
  nor _56999_ (_06294_, _06177_, _00254_);
  nor _57000_ (_06295_, _06153_, _00213_);
  nor _57001_ (_06296_, _06295_, _06294_);
  nor _57002_ (_06297_, _06147_, _00059_);
  nor _57003_ (_06298_, _06133_, _00018_);
  nor _57004_ (_06299_, _06298_, _06297_);
  and _57005_ (_06300_, _06299_, _06296_);
  and _57006_ (_06301_, _06300_, _06293_);
  nor _57007_ (_06302_, _06137_, _00459_);
  nor _57008_ (_06303_, _06166_, _00418_);
  nor _57009_ (_06304_, _06303_, _06302_);
  nor _57010_ (_06305_, _06126_, _00642_);
  nor _57011_ (_06306_, _06172_, _00336_);
  nor _57012_ (_06307_, _06306_, _06305_);
  and _57013_ (_06308_, _06307_, _06304_);
  nor _57014_ (_06309_, _06159_, _00155_);
  nor _57015_ (_06310_, _06161_, _43510_);
  nor _57016_ (_06311_, _06310_, _06309_);
  nor _57017_ (_06312_, _06164_, _00601_);
  nor _57018_ (_06313_, _06143_, _00377_);
  nor _57019_ (_06314_, _06313_, _06312_);
  and _57020_ (_06315_, _06314_, _06311_);
  and _57021_ (_06316_, _06315_, _06308_);
  and _57022_ (_06317_, _06316_, _06301_);
  and _57023_ (_06318_, _06317_, _06286_);
  and _57024_ (_06319_, _06213_, _06182_);
  nor _57025_ (_06320_, _06319_, _06318_);
  not _57026_ (_06321_, _05951_);
  and _57027_ (_06322_, _06256_, _06321_);
  and _57028_ (_06323_, _06256_, _05944_);
  nor _57029_ (_06324_, _06323_, _06322_);
  nor _57030_ (_06325_, _06324_, _06320_);
  not _57031_ (_06326_, _05981_);
  and _57032_ (_06327_, _05923_, _05892_);
  and _57033_ (_06328_, _06327_, _06255_);
  nor _57034_ (_06329_, _06328_, _06326_);
  nor _57035_ (_06330_, _06329_, _06006_);
  not _57036_ (_06331_, _05933_);
  and _57037_ (_06332_, _06327_, _06331_);
  not _57038_ (_06333_, _06332_);
  not _57039_ (_06334_, _05972_);
  and _57040_ (_06335_, _06327_, _06334_);
  and _57041_ (_06336_, _05923_, _05979_);
  and _57042_ (_06337_, _06336_, _05852_);
  nor _57043_ (_06338_, _06337_, _06335_);
  and _57044_ (_06339_, _06338_, _06333_);
  or _57045_ (_06340_, _06339_, _06006_);
  nor _57046_ (_06341_, _06009_, _05981_);
  not _57047_ (_06342_, _05980_);
  and _57048_ (_06343_, _06255_, _06342_);
  and _57049_ (_06344_, _06343_, _06260_);
  nor _57050_ (_06345_, _05980_, _05972_);
  and _57051_ (_06346_, _06345_, _06260_);
  or _57052_ (_06347_, _06346_, _06344_);
  nor _57053_ (_06348_, _06347_, _06341_);
  and _57054_ (_06349_, _06348_, _06340_);
  and _57055_ (_06350_, _06336_, _06331_);
  and _57056_ (_06351_, _06350_, _06260_);
  not _57057_ (_06352_, _06351_);
  and _57058_ (_06353_, _06327_, _05852_);
  and _57059_ (_06354_, _06353_, _06260_);
  nand _57060_ (_06355_, _06336_, _05850_);
  nor _57061_ (_06356_, _06355_, _06006_);
  nor _57062_ (_06357_, _06356_, _06354_);
  and _57063_ (_06358_, _06357_, _06352_);
  nand _57064_ (_06359_, _06358_, _06349_);
  nor _57065_ (_06360_, _06359_, _06330_);
  and _57066_ (_06361_, _06256_, _05779_);
  and _57067_ (_06362_, _06280_, _05926_);
  nor _57068_ (_06363_, _06362_, _06361_);
  not _57069_ (_06364_, _05958_);
  and _57070_ (_06365_, _06364_, _05926_);
  nor _57071_ (_06366_, _05973_, _05965_);
  nor _57072_ (_06367_, _06366_, _06365_);
  and _57073_ (_06368_, _06367_, _06363_);
  nor _57074_ (_06369_, _05973_, _05954_);
  and _57075_ (_06370_, _06342_, _05852_);
  and _57076_ (_06371_, _06370_, _06260_);
  nor _57077_ (_06372_, _06371_, _06369_);
  and _57078_ (_06373_, _05976_, _05926_);
  not _57079_ (_06374_, _06373_);
  nor _57080_ (_06375_, _05973_, _05960_);
  nor _57081_ (_06376_, _06375_, _06218_);
  and _57082_ (_06377_, _06376_, _06374_);
  and _57083_ (_06378_, _06377_, _06372_);
  and _57084_ (_06379_, _06256_, _05938_);
  nor _57085_ (_06380_, _06379_, _05927_);
  and _57086_ (_06381_, _06380_, _06378_);
  and _57087_ (_06382_, _06381_, _06368_);
  and _57088_ (_06383_, _06382_, _06360_);
  and _57089_ (_06384_, _06383_, _05630_);
  nor _57090_ (_06385_, _06384_, _05597_);
  and _57091_ (_06386_, _06384_, _05597_);
  nor _57092_ (_06387_, _06386_, _06385_);
  nor _57093_ (_06388_, _06383_, _05630_);
  nor _57094_ (_06389_, _06388_, _06384_);
  and _57095_ (_06390_, _06389_, _06387_);
  nor _57096_ (_06391_, _06383_, _06085_);
  and _57097_ (_06392_, _06383_, _06040_);
  nor _57098_ (_06393_, _06392_, _06391_);
  nor _57099_ (_06394_, _06383_, _06033_);
  and _57100_ (_06395_, _06383_, _06028_);
  nor _57101_ (_06396_, _06395_, _06394_);
  and _57102_ (_06397_, _06396_, _06393_);
  and _57103_ (_06398_, _06397_, _06390_);
  and _57104_ (_06399_, _06398_, _04719_);
  nor _57105_ (_06400_, _06389_, _06387_);
  and _57106_ (_06401_, _06400_, _06397_);
  and _57107_ (_06402_, _06401_, _04680_);
  nor _57108_ (_06403_, _06402_, _06399_);
  nor _57109_ (_06404_, _06396_, _06393_);
  not _57110_ (_06405_, _06387_);
  nor _57111_ (_06406_, _06389_, _06405_);
  and _57112_ (_06407_, _06406_, _06404_);
  and _57113_ (_06408_, _06407_, _04699_);
  not _57114_ (_06409_, _06393_);
  nor _57115_ (_06410_, _06396_, _06409_);
  and _57116_ (_06411_, _06410_, _06406_);
  and _57117_ (_06412_, _06411_, _04697_);
  nor _57118_ (_06413_, _06412_, _06408_);
  and _57119_ (_06414_, _06413_, _06403_);
  and _57120_ (_06415_, _06410_, _06390_);
  and _57121_ (_06416_, _06415_, _04678_);
  and _57122_ (_06417_, _06410_, _06400_);
  and _57123_ (_06418_, _06417_, _04717_);
  nor _57124_ (_06419_, _06418_, _06416_);
  and _57125_ (_06420_, _06404_, _06400_);
  and _57126_ (_06421_, _06420_, _04689_);
  and _57127_ (_06422_, _06389_, _06405_);
  and _57128_ (_06423_, _06422_, _06404_);
  and _57129_ (_06424_, _06423_, _04691_);
  nor _57130_ (_06425_, _06424_, _06421_);
  and _57131_ (_06426_, _06425_, _06419_);
  and _57132_ (_06427_, _06426_, _06414_);
  and _57133_ (_06428_, _06396_, _06409_);
  and _57134_ (_06429_, _06428_, _06422_);
  and _57135_ (_06430_, _06429_, _04713_);
  and _57136_ (_06431_, _06406_, _06397_);
  and _57137_ (_06432_, _06431_, _04693_);
  nor _57138_ (_06433_, _06432_, _06430_);
  and _57139_ (_06434_, _06428_, _06390_);
  and _57140_ (_06435_, _06434_, _04701_);
  and _57141_ (_06436_, _06422_, _06397_);
  and _57142_ (_06437_, _06436_, _04685_);
  nor _57143_ (_06438_, _06437_, _06435_);
  and _57144_ (_06439_, _06438_, _06433_);
  and _57145_ (_06440_, _06404_, _06390_);
  and _57146_ (_06441_, _06440_, _04704_);
  and _57147_ (_06442_, _06422_, _06410_);
  and _57148_ (_06443_, _06442_, _04683_);
  nor _57149_ (_06444_, _06443_, _06441_);
  and _57150_ (_06445_, _06428_, _06406_);
  and _57151_ (_06446_, _06445_, _04706_);
  and _57152_ (_06447_, _06428_, _06400_);
  and _57153_ (_06448_, _06447_, _04711_);
  nor _57154_ (_06449_, _06448_, _06446_);
  and _57155_ (_06450_, _06449_, _06444_);
  and _57156_ (_06451_, _06450_, _06439_);
  and _57157_ (_06452_, _06451_, _06427_);
  nor _57158_ (_06453_, _06452_, _05982_);
  not _57159_ (_06454_, _06324_);
  and _57160_ (_06455_, _06260_, _05926_);
  nor _57161_ (_06456_, _06455_, _06261_);
  not _57162_ (_06457_, _06456_);
  and _57163_ (_06458_, _06457_, _06320_);
  nor _57164_ (_06459_, _06320_, _06273_);
  not _57165_ (_06460_, \oc8051_golden_model_1.SP [3]);
  and _57166_ (_06461_, _06271_, _05926_);
  and _57167_ (_06462_, _06461_, _06460_);
  nor _57168_ (_06463_, _06462_, _06459_);
  nor _57169_ (_06464_, _06012_, _05981_);
  not _57170_ (_06465_, _06464_);
  nor _57171_ (_06466_, _06461_, _06272_);
  not _57172_ (_06467_, _06466_);
  nor _57173_ (_06468_, _06014_, _05981_);
  nor _57174_ (_06469_, _06468_, _06341_);
  and _57175_ (_06470_, _06469_, \oc8051_golden_model_1.PSW [3]);
  or _57176_ (_06471_, _06470_, _06467_);
  and _57177_ (_06472_, _06471_, _06465_);
  not _57178_ (_06473_, _06213_);
  nand _57179_ (_06474_, _06469_, _06465_);
  and _57180_ (_06475_, _06474_, _06473_);
  or _57181_ (_06476_, _06475_, _06472_);
  and _57182_ (_06477_, _06476_, _06269_);
  and _57183_ (_06478_, _06477_, _06463_);
  and _57184_ (_06479_, _06320_, _06268_);
  nor _57185_ (_06480_, _06006_, _05981_);
  nor _57186_ (_06481_, _06480_, _06267_);
  not _57187_ (_06482_, _06481_);
  nor _57188_ (_06483_, _06482_, _06479_);
  not _57189_ (_06484_, _06483_);
  nor _57190_ (_06485_, _06484_, _06478_);
  and _57191_ (_06486_, _06482_, _06213_);
  nor _57192_ (_06487_, _06486_, _06457_);
  not _57193_ (_06488_, _06487_);
  nor _57194_ (_06489_, _06488_, _06485_);
  nor _57195_ (_06490_, _06489_, _06458_);
  not _57196_ (_06491_, _06019_);
  and _57197_ (_06492_, _06328_, _06491_);
  and _57198_ (_06493_, _06353_, _06491_);
  nor _57199_ (_06494_, _06493_, _06492_);
  and _57200_ (_06495_, _06335_, _06491_);
  and _57201_ (_06496_, _06332_, _06491_);
  nor _57202_ (_06497_, _06496_, _06495_);
  and _57203_ (_06498_, _06336_, _06491_);
  not _57204_ (_06499_, _06498_);
  and _57205_ (_06500_, _06499_, _06497_);
  and _57206_ (_06501_, _06500_, _06494_);
  not _57207_ (_06502_, _06501_);
  nor _57208_ (_06503_, _06502_, _06490_);
  and _57209_ (_06504_, _06491_, _05926_);
  and _57210_ (_06505_, _06256_, _06491_);
  nor _57211_ (_06506_, _06505_, _06504_);
  not _57212_ (_06507_, _06506_);
  nor _57213_ (_06508_, _06501_, _06213_);
  nor _57214_ (_06509_, _06508_, _06507_);
  not _57215_ (_06510_, _06509_);
  nor _57216_ (_06511_, _06510_, _06503_);
  nor _57217_ (_06512_, _05981_, _05977_);
  nor _57218_ (_06513_, _06506_, _06320_);
  nor _57219_ (_06514_, _06513_, _06512_);
  not _57220_ (_06515_, _06514_);
  nor _57221_ (_06516_, _06515_, _06511_);
  not _57222_ (_06517_, _06512_);
  nor _57223_ (_06518_, _06517_, _06213_);
  or _57224_ (_06519_, _06518_, _06516_);
  and _57225_ (_06520_, _06519_, _06258_);
  and _57226_ (_06521_, _06320_, _06257_);
  or _57227_ (_06522_, _06521_, _06520_);
  and _57228_ (_06523_, _06522_, _05982_);
  or _57229_ (_06524_, _06523_, _06454_);
  nor _57230_ (_06525_, _06524_, _06453_);
  or _57231_ (_06526_, _06525_, _06325_);
  not _57232_ (_06527_, _05965_);
  and _57233_ (_06528_, _06256_, _06527_);
  nor _57234_ (_06529_, _06528_, _06366_);
  nor _57235_ (_06530_, _05981_, _05965_);
  not _57236_ (_06531_, _06530_);
  and _57237_ (_06532_, _06531_, _06529_);
  nor _57238_ (_06533_, _05981_, _05954_);
  not _57239_ (_06534_, _06533_);
  not _57240_ (_06535_, _05954_);
  and _57241_ (_06536_, _06256_, _06535_);
  nor _57242_ (_06537_, _06536_, _06369_);
  and _57243_ (_06538_, _06537_, _06534_);
  and _57244_ (_06539_, _06538_, _06532_);
  nor _57245_ (_06540_, _05981_, _05958_);
  not _57246_ (_06541_, _06540_);
  nor _57247_ (_06542_, _05981_, _05960_);
  not _57248_ (_06543_, _06542_);
  not _57249_ (_06544_, _05960_);
  and _57250_ (_06545_, _06256_, _06544_);
  nor _57251_ (_06546_, _06545_, _06375_);
  and _57252_ (_06547_, _06546_, _06543_);
  and _57253_ (_06548_, _06547_, _06541_);
  and _57254_ (_06549_, _06548_, _06539_);
  nand _57255_ (_06550_, _06549_, _06526_);
  and _57256_ (_06551_, _06256_, _06364_);
  nor _57257_ (_06552_, _06549_, _06473_);
  nor _57258_ (_06553_, _06552_, _06551_);
  and _57259_ (_06554_, _06553_, _06550_);
  and _57260_ (_06555_, _06551_, \oc8051_golden_model_1.SP [3]);
  or _57261_ (_06556_, _06555_, _06365_);
  nor _57262_ (_06557_, _06556_, _06554_);
  not _57263_ (_06558_, _06365_);
  nor _57264_ (_06559_, _06320_, _06558_);
  or _57265_ (_06560_, _06559_, _06557_);
  and _57266_ (_06561_, _06560_, _06285_);
  or _57267_ (_06562_, _06561_, _06284_);
  nand _57268_ (_06563_, _06562_, _06282_);
  and _57269_ (_06564_, _06281_, _06460_);
  nor _57270_ (_06565_, _06564_, _06362_);
  nand _57271_ (_06566_, _06565_, _06563_);
  not _57272_ (_06567_, _05779_);
  nor _57273_ (_06568_, _05981_, _06567_);
  and _57274_ (_06569_, _06362_, _06320_);
  nor _57275_ (_06570_, _06569_, _06568_);
  nand _57276_ (_06571_, _06570_, _06566_);
  and _57277_ (_06572_, _06568_, _06213_);
  nor _57278_ (_06573_, _06572_, _05927_);
  and _57279_ (_06574_, _06573_, _06571_);
  and _57280_ (_06575_, _06320_, _05927_);
  or _57281_ (_06576_, _06575_, _06574_);
  nand _57282_ (_06577_, _06576_, _06279_);
  nor _57283_ (_06578_, _06279_, _06213_);
  not _57284_ (_06579_, _06578_);
  and _57285_ (_06580_, _06579_, _06577_);
  nor _57286_ (_06581_, _06133_, _00013_);
  nor _57287_ (_06582_, _06147_, _00054_);
  nor _57288_ (_06583_, _06582_, _06581_);
  nor _57289_ (_06584_, _06164_, _00596_);
  nor _57290_ (_06585_, _06177_, _00249_);
  nor _57291_ (_06586_, _06585_, _06584_);
  and _57292_ (_06587_, _06586_, _06583_);
  nor _57293_ (_06588_, _06137_, _00454_);
  nor _57294_ (_06589_, _06143_, _00372_);
  nor _57295_ (_06590_, _06589_, _06588_);
  nor _57296_ (_06591_, _06153_, _00208_);
  nor _57297_ (_06592_, _06161_, _43505_);
  nor _57298_ (_06593_, _06592_, _06591_);
  and _57299_ (_06594_, _06593_, _06590_);
  and _57300_ (_06595_, _06594_, _06587_);
  nor _57301_ (_06596_, _06175_, _00495_);
  nor _57302_ (_06597_, _06172_, _00331_);
  nor _57303_ (_06598_, _06597_, _06596_);
  nor _57304_ (_06599_, _06126_, _00637_);
  nor _57305_ (_06600_, _06170_, _00536_);
  nor _57306_ (_06601_, _06600_, _06599_);
  and _57307_ (_06602_, _06601_, _06598_);
  nor _57308_ (_06603_, _06166_, _00413_);
  nor _57309_ (_06604_, _06139_, _00095_);
  nor _57310_ (_06605_, _06604_, _06603_);
  nor _57311_ (_06606_, _06151_, _00290_);
  nor _57312_ (_06607_, _06159_, _00144_);
  nor _57313_ (_06608_, _06607_, _06606_);
  and _57314_ (_06609_, _06608_, _06605_);
  and _57315_ (_06610_, _06609_, _06602_);
  and _57316_ (_06611_, _06610_, _06595_);
  nor _57317_ (_06612_, _06611_, _06182_);
  not _57318_ (_06613_, _06612_);
  nor _57319_ (_06614_, _06362_, _06257_);
  and _57320_ (_06615_, _06614_, _06558_);
  and _57321_ (_06616_, _06506_, _06456_);
  nor _57322_ (_06617_, _06268_, _05927_);
  and _57323_ (_06618_, _06617_, _06324_);
  and _57324_ (_06619_, _06618_, _06616_);
  and _57325_ (_06620_, _06619_, _06615_);
  nor _57326_ (_06621_, _06620_, _06613_);
  not _57327_ (_06622_, _06621_);
  and _57328_ (_06623_, _06612_, _06272_);
  not _57329_ (_06624_, _06623_);
  nor _57330_ (_06625_, _06151_, _00275_);
  nor _57331_ (_06627_, _06139_, _00080_);
  nor _57332_ (_06628_, _06627_, _06625_);
  nor _57333_ (_06629_, _06175_, _00480_);
  nor _57334_ (_06630_, _06143_, _00357_);
  nor _57335_ (_06631_, _06630_, _06629_);
  and _57336_ (_06632_, _06631_, _06628_);
  nor _57337_ (_06633_, _06177_, _00234_);
  nor _57338_ (_06634_, _06153_, _00193_);
  nor _57339_ (_06635_, _06634_, _06633_);
  nor _57340_ (_06636_, _06161_, _43490_);
  nor _57341_ (_06637_, _06147_, _00039_);
  nor _57342_ (_06638_, _06637_, _06636_);
  and _57343_ (_06639_, _06638_, _06635_);
  and _57344_ (_06640_, _06639_, _06632_);
  nor _57345_ (_06641_, _06126_, _00622_);
  nor _57346_ (_06642_, _06164_, _00574_);
  nor _57347_ (_06643_, _06642_, _06641_);
  nor _57348_ (_06644_, _06170_, _00521_);
  nor _57349_ (_06645_, _06137_, _00439_);
  nor _57350_ (_06646_, _06645_, _06644_);
  and _57351_ (_06647_, _06646_, _06643_);
  nor _57352_ (_06648_, _06159_, _00121_);
  nor _57353_ (_06649_, _06133_, _43531_);
  nor _57354_ (_06650_, _06649_, _06648_);
  nor _57355_ (_06651_, _06166_, _00398_);
  nor _57356_ (_06652_, _06172_, _00316_);
  nor _57357_ (_06653_, _06652_, _06651_);
  and _57358_ (_06654_, _06653_, _06650_);
  and _57359_ (_06655_, _06654_, _06647_);
  and _57360_ (_06656_, _06655_, _06640_);
  not _57361_ (_06657_, _06656_);
  nand _57362_ (_06658_, _06517_, _06481_);
  nor _57363_ (_06659_, _06658_, _06474_);
  nand _57364_ (_06660_, _06659_, _06501_);
  nor _57365_ (_06661_, _06568_, _06278_);
  and _57366_ (_06662_, _06661_, _06285_);
  nand _57367_ (_06663_, _06662_, _06549_);
  or _57368_ (_06664_, _06663_, _06660_);
  and _57369_ (_06665_, _06664_, _06657_);
  not _57370_ (_06666_, _06665_);
  and _57371_ (_06667_, _06440_, _04653_);
  and _57372_ (_06668_, _06420_, _04645_);
  nor _57373_ (_06669_, _06668_, _06667_);
  and _57374_ (_06670_, _06429_, _04643_);
  and _57375_ (_06671_, _06431_, _04647_);
  nor _57376_ (_06672_, _06671_, _06670_);
  and _57377_ (_06673_, _06672_, _06669_);
  and _57378_ (_06674_, _06434_, _04660_);
  and _57379_ (_06675_, _06447_, _04667_);
  nor _57380_ (_06676_, _06675_, _06674_);
  and _57381_ (_06677_, _06398_, _04673_);
  and _57382_ (_06678_, _06401_, _04634_);
  nor _57383_ (_06679_, _06678_, _06677_);
  and _57384_ (_06680_, _06679_, _06676_);
  and _57385_ (_06681_, _06680_, _06673_);
  and _57386_ (_06682_, _06415_, _04671_);
  and _57387_ (_06683_, _06442_, _04632_);
  nor _57388_ (_06684_, _06683_, _06682_);
  and _57389_ (_06685_, _06407_, _04658_);
  and _57390_ (_06686_, _06423_, _04665_);
  nor _57391_ (_06687_, _06686_, _06685_);
  and _57392_ (_06688_, _06687_, _06684_);
  and _57393_ (_06689_, _06445_, _04655_);
  and _57394_ (_06690_, _06436_, _04639_);
  nor _57395_ (_06691_, _06690_, _06689_);
  and _57396_ (_06692_, _06411_, _04651_);
  and _57397_ (_06693_, _06417_, _04637_);
  nor _57398_ (_06694_, _06693_, _06692_);
  and _57399_ (_06695_, _06694_, _06691_);
  and _57400_ (_06696_, _06695_, _06688_);
  and _57401_ (_06697_, _06696_, _06681_);
  nor _57402_ (_06698_, _06697_, _05982_);
  nor _57403_ (_06699_, _06335_, _06328_);
  nor _57404_ (_06700_, _06699_, _06012_);
  nor _57405_ (_06701_, _06699_, _06567_);
  nor _57406_ (_06702_, _06701_, _06700_);
  and _57407_ (_06703_, _06353_, _06535_);
  not _57408_ (_06704_, _06703_);
  and _57409_ (_06705_, _06353_, _05976_);
  not _57410_ (_06706_, _06014_);
  and _57411_ (_06707_, _06353_, _06706_);
  nor _57412_ (_06708_, _06707_, _06705_);
  and _57413_ (_06709_, _06708_, _06704_);
  and _57414_ (_06710_, _06709_, _06702_);
  nor _57415_ (_06711_, _06699_, _05965_);
  nor _57416_ (_06712_, _06699_, _05960_);
  nor _57417_ (_06713_, _06712_, _06711_);
  not _57418_ (_06714_, _06713_);
  not _57419_ (_06715_, \oc8051_golden_model_1.SP [2]);
  not _57420_ (_06716_, _06551_);
  nor _57421_ (_06717_, _06461_, _06281_);
  and _57422_ (_06718_, _06717_, _06716_);
  nor _57423_ (_06719_, _06718_, _06715_);
  nor _57424_ (_06720_, _06719_, _06714_);
  and _57425_ (_06721_, _06720_, _06710_);
  or _57426_ (_06722_, _05777_, _05942_);
  nor _57427_ (_06723_, _06722_, _06699_);
  and _57428_ (_06724_, _05945_, _05954_);
  nor _57429_ (_06725_, _05936_, _05699_);
  not _57430_ (_06726_, _06725_);
  and _57431_ (_06727_, _06726_, _06724_);
  nor _57432_ (_06728_, _06727_, _06699_);
  nor _57433_ (_06729_, _06728_, _06723_);
  not _57434_ (_06730_, _06699_);
  nand _57435_ (_06731_, _06006_, _05958_);
  or _57436_ (_06732_, _06731_, _06706_);
  and _57437_ (_06733_, _06732_, _06730_);
  and _57438_ (_06734_, _06327_, _05851_);
  not _57439_ (_06735_, _06734_);
  and _57440_ (_06736_, _06006_, _05960_);
  and _57441_ (_06737_, _06736_, _05963_);
  nor _57442_ (_06738_, _06737_, _06735_);
  nor _57443_ (_06739_, _06738_, _06733_);
  and _57444_ (_06740_, _06739_, _06729_);
  and _57445_ (_06741_, _06734_, _06266_);
  and _57446_ (_06742_, _06734_, _06271_);
  nor _57447_ (_06743_, _06742_, _06741_);
  and _57448_ (_06744_, _06332_, _06535_);
  not _57449_ (_06745_, _06744_);
  and _57450_ (_06746_, _06745_, _06743_);
  and _57451_ (_06747_, _06734_, _05938_);
  or _57452_ (_06748_, _05976_, _05944_);
  and _57453_ (_06749_, _06748_, _06332_);
  nor _57454_ (_06750_, _06749_, _06747_);
  and _57455_ (_06751_, _06750_, _06746_);
  and _57456_ (_06752_, _06734_, _06364_);
  not _57457_ (_06753_, _06752_);
  and _57458_ (_06754_, _06734_, _05779_);
  and _57459_ (_06755_, _06734_, _06527_);
  nor _57460_ (_06756_, _06755_, _06754_);
  and _57461_ (_06757_, _06756_, _06753_);
  and _57462_ (_06758_, _06332_, _06706_);
  and _57463_ (_06759_, _06353_, _05944_);
  nor _57464_ (_06760_, _06759_, _06758_);
  and _57465_ (_06761_, _06760_, _06757_);
  and _57466_ (_06762_, _06761_, _06751_);
  and _57467_ (_06763_, _06762_, _06740_);
  and _57468_ (_06764_, _06763_, _06721_);
  not _57469_ (_06765_, _06764_);
  nor _57470_ (_06766_, _06765_, _06698_);
  and _57471_ (_06767_, _06766_, _06666_);
  and _57472_ (_06768_, _06767_, _06624_);
  and _57473_ (_06769_, _06768_, _06622_);
  not _57474_ (_06770_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor _57475_ (_06771_, _06279_, _06251_);
  not _57476_ (_06772_, _06771_);
  nor _57477_ (_06773_, _06506_, _06214_);
  not _57478_ (_06774_, _06480_);
  nor _57479_ (_06775_, _06774_, _06251_);
  or _57480_ (_06776_, _06465_, _06251_);
  nor _57481_ (_06777_, _06469_, _06251_);
  not _57482_ (_06778_, _06017_);
  and _57483_ (_06779_, _06343_, _06778_);
  nor _57484_ (_06780_, _06779_, _06707_);
  and _57485_ (_06781_, _06328_, _06706_);
  not _57486_ (_06782_, _06781_);
  and _57487_ (_06783_, _06343_, _06706_);
  nor _57488_ (_06784_, _06783_, _06468_);
  and _57489_ (_06785_, _06336_, _05814_);
  nand _57490_ (_06786_, _06785_, _06706_);
  and _57491_ (_06787_, _06786_, _06784_);
  and _57492_ (_06788_, _06787_, _06782_);
  and _57493_ (_06789_, _06788_, _06780_);
  and _57494_ (_06790_, _06327_, _05814_);
  not _57495_ (_06791_, _06790_);
  nor _57496_ (_06792_, _06343_, _06785_);
  and _57497_ (_06793_, _06792_, _06791_);
  nor _57498_ (_06794_, _06793_, _06009_);
  nor _57499_ (_06795_, _06794_, _06341_);
  and _57500_ (_06796_, _06795_, _06789_);
  or _57501_ (_06797_, _06796_, _06777_);
  nand _57502_ (_06798_, _06797_, _06273_);
  nand _57503_ (_06799_, _06274_, _06798_);
  not _57504_ (_06800_, \oc8051_golden_model_1.SP [0]);
  and _57505_ (_06801_, _06461_, _06800_);
  nor _57506_ (_06802_, _06801_, _06464_);
  nor _57507_ (_06803_, _06792_, _06012_);
  and _57508_ (_06804_, _06790_, _06266_);
  nor _57509_ (_06805_, _06804_, _06803_);
  and _57510_ (_06806_, _06805_, _06802_);
  nand _57511_ (_06807_, _06806_, _06799_);
  nand _57512_ (_06808_, _06807_, _06776_);
  and _57513_ (_06809_, _06808_, _06269_);
  or _57514_ (_06810_, _06270_, _06809_);
  and _57515_ (_06811_, _06267_, _06251_);
  nor _57516_ (_06812_, _06792_, _06006_);
  not _57517_ (_06813_, _06812_);
  nor _57518_ (_06814_, _06354_, _06330_);
  and _57519_ (_06815_, _06814_, _06813_);
  not _57520_ (_06816_, _06815_);
  nor _57521_ (_06817_, _06816_, _06811_);
  and _57522_ (_06818_, _06817_, _06810_);
  or _57523_ (_06819_, _06818_, _06775_);
  nand _57524_ (_06820_, _06819_, _06456_);
  nor _57525_ (_06821_, _06456_, _06214_);
  nor _57526_ (_06822_, _06821_, _06502_);
  nand _57527_ (_06823_, _06822_, _06820_);
  and _57528_ (_06824_, _06502_, _06251_);
  and _57529_ (_06825_, _06343_, _06491_);
  nor _57530_ (_06826_, _06825_, _06507_);
  not _57531_ (_06827_, _06826_);
  nor _57532_ (_06828_, _06827_, _06824_);
  and _57533_ (_06829_, _06828_, _06823_);
  nor _57534_ (_06830_, _06829_, _06773_);
  not _57535_ (_06831_, _06353_);
  and _57536_ (_06832_, _06329_, _06831_);
  and _57537_ (_06833_, _06832_, _06792_);
  nor _57538_ (_06834_, _06833_, _05977_);
  nor _57539_ (_06835_, _06834_, _06830_);
  nor _57540_ (_06836_, _06517_, _06251_);
  or _57541_ (_06837_, _06836_, _06835_);
  and _57542_ (_06838_, _06837_, _06258_);
  nor _57543_ (_06839_, _06838_, _06259_);
  nor _57544_ (_06840_, _06833_, _05945_);
  nor _57545_ (_06841_, _06840_, _06839_);
  and _57546_ (_06842_, _06401_, _04578_);
  and _57547_ (_06843_, _06398_, _04539_);
  nor _57548_ (_06844_, _06843_, _06842_);
  and _57549_ (_06845_, _06440_, _04572_);
  and _57550_ (_06846_, _06434_, _04570_);
  nor _57551_ (_06847_, _06846_, _06845_);
  and _57552_ (_06848_, _06847_, _06844_);
  and _57553_ (_06849_, _06411_, _04563_);
  and _57554_ (_06850_, _06417_, _04580_);
  nor _57555_ (_06851_, _06850_, _06849_);
  and _57556_ (_06852_, _06447_, _04552_);
  and _57557_ (_06853_, _06436_, _04544_);
  nor _57558_ (_06854_, _06853_, _06852_);
  and _57559_ (_06855_, _06854_, _06851_);
  and _57560_ (_06856_, _06855_, _06848_);
  and _57561_ (_06857_, _06423_, _04550_);
  and _57562_ (_06858_, _06442_, _04546_);
  nor _57563_ (_06859_, _06858_, _06857_);
  and _57564_ (_06860_, _06407_, _04565_);
  and _57565_ (_06861_, _06420_, _04554_);
  nor _57566_ (_06862_, _06861_, _06860_);
  and _57567_ (_06863_, _06862_, _06859_);
  and _57568_ (_06864_, _06415_, _04541_);
  and _57569_ (_06865_, _06431_, _04558_);
  nor _57570_ (_06866_, _06865_, _06864_);
  and _57571_ (_06867_, _06445_, _04567_);
  and _57572_ (_06868_, _06429_, _04560_);
  nor _57573_ (_06869_, _06868_, _06867_);
  and _57574_ (_06870_, _06869_, _06866_);
  and _57575_ (_06871_, _06870_, _06863_);
  and _57576_ (_06872_, _06871_, _06856_);
  nor _57577_ (_06873_, _06872_, _05982_);
  or _57578_ (_06874_, _06873_, _06841_);
  and _57579_ (_06875_, _06323_, _06214_);
  and _57580_ (_06876_, _06343_, _06321_);
  nor _57581_ (_06877_, _06876_, _06322_);
  not _57582_ (_06878_, _06877_);
  nor _57583_ (_06879_, _06878_, _06875_);
  and _57584_ (_06880_, _06879_, _06874_);
  not _57585_ (_06881_, _06322_);
  nor _57586_ (_06882_, _06881_, _06214_);
  or _57587_ (_06883_, _06882_, _06880_);
  and _57588_ (_06884_, _06343_, _06535_);
  not _57589_ (_06885_, _06884_);
  and _57590_ (_06886_, _06336_, _06255_);
  and _57591_ (_06887_, _06886_, _06535_);
  and _57592_ (_06888_, _06337_, _06535_);
  nor _57593_ (_06889_, _06888_, _06887_);
  and _57594_ (_06890_, _06889_, _06885_);
  and _57595_ (_06891_, _06328_, _06535_);
  nor _57596_ (_06892_, _06891_, _06703_);
  and _57597_ (_06893_, _06892_, _06890_);
  and _57598_ (_06894_, _06893_, _06883_);
  nor _57599_ (_06895_, _06538_, _06252_);
  nor _57600_ (_06896_, _06793_, _05960_);
  nor _57601_ (_06897_, _06896_, _06895_);
  and _57602_ (_06898_, _06897_, _06894_);
  nor _57603_ (_06899_, _06547_, _06252_);
  nor _57604_ (_06900_, _06793_, _05965_);
  nor _57605_ (_06901_, _06900_, _06899_);
  and _57606_ (_06902_, _06901_, _06898_);
  nor _57607_ (_06903_, _06532_, _06252_);
  nor _57608_ (_06904_, _06833_, _05958_);
  nor _57609_ (_06905_, _06904_, _06903_);
  and _57610_ (_06906_, _06905_, _06902_);
  nor _57611_ (_06907_, _06541_, _06251_);
  or _57612_ (_06908_, _06907_, _06906_);
  and _57613_ (_06909_, _06551_, _06800_);
  nor _57614_ (_06910_, _06909_, _06365_);
  and _57615_ (_06911_, _06910_, _06908_);
  nor _57616_ (_06912_, _06558_, _06214_);
  nor _57617_ (_06913_, _06912_, _06911_);
  nor _57618_ (_06914_, _06833_, _05963_);
  nor _57619_ (_06915_, _06914_, _06913_);
  nor _57620_ (_06916_, _06285_, _06251_);
  or _57621_ (_06917_, _06916_, _06915_);
  and _57622_ (_06918_, _06281_, _06800_);
  nor _57623_ (_06919_, _06918_, _06362_);
  and _57624_ (_06920_, _06919_, _06917_);
  not _57625_ (_06921_, _06362_);
  nor _57626_ (_06922_, _06921_, _06214_);
  nor _57627_ (_06923_, _06922_, _06920_);
  nor _57628_ (_06924_, _06833_, _06567_);
  nor _57629_ (_06925_, _06924_, _06923_);
  not _57630_ (_06926_, _06568_);
  nor _57631_ (_06927_, _06926_, _06251_);
  or _57632_ (_06928_, _06927_, _06925_);
  and _57633_ (_06929_, _06928_, _05928_);
  or _57634_ (_06930_, _06929_, _06215_);
  and _57635_ (_06931_, _06353_, _05938_);
  and _57636_ (_06932_, _06792_, _06329_);
  nor _57637_ (_06933_, _06932_, _06277_);
  nor _57638_ (_06934_, _06933_, _06931_);
  nand _57639_ (_06935_, _06934_, _06930_);
  nand _57640_ (_06936_, _06935_, _06772_);
  or _57641_ (_06937_, _06936_, _06770_);
  nor _57642_ (_06938_, _06126_, _00632_);
  nor _57643_ (_06939_, _06133_, _00008_);
  nor _57644_ (_06940_, _06939_, _06938_);
  nor _57645_ (_06941_, _06137_, _00449_);
  nor _57646_ (_06942_, _06161_, _43500_);
  nor _57647_ (_06943_, _06942_, _06941_);
  and _57648_ (_06944_, _06943_, _06940_);
  nor _57649_ (_06945_, _06143_, _00367_);
  nor _57650_ (_06946_, _06147_, _00049_);
  nor _57651_ (_06947_, _06946_, _06945_);
  nor _57652_ (_06948_, _06177_, _00244_);
  nor _57653_ (_06949_, _06159_, _00133_);
  nor _57654_ (_06950_, _06949_, _06948_);
  and _57655_ (_06951_, _06950_, _06947_);
  and _57656_ (_06952_, _06951_, _06944_);
  nor _57657_ (_06953_, _06153_, _00203_);
  nor _57658_ (_06954_, _06139_, _00090_);
  nor _57659_ (_06955_, _06954_, _06953_);
  nor _57660_ (_06956_, _06170_, _00531_);
  nor _57661_ (_06957_, _06166_, _00408_);
  nor _57662_ (_06958_, _06957_, _06956_);
  and _57663_ (_06959_, _06958_, _06955_);
  nor _57664_ (_06960_, _06164_, _00590_);
  nor _57665_ (_06961_, _06172_, _00326_);
  nor _57666_ (_06962_, _06961_, _06960_);
  nor _57667_ (_06963_, _06175_, _00490_);
  nor _57668_ (_06964_, _06151_, _00285_);
  nor _57669_ (_06965_, _06964_, _06963_);
  and _57670_ (_06966_, _06965_, _06962_);
  and _57671_ (_06967_, _06966_, _06959_);
  and _57672_ (_06968_, _06967_, _06952_);
  nor _57673_ (_06969_, _06968_, _06182_);
  and _57674_ (_06970_, _06620_, _06273_);
  not _57675_ (_06971_, _06970_);
  and _57676_ (_06972_, _06971_, _06969_);
  not _57677_ (_06973_, _06972_);
  nor _57678_ (_06974_, _06137_, _00434_);
  nor _57679_ (_06975_, _06166_, _00393_);
  nor _57680_ (_06976_, _06975_, _06974_);
  nor _57681_ (_06977_, _06175_, _00475_);
  nor _57682_ (_06978_, _06143_, _00352_);
  nor _57683_ (_06979_, _06978_, _06977_);
  and _57684_ (_06980_, _06979_, _06976_);
  nor _57685_ (_06981_, _06159_, _00116_);
  nor _57686_ (_06982_, _06147_, _00034_);
  nor _57687_ (_06983_, _06982_, _06981_);
  nor _57688_ (_06984_, _06151_, _00270_);
  nor _57689_ (_06985_, _06153_, _00188_);
  nor _57690_ (_06986_, _06985_, _06984_);
  and _57691_ (_06987_, _06986_, _06983_);
  and _57692_ (_06988_, _06987_, _06980_);
  nor _57693_ (_06989_, _06170_, _00516_);
  nor _57694_ (_06990_, _06161_, _43485_);
  nor _57695_ (_06991_, _06990_, _06989_);
  nor _57696_ (_06992_, _06172_, _00311_);
  nor _57697_ (_06993_, _06139_, _00075_);
  nor _57698_ (_06994_, _06993_, _06992_);
  and _57699_ (_06995_, _06994_, _06991_);
  nor _57700_ (_06996_, _06126_, _00617_);
  nor _57701_ (_06997_, _06133_, _43526_);
  nor _57702_ (_06998_, _06997_, _06996_);
  nor _57703_ (_06999_, _06164_, _00566_);
  nor _57704_ (_07000_, _06177_, _00229_);
  nor _57705_ (_07001_, _07000_, _06999_);
  and _57706_ (_07002_, _07001_, _06998_);
  and _57707_ (_07003_, _07002_, _06995_);
  and _57708_ (_07004_, _07003_, _06988_);
  not _57709_ (_07005_, _07004_);
  and _57710_ (_07006_, _07005_, _06664_);
  not _57711_ (_07007_, _07006_);
  and _57712_ (_07008_, _06407_, _04612_);
  and _57713_ (_07009_, _06440_, _04619_);
  nor _57714_ (_07010_, _07009_, _07008_);
  and _57715_ (_07011_, _06420_, _04596_);
  and _57716_ (_07012_, _06411_, _04609_);
  nor _57717_ (_07013_, _07012_, _07011_);
  and _57718_ (_07014_, _07013_, _07010_);
  and _57719_ (_07015_, _06429_, _04626_);
  and _57720_ (_07016_, _06398_, _04606_);
  nor _57721_ (_07017_, _07016_, _07015_);
  and _57722_ (_07018_, _06445_, _04614_);
  and _57723_ (_07019_, _06447_, _04624_);
  nor _57724_ (_07020_, _07019_, _07018_);
  and _57725_ (_07021_, _07020_, _07017_);
  and _57726_ (_07022_, _07021_, _07014_);
  and _57727_ (_07023_, _06442_, _04587_);
  and _57728_ (_07024_, _06436_, _04590_);
  nor _57729_ (_07025_, _07024_, _07023_);
  and _57730_ (_07026_, _06417_, _04585_);
  and _57731_ (_07027_, _06431_, _04598_);
  nor _57732_ (_07028_, _07027_, _07026_);
  and _57733_ (_07029_, _07028_, _07025_);
  and _57734_ (_07030_, _06423_, _04600_);
  and _57735_ (_07031_, _06401_, _04604_);
  nor _57736_ (_07032_, _07031_, _07030_);
  and _57737_ (_07033_, _06415_, _04592_);
  and _57738_ (_07034_, _06434_, _04617_);
  nor _57739_ (_07035_, _07034_, _07033_);
  and _57740_ (_07036_, _07035_, _07032_);
  and _57741_ (_07037_, _07036_, _07029_);
  and _57742_ (_07038_, _07037_, _07022_);
  nor _57743_ (_07039_, _07038_, _05982_);
  and _57744_ (_07040_, _06886_, _06527_);
  and _57745_ (_07041_, _06336_, _06334_);
  and _57746_ (_07042_, _07041_, _06527_);
  nor _57747_ (_07043_, _07042_, _07040_);
  and _57748_ (_07044_, _06551_, \oc8051_golden_model_1.SP [1]);
  nor _57749_ (_07045_, _06355_, _05963_);
  nor _57750_ (_07046_, _07045_, _07044_);
  nand _57751_ (_07047_, _07046_, _07043_);
  and _57752_ (_07048_, _06012_, _06009_);
  nor _57753_ (_07049_, _07048_, _06355_);
  nor _57754_ (_07050_, _06355_, _05960_);
  or _57755_ (_07051_, _07050_, _06356_);
  or _57756_ (_07052_, _07051_, _07049_);
  or _57757_ (_07053_, _07052_, _06728_);
  or _57758_ (_07054_, _07053_, _07047_);
  or _57759_ (_07055_, _05976_, _06364_);
  nor _57760_ (_07056_, _07055_, _06706_);
  and _57761_ (_07057_, _07056_, _06724_);
  nor _57762_ (_07058_, _07057_, _06355_);
  or _57763_ (_07059_, _07058_, _06714_);
  nor _57764_ (_07060_, _07059_, _07054_);
  nor _57765_ (_07061_, _06355_, _06567_);
  not _57766_ (_07062_, _07061_);
  or _57767_ (_07063_, _06355_, _06277_);
  and _57768_ (_07064_, _07063_, _07062_);
  and _57769_ (_07065_, _07064_, _06702_);
  nor _57770_ (_07066_, _06733_, _06723_);
  not _57771_ (_07067_, \oc8051_golden_model_1.SP [1]);
  nor _57772_ (_07068_, _06717_, _07067_);
  not _57773_ (_07069_, _07068_);
  and _57774_ (_07070_, _07069_, _07066_);
  and _57775_ (_07071_, _07070_, _07065_);
  and _57776_ (_07072_, _07071_, _07060_);
  not _57777_ (_07073_, _07072_);
  nor _57778_ (_07074_, _07073_, _07039_);
  and _57779_ (_07075_, _07074_, _07007_);
  and _57780_ (_07076_, _07075_, _06973_);
  not _57781_ (_07077_, \oc8051_golden_model_1.IRAM[1] [0]);
  and _57782_ (_07078_, _06935_, _06772_);
  or _57783_ (_07079_, _07078_, _07077_);
  and _57784_ (_07080_, _07079_, _07076_);
  nand _57785_ (_07081_, _07080_, _06937_);
  not _57786_ (_07082_, \oc8051_golden_model_1.IRAM[3] [0]);
  or _57787_ (_07083_, _07078_, _07082_);
  not _57788_ (_07084_, _07076_);
  not _57789_ (_07085_, \oc8051_golden_model_1.IRAM[2] [0]);
  or _57790_ (_07086_, _06936_, _07085_);
  and _57791_ (_07087_, _07086_, _07084_);
  nand _57792_ (_07088_, _07087_, _07083_);
  nand _57793_ (_07089_, _07088_, _07081_);
  nand _57794_ (_07090_, _07089_, _06769_);
  not _57795_ (_07091_, _06769_);
  not _57796_ (_07092_, \oc8051_golden_model_1.IRAM[7] [0]);
  or _57797_ (_07093_, _07078_, _07092_);
  not _57798_ (_07094_, \oc8051_golden_model_1.IRAM[6] [0]);
  or _57799_ (_07095_, _06936_, _07094_);
  and _57800_ (_07096_, _07095_, _07084_);
  nand _57801_ (_07097_, _07096_, _07093_);
  not _57802_ (_07098_, \oc8051_golden_model_1.IRAM[4] [0]);
  or _57803_ (_07099_, _06936_, _07098_);
  not _57804_ (_07100_, \oc8051_golden_model_1.IRAM[5] [0]);
  or _57805_ (_07101_, _07078_, _07100_);
  and _57806_ (_07102_, _07101_, _07076_);
  nand _57807_ (_07103_, _07102_, _07099_);
  nand _57808_ (_07104_, _07103_, _07097_);
  nand _57809_ (_07105_, _07104_, _07091_);
  nand _57810_ (_07106_, _07105_, _07090_);
  nand _57811_ (_07107_, _07106_, _06580_);
  not _57812_ (_07108_, _06580_);
  nand _57813_ (_07109_, _06936_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _57814_ (_07110_, _07078_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _57815_ (_07111_, _07110_, _07084_);
  nand _57816_ (_07112_, _07111_, _07109_);
  nand _57817_ (_07113_, _07078_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand _57818_ (_07114_, _06936_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _57819_ (_07115_, _07114_, _07076_);
  nand _57820_ (_07116_, _07115_, _07113_);
  nand _57821_ (_07117_, _07116_, _07112_);
  nand _57822_ (_07118_, _07117_, _06769_);
  not _57823_ (_07119_, \oc8051_golden_model_1.IRAM[15] [0]);
  or _57824_ (_07120_, _07078_, _07119_);
  nand _57825_ (_07121_, _07078_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _57826_ (_07122_, _07121_, _07084_);
  nand _57827_ (_07123_, _07122_, _07120_);
  not _57828_ (_07124_, \oc8051_golden_model_1.IRAM[12] [0]);
  or _57829_ (_07125_, _06936_, _07124_);
  nand _57830_ (_07126_, _06936_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _57831_ (_07127_, _07126_, _07076_);
  nand _57832_ (_07128_, _07127_, _07125_);
  nand _57833_ (_07129_, _07128_, _07123_);
  nand _57834_ (_07130_, _07129_, _07091_);
  nand _57835_ (_07131_, _07130_, _07118_);
  nand _57836_ (_07132_, _07131_, _07108_);
  and _57837_ (_07133_, _07132_, _07107_);
  and _57838_ (_07134_, _07133_, _06276_);
  nor _57839_ (_07135_, _06343_, _06337_);
  nor _57840_ (_07136_, _06370_, _05935_);
  and _57841_ (_07137_, _07136_, _07135_);
  nor _57842_ (_07138_, _07137_, _06017_);
  not _57843_ (_07139_, _07138_);
  nor _57844_ (_07140_, _07139_, _07134_);
  and _57845_ (_07141_, _06335_, _06706_);
  not _57846_ (_07142_, _07141_);
  nor _57847_ (_07143_, _07142_, _06182_);
  and _57848_ (_07144_, _07143_, _06251_);
  nor _57849_ (_07145_, _07144_, _07140_);
  and _57850_ (_07146_, _06758_, \oc8051_golden_model_1.SP [0]);
  and _57851_ (_07147_, _05923_, _05814_);
  and _57852_ (_07148_, _07147_, _06271_);
  nor _57853_ (_07149_, _07148_, _07146_);
  and _57854_ (_07150_, _07149_, _07145_);
  not _57855_ (_07151_, _06341_);
  nor _57856_ (_07152_, _07151_, _06182_);
  nor _57857_ (_07153_, _06343_, _06345_);
  nor _57858_ (_07154_, _07153_, _06009_);
  not _57859_ (_07155_, _07154_);
  nor _57860_ (_07156_, _07155_, _07133_);
  nor _57861_ (_07157_, _07156_, _07152_);
  and _57862_ (_07158_, _07157_, _07150_);
  and _57863_ (_07159_, _07152_, _06252_);
  nor _57864_ (_07160_, _07159_, _07158_);
  nor _57865_ (_07161_, _07160_, _06275_);
  not _57866_ (_07162_, _07161_);
  and _57867_ (_07163_, _07162_, _06274_);
  nor _57868_ (_07164_, _06010_, _06800_);
  nor _57869_ (_07165_, _07164_, _07163_);
  not _57870_ (_07166_, _06461_);
  nor _57871_ (_07167_, _07166_, _06182_);
  and _57872_ (_07168_, _07167_, _06251_);
  and _57873_ (_07169_, _06785_, _06266_);
  nor _57874_ (_07170_, _07169_, _06804_);
  not _57875_ (_07171_, _07170_);
  nor _57876_ (_07172_, _07171_, _07168_);
  and _57877_ (_07173_, _07172_, _07165_);
  nor _57878_ (_07174_, _07153_, _06012_);
  not _57879_ (_07175_, _07174_);
  nor _57880_ (_07176_, _07175_, _07133_);
  not _57881_ (_07177_, _07176_);
  and _57882_ (_07178_, _07177_, _07173_);
  nor _57883_ (_07179_, _06269_, _06182_);
  nor _57884_ (_07180_, _06465_, _06182_);
  and _57885_ (_07181_, _07180_, _06251_);
  nor _57886_ (_07182_, _07181_, _07179_);
  and _57887_ (_07183_, _07182_, _07178_);
  nor _57888_ (_07184_, _07183_, _06270_);
  or _57889_ (_07185_, _07184_, _06267_);
  nand _57890_ (_07186_, _06267_, _06800_);
  nand _57891_ (_07187_, _07186_, _07185_);
  and _57892_ (_07188_, _07187_, _06265_);
  nor _57893_ (_07189_, _07188_, _06263_);
  and _57894_ (_07190_, _06785_, _06491_);
  nor _57895_ (_07191_, _06007_, _06800_);
  nor _57896_ (_07192_, _07191_, _07190_);
  and _57897_ (_07193_, _07192_, _06494_);
  not _57898_ (_07194_, _07193_);
  nor _57899_ (_07195_, _07194_, _07189_);
  nor _57900_ (_07196_, _06258_, _06182_);
  nor _57901_ (_07197_, _07153_, _06019_);
  not _57902_ (_07198_, _07197_);
  nor _57903_ (_07199_, _07198_, _07133_);
  nor _57904_ (_07200_, _07199_, _07196_);
  and _57905_ (_07201_, _07200_, _07195_);
  nor _57906_ (_07202_, _07201_, _06259_);
  nor _57907_ (_07203_, _07202_, _06254_);
  nor _57908_ (_07204_, _05978_, \oc8051_golden_model_1.SP [0]);
  nor _57909_ (_07205_, _07204_, _07203_);
  and _57910_ (_07206_, _06343_, _05944_);
  and _57911_ (_07207_, _06345_, _05944_);
  nor _57912_ (_07208_, _07207_, _07206_);
  and _57913_ (_07209_, _06336_, _05851_);
  and _57914_ (_07210_, _07209_, _05944_);
  and _57915_ (_07211_, _06699_, _06333_);
  and _57916_ (_07212_, _06355_, _06831_);
  and _57917_ (_07213_, _07212_, _07211_);
  nor _57918_ (_07214_, _07213_, _05945_);
  nor _57919_ (_07215_, _07214_, _07210_);
  and _57920_ (_07216_, _07215_, _07208_);
  and _57921_ (_07217_, _07216_, _05982_);
  nor _57922_ (_07218_, _07217_, _06182_);
  and _57923_ (_07219_, _07218_, _06251_);
  and _57924_ (_07220_, _07147_, _06321_);
  nor _57925_ (_07221_, _07220_, _07219_);
  not _57926_ (_07222_, _07221_);
  nor _57927_ (_07223_, _07222_, _07205_);
  nor _57928_ (_07224_, _07153_, _05951_);
  not _57929_ (_07225_, _07224_);
  nor _57930_ (_07226_, _07225_, _07133_);
  nor _57931_ (_07227_, _07226_, _06220_);
  and _57932_ (_07228_, _07227_, _07223_);
  nor _57933_ (_07229_, _07228_, _06253_);
  nor _57934_ (_07230_, _07229_, _06217_);
  nor _57935_ (_07231_, _05952_, \oc8051_golden_model_1.SP [0]);
  nor _57936_ (_07232_, _07231_, _07230_);
  not _57937_ (_07233_, _05961_);
  not _57938_ (_07234_, _06545_);
  nor _57939_ (_07235_, _07234_, _06182_);
  not _57940_ (_07236_, _07235_);
  not _57941_ (_07237_, _06369_);
  nor _57942_ (_07238_, _07237_, _06182_);
  not _57943_ (_07239_, _07238_);
  not _57944_ (_07240_, _06536_);
  nor _57945_ (_07241_, _07240_, _06182_);
  not _57946_ (_07242_, _06375_);
  nor _57947_ (_07243_, _07242_, _06182_);
  nor _57948_ (_07244_, _07243_, _07241_);
  and _57949_ (_07245_, _07244_, _07239_);
  and _57950_ (_07246_, _07245_, _07236_);
  nor _57951_ (_07247_, _07246_, _06252_);
  nor _57952_ (_07248_, _07247_, _07233_);
  not _57953_ (_07249_, _07248_);
  nor _57954_ (_07250_, _07249_, _07232_);
  nor _57955_ (_07251_, _05961_, \oc8051_golden_model_1.SP [0]);
  nor _57956_ (_07252_, _07251_, _07250_);
  not _57957_ (_07253_, _05959_);
  nor _57958_ (_07254_, _06529_, _06182_);
  and _57959_ (_07255_, _07254_, _06251_);
  or _57960_ (_07256_, _07255_, _07253_);
  nor _57961_ (_07257_, _07256_, _07252_);
  nor _57962_ (_07258_, _07257_, _06216_);
  and _57963_ (_07259_, _07147_, _05779_);
  nor _57964_ (_07260_, _07259_, _07258_);
  nor _57965_ (_07261_, _06926_, _06182_);
  and _57966_ (_07262_, _06343_, _05779_);
  and _57967_ (_07263_, _06345_, _05779_);
  nor _57968_ (_07264_, _07263_, _07262_);
  nor _57969_ (_07265_, _07264_, _07133_);
  nor _57970_ (_07266_, _07265_, _07261_);
  and _57971_ (_07267_, _07266_, _07260_);
  and _57972_ (_07268_, _07261_, _06252_);
  nor _57973_ (_07269_, _07268_, _07267_);
  nor _57974_ (_07270_, _06182_, _05928_);
  nor _57975_ (_07271_, _06361_, _05940_);
  nor _57976_ (_07272_, _07271_, _06800_);
  nor _57977_ (_07273_, _07272_, _07270_);
  not _57978_ (_07274_, _07273_);
  nor _57979_ (_07275_, _07274_, _07269_);
  nor _57980_ (_07276_, _07275_, _06215_);
  and _57981_ (_07277_, _07147_, _05938_);
  nor _57982_ (_07278_, _07277_, _07276_);
  and _57983_ (_07279_, _06343_, _05938_);
  and _57984_ (_07280_, _06345_, _05938_);
  or _57985_ (_07281_, _07280_, _07279_);
  not _57986_ (_07282_, _07281_);
  nor _57987_ (_07283_, _07282_, _07133_);
  not _57988_ (_07284_, _07283_);
  and _57989_ (_07285_, _07284_, _07278_);
  nor _57990_ (_07286_, _06279_, _06182_);
  and _57991_ (_07287_, _07286_, _06251_);
  not _57992_ (_07288_, _07287_);
  and _57993_ (_07289_, _07288_, _07285_);
  and _57994_ (_07290_, _07286_, _07005_);
  and _57995_ (_07291_, _06969_, _05927_);
  and _57996_ (_07292_, _07209_, _05779_);
  nor _57997_ (_07293_, _07292_, _06754_);
  not _57998_ (_07294_, _07293_);
  and _57999_ (_07295_, _07067_, \oc8051_golden_model_1.SP [0]);
  and _58000_ (_07296_, \oc8051_golden_model_1.SP [1], _06800_);
  nor _58001_ (_07297_, _07296_, _07295_);
  nor _58002_ (_07298_, _07297_, _05959_);
  and _58003_ (_07299_, _07005_, _06220_);
  and _58004_ (_07300_, _06969_, _06257_);
  not _58005_ (_07301_, _07297_);
  and _58006_ (_07302_, _07301_, _06267_);
  not _58007_ (_07303_, _06267_);
  nor _58008_ (_07304_, _07153_, _06017_);
  not _58009_ (_07305_, \oc8051_golden_model_1.IRAM[0] [1]);
  or _58010_ (_07306_, _06936_, _07305_);
  not _58011_ (_07307_, \oc8051_golden_model_1.IRAM[1] [1]);
  or _58012_ (_07308_, _07078_, _07307_);
  and _58013_ (_07309_, _07308_, _07076_);
  nand _58014_ (_07310_, _07309_, _07306_);
  not _58015_ (_07311_, \oc8051_golden_model_1.IRAM[3] [1]);
  or _58016_ (_07312_, _07078_, _07311_);
  not _58017_ (_07313_, \oc8051_golden_model_1.IRAM[2] [1]);
  or _58018_ (_07314_, _06936_, _07313_);
  and _58019_ (_07315_, _07314_, _07084_);
  nand _58020_ (_07316_, _07315_, _07312_);
  nand _58021_ (_07317_, _07316_, _07310_);
  nand _58022_ (_07318_, _07317_, _06769_);
  not _58023_ (_07319_, \oc8051_golden_model_1.IRAM[7] [1]);
  or _58024_ (_07320_, _07078_, _07319_);
  not _58025_ (_07321_, \oc8051_golden_model_1.IRAM[6] [1]);
  or _58026_ (_07322_, _06936_, _07321_);
  and _58027_ (_07323_, _07322_, _07084_);
  nand _58028_ (_07324_, _07323_, _07320_);
  not _58029_ (_07325_, \oc8051_golden_model_1.IRAM[4] [1]);
  or _58030_ (_07326_, _06936_, _07325_);
  not _58031_ (_07327_, \oc8051_golden_model_1.IRAM[5] [1]);
  or _58032_ (_07328_, _07078_, _07327_);
  and _58033_ (_07329_, _07328_, _07076_);
  nand _58034_ (_07330_, _07329_, _07326_);
  nand _58035_ (_07331_, _07330_, _07324_);
  nand _58036_ (_07332_, _07331_, _07091_);
  nand _58037_ (_07333_, _07332_, _07318_);
  nand _58038_ (_07334_, _07333_, _06580_);
  nand _58039_ (_07335_, _06936_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _58040_ (_07336_, _07078_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _58041_ (_07337_, _07336_, _07084_);
  nand _58042_ (_07338_, _07337_, _07335_);
  nand _58043_ (_07339_, _07078_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand _58044_ (_07340_, _06936_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _58045_ (_07341_, _07340_, _07076_);
  nand _58046_ (_07342_, _07341_, _07339_);
  nand _58047_ (_07343_, _07342_, _07338_);
  nand _58048_ (_07344_, _07343_, _06769_);
  nand _58049_ (_07345_, _06936_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _58050_ (_07346_, _07078_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _58051_ (_07347_, _07346_, _07084_);
  nand _58052_ (_07348_, _07347_, _07345_);
  nand _58053_ (_07349_, _07078_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand _58054_ (_07350_, _06936_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _58055_ (_07351_, _07350_, _07076_);
  nand _58056_ (_07352_, _07351_, _07349_);
  nand _58057_ (_07353_, _07352_, _07348_);
  nand _58058_ (_07354_, _07353_, _07091_);
  nand _58059_ (_07355_, _07354_, _07344_);
  nand _58060_ (_07356_, _07355_, _07108_);
  nand _58061_ (_07357_, _07356_, _07334_);
  and _58062_ (_07358_, _07357_, _06276_);
  or _58063_ (_07359_, _07358_, _07304_);
  and _58064_ (_07360_, _07143_, _07004_);
  or _58065_ (_07361_, _07360_, _07359_);
  and _58066_ (_07362_, _07297_, _06758_);
  not _58067_ (_07363_, _07362_);
  and _58068_ (_07364_, _07209_, _06271_);
  nor _58069_ (_07365_, _07364_, _06742_);
  and _58070_ (_07366_, _07365_, _07363_);
  not _58071_ (_07367_, _07366_);
  nor _58072_ (_07368_, _07367_, _07361_);
  and _58073_ (_07369_, _07357_, _07154_);
  nor _58074_ (_07370_, _07369_, _07152_);
  and _58075_ (_07371_, _07370_, _07368_);
  and _58076_ (_07372_, _07152_, _07005_);
  nor _58077_ (_07373_, _07372_, _07371_);
  and _58078_ (_07374_, _06968_, _06275_);
  nor _58079_ (_07375_, _07374_, _07373_);
  or _58080_ (_07376_, _07301_, _06010_);
  nand _58081_ (_07377_, _07376_, _07375_);
  and _58082_ (_07378_, _07167_, _07004_);
  and _58083_ (_07379_, _07209_, _06266_);
  nor _58084_ (_07380_, _07379_, _06741_);
  not _58085_ (_07381_, _07380_);
  nor _58086_ (_07382_, _07381_, _07378_);
  not _58087_ (_07383_, _07382_);
  nor _58088_ (_07384_, _07383_, _07377_);
  and _58089_ (_07385_, _07357_, _07174_);
  nor _58090_ (_07386_, _07385_, _07180_);
  and _58091_ (_07387_, _07386_, _07384_);
  and _58092_ (_07388_, _07180_, _07005_);
  nor _58093_ (_07389_, _07388_, _07387_);
  and _58094_ (_07390_, _06968_, _07179_);
  nor _58095_ (_07391_, _07390_, _07389_);
  and _58096_ (_07392_, _07391_, _07303_);
  nor _58097_ (_07393_, _07392_, _07302_);
  and _58098_ (_07394_, _06968_, _06264_);
  or _58099_ (_07395_, _07394_, _07393_);
  nor _58100_ (_07396_, _07301_, _06007_);
  not _58101_ (_07397_, _07396_);
  and _58102_ (_07398_, _07209_, _06491_);
  and _58103_ (_07399_, _06734_, _06491_);
  nor _58104_ (_07400_, _07399_, _07398_);
  and _58105_ (_07401_, _07400_, _07397_);
  not _58106_ (_07402_, _07401_);
  nor _58107_ (_07403_, _07402_, _07395_);
  and _58108_ (_07404_, _07357_, _07197_);
  nor _58109_ (_07405_, _07404_, _07196_);
  and _58110_ (_07406_, _07405_, _07403_);
  nor _58111_ (_07407_, _07406_, _07300_);
  nor _58112_ (_07408_, _07407_, _06254_);
  nor _58113_ (_07409_, _07297_, _05978_);
  nor _58114_ (_07410_, _07409_, _07408_);
  and _58115_ (_07411_, _07218_, _07004_);
  nor _58116_ (_07412_, _05951_, _05850_);
  and _58117_ (_07413_, _07412_, _05923_);
  nor _58118_ (_07414_, _07413_, _07411_);
  not _58119_ (_07415_, _07414_);
  nor _58120_ (_07416_, _07415_, _07410_);
  and _58121_ (_07417_, _07357_, _07224_);
  nor _58122_ (_07418_, _07417_, _06220_);
  and _58123_ (_07419_, _07418_, _07416_);
  nor _58124_ (_07420_, _07419_, _07299_);
  nor _58125_ (_07421_, _07420_, _06217_);
  nor _58126_ (_07422_, _07297_, _05952_);
  nor _58127_ (_07423_, _07422_, _07421_);
  nor _58128_ (_07424_, _07246_, _07005_);
  nor _58129_ (_07425_, _07424_, _07233_);
  not _58130_ (_07426_, _07425_);
  nor _58131_ (_07427_, _07426_, _07423_);
  nor _58132_ (_07428_, _07297_, _05961_);
  nor _58133_ (_07429_, _07428_, _07427_);
  and _58134_ (_07430_, _07254_, _07004_);
  or _58135_ (_07431_, _07430_, _07253_);
  nor _58136_ (_07432_, _07431_, _07429_);
  nor _58137_ (_07433_, _07432_, _07298_);
  nor _58138_ (_07434_, _07433_, _07294_);
  not _58139_ (_07435_, _07264_);
  and _58140_ (_07436_, _07357_, _07435_);
  nor _58141_ (_07437_, _07436_, _07261_);
  and _58142_ (_07438_, _07437_, _07434_);
  and _58143_ (_07439_, _07261_, _07005_);
  nor _58144_ (_07440_, _07439_, _07438_);
  nor _58145_ (_07441_, _07301_, _07271_);
  nor _58146_ (_07442_, _07441_, _07270_);
  not _58147_ (_07443_, _07442_);
  nor _58148_ (_07444_, _07443_, _07440_);
  nor _58149_ (_07445_, _07444_, _07291_);
  and _58150_ (_07446_, _07209_, _05938_);
  nor _58151_ (_07447_, _07446_, _06747_);
  not _58152_ (_07448_, _07447_);
  nor _58153_ (_07449_, _07448_, _07445_);
  and _58154_ (_07450_, _07357_, _07281_);
  nor _58155_ (_07451_, _07450_, _07286_);
  and _58156_ (_07452_, _07451_, _07449_);
  nor _58157_ (_07453_, _07452_, _07290_);
  not _58158_ (_07454_, _01354_);
  nor _58159_ (_07455_, _07211_, _05945_);
  not _58160_ (_07456_, _07455_);
  not _58161_ (_07457_, _06759_);
  nor _58162_ (_07458_, _07210_, _07141_);
  and _58163_ (_07459_, _07458_, _07457_);
  not _58164_ (_07460_, _07208_);
  nor _58165_ (_07461_, _06355_, _05945_);
  nor _58166_ (_07462_, _07461_, _07460_);
  and _58167_ (_07463_, _07462_, _07459_);
  and _58168_ (_07464_, _07463_, _07456_);
  nor _58169_ (_07465_, _07464_, _06182_);
  nor _58170_ (_07466_, _07465_, _07235_);
  nor _58171_ (_07467_, _07167_, _06264_);
  and _58172_ (_07468_, _07467_, _07466_);
  nor _58173_ (_07469_, _07180_, _07179_);
  nor _58174_ (_07470_, _06182_, _05982_);
  not _58175_ (_07471_, _07470_);
  and _58176_ (_07472_, _07412_, _06785_);
  nor _58177_ (_07473_, _07472_, _06492_);
  and _58178_ (_07474_, _07264_, _07175_);
  and _58179_ (_07475_, _07474_, _07473_);
  not _58180_ (_07476_, _07049_);
  and _58181_ (_07477_, _07476_, _06743_);
  nor _58182_ (_07478_, _07281_, _07154_);
  and _58183_ (_07479_, _07478_, _07477_);
  and _58184_ (_07480_, _07479_, _07475_);
  not _58185_ (_07481_, _07209_);
  and _58186_ (_07482_, _07153_, _07481_);
  nor _58187_ (_07483_, _07482_, _06017_);
  nand _58188_ (_07484_, _07136_, _05981_);
  and _58189_ (_07485_, _07484_, _06778_);
  or _58190_ (_07486_, _07485_, _07483_);
  not _58191_ (_07487_, _07486_);
  nor _58192_ (_07488_, _07197_, _06493_);
  and _58193_ (_07489_, _07488_, _07225_);
  and _58194_ (_07490_, _07489_, _07487_);
  and _58195_ (_07491_, _07490_, _07480_);
  and _58196_ (_07492_, _06350_, _06321_);
  not _58197_ (_07493_, _07492_);
  and _58198_ (_07494_, _06007_, _05978_);
  and _58199_ (_07495_, _06010_, _05952_);
  and _58200_ (_07496_, _07495_, _07494_);
  and _58201_ (_07497_, _07496_, _07493_);
  nor _58202_ (_07498_, _06699_, _06009_);
  not _58203_ (_07499_, _07498_);
  and _58204_ (_07500_, _07499_, _06497_);
  and _58205_ (_07501_, _07500_, _07497_);
  nor _58206_ (_07502_, _07364_, _07398_);
  and _58207_ (_07503_, _07502_, _07293_);
  not _58208_ (_07504_, _06758_);
  and _58209_ (_07505_, _07041_, _06491_);
  nor _58210_ (_07506_, _07446_, _07505_);
  and _58211_ (_07507_, _07506_, _07504_);
  and _58212_ (_07508_, _07507_, _07503_);
  and _58213_ (_07509_, _07271_, _05962_);
  and _58214_ (_07510_, _06327_, _05938_);
  nor _58215_ (_07511_, _07510_, _06267_);
  and _58216_ (_07512_, _06886_, _06491_);
  nor _58217_ (_07513_, _07379_, _07512_);
  and _58218_ (_07514_, _07513_, _07511_);
  and _58219_ (_07515_, _07514_, _07509_);
  and _58220_ (_07516_, _07515_, _07508_);
  and _58221_ (_07517_, _07516_, _07501_);
  nor _58222_ (_07518_, _07213_, _05951_);
  not _58223_ (_07519_, _07518_);
  and _58224_ (_07520_, _07519_, _07065_);
  and _58225_ (_07521_, _07520_, _07517_);
  and _58226_ (_07522_, _07521_, _07491_);
  and _58227_ (_07523_, _07522_, _07471_);
  and _58228_ (_07524_, _07523_, _07469_);
  and _58229_ (_07525_, _07524_, _07468_);
  nor _58230_ (_07526_, _07261_, _06220_);
  nor _58231_ (_07527_, _07254_, _07196_);
  and _58232_ (_07528_, _07527_, _07526_);
  nor _58233_ (_07529_, _07286_, _07270_);
  nor _58234_ (_07530_, _07152_, _06275_);
  and _58235_ (_07531_, _07530_, _07529_);
  and _58236_ (_07532_, _07531_, _07528_);
  and _58237_ (_07533_, _07532_, _07245_);
  and _58238_ (_07534_, _07533_, _07525_);
  nor _58239_ (_07535_, _07534_, _07454_);
  not _58240_ (_07536_, _07535_);
  nor _58241_ (_07537_, _07536_, _07453_);
  and _58242_ (_07538_, _07537_, _07289_);
  not _58243_ (_07539_, _07270_);
  or _58244_ (_07540_, _07539_, _06318_);
  or _58245_ (_07541_, _07153_, _06567_);
  not _58246_ (_07542_, \oc8051_golden_model_1.IRAM[0] [3]);
  or _58247_ (_07543_, _06936_, _07542_);
  not _58248_ (_07544_, \oc8051_golden_model_1.IRAM[1] [3]);
  or _58249_ (_07545_, _07078_, _07544_);
  and _58250_ (_07546_, _07545_, _07076_);
  nand _58251_ (_07547_, _07546_, _07543_);
  not _58252_ (_07548_, \oc8051_golden_model_1.IRAM[3] [3]);
  or _58253_ (_07549_, _07078_, _07548_);
  not _58254_ (_07550_, \oc8051_golden_model_1.IRAM[2] [3]);
  or _58255_ (_07551_, _06936_, _07550_);
  and _58256_ (_07552_, _07551_, _07084_);
  nand _58257_ (_07553_, _07552_, _07549_);
  nand _58258_ (_07554_, _07553_, _07547_);
  nand _58259_ (_07555_, _07554_, _06769_);
  not _58260_ (_07556_, \oc8051_golden_model_1.IRAM[7] [3]);
  or _58261_ (_07557_, _07078_, _07556_);
  not _58262_ (_07558_, \oc8051_golden_model_1.IRAM[6] [3]);
  or _58263_ (_07559_, _06936_, _07558_);
  and _58264_ (_07560_, _07559_, _07084_);
  nand _58265_ (_07561_, _07560_, _07557_);
  not _58266_ (_07562_, \oc8051_golden_model_1.IRAM[4] [3]);
  or _58267_ (_07563_, _06936_, _07562_);
  not _58268_ (_07564_, \oc8051_golden_model_1.IRAM[5] [3]);
  or _58269_ (_07565_, _07078_, _07564_);
  and _58270_ (_07566_, _07565_, _07076_);
  nand _58271_ (_07567_, _07566_, _07563_);
  nand _58272_ (_07568_, _07567_, _07561_);
  nand _58273_ (_07569_, _07568_, _07091_);
  nand _58274_ (_07570_, _07569_, _07555_);
  nand _58275_ (_07571_, _07570_, _06580_);
  nand _58276_ (_07572_, _06936_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _58277_ (_07573_, _07078_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _58278_ (_07574_, _07573_, _07084_);
  nand _58279_ (_07575_, _07574_, _07572_);
  nand _58280_ (_07576_, _07078_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand _58281_ (_07577_, _06936_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _58282_ (_07578_, _07577_, _07076_);
  nand _58283_ (_07579_, _07578_, _07576_);
  nand _58284_ (_07580_, _07579_, _07575_);
  nand _58285_ (_07581_, _07580_, _06769_);
  nand _58286_ (_07582_, _06936_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _58287_ (_07583_, _07078_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _58288_ (_07584_, _07583_, _07084_);
  nand _58289_ (_07585_, _07584_, _07582_);
  nand _58290_ (_07586_, _07078_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand _58291_ (_07587_, _06936_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _58292_ (_07588_, _07587_, _07076_);
  nand _58293_ (_07589_, _07588_, _07586_);
  nand _58294_ (_07590_, _07589_, _07585_);
  nand _58295_ (_07591_, _07590_, _07091_);
  nand _58296_ (_07592_, _07591_, _07581_);
  nand _58297_ (_07593_, _07592_, _07108_);
  nand _58298_ (_07594_, _07593_, _07571_);
  not _58299_ (_07595_, _07594_);
  or _58300_ (_07596_, _07595_, _07541_);
  and _58301_ (_07597_, _07594_, _07224_);
  and _58302_ (_07598_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _58303_ (_07599_, _07598_, \oc8051_golden_model_1.SP [2]);
  nor _58304_ (_07600_, _07599_, \oc8051_golden_model_1.SP [3]);
  and _58305_ (_07601_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _58306_ (_07602_, _07601_, \oc8051_golden_model_1.SP [3]);
  and _58307_ (_07603_, _07602_, \oc8051_golden_model_1.SP [0]);
  nor _58308_ (_07604_, _07603_, _07600_);
  not _58309_ (_07605_, _07604_);
  nor _58310_ (_07606_, _07605_, _05978_);
  not _58311_ (_07607_, _06317_);
  and _58312_ (_07608_, _07607_, _07196_);
  and _58313_ (_07609_, _07594_, _07197_);
  nor _58314_ (_07610_, _07605_, _06007_);
  not _58315_ (_07611_, _06010_);
  and _58316_ (_07612_, _07594_, _07154_);
  and _58317_ (_07613_, _07604_, _06758_);
  and _58318_ (_07614_, _07594_, _06276_);
  not _58319_ (_07615_, \oc8051_golden_model_1.PSW [3]);
  and _58320_ (_07616_, _06018_, _07615_);
  nor _58321_ (_07617_, _07616_, _07614_);
  nor _58322_ (_07618_, _07617_, _07143_);
  and _58323_ (_07619_, _07143_, _06213_);
  nor _58324_ (_07620_, _07619_, _06758_);
  not _58325_ (_07621_, _07620_);
  nor _58326_ (_07622_, _07621_, _07618_);
  or _58327_ (_07623_, _07622_, _07154_);
  nor _58328_ (_07624_, _07623_, _07613_);
  or _58329_ (_07625_, _07624_, _07152_);
  nor _58330_ (_07626_, _07625_, _07612_);
  and _58331_ (_07627_, _07152_, _06473_);
  or _58332_ (_07628_, _07627_, _06275_);
  nor _58333_ (_07629_, _07628_, _07626_);
  and _58334_ (_07630_, _06318_, _06272_);
  nor _58335_ (_07631_, _07630_, _07629_);
  nor _58336_ (_07632_, _07631_, _07611_);
  nor _58337_ (_07633_, _07604_, _06010_);
  nor _58338_ (_07634_, _07633_, _07167_);
  not _58339_ (_07635_, _07634_);
  nor _58340_ (_07636_, _07635_, _07632_);
  and _58341_ (_07637_, _07167_, _06473_);
  nor _58342_ (_07638_, _07637_, _07174_);
  not _58343_ (_07639_, _07638_);
  nor _58344_ (_07640_, _07639_, _07636_);
  and _58345_ (_07641_, _07594_, _07174_);
  nor _58346_ (_07642_, _07641_, _07180_);
  not _58347_ (_07643_, _07642_);
  nor _58348_ (_07644_, _07643_, _07640_);
  and _58349_ (_07645_, _07180_, _06473_);
  nor _58350_ (_07646_, _07645_, _07179_);
  not _58351_ (_07647_, _07646_);
  nor _58352_ (_07648_, _07647_, _07644_);
  and _58353_ (_07649_, _06318_, _07179_);
  nor _58354_ (_07650_, _07649_, _07648_);
  and _58355_ (_07651_, _07650_, _07303_);
  and _58356_ (_07652_, _07604_, _06267_);
  nor _58357_ (_07653_, _07652_, _07651_);
  nor _58358_ (_07654_, _07653_, _06264_);
  and _58359_ (_07655_, _06264_, _06320_);
  or _58360_ (_07656_, _07655_, _07654_);
  and _58361_ (_07657_, _07656_, _06007_);
  or _58362_ (_07658_, _07657_, _07197_);
  nor _58363_ (_07659_, _07658_, _07610_);
  or _58364_ (_07660_, _07659_, _07196_);
  nor _58365_ (_07661_, _07660_, _07609_);
  nor _58366_ (_07662_, _07661_, _07608_);
  nor _58367_ (_07663_, _07662_, _06254_);
  nor _58368_ (_07664_, _07663_, _07606_);
  or _58369_ (_07665_, _07664_, _07218_);
  nand _58370_ (_07666_, _07218_, _06473_);
  and _58371_ (_07667_, _07666_, _07225_);
  and _58372_ (_07668_, _07667_, _07665_);
  or _58373_ (_07669_, _07668_, _06220_);
  nor _58374_ (_07670_, _07669_, _07597_);
  nor _58375_ (_07671_, _06219_, _06214_);
  nor _58376_ (_07672_, _07671_, _07670_);
  nor _58377_ (_07673_, _07672_, _06217_);
  nor _58378_ (_07674_, _07605_, _05952_);
  not _58379_ (_07675_, _07674_);
  and _58380_ (_07676_, _07675_, _07246_);
  not _58381_ (_07677_, _07676_);
  nor _58382_ (_07678_, _07677_, _07673_);
  nor _58383_ (_07679_, _07246_, _06473_);
  nor _58384_ (_07680_, _07679_, _07233_);
  not _58385_ (_07681_, _07680_);
  nor _58386_ (_07682_, _07681_, _07678_);
  nor _58387_ (_07683_, _07605_, _05961_);
  or _58388_ (_07684_, _07683_, _07254_);
  nor _58389_ (_07685_, _07684_, _07682_);
  and _58390_ (_07686_, _07254_, _06213_);
  or _58391_ (_07687_, _07686_, _07253_);
  nor _58392_ (_07688_, _07687_, _07685_);
  nor _58393_ (_07689_, _07605_, _05959_);
  nor _58394_ (_07690_, _07689_, _07435_);
  not _58395_ (_07691_, _07690_);
  nor _58396_ (_07692_, _07691_, _07688_);
  nor _58397_ (_07693_, _07692_, _07261_);
  and _58398_ (_07694_, _07693_, _07596_);
  not _58399_ (_07695_, _07271_);
  and _58400_ (_07696_, _07261_, _06473_);
  nor _58401_ (_07697_, _07696_, _07695_);
  not _58402_ (_07698_, _07697_);
  nor _58403_ (_07699_, _07698_, _07694_);
  nor _58404_ (_07700_, _07604_, _07271_);
  nor _58405_ (_07701_, _07700_, _07270_);
  not _58406_ (_07702_, _07701_);
  nor _58407_ (_07703_, _07702_, _07699_);
  nor _58408_ (_07704_, _07703_, _07281_);
  and _58409_ (_07705_, _07704_, _07540_);
  and _58410_ (_07706_, _07594_, _07281_);
  nor _58411_ (_07707_, _07706_, _07286_);
  not _58412_ (_07708_, _07707_);
  nor _58413_ (_07709_, _07708_, _07705_);
  nor _58414_ (_07710_, _06279_, _06214_);
  nor _58415_ (_07711_, _07710_, _07709_);
  and _58416_ (_07712_, _07286_, _06657_);
  and _58417_ (_07713_, _06612_, _05927_);
  nor _58418_ (_07714_, _07598_, \oc8051_golden_model_1.SP [2]);
  nor _58419_ (_07715_, _07714_, _07599_);
  not _58420_ (_07716_, _07715_);
  nor _58421_ (_07717_, _07716_, _05959_);
  and _58422_ (_07718_, _06657_, _06220_);
  and _58423_ (_07719_, _06612_, _06257_);
  and _58424_ (_07720_, _07715_, _06267_);
  and _58425_ (_07721_, _07152_, _06657_);
  not _58426_ (_07722_, \oc8051_golden_model_1.IRAM[0] [2]);
  or _58427_ (_07723_, _06936_, _07722_);
  not _58428_ (_07724_, \oc8051_golden_model_1.IRAM[1] [2]);
  or _58429_ (_07725_, _07078_, _07724_);
  and _58430_ (_07726_, _07725_, _07076_);
  nand _58431_ (_07727_, _07726_, _07723_);
  not _58432_ (_07728_, \oc8051_golden_model_1.IRAM[3] [2]);
  or _58433_ (_07729_, _07078_, _07728_);
  not _58434_ (_07730_, \oc8051_golden_model_1.IRAM[2] [2]);
  or _58435_ (_07731_, _06936_, _07730_);
  and _58436_ (_07732_, _07731_, _07084_);
  nand _58437_ (_07733_, _07732_, _07729_);
  nand _58438_ (_07734_, _07733_, _07727_);
  nand _58439_ (_07735_, _07734_, _06769_);
  not _58440_ (_07736_, \oc8051_golden_model_1.IRAM[7] [2]);
  or _58441_ (_07737_, _07078_, _07736_);
  not _58442_ (_07738_, \oc8051_golden_model_1.IRAM[6] [2]);
  or _58443_ (_07739_, _06936_, _07738_);
  and _58444_ (_07740_, _07739_, _07084_);
  nand _58445_ (_07741_, _07740_, _07737_);
  not _58446_ (_07742_, \oc8051_golden_model_1.IRAM[4] [2]);
  or _58447_ (_07743_, _06936_, _07742_);
  not _58448_ (_07744_, \oc8051_golden_model_1.IRAM[5] [2]);
  or _58449_ (_07745_, _07078_, _07744_);
  and _58450_ (_07746_, _07745_, _07076_);
  nand _58451_ (_07747_, _07746_, _07743_);
  nand _58452_ (_07748_, _07747_, _07741_);
  nand _58453_ (_07749_, _07748_, _07091_);
  nand _58454_ (_07750_, _07749_, _07735_);
  nand _58455_ (_07751_, _07750_, _06580_);
  nand _58456_ (_07752_, _06936_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _58457_ (_07753_, _07078_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _58458_ (_07754_, _07753_, _07084_);
  nand _58459_ (_07755_, _07754_, _07752_);
  nand _58460_ (_07756_, _07078_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand _58461_ (_07757_, _06936_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _58462_ (_07758_, _07757_, _07076_);
  nand _58463_ (_07759_, _07758_, _07756_);
  nand _58464_ (_07760_, _07759_, _07755_);
  nand _58465_ (_07761_, _07760_, _06769_);
  not _58466_ (_07762_, \oc8051_golden_model_1.IRAM[15] [2]);
  or _58467_ (_07763_, _07078_, _07762_);
  not _58468_ (_07764_, \oc8051_golden_model_1.IRAM[14] [2]);
  or _58469_ (_07765_, _06936_, _07764_);
  and _58470_ (_07766_, _07765_, _07084_);
  nand _58471_ (_07767_, _07766_, _07763_);
  nand _58472_ (_07768_, _07078_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand _58473_ (_07769_, _06936_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _58474_ (_07770_, _07769_, _07076_);
  nand _58475_ (_07771_, _07770_, _07768_);
  nand _58476_ (_07772_, _07771_, _07767_);
  nand _58477_ (_07773_, _07772_, _07091_);
  nand _58478_ (_07774_, _07773_, _07761_);
  nand _58479_ (_07775_, _07774_, _07108_);
  nand _58480_ (_07776_, _07775_, _07751_);
  or _58481_ (_07777_, _07776_, _05934_);
  and _58482_ (_07778_, _07777_, _07485_);
  and _58483_ (_07779_, _07143_, _06656_);
  nor _58484_ (_07780_, _07779_, _07778_);
  and _58485_ (_07781_, _07716_, _06758_);
  and _58486_ (_07782_, _06336_, _06271_);
  nor _58487_ (_07783_, _07782_, _07781_);
  and _58488_ (_07784_, _07783_, _07780_);
  and _58489_ (_07785_, _07776_, _07154_);
  nor _58490_ (_07786_, _07785_, _07152_);
  and _58491_ (_07787_, _07786_, _07784_);
  nor _58492_ (_07788_, _07787_, _07721_);
  nor _58493_ (_07789_, _07788_, _06275_);
  nor _58494_ (_07790_, _07789_, _06623_);
  nor _58495_ (_07791_, _07715_, _06010_);
  nor _58496_ (_07792_, _07791_, _07790_);
  and _58497_ (_07793_, _07167_, _06656_);
  and _58498_ (_07794_, _06336_, _06266_);
  nor _58499_ (_07795_, _07794_, _07793_);
  and _58500_ (_07796_, _07795_, _07792_);
  and _58501_ (_07797_, _07776_, _07174_);
  nor _58502_ (_07798_, _07797_, _07180_);
  and _58503_ (_07799_, _07798_, _07796_);
  and _58504_ (_07800_, _07180_, _06657_);
  nor _58505_ (_07801_, _07800_, _07799_);
  and _58506_ (_07802_, _06611_, _07179_);
  nor _58507_ (_07803_, _07802_, _07801_);
  and _58508_ (_07804_, _07803_, _07303_);
  nor _58509_ (_07805_, _07804_, _07720_);
  and _58510_ (_07806_, _06264_, _06611_);
  or _58511_ (_07807_, _07806_, _07805_);
  nor _58512_ (_07808_, _07715_, _06007_);
  nor _58513_ (_07809_, _07808_, _06498_);
  not _58514_ (_07810_, _07809_);
  nor _58515_ (_07811_, _07810_, _07807_);
  and _58516_ (_07812_, _07776_, _07197_);
  nor _58517_ (_07813_, _07812_, _07196_);
  and _58518_ (_07814_, _07813_, _07811_);
  nor _58519_ (_07815_, _07814_, _07719_);
  nor _58520_ (_07816_, _07815_, _06254_);
  nor _58521_ (_07817_, _07716_, _05978_);
  nor _58522_ (_07818_, _07817_, _07816_);
  and _58523_ (_07819_, _07218_, _06656_);
  and _58524_ (_07820_, _06336_, _06321_);
  nor _58525_ (_07821_, _07820_, _07819_);
  not _58526_ (_07822_, _07821_);
  nor _58527_ (_07823_, _07822_, _07818_);
  and _58528_ (_07824_, _07776_, _07224_);
  nor _58529_ (_07825_, _07824_, _06220_);
  and _58530_ (_07826_, _07825_, _07823_);
  nor _58531_ (_07827_, _07826_, _07718_);
  nor _58532_ (_07828_, _07827_, _06217_);
  nor _58533_ (_07829_, _07716_, _05952_);
  nor _58534_ (_07830_, _07829_, _07828_);
  nor _58535_ (_07831_, _07246_, _06657_);
  nor _58536_ (_07832_, _07831_, _07233_);
  not _58537_ (_07833_, _07832_);
  nor _58538_ (_07834_, _07833_, _07830_);
  nor _58539_ (_07835_, _07716_, _05961_);
  nor _58540_ (_07836_, _07835_, _07834_);
  and _58541_ (_07837_, _07254_, _06656_);
  or _58542_ (_07838_, _07837_, _07253_);
  nor _58543_ (_07839_, _07838_, _07836_);
  nor _58544_ (_07840_, _07839_, _07717_);
  and _58545_ (_07841_, _06336_, _05779_);
  nor _58546_ (_07842_, _07841_, _07840_);
  and _58547_ (_07843_, _07776_, _07435_);
  nor _58548_ (_07844_, _07843_, _07261_);
  and _58549_ (_07845_, _07844_, _07842_);
  and _58550_ (_07846_, _07261_, _06657_);
  nor _58551_ (_07847_, _07846_, _07845_);
  nor _58552_ (_07848_, _07715_, _07271_);
  nor _58553_ (_07849_, _07848_, _07270_);
  not _58554_ (_07850_, _07849_);
  nor _58555_ (_07851_, _07850_, _07847_);
  nor _58556_ (_07852_, _07851_, _07713_);
  and _58557_ (_07853_, _06336_, _05938_);
  nor _58558_ (_07854_, _07853_, _07852_);
  and _58559_ (_07855_, _07776_, _07281_);
  nor _58560_ (_07856_, _07855_, _07286_);
  and _58561_ (_07857_, _07856_, _07854_);
  nor _58562_ (_07858_, _07857_, _07712_);
  nor _58563_ (_07859_, _07858_, _07536_);
  not _58564_ (_07860_, _07859_);
  nor _58565_ (_07861_, _07860_, _07711_);
  and _58566_ (_07862_, _07861_, _07538_);
  or _58567_ (_07863_, _07862_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand _58568_ (_07864_, _07601_, _06800_);
  or _58569_ (_07865_, _07715_, _07296_);
  and _58570_ (_07866_, _07865_, _07864_);
  and _58571_ (_07867_, _07602_, _06800_);
  and _58572_ (_07868_, _07864_, _07605_);
  nor _58573_ (_07869_, _07868_, _07867_);
  and _58574_ (_07870_, _07509_, _07504_);
  and _58575_ (_07871_, _07870_, _07496_);
  nor _58576_ (_07872_, _07871_, _07454_);
  and _58577_ (_07873_, _07872_, _07869_);
  and _58578_ (_07874_, _07873_, _07866_);
  and _58579_ (_07875_, _07874_, _07295_);
  not _58580_ (_07876_, _07875_);
  and _58581_ (_07877_, _07876_, _07863_);
  not _58582_ (_07878_, _07862_);
  and _58583_ (_07879_, _06656_, _06473_);
  and _58584_ (_07880_, _07004_, _06252_);
  and _58585_ (_07881_, _07880_, _07879_);
  and _58586_ (_07882_, _06317_, _06182_);
  not _58587_ (_07883_, _06968_);
  and _58588_ (_07884_, _07883_, _06611_);
  and _58589_ (_07885_, _07884_, _07882_);
  and _58590_ (_07886_, _07885_, _07881_);
  and _58591_ (_07887_, _07886_, \oc8051_golden_model_1.SBUF [7]);
  not _58592_ (_07888_, _07887_);
  and _58593_ (_07889_, _07004_, _06251_);
  and _58594_ (_07890_, _06656_, _06213_);
  and _58595_ (_07891_, _07890_, _07889_);
  nor _58596_ (_07892_, _06968_, _06611_);
  and _58597_ (_07893_, _07892_, _07882_);
  and _58598_ (_07894_, _07893_, _07891_);
  and _58599_ (_07895_, _07894_, \oc8051_golden_model_1.P3 [7]);
  not _58600_ (_07896_, _06611_);
  and _58601_ (_07897_, _06968_, _07896_);
  and _58602_ (_07898_, _07897_, _07882_);
  and _58603_ (_07899_, _07889_, _07879_);
  and _58604_ (_07900_, _07899_, _07898_);
  and _58605_ (_07901_, _07900_, \oc8051_golden_model_1.IE [7]);
  nor _58606_ (_07902_, _07901_, _07895_);
  and _58607_ (_07903_, _07902_, _07888_);
  and _58608_ (_07904_, _07898_, _07891_);
  and _58609_ (_07905_, _07904_, \oc8051_golden_model_1.P2 [7]);
  and _58610_ (_07906_, _06968_, _06611_);
  and _58611_ (_07907_, _07906_, _07882_);
  nor _58612_ (_07908_, _06656_, _06213_);
  and _58613_ (_07909_, _07880_, _07908_);
  and _58614_ (_07910_, _07909_, _07907_);
  and _58615_ (_07911_, _07910_, \oc8051_golden_model_1.TH1 [7]);
  nor _58616_ (_07912_, _07911_, _07905_);
  and _58617_ (_07913_, _07912_, _07903_);
  and _58618_ (_07914_, _07881_, _07907_);
  and _58619_ (_07915_, _07914_, \oc8051_golden_model_1.TMOD [7]);
  not _58620_ (_07916_, _07915_);
  nor _58621_ (_07917_, _07004_, _06252_);
  and _58622_ (_07918_, _07879_, _07917_);
  and _58623_ (_07919_, _07918_, _07907_);
  and _58624_ (_07920_, _07919_, \oc8051_golden_model_1.TL0 [7]);
  and _58625_ (_07921_, _07908_, _07889_);
  and _58626_ (_07922_, _07921_, _07907_);
  and _58627_ (_07923_, _07922_, \oc8051_golden_model_1.TH0 [7]);
  nor _58628_ (_07924_, _07923_, _07920_);
  and _58629_ (_07925_, _07924_, _07916_);
  and _58630_ (_07926_, _07891_, _07907_);
  and _58631_ (_07927_, _07926_, \oc8051_golden_model_1.P0 [7]);
  and _58632_ (_07928_, _07899_, _07907_);
  and _58633_ (_07929_, _07928_, \oc8051_golden_model_1.TCON [7]);
  nor _58634_ (_07930_, _07929_, _07927_);
  and _58635_ (_07931_, _07930_, _07925_);
  and _58636_ (_07932_, _07931_, _07913_);
  nor _58637_ (_07933_, _06317_, _06286_);
  and _58638_ (_07934_, _07933_, _07884_);
  and _58639_ (_07935_, _07934_, _07891_);
  and _58640_ (_07936_, _07935_, \oc8051_golden_model_1.PSW [7]);
  not _58641_ (_07937_, _07936_);
  and _58642_ (_07938_, _07933_, _07897_);
  and _58643_ (_07939_, _07938_, _07891_);
  and _58644_ (_07940_, _07939_, \oc8051_golden_model_1.ACC [7]);
  and _58645_ (_07941_, _07933_, _07892_);
  and _58646_ (_07942_, _07941_, _07891_);
  and _58647_ (_07943_, _07942_, \oc8051_golden_model_1.B [7]);
  nor _58648_ (_07944_, _07943_, _07940_);
  and _58649_ (_07945_, _07944_, _07937_);
  and _58650_ (_07946_, _07899_, _07893_);
  and _58651_ (_07947_, _07946_, \oc8051_golden_model_1.IP [7]);
  and _58652_ (_07948_, _07907_, _06213_);
  nor _58653_ (_07949_, _07004_, _06251_);
  and _58654_ (_07950_, _07949_, _06657_);
  and _58655_ (_07951_, _07950_, _07948_);
  and _58656_ (_07952_, _07951_, \oc8051_golden_model_1.PCON [7]);
  nor _58657_ (_07953_, _07952_, _07947_);
  and _58658_ (_07954_, _07953_, _07945_);
  and _58659_ (_07955_, _07880_, _07890_);
  and _58660_ (_07956_, _07955_, _07907_);
  and _58661_ (_07957_, _07956_, \oc8051_golden_model_1.SP [7]);
  not _58662_ (_07958_, _07957_);
  and _58663_ (_07959_, _07917_, _06656_);
  and _58664_ (_07960_, _07959_, _07948_);
  and _58665_ (_07961_, _07960_, \oc8051_golden_model_1.DPL [7]);
  and _58666_ (_07962_, _07949_, _07890_);
  and _58667_ (_07963_, _07962_, _07907_);
  and _58668_ (_07964_, _07963_, \oc8051_golden_model_1.DPH [7]);
  nor _58669_ (_07965_, _07964_, _07961_);
  and _58670_ (_07966_, _07965_, _07958_);
  and _58671_ (_07967_, _07949_, _07879_);
  and _58672_ (_07968_, _07967_, _07907_);
  and _58673_ (_07969_, _07968_, \oc8051_golden_model_1.TL1 [7]);
  not _58674_ (_07970_, _07969_);
  and _58675_ (_07971_, _07885_, _07891_);
  and _58676_ (_07972_, _07971_, \oc8051_golden_model_1.P1 [7]);
  and _58677_ (_07973_, _07899_, _07885_);
  and _58678_ (_07974_, _07973_, \oc8051_golden_model_1.SCON [7]);
  nor _58679_ (_07975_, _07974_, _07972_);
  and _58680_ (_07976_, _07975_, _07970_);
  and _58681_ (_07977_, _07976_, _07966_);
  and _58682_ (_07978_, _07977_, _07954_);
  and _58683_ (_07979_, _07978_, _07932_);
  not _58684_ (_07980_, \oc8051_golden_model_1.IRAM[0] [7]);
  or _58685_ (_07981_, _06936_, _07980_);
  not _58686_ (_07982_, \oc8051_golden_model_1.IRAM[1] [7]);
  or _58687_ (_07983_, _07078_, _07982_);
  and _58688_ (_07984_, _07983_, _07076_);
  nand _58689_ (_07985_, _07984_, _07981_);
  not _58690_ (_07986_, \oc8051_golden_model_1.IRAM[3] [7]);
  or _58691_ (_07987_, _07078_, _07986_);
  not _58692_ (_07988_, \oc8051_golden_model_1.IRAM[2] [7]);
  or _58693_ (_07989_, _06936_, _07988_);
  and _58694_ (_07990_, _07989_, _07084_);
  nand _58695_ (_07991_, _07990_, _07987_);
  nand _58696_ (_07992_, _07991_, _07985_);
  nand _58697_ (_07993_, _07992_, _06769_);
  not _58698_ (_07994_, \oc8051_golden_model_1.IRAM[7] [7]);
  or _58699_ (_07995_, _07078_, _07994_);
  not _58700_ (_07996_, \oc8051_golden_model_1.IRAM[6] [7]);
  or _58701_ (_07997_, _06936_, _07996_);
  and _58702_ (_07998_, _07997_, _07084_);
  nand _58703_ (_07999_, _07998_, _07995_);
  not _58704_ (_08000_, \oc8051_golden_model_1.IRAM[4] [7]);
  or _58705_ (_08001_, _06936_, _08000_);
  not _58706_ (_08002_, \oc8051_golden_model_1.IRAM[5] [7]);
  or _58707_ (_08003_, _07078_, _08002_);
  and _58708_ (_08004_, _08003_, _07076_);
  nand _58709_ (_08005_, _08004_, _08001_);
  nand _58710_ (_08006_, _08005_, _07999_);
  nand _58711_ (_08007_, _08006_, _07091_);
  nand _58712_ (_08008_, _08007_, _07993_);
  nand _58713_ (_08009_, _08008_, _06580_);
  not _58714_ (_08010_, \oc8051_golden_model_1.IRAM[11] [7]);
  or _58715_ (_08011_, _07078_, _08010_);
  not _58716_ (_08012_, \oc8051_golden_model_1.IRAM[10] [7]);
  or _58717_ (_08013_, _06936_, _08012_);
  and _58718_ (_08014_, _08013_, _07084_);
  nand _58719_ (_08015_, _08014_, _08011_);
  not _58720_ (_08016_, \oc8051_golden_model_1.IRAM[8] [7]);
  or _58721_ (_08017_, _06936_, _08016_);
  not _58722_ (_08018_, \oc8051_golden_model_1.IRAM[9] [7]);
  or _58723_ (_08019_, _07078_, _08018_);
  and _58724_ (_08020_, _08019_, _07076_);
  nand _58725_ (_08021_, _08020_, _08017_);
  nand _58726_ (_08022_, _08021_, _08015_);
  nand _58727_ (_08023_, _08022_, _06769_);
  not _58728_ (_08024_, \oc8051_golden_model_1.IRAM[15] [7]);
  or _58729_ (_08025_, _07078_, _08024_);
  not _58730_ (_08026_, \oc8051_golden_model_1.IRAM[14] [7]);
  or _58731_ (_08027_, _06936_, _08026_);
  and _58732_ (_08028_, _08027_, _07084_);
  nand _58733_ (_08029_, _08028_, _08025_);
  not _58734_ (_08030_, \oc8051_golden_model_1.IRAM[12] [7]);
  or _58735_ (_08031_, _06936_, _08030_);
  not _58736_ (_08032_, \oc8051_golden_model_1.IRAM[13] [7]);
  or _58737_ (_08033_, _07078_, _08032_);
  and _58738_ (_08034_, _08033_, _07076_);
  nand _58739_ (_08035_, _08034_, _08031_);
  nand _58740_ (_08036_, _08035_, _08029_);
  nand _58741_ (_08037_, _08036_, _07091_);
  nand _58742_ (_08038_, _08037_, _08023_);
  nand _58743_ (_08039_, _08038_, _07108_);
  nand _58744_ (_08040_, _08039_, _08009_);
  or _58745_ (_08041_, _08040_, _06182_);
  and _58746_ (_08042_, _08041_, _07979_);
  not _58747_ (_08043_, _08042_);
  and _58748_ (_08044_, _07904_, \oc8051_golden_model_1.P2 [6]);
  not _58749_ (_08045_, _08044_);
  and _58750_ (_08046_, _07886_, \oc8051_golden_model_1.SBUF [6]);
  not _58751_ (_08047_, _08046_);
  and _58752_ (_08048_, _07894_, \oc8051_golden_model_1.P3 [6]);
  and _58753_ (_08049_, _07900_, \oc8051_golden_model_1.IE [6]);
  nor _58754_ (_08050_, _08049_, _08048_);
  and _58755_ (_08051_, _08050_, _08047_);
  and _58756_ (_08052_, _08051_, _08045_);
  and _58757_ (_08053_, _07926_, \oc8051_golden_model_1.P0 [6]);
  not _58758_ (_08054_, _08053_);
  and _58759_ (_08055_, _07960_, \oc8051_golden_model_1.DPL [6]);
  and _58760_ (_08056_, _07963_, \oc8051_golden_model_1.DPH [6]);
  nor _58761_ (_08057_, _08056_, _08055_);
  and _58762_ (_08058_, _08057_, _08054_);
  and _58763_ (_08059_, _07971_, \oc8051_golden_model_1.P1 [6]);
  and _58764_ (_08060_, _07973_, \oc8051_golden_model_1.SCON [6]);
  nor _58765_ (_08061_, _08060_, _08059_);
  and _58766_ (_08062_, _07968_, \oc8051_golden_model_1.TL1 [6]);
  and _58767_ (_08063_, _07910_, \oc8051_golden_model_1.TH1 [6]);
  nor _58768_ (_08064_, _08063_, _08062_);
  and _58769_ (_08065_, _08064_, _08061_);
  and _58770_ (_08066_, _08065_, _08058_);
  and _58771_ (_08067_, _08066_, _08052_);
  and _58772_ (_08068_, _07935_, \oc8051_golden_model_1.PSW [6]);
  not _58773_ (_08069_, _08068_);
  and _58774_ (_08070_, _07942_, \oc8051_golden_model_1.B [6]);
  and _58775_ (_08071_, _07939_, \oc8051_golden_model_1.ACC [6]);
  nor _58776_ (_08072_, _08071_, _08070_);
  and _58777_ (_08073_, _08072_, _08069_);
  and _58778_ (_08074_, _07946_, \oc8051_golden_model_1.IP [6]);
  and _58779_ (_08075_, _07951_, \oc8051_golden_model_1.PCON [6]);
  nor _58780_ (_08076_, _08075_, _08074_);
  and _58781_ (_08077_, _08076_, _08073_);
  and _58782_ (_08078_, _07928_, \oc8051_golden_model_1.TCON [6]);
  not _58783_ (_08079_, _08078_);
  and _58784_ (_08080_, _07922_, \oc8051_golden_model_1.TH0 [6]);
  and _58785_ (_08081_, _07919_, \oc8051_golden_model_1.TL0 [6]);
  nor _58786_ (_08082_, _08081_, _08080_);
  and _58787_ (_08083_, _08082_, _08079_);
  and _58788_ (_08084_, _07914_, \oc8051_golden_model_1.TMOD [6]);
  and _58789_ (_08085_, _07956_, \oc8051_golden_model_1.SP [6]);
  nor _58790_ (_08086_, _08085_, _08084_);
  and _58791_ (_08087_, _08086_, _08083_);
  and _58792_ (_08088_, _08087_, _08077_);
  and _58793_ (_08089_, _08088_, _08067_);
  not _58794_ (_08090_, \oc8051_golden_model_1.IRAM[0] [6]);
  or _58795_ (_08091_, _06936_, _08090_);
  not _58796_ (_08092_, \oc8051_golden_model_1.IRAM[1] [6]);
  or _58797_ (_08093_, _07078_, _08092_);
  and _58798_ (_08094_, _08093_, _07076_);
  nand _58799_ (_08095_, _08094_, _08091_);
  not _58800_ (_08096_, \oc8051_golden_model_1.IRAM[3] [6]);
  or _58801_ (_08097_, _07078_, _08096_);
  not _58802_ (_08098_, \oc8051_golden_model_1.IRAM[2] [6]);
  or _58803_ (_08099_, _06936_, _08098_);
  and _58804_ (_08100_, _08099_, _07084_);
  nand _58805_ (_08101_, _08100_, _08097_);
  nand _58806_ (_08102_, _08101_, _08095_);
  nand _58807_ (_08103_, _08102_, _06769_);
  not _58808_ (_08104_, \oc8051_golden_model_1.IRAM[7] [6]);
  or _58809_ (_08105_, _07078_, _08104_);
  not _58810_ (_08106_, \oc8051_golden_model_1.IRAM[6] [6]);
  or _58811_ (_08107_, _06936_, _08106_);
  and _58812_ (_08108_, _08107_, _07084_);
  nand _58813_ (_08109_, _08108_, _08105_);
  not _58814_ (_08110_, \oc8051_golden_model_1.IRAM[4] [6]);
  or _58815_ (_08111_, _06936_, _08110_);
  not _58816_ (_08112_, \oc8051_golden_model_1.IRAM[5] [6]);
  or _58817_ (_08113_, _07078_, _08112_);
  and _58818_ (_08114_, _08113_, _07076_);
  nand _58819_ (_08115_, _08114_, _08111_);
  nand _58820_ (_08116_, _08115_, _08109_);
  nand _58821_ (_08117_, _08116_, _07091_);
  nand _58822_ (_08118_, _08117_, _08103_);
  nand _58823_ (_08119_, _08118_, _06580_);
  nand _58824_ (_08120_, _06936_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _58825_ (_08121_, _07078_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _58826_ (_08122_, _08121_, _07084_);
  nand _58827_ (_08123_, _08122_, _08120_);
  nand _58828_ (_08124_, _07078_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand _58829_ (_08125_, _06936_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _58830_ (_08126_, _08125_, _07076_);
  nand _58831_ (_08127_, _08126_, _08124_);
  nand _58832_ (_08128_, _08127_, _08123_);
  nand _58833_ (_08129_, _08128_, _06769_);
  nand _58834_ (_08130_, _06936_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _58835_ (_08131_, _07078_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _58836_ (_08132_, _08131_, _07084_);
  nand _58837_ (_08133_, _08132_, _08130_);
  nand _58838_ (_08134_, _07078_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand _58839_ (_08135_, _06936_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _58840_ (_08136_, _08135_, _07076_);
  nand _58841_ (_08137_, _08136_, _08134_);
  nand _58842_ (_08138_, _08137_, _08133_);
  nand _58843_ (_08139_, _08138_, _07091_);
  nand _58844_ (_08140_, _08139_, _08129_);
  nand _58845_ (_08141_, _08140_, _07108_);
  nand _58846_ (_08142_, _08141_, _08119_);
  or _58847_ (_08143_, _08142_, _06182_);
  and _58848_ (_08144_, _08143_, _08089_);
  not _58849_ (_08145_, _08144_);
  and _58850_ (_08146_, _07935_, \oc8051_golden_model_1.PSW [5]);
  and _58851_ (_08147_, _07942_, \oc8051_golden_model_1.B [5]);
  nor _58852_ (_08148_, _08147_, _08146_);
  and _58853_ (_08149_, _07973_, \oc8051_golden_model_1.SCON [5]);
  and _58854_ (_08150_, _07894_, \oc8051_golden_model_1.P3 [5]);
  nor _58855_ (_08151_, _08150_, _08149_);
  and _58856_ (_08152_, _08151_, _08148_);
  and _58857_ (_08153_, _07919_, \oc8051_golden_model_1.TL0 [5]);
  and _58858_ (_08154_, _07939_, \oc8051_golden_model_1.ACC [5]);
  nor _58859_ (_08155_, _08154_, _08153_);
  and _58860_ (_08156_, _07922_, \oc8051_golden_model_1.TH0 [5]);
  and _58861_ (_08157_, _07904_, \oc8051_golden_model_1.P2 [5]);
  nor _58862_ (_08158_, _08157_, _08156_);
  and _58863_ (_08159_, _08158_, _08155_);
  and _58864_ (_08160_, _07971_, \oc8051_golden_model_1.P1 [5]);
  and _58865_ (_08161_, _07900_, \oc8051_golden_model_1.IE [5]);
  nor _58866_ (_08162_, _08161_, _08160_);
  and _58867_ (_08163_, _07886_, \oc8051_golden_model_1.SBUF [5]);
  and _58868_ (_08164_, _07946_, \oc8051_golden_model_1.IP [5]);
  nor _58869_ (_08165_, _08164_, _08163_);
  and _58870_ (_08166_, _08165_, _08162_);
  and _58871_ (_08167_, _08166_, _08159_);
  and _58872_ (_08168_, _08167_, _08152_);
  and _58873_ (_08169_, _07926_, \oc8051_golden_model_1.P0 [5]);
  not _58874_ (_08170_, _08169_);
  and _58875_ (_08171_, _07960_, \oc8051_golden_model_1.DPL [5]);
  and _58876_ (_08172_, _07880_, _06656_);
  and _58877_ (_08173_, _07948_, _08172_);
  and _58878_ (_08174_, _08173_, \oc8051_golden_model_1.SP [5]);
  nor _58879_ (_08175_, _08174_, _08171_);
  and _58880_ (_08176_, _08175_, _08170_);
  and _58881_ (_08177_, _07928_, \oc8051_golden_model_1.TCON [5]);
  and _58882_ (_08178_, _07914_, \oc8051_golden_model_1.TMOD [5]);
  nor _58883_ (_08179_, _08178_, _08177_);
  and _58884_ (_08180_, _07968_, \oc8051_golden_model_1.TL1 [5]);
  and _58885_ (_08181_, _07910_, \oc8051_golden_model_1.TH1 [5]);
  nor _58886_ (_08182_, _08181_, _08180_);
  and _58887_ (_08183_, _08182_, _08179_);
  and _58888_ (_08184_, _07951_, \oc8051_golden_model_1.PCON [5]);
  and _58889_ (_08185_, _07949_, _06656_);
  and _58890_ (_08186_, _08185_, _07948_);
  and _58891_ (_08187_, _08186_, \oc8051_golden_model_1.DPH [5]);
  nor _58892_ (_08188_, _08187_, _08184_);
  and _58893_ (_08189_, _08188_, _08183_);
  and _58894_ (_08190_, _08189_, _08176_);
  and _58895_ (_08191_, _08190_, _08168_);
  not _58896_ (_08192_, \oc8051_golden_model_1.IRAM[0] [5]);
  or _58897_ (_08193_, _06936_, _08192_);
  not _58898_ (_08194_, \oc8051_golden_model_1.IRAM[1] [5]);
  or _58899_ (_08195_, _07078_, _08194_);
  and _58900_ (_08196_, _08195_, _07076_);
  nand _58901_ (_08197_, _08196_, _08193_);
  not _58902_ (_08198_, \oc8051_golden_model_1.IRAM[3] [5]);
  or _58903_ (_08199_, _07078_, _08198_);
  not _58904_ (_08200_, \oc8051_golden_model_1.IRAM[2] [5]);
  or _58905_ (_08201_, _06936_, _08200_);
  and _58906_ (_08202_, _08201_, _07084_);
  nand _58907_ (_08203_, _08202_, _08199_);
  nand _58908_ (_08204_, _08203_, _08197_);
  nand _58909_ (_08205_, _08204_, _06769_);
  not _58910_ (_08206_, \oc8051_golden_model_1.IRAM[7] [5]);
  or _58911_ (_08207_, _07078_, _08206_);
  not _58912_ (_08208_, \oc8051_golden_model_1.IRAM[6] [5]);
  or _58913_ (_08209_, _06936_, _08208_);
  and _58914_ (_08210_, _08209_, _07084_);
  nand _58915_ (_08211_, _08210_, _08207_);
  not _58916_ (_08212_, \oc8051_golden_model_1.IRAM[4] [5]);
  or _58917_ (_08213_, _06936_, _08212_);
  not _58918_ (_08214_, \oc8051_golden_model_1.IRAM[5] [5]);
  or _58919_ (_08215_, _07078_, _08214_);
  and _58920_ (_08216_, _08215_, _07076_);
  nand _58921_ (_08217_, _08216_, _08213_);
  nand _58922_ (_08218_, _08217_, _08211_);
  nand _58923_ (_08219_, _08218_, _07091_);
  nand _58924_ (_08220_, _08219_, _08205_);
  nand _58925_ (_08221_, _08220_, _06580_);
  nand _58926_ (_08222_, _06936_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _58927_ (_08223_, _07078_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _58928_ (_08224_, _08223_, _07084_);
  nand _58929_ (_08225_, _08224_, _08222_);
  nand _58930_ (_08226_, _07078_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand _58931_ (_08227_, _06936_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _58932_ (_08228_, _08227_, _07076_);
  nand _58933_ (_08229_, _08228_, _08226_);
  nand _58934_ (_08230_, _08229_, _08225_);
  nand _58935_ (_08231_, _08230_, _06769_);
  nand _58936_ (_08232_, _06936_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _58937_ (_08233_, _07078_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _58938_ (_08234_, _08233_, _07084_);
  nand _58939_ (_08235_, _08234_, _08232_);
  nand _58940_ (_08236_, _07078_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand _58941_ (_08237_, _06936_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _58942_ (_08238_, _08237_, _07076_);
  nand _58943_ (_08239_, _08238_, _08236_);
  nand _58944_ (_08240_, _08239_, _08235_);
  nand _58945_ (_08241_, _08240_, _07091_);
  nand _58946_ (_08242_, _08241_, _08231_);
  nand _58947_ (_08243_, _08242_, _07108_);
  nand _58948_ (_08244_, _08243_, _08221_);
  or _58949_ (_08245_, _08244_, _06182_);
  and _58950_ (_08246_, _08245_, _08191_);
  not _58951_ (_08247_, _08246_);
  and _58952_ (_08248_, _07900_, \oc8051_golden_model_1.IE [3]);
  and _58953_ (_08249_, _07946_, \oc8051_golden_model_1.IP [3]);
  nor _58954_ (_08250_, _08249_, _08248_);
  and _58955_ (_08251_, _07886_, \oc8051_golden_model_1.SBUF [3]);
  and _58956_ (_08252_, _07904_, \oc8051_golden_model_1.P2 [3]);
  nor _58957_ (_08253_, _08252_, _08251_);
  and _58958_ (_08254_, _08253_, _08250_);
  and _58959_ (_08255_, _07894_, \oc8051_golden_model_1.P3 [3]);
  and _58960_ (_08256_, _07939_, \oc8051_golden_model_1.ACC [3]);
  nor _58961_ (_08257_, _08256_, _08255_);
  and _58962_ (_08258_, _07935_, \oc8051_golden_model_1.PSW [3]);
  and _58963_ (_08259_, _07942_, \oc8051_golden_model_1.B [3]);
  nor _58964_ (_08260_, _08259_, _08258_);
  and _58965_ (_08261_, _08260_, _08257_);
  and _58966_ (_08262_, _07971_, \oc8051_golden_model_1.P1 [3]);
  and _58967_ (_08263_, _07973_, \oc8051_golden_model_1.SCON [3]);
  nor _58968_ (_08264_, _08263_, _08262_);
  and _58969_ (_08265_, _07919_, \oc8051_golden_model_1.TL0 [3]);
  and _58970_ (_08266_, _07922_, \oc8051_golden_model_1.TH0 [3]);
  nor _58971_ (_08267_, _08266_, _08265_);
  and _58972_ (_08268_, _08267_, _08264_);
  and _58973_ (_08269_, _08268_, _08261_);
  and _58974_ (_08270_, _08269_, _08254_);
  and _58975_ (_08271_, _07926_, \oc8051_golden_model_1.P0 [3]);
  not _58976_ (_08272_, _08271_);
  and _58977_ (_08273_, _07960_, \oc8051_golden_model_1.DPL [3]);
  and _58978_ (_08274_, _08173_, \oc8051_golden_model_1.SP [3]);
  nor _58979_ (_08275_, _08274_, _08273_);
  and _58980_ (_08276_, _08275_, _08272_);
  and _58981_ (_08277_, _07928_, \oc8051_golden_model_1.TCON [3]);
  and _58982_ (_08278_, _07914_, \oc8051_golden_model_1.TMOD [3]);
  nor _58983_ (_08279_, _08278_, _08277_);
  and _58984_ (_08280_, _07968_, \oc8051_golden_model_1.TL1 [3]);
  and _58985_ (_08281_, _07910_, \oc8051_golden_model_1.TH1 [3]);
  nor _58986_ (_08282_, _08281_, _08280_);
  and _58987_ (_08283_, _08282_, _08279_);
  and _58988_ (_08284_, _07951_, \oc8051_golden_model_1.PCON [3]);
  and _58989_ (_08285_, _08186_, \oc8051_golden_model_1.DPH [3]);
  nor _58990_ (_08286_, _08285_, _08284_);
  and _58991_ (_08287_, _08286_, _08283_);
  and _58992_ (_08288_, _08287_, _08276_);
  and _58993_ (_08289_, _08288_, _08270_);
  or _58994_ (_08290_, _07594_, _06182_);
  and _58995_ (_08291_, _08290_, _08289_);
  not _58996_ (_08292_, _08291_);
  and _58997_ (_08293_, _07886_, \oc8051_golden_model_1.SBUF [1]);
  not _58998_ (_08294_, _08293_);
  and _58999_ (_08295_, _07900_, \oc8051_golden_model_1.IE [1]);
  and _59000_ (_08296_, _07894_, \oc8051_golden_model_1.P3 [1]);
  nor _59001_ (_08297_, _08296_, _08295_);
  and _59002_ (_08298_, _08297_, _08294_);
  and _59003_ (_08299_, _07904_, \oc8051_golden_model_1.P2 [1]);
  and _59004_ (_08300_, _07968_, \oc8051_golden_model_1.TL1 [1]);
  nor _59005_ (_08301_, _08300_, _08299_);
  and _59006_ (_08302_, _08301_, _08298_);
  and _59007_ (_08303_, _07914_, \oc8051_golden_model_1.TMOD [1]);
  not _59008_ (_08304_, _08303_);
  and _59009_ (_08305_, _07919_, \oc8051_golden_model_1.TL0 [1]);
  and _59010_ (_08306_, _07922_, \oc8051_golden_model_1.TH0 [1]);
  nor _59011_ (_08307_, _08306_, _08305_);
  and _59012_ (_08308_, _08307_, _08304_);
  and _59013_ (_08309_, _07928_, \oc8051_golden_model_1.TCON [1]);
  and _59014_ (_08310_, _07956_, \oc8051_golden_model_1.SP [1]);
  nor _59015_ (_08311_, _08310_, _08309_);
  and _59016_ (_08312_, _08311_, _08308_);
  and _59017_ (_08313_, _08312_, _08302_);
  and _59018_ (_08314_, _07939_, \oc8051_golden_model_1.ACC [1]);
  and _59019_ (_08315_, _07942_, \oc8051_golden_model_1.B [1]);
  nor _59020_ (_08316_, _08315_, _08314_);
  and _59021_ (_08317_, _07935_, \oc8051_golden_model_1.PSW [1]);
  not _59022_ (_08318_, _08317_);
  and _59023_ (_08319_, _08318_, _08316_);
  and _59024_ (_08320_, _07946_, \oc8051_golden_model_1.IP [1]);
  and _59025_ (_08321_, _07951_, \oc8051_golden_model_1.PCON [1]);
  nor _59026_ (_08322_, _08321_, _08320_);
  and _59027_ (_08323_, _08322_, _08319_);
  and _59028_ (_08324_, _07926_, \oc8051_golden_model_1.P0 [1]);
  not _59029_ (_08325_, _08324_);
  and _59030_ (_08326_, _07960_, \oc8051_golden_model_1.DPL [1]);
  and _59031_ (_08327_, _07963_, \oc8051_golden_model_1.DPH [1]);
  nor _59032_ (_08328_, _08327_, _08326_);
  and _59033_ (_08329_, _08328_, _08325_);
  and _59034_ (_08330_, _07910_, \oc8051_golden_model_1.TH1 [1]);
  not _59035_ (_08331_, _08330_);
  and _59036_ (_08332_, _07973_, \oc8051_golden_model_1.SCON [1]);
  and _59037_ (_08333_, _07971_, \oc8051_golden_model_1.P1 [1]);
  nor _59038_ (_08334_, _08333_, _08332_);
  and _59039_ (_08335_, _08334_, _08331_);
  and _59040_ (_08336_, _08335_, _08329_);
  and _59041_ (_08337_, _08336_, _08323_);
  and _59042_ (_08338_, _08337_, _08313_);
  or _59043_ (_08339_, _07357_, _06182_);
  and _59044_ (_08340_, _08339_, _08338_);
  not _59045_ (_08341_, _08340_);
  and _59046_ (_08342_, _07904_, \oc8051_golden_model_1.P2 [0]);
  not _59047_ (_08343_, _08342_);
  and _59048_ (_08344_, _07886_, \oc8051_golden_model_1.SBUF [0]);
  not _59049_ (_08345_, _08344_);
  and _59050_ (_08346_, _07900_, \oc8051_golden_model_1.IE [0]);
  and _59051_ (_08347_, _07894_, \oc8051_golden_model_1.P3 [0]);
  nor _59052_ (_08348_, _08347_, _08346_);
  and _59053_ (_08349_, _08348_, _08345_);
  and _59054_ (_08350_, _08349_, _08343_);
  and _59055_ (_08351_, _07960_, \oc8051_golden_model_1.DPL [0]);
  and _59056_ (_08352_, _07963_, \oc8051_golden_model_1.DPH [0]);
  nor _59057_ (_08353_, _08352_, _08351_);
  and _59058_ (_08354_, _07926_, \oc8051_golden_model_1.P0 [0]);
  not _59059_ (_08355_, _08354_);
  and _59060_ (_08356_, _08355_, _08353_);
  and _59061_ (_08357_, _07968_, \oc8051_golden_model_1.TL1 [0]);
  and _59062_ (_08358_, _07910_, \oc8051_golden_model_1.TH1 [0]);
  nor _59063_ (_08359_, _08358_, _08357_);
  and _59064_ (_08360_, _07973_, \oc8051_golden_model_1.SCON [0]);
  and _59065_ (_08361_, _07971_, \oc8051_golden_model_1.P1 [0]);
  nor _59066_ (_08362_, _08361_, _08360_);
  and _59067_ (_08363_, _08362_, _08359_);
  and _59068_ (_08364_, _08363_, _08356_);
  and _59069_ (_08365_, _08364_, _08350_);
  and _59070_ (_08366_, _07935_, \oc8051_golden_model_1.PSW [0]);
  not _59071_ (_08367_, _08366_);
  and _59072_ (_08368_, _07939_, \oc8051_golden_model_1.ACC [0]);
  and _59073_ (_08369_, _07942_, \oc8051_golden_model_1.B [0]);
  nor _59074_ (_08370_, _08369_, _08368_);
  and _59075_ (_08371_, _08370_, _08367_);
  and _59076_ (_08372_, _07946_, \oc8051_golden_model_1.IP [0]);
  and _59077_ (_08373_, _07951_, \oc8051_golden_model_1.PCON [0]);
  nor _59078_ (_08374_, _08373_, _08372_);
  and _59079_ (_08375_, _08374_, _08371_);
  and _59080_ (_08376_, _07914_, \oc8051_golden_model_1.TMOD [0]);
  not _59081_ (_08377_, _08376_);
  and _59082_ (_08378_, _07919_, \oc8051_golden_model_1.TL0 [0]);
  and _59083_ (_08379_, _07922_, \oc8051_golden_model_1.TH0 [0]);
  nor _59084_ (_08380_, _08379_, _08378_);
  and _59085_ (_08381_, _08380_, _08377_);
  and _59086_ (_08382_, _07928_, \oc8051_golden_model_1.TCON [0]);
  and _59087_ (_08383_, _07956_, \oc8051_golden_model_1.SP [0]);
  nor _59088_ (_08384_, _08383_, _08382_);
  and _59089_ (_08385_, _08384_, _08381_);
  and _59090_ (_08386_, _08385_, _08375_);
  and _59091_ (_08387_, _08386_, _08365_);
  not _59092_ (_08388_, _08387_);
  and _59093_ (_08389_, _07133_, _06286_);
  or _59094_ (_08390_, _08389_, _08388_);
  and _59095_ (_08391_, _08390_, _08341_);
  and _59096_ (_08392_, _07886_, \oc8051_golden_model_1.SBUF [2]);
  not _59097_ (_08393_, _08392_);
  and _59098_ (_08394_, _07900_, \oc8051_golden_model_1.IE [2]);
  and _59099_ (_08395_, _07894_, \oc8051_golden_model_1.P3 [2]);
  nor _59100_ (_08396_, _08395_, _08394_);
  and _59101_ (_08397_, _08396_, _08393_);
  and _59102_ (_08398_, _07904_, \oc8051_golden_model_1.P2 [2]);
  and _59103_ (_08399_, _07968_, \oc8051_golden_model_1.TL1 [2]);
  nor _59104_ (_08400_, _08399_, _08398_);
  and _59105_ (_08401_, _08400_, _08397_);
  and _59106_ (_08402_, _07928_, \oc8051_golden_model_1.TCON [2]);
  not _59107_ (_08403_, _08402_);
  and _59108_ (_08404_, _07922_, \oc8051_golden_model_1.TH0 [2]);
  and _59109_ (_08405_, _07919_, \oc8051_golden_model_1.TL0 [2]);
  nor _59110_ (_08406_, _08405_, _08404_);
  and _59111_ (_08407_, _08406_, _08403_);
  and _59112_ (_08408_, _07914_, \oc8051_golden_model_1.TMOD [2]);
  and _59113_ (_08409_, _07926_, \oc8051_golden_model_1.P0 [2]);
  nor _59114_ (_08410_, _08409_, _08408_);
  and _59115_ (_08411_, _08410_, _08407_);
  and _59116_ (_08412_, _08411_, _08401_);
  and _59117_ (_08413_, _07935_, \oc8051_golden_model_1.PSW [2]);
  not _59118_ (_08414_, _08413_);
  and _59119_ (_08415_, _07939_, \oc8051_golden_model_1.ACC [2]);
  and _59120_ (_08416_, _07942_, \oc8051_golden_model_1.B [2]);
  nor _59121_ (_08417_, _08416_, _08415_);
  and _59122_ (_08418_, _08417_, _08414_);
  and _59123_ (_08419_, _07946_, \oc8051_golden_model_1.IP [2]);
  and _59124_ (_08420_, _07951_, \oc8051_golden_model_1.PCON [2]);
  nor _59125_ (_08421_, _08420_, _08419_);
  and _59126_ (_08422_, _08421_, _08418_);
  and _59127_ (_08423_, _07956_, \oc8051_golden_model_1.SP [2]);
  not _59128_ (_08424_, _08423_);
  and _59129_ (_08425_, _07960_, \oc8051_golden_model_1.DPL [2]);
  and _59130_ (_08426_, _07963_, \oc8051_golden_model_1.DPH [2]);
  nor _59131_ (_08427_, _08426_, _08425_);
  and _59132_ (_08428_, _08427_, _08424_);
  and _59133_ (_08429_, _07910_, \oc8051_golden_model_1.TH1 [2]);
  not _59134_ (_08430_, _08429_);
  and _59135_ (_08431_, _07973_, \oc8051_golden_model_1.SCON [2]);
  and _59136_ (_08432_, _07971_, \oc8051_golden_model_1.P1 [2]);
  nor _59137_ (_08433_, _08432_, _08431_);
  and _59138_ (_08434_, _08433_, _08430_);
  and _59139_ (_08435_, _08434_, _08428_);
  and _59140_ (_08436_, _08435_, _08422_);
  and _59141_ (_08437_, _08436_, _08412_);
  or _59142_ (_08438_, _07776_, _06182_);
  and _59143_ (_08439_, _08438_, _08437_);
  not _59144_ (_08440_, _08439_);
  and _59145_ (_08441_, _08440_, _08391_);
  and _59146_ (_08442_, _08441_, _08292_);
  and _59147_ (_08443_, _07904_, \oc8051_golden_model_1.P2 [4]);
  not _59148_ (_08444_, _08443_);
  and _59149_ (_08445_, _07886_, \oc8051_golden_model_1.SBUF [4]);
  not _59150_ (_08446_, _08445_);
  and _59151_ (_08447_, _07894_, \oc8051_golden_model_1.P3 [4]);
  and _59152_ (_08448_, _07900_, \oc8051_golden_model_1.IE [4]);
  nor _59153_ (_08449_, _08448_, _08447_);
  and _59154_ (_08450_, _08449_, _08446_);
  and _59155_ (_08451_, _08450_, _08444_);
  and _59156_ (_08452_, _07956_, \oc8051_golden_model_1.SP [4]);
  not _59157_ (_08453_, _08452_);
  and _59158_ (_08454_, _07960_, \oc8051_golden_model_1.DPL [4]);
  and _59159_ (_08455_, _07963_, \oc8051_golden_model_1.DPH [4]);
  nor _59160_ (_08456_, _08455_, _08454_);
  and _59161_ (_08457_, _08456_, _08453_);
  and _59162_ (_08458_, _07971_, \oc8051_golden_model_1.P1 [4]);
  and _59163_ (_08459_, _07973_, \oc8051_golden_model_1.SCON [4]);
  nor _59164_ (_08460_, _08459_, _08458_);
  and _59165_ (_08461_, _07910_, \oc8051_golden_model_1.TH1 [4]);
  and _59166_ (_08462_, _07968_, \oc8051_golden_model_1.TL1 [4]);
  nor _59167_ (_08463_, _08462_, _08461_);
  and _59168_ (_08464_, _08463_, _08460_);
  and _59169_ (_08465_, _08464_, _08457_);
  and _59170_ (_08466_, _08465_, _08451_);
  and _59171_ (_08467_, _07935_, \oc8051_golden_model_1.PSW [4]);
  not _59172_ (_08468_, _08467_);
  and _59173_ (_08469_, _07939_, \oc8051_golden_model_1.ACC [4]);
  and _59174_ (_08470_, _07942_, \oc8051_golden_model_1.B [4]);
  nor _59175_ (_08471_, _08470_, _08469_);
  and _59176_ (_08472_, _08471_, _08468_);
  and _59177_ (_08473_, _07946_, \oc8051_golden_model_1.IP [4]);
  and _59178_ (_08474_, _07951_, \oc8051_golden_model_1.PCON [4]);
  nor _59179_ (_08475_, _08474_, _08473_);
  and _59180_ (_08476_, _08475_, _08472_);
  and _59181_ (_08477_, _07928_, \oc8051_golden_model_1.TCON [4]);
  not _59182_ (_08478_, _08477_);
  and _59183_ (_08479_, _07919_, \oc8051_golden_model_1.TL0 [4]);
  and _59184_ (_08480_, _07922_, \oc8051_golden_model_1.TH0 [4]);
  nor _59185_ (_08481_, _08480_, _08479_);
  and _59186_ (_08482_, _08481_, _08478_);
  and _59187_ (_08483_, _07914_, \oc8051_golden_model_1.TMOD [4]);
  and _59188_ (_08484_, _07926_, \oc8051_golden_model_1.P0 [4]);
  nor _59189_ (_08485_, _08484_, _08483_);
  and _59190_ (_08486_, _08485_, _08482_);
  and _59191_ (_08487_, _08486_, _08476_);
  and _59192_ (_08488_, _08487_, _08466_);
  not _59193_ (_08489_, \oc8051_golden_model_1.IRAM[0] [4]);
  or _59194_ (_08490_, _06936_, _08489_);
  not _59195_ (_08491_, \oc8051_golden_model_1.IRAM[1] [4]);
  or _59196_ (_08492_, _07078_, _08491_);
  and _59197_ (_08493_, _08492_, _07076_);
  nand _59198_ (_08494_, _08493_, _08490_);
  not _59199_ (_08495_, \oc8051_golden_model_1.IRAM[3] [4]);
  or _59200_ (_08496_, _07078_, _08495_);
  not _59201_ (_08497_, \oc8051_golden_model_1.IRAM[2] [4]);
  or _59202_ (_08498_, _06936_, _08497_);
  and _59203_ (_08499_, _08498_, _07084_);
  nand _59204_ (_08500_, _08499_, _08496_);
  nand _59205_ (_08501_, _08500_, _08494_);
  nand _59206_ (_08502_, _08501_, _06769_);
  not _59207_ (_08503_, \oc8051_golden_model_1.IRAM[7] [4]);
  or _59208_ (_08504_, _07078_, _08503_);
  not _59209_ (_08505_, \oc8051_golden_model_1.IRAM[6] [4]);
  or _59210_ (_08506_, _06936_, _08505_);
  and _59211_ (_08507_, _08506_, _07084_);
  nand _59212_ (_08508_, _08507_, _08504_);
  not _59213_ (_08509_, \oc8051_golden_model_1.IRAM[4] [4]);
  or _59214_ (_08510_, _06936_, _08509_);
  not _59215_ (_08511_, \oc8051_golden_model_1.IRAM[5] [4]);
  or _59216_ (_08512_, _07078_, _08511_);
  and _59217_ (_08513_, _08512_, _07076_);
  nand _59218_ (_08514_, _08513_, _08510_);
  nand _59219_ (_08515_, _08514_, _08508_);
  nand _59220_ (_08516_, _08515_, _07091_);
  nand _59221_ (_08517_, _08516_, _08502_);
  nand _59222_ (_08518_, _08517_, _06580_);
  nand _59223_ (_08519_, _06936_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _59224_ (_08520_, _07078_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _59225_ (_08521_, _08520_, _07084_);
  nand _59226_ (_08522_, _08521_, _08519_);
  nand _59227_ (_08523_, _07078_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand _59228_ (_08524_, _06936_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _59229_ (_08525_, _08524_, _07076_);
  nand _59230_ (_08526_, _08525_, _08523_);
  nand _59231_ (_08527_, _08526_, _08522_);
  nand _59232_ (_08528_, _08527_, _06769_);
  nand _59233_ (_08529_, _06936_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _59234_ (_08530_, _07078_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _59235_ (_08531_, _08530_, _07084_);
  nand _59236_ (_08532_, _08531_, _08529_);
  nand _59237_ (_08533_, _07078_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand _59238_ (_08534_, _06936_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _59239_ (_08535_, _08534_, _07076_);
  nand _59240_ (_08536_, _08535_, _08533_);
  nand _59241_ (_08537_, _08536_, _08532_);
  nand _59242_ (_08538_, _08537_, _07091_);
  nand _59243_ (_08539_, _08538_, _08528_);
  nand _59244_ (_08540_, _08539_, _07108_);
  nand _59245_ (_08541_, _08540_, _08518_);
  or _59246_ (_08542_, _08541_, _06182_);
  and _59247_ (_08543_, _08542_, _08488_);
  not _59248_ (_08544_, _08543_);
  and _59249_ (_08545_, _08544_, _08442_);
  and _59250_ (_08546_, _08545_, _08247_);
  and _59251_ (_08547_, _08546_, _08145_);
  or _59252_ (_08548_, _08547_, _08043_);
  nand _59253_ (_08549_, _08547_, _08043_);
  and _59254_ (_08550_, _08549_, _08548_);
  and _59255_ (_08551_, _08550_, _07286_);
  not _59256_ (_08552_, _08040_);
  and _59257_ (_08553_, _08541_, _08244_);
  and _59258_ (_08554_, _07776_, _07594_);
  not _59259_ (_08555_, _07133_);
  and _59260_ (_08556_, _07357_, _08555_);
  and _59261_ (_08557_, _08556_, _08554_);
  and _59262_ (_08558_, _08557_, _08553_);
  and _59263_ (_08559_, _08558_, _08142_);
  or _59264_ (_08560_, _08559_, _08552_);
  nand _59265_ (_08561_, _08559_, _08552_);
  and _59266_ (_08562_, _08561_, _08560_);
  and _59267_ (_08563_, _06337_, _05779_);
  and _59268_ (_08564_, _06350_, _05779_);
  nor _59269_ (_08565_, _08564_, _08563_);
  nor _59270_ (_08566_, _07211_, _06567_);
  nor _59271_ (_08567_, _07212_, _06567_);
  nor _59272_ (_08568_, _08567_, _08566_);
  and _59273_ (_08569_, _08568_, _08565_);
  or _59274_ (_08570_, _08569_, _08562_);
  not _59275_ (_08571_, _07243_);
  not _59276_ (_08572_, \oc8051_golden_model_1.ACC [7]);
  and _59277_ (_08573_, _08042_, _08572_);
  nor _59278_ (_08574_, _08042_, _08572_);
  nor _59279_ (_08575_, _08574_, _08573_);
  and _59280_ (_08576_, _08575_, _07241_);
  not _59281_ (_08577_, _07241_);
  and _59282_ (_08578_, _06420_, _04431_);
  and _59283_ (_08579_, _06445_, _04415_);
  nor _59284_ (_08580_, _08579_, _08578_);
  and _59285_ (_08581_, _06434_, _04434_);
  and _59286_ (_08582_, _06436_, _04419_);
  nor _59287_ (_08583_, _08582_, _08581_);
  and _59288_ (_08584_, _08583_, _08580_);
  and _59289_ (_08585_, _06417_, _04355_);
  and _59290_ (_08586_, _06415_, _04439_);
  nor _59291_ (_08587_, _08586_, _08585_);
  and _59292_ (_08588_, _06411_, _04387_);
  and _59293_ (_08589_, _06431_, _04392_);
  nor _59294_ (_08590_, _08589_, _08588_);
  and _59295_ (_08591_, _08590_, _08587_);
  and _59296_ (_08592_, _08591_, _08584_);
  and _59297_ (_08593_, _06447_, _04397_);
  and _59298_ (_08594_, _06429_, _04406_);
  nor _59299_ (_08595_, _08594_, _08593_);
  and _59300_ (_08596_, _06440_, _04401_);
  and _59301_ (_08597_, _06401_, _04381_);
  nor _59302_ (_08598_, _08597_, _08596_);
  and _59303_ (_08599_, _08598_, _08595_);
  and _59304_ (_08600_, _06407_, _04423_);
  and _59305_ (_08601_, _06398_, _04442_);
  nor _59306_ (_08602_, _08601_, _08600_);
  and _59307_ (_08603_, _06423_, _04411_);
  and _59308_ (_08604_, _06442_, _04426_);
  nor _59309_ (_08605_, _08604_, _08603_);
  and _59310_ (_08606_, _08605_, _08602_);
  and _59311_ (_08607_, _08606_, _08599_);
  and _59312_ (_08608_, _08607_, _08592_);
  nand _59313_ (_08609_, _08608_, _06220_);
  not _59314_ (_08610_, _07179_);
  and _59315_ (_08611_, _07948_, \oc8051_golden_model_1.P0 [7]);
  not _59316_ (_08612_, _06214_);
  nor _59317_ (_08613_, _06969_, _08612_);
  and _59318_ (_08614_, _06613_, _06320_);
  and _59319_ (_08615_, _08614_, _08613_);
  and _59320_ (_08616_, _08615_, _07907_);
  and _59321_ (_08617_, _08616_, \oc8051_golden_model_1.TCON [7]);
  nor _59322_ (_08618_, _06612_, _06320_);
  and _59323_ (_08619_, _08618_, _08613_);
  and _59324_ (_08620_, _08619_, _07885_);
  and _59325_ (_08621_, _08620_, \oc8051_golden_model_1.P1 [7]);
  and _59326_ (_08622_, _08615_, _07885_);
  and _59327_ (_08623_, _08622_, \oc8051_golden_model_1.SCON [7]);
  and _59328_ (_08624_, _08619_, _07898_);
  and _59329_ (_08625_, _08624_, \oc8051_golden_model_1.P2 [7]);
  and _59330_ (_08626_, _08615_, _07898_);
  and _59331_ (_08627_, _08626_, \oc8051_golden_model_1.IE [7]);
  and _59332_ (_08628_, _08619_, _07893_);
  and _59333_ (_08629_, _08628_, \oc8051_golden_model_1.P3 [7]);
  and _59334_ (_08630_, _08619_, _07934_);
  and _59335_ (_08631_, _08630_, \oc8051_golden_model_1.PSW [7]);
  and _59336_ (_08632_, _08615_, _07893_);
  and _59337_ (_08633_, _08632_, \oc8051_golden_model_1.IP [7]);
  and _59338_ (_08634_, _07941_, _08619_);
  and _59339_ (_08635_, _08634_, \oc8051_golden_model_1.B [7]);
  and _59340_ (_08636_, _08619_, _07938_);
  and _59341_ (_08637_, _08636_, \oc8051_golden_model_1.ACC [7]);
  or _59342_ (_08638_, _08637_, _08635_);
  or _59343_ (_08639_, _08638_, _08633_);
  or _59344_ (_08640_, _08639_, _08631_);
  or _59345_ (_08641_, _08640_, _08629_);
  or _59346_ (_08642_, _08641_, _08627_);
  or _59347_ (_08643_, _08642_, _08625_);
  or _59348_ (_08644_, _08643_, _08623_);
  or _59349_ (_08645_, _08644_, _08621_);
  or _59350_ (_08646_, _08645_, _08617_);
  nor _59351_ (_08647_, _08646_, _08611_);
  and _59352_ (_08648_, _08647_, _08041_);
  nor _59353_ (_08649_, _08648_, _07950_);
  or _59354_ (_08650_, _08649_, _08610_);
  not _59355_ (_08651_, _06275_);
  not _59356_ (_08652_, _07152_);
  nor _59357_ (_08653_, _07213_, _06009_);
  nor _59358_ (_08654_, _08653_, _07364_);
  or _59359_ (_08655_, _08654_, _08562_);
  and _59360_ (_08656_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and _59361_ (_08657_, _08656_, \oc8051_golden_model_1.PC [6]);
  and _59362_ (_08658_, _08657_, _05929_);
  and _59363_ (_08659_, _08658_, \oc8051_golden_model_1.PC [7]);
  nor _59364_ (_08660_, _08658_, \oc8051_golden_model_1.PC [7]);
  nor _59365_ (_08661_, _08660_, _08659_);
  and _59366_ (_08662_, _08661_, _06758_);
  nor _59367_ (_08663_, _06758_, _08572_);
  nor _59368_ (_08664_, _08663_, _08662_);
  nand _59369_ (_08665_, _08664_, _08654_);
  and _59370_ (_08666_, _08665_, _08655_);
  or _59371_ (_08667_, _08666_, _07154_);
  nor _59372_ (_08668_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _59373_ (_08669_, _08668_, _06715_);
  nor _59374_ (_08670_, _08669_, _06460_);
  nor _59375_ (_08671_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _59376_ (_08672_, _08671_, _06460_);
  and _59377_ (_08673_, _08672_, _06800_);
  nor _59378_ (_08674_, _08673_, _08670_);
  nor _59379_ (_08675_, _06551_, _06281_);
  nor _59380_ (_08676_, _08675_, _08674_);
  and _59381_ (_08677_, _07594_, _07198_);
  and _59382_ (_08678_, _07197_, _06213_);
  not _59383_ (_08679_, _08678_);
  nand _59384_ (_08680_, _08679_, _08675_);
  nor _59385_ (_08681_, _08680_, _08677_);
  nor _59386_ (_08682_, _08681_, _08676_);
  nor _59387_ (_08683_, _08668_, _06715_);
  nor _59388_ (_08684_, _08683_, _08669_);
  nor _59389_ (_08685_, _08684_, _08675_);
  not _59390_ (_08686_, _08685_);
  nand _59391_ (_08687_, _07776_, _07198_);
  and _59392_ (_08688_, _07197_, _06656_);
  not _59393_ (_08689_, _08688_);
  and _59394_ (_08690_, _08689_, _08675_);
  nand _59395_ (_08691_, _08690_, _08687_);
  and _59396_ (_08692_, _08691_, _08686_);
  or _59397_ (_08693_, _07197_, _07133_);
  and _59398_ (_08694_, _07197_, _06251_);
  not _59399_ (_08695_, _08694_);
  and _59400_ (_08696_, _08695_, _08675_);
  nand _59401_ (_08697_, _08696_, _08693_);
  nor _59402_ (_08698_, _08675_, \oc8051_golden_model_1.SP [0]);
  not _59403_ (_08699_, _08698_);
  and _59404_ (_08700_, _08699_, _08697_);
  nand _59405_ (_08701_, _08700_, \oc8051_golden_model_1.IRAM[0] [7]);
  nor _59406_ (_08702_, _08675_, _07297_);
  not _59407_ (_08703_, _08702_);
  or _59408_ (_08704_, _07357_, _07197_);
  or _59409_ (_08705_, _07198_, _07004_);
  and _59410_ (_08706_, _08705_, _08675_);
  nand _59411_ (_08707_, _08706_, _08704_);
  and _59412_ (_08708_, _08707_, _08703_);
  not _59413_ (_08709_, _08708_);
  or _59414_ (_08710_, _08700_, _07982_);
  and _59415_ (_08711_, _08710_, _08709_);
  nand _59416_ (_08712_, _08711_, _08701_);
  nand _59417_ (_08713_, _08700_, \oc8051_golden_model_1.IRAM[2] [7]);
  or _59418_ (_08714_, _08700_, _07986_);
  and _59419_ (_08715_, _08714_, _08708_);
  nand _59420_ (_08716_, _08715_, _08713_);
  nand _59421_ (_08717_, _08716_, _08712_);
  nand _59422_ (_08718_, _08717_, _08692_);
  not _59423_ (_08719_, _08692_);
  nand _59424_ (_08720_, _08700_, \oc8051_golden_model_1.IRAM[4] [7]);
  or _59425_ (_08721_, _08700_, _08002_);
  and _59426_ (_08722_, _08721_, _08709_);
  nand _59427_ (_08723_, _08722_, _08720_);
  nand _59428_ (_08724_, _08700_, \oc8051_golden_model_1.IRAM[6] [7]);
  or _59429_ (_08725_, _08700_, _07994_);
  and _59430_ (_08726_, _08725_, _08708_);
  nand _59431_ (_08727_, _08726_, _08724_);
  nand _59432_ (_08728_, _08727_, _08723_);
  nand _59433_ (_08729_, _08728_, _08719_);
  nand _59434_ (_08730_, _08729_, _08718_);
  nand _59435_ (_08731_, _08730_, _08682_);
  not _59436_ (_08732_, _08682_);
  nand _59437_ (_08733_, _08700_, \oc8051_golden_model_1.IRAM[10] [7]);
  or _59438_ (_08734_, _08700_, _08010_);
  and _59439_ (_08735_, _08734_, _08708_);
  nand _59440_ (_08736_, _08735_, _08733_);
  nand _59441_ (_08737_, _08700_, \oc8051_golden_model_1.IRAM[8] [7]);
  or _59442_ (_08738_, _08700_, _08018_);
  and _59443_ (_08739_, _08738_, _08709_);
  nand _59444_ (_08740_, _08739_, _08737_);
  nand _59445_ (_08741_, _08740_, _08736_);
  nand _59446_ (_08742_, _08741_, _08692_);
  nand _59447_ (_08743_, _08700_, \oc8051_golden_model_1.IRAM[12] [7]);
  or _59448_ (_08744_, _08700_, _08032_);
  and _59449_ (_08745_, _08744_, _08709_);
  nand _59450_ (_08746_, _08745_, _08743_);
  nand _59451_ (_08747_, _08700_, \oc8051_golden_model_1.IRAM[14] [7]);
  or _59452_ (_08748_, _08700_, _08024_);
  and _59453_ (_08749_, _08748_, _08708_);
  nand _59454_ (_08750_, _08749_, _08747_);
  nand _59455_ (_08751_, _08750_, _08746_);
  nand _59456_ (_08752_, _08751_, _08719_);
  nand _59457_ (_08753_, _08752_, _08742_);
  nand _59458_ (_08754_, _08753_, _08732_);
  and _59459_ (_08755_, _08754_, _08731_);
  or _59460_ (_08756_, _08755_, _07155_);
  and _59461_ (_08757_, _08756_, _08667_);
  and _59462_ (_08758_, _08757_, _08652_);
  and _59463_ (_08759_, _08543_, _08246_);
  not _59464_ (_08760_, _08390_);
  and _59465_ (_08761_, _08760_, _08340_);
  and _59466_ (_08762_, _08439_, _08291_);
  and _59467_ (_08763_, _08762_, _08761_);
  and _59468_ (_08764_, _08763_, _08759_);
  and _59469_ (_08765_, _08764_, _08144_);
  or _59470_ (_08766_, _08765_, _08043_);
  nand _59471_ (_08767_, _08765_, _08043_);
  and _59472_ (_08768_, _08767_, _08766_);
  and _59473_ (_08769_, _08768_, _07152_);
  or _59474_ (_08770_, _08769_, _08758_);
  and _59475_ (_08771_, _08770_, _08651_);
  not _59476_ (_08772_, _07950_);
  nand _59477_ (_08773_, _08648_, _08772_);
  and _59478_ (_08774_, _08773_, _06275_);
  or _59479_ (_08775_, _08774_, _07611_);
  or _59480_ (_08776_, _08775_, _08771_);
  nor _59481_ (_08777_, _08661_, _06010_);
  nor _59482_ (_08778_, _08777_, _07167_);
  and _59483_ (_08779_, _08778_, _08776_);
  and _59484_ (_08780_, _08552_, _07167_);
  or _59485_ (_08781_, _08780_, _07179_);
  or _59486_ (_08782_, _08781_, _08779_);
  and _59487_ (_08783_, _08782_, _08650_);
  or _59488_ (_08784_, _08783_, _06267_);
  nand _59489_ (_08785_, _08042_, _06267_);
  and _59490_ (_08786_, _08785_, _06265_);
  and _59491_ (_08787_, _08786_, _08784_);
  nor _59492_ (_08788_, _08648_, _08772_);
  not _59493_ (_08789_, _08788_);
  and _59494_ (_08790_, _08789_, _08773_);
  and _59495_ (_08791_, _08790_, _06264_);
  or _59496_ (_08792_, _08791_, _08787_);
  and _59497_ (_08793_, _08792_, _06007_);
  not _59498_ (_08794_, _08661_);
  or _59499_ (_08795_, _08794_, _06007_);
  nand _59500_ (_08796_, _08795_, _06501_);
  or _59501_ (_08797_, _08796_, _08793_);
  nand _59502_ (_08798_, _08042_, _06502_);
  and _59503_ (_08799_, _08798_, _08797_);
  or _59504_ (_08800_, _08799_, _07197_);
  not _59505_ (_08801_, _07196_);
  and _59506_ (_08802_, _08755_, _06286_);
  nand _59507_ (_08803_, _07979_, _07197_);
  or _59508_ (_08804_, _08803_, _08802_);
  and _59509_ (_08805_, _08804_, _08801_);
  and _59510_ (_08806_, _08805_, _08800_);
  and _59511_ (_08807_, _07950_, \oc8051_golden_model_1.PSW [7]);
  or _59512_ (_08808_, _08807_, _08649_);
  and _59513_ (_08809_, _08808_, _07196_);
  or _59514_ (_08810_, _08809_, _06254_);
  or _59515_ (_08811_, _08810_, _08806_);
  nor _59516_ (_08812_, _07215_, _06182_);
  nor _59517_ (_08813_, _08661_, _05978_);
  nor _59518_ (_08814_, _08813_, _08812_);
  and _59519_ (_08815_, _08814_, _08811_);
  nor _59520_ (_08816_, _07208_, _06182_);
  not _59521_ (_08817_, _08812_);
  nor _59522_ (_08818_, _08040_, _08817_);
  or _59523_ (_08819_, _08818_, _08816_);
  or _59524_ (_08820_, _08819_, _08815_);
  not _59525_ (_08821_, _08816_);
  or _59526_ (_08822_, _08755_, _08821_);
  and _59527_ (_08823_, _08822_, _07471_);
  and _59528_ (_08824_, _08823_, _08820_);
  not _59529_ (_08825_, _08608_);
  nor _59530_ (_08826_, _08825_, _08040_);
  and _59531_ (_08827_, _06423_, _04849_);
  and _59532_ (_08828_, _06445_, _04839_);
  nor _59533_ (_08829_, _08828_, _08827_);
  and _59534_ (_08830_, _06447_, _04851_);
  and _59535_ (_08831_, _06436_, _04823_);
  nor _59536_ (_08832_, _08831_, _08830_);
  and _59537_ (_08833_, _08832_, _08829_);
  and _59538_ (_08834_, _06411_, _04835_);
  and _59539_ (_08835_, _06431_, _04831_);
  nor _59540_ (_08836_, _08835_, _08834_);
  and _59541_ (_08837_, _06415_, _04855_);
  and _59542_ (_08838_, _06442_, _04816_);
  nor _59543_ (_08839_, _08838_, _08837_);
  and _59544_ (_08840_, _08839_, _08836_);
  and _59545_ (_08841_, _08840_, _08833_);
  and _59546_ (_08842_, _06434_, _04844_);
  and _59547_ (_08843_, _06429_, _04827_);
  nor _59548_ (_08844_, _08843_, _08842_);
  and _59549_ (_08845_, _06440_, _04837_);
  and _59550_ (_08846_, _06401_, _04818_);
  nor _59551_ (_08847_, _08846_, _08845_);
  and _59552_ (_08848_, _08847_, _08844_);
  and _59553_ (_08849_, _06407_, _04842_);
  and _59554_ (_08850_, _06398_, _04857_);
  nor _59555_ (_08851_, _08850_, _08849_);
  and _59556_ (_08852_, _06420_, _04829_);
  and _59557_ (_08853_, _06417_, _04821_);
  nor _59558_ (_08854_, _08853_, _08852_);
  and _59559_ (_08855_, _08854_, _08851_);
  and _59560_ (_08856_, _08855_, _08848_);
  and _59561_ (_08857_, _08856_, _08841_);
  and _59562_ (_08858_, _08857_, _08825_);
  and _59563_ (_08859_, _06407_, _04750_);
  and _59564_ (_08860_, _06442_, _04724_);
  nor _59565_ (_08861_, _08860_, _08859_);
  and _59566_ (_08862_, _06411_, _04743_);
  and _59567_ (_08863_, _06431_, _04739_);
  nor _59568_ (_08864_, _08863_, _08862_);
  and _59569_ (_08865_, _08864_, _08861_);
  and _59570_ (_08866_, _06445_, _04747_);
  and _59571_ (_08868_, _06429_, _04735_);
  nor _59572_ (_08869_, _08868_, _08866_);
  and _59573_ (_08870_, _06440_, _04745_);
  and _59574_ (_08871_, _06423_, _04757_);
  nor _59575_ (_08872_, _08871_, _08870_);
  and _59576_ (_08873_, _08872_, _08869_);
  and _59577_ (_08874_, _08873_, _08865_);
  and _59578_ (_08875_, _06447_, _04759_);
  and _59579_ (_08876_, _06398_, _04765_);
  nor _59580_ (_08877_, _08876_, _08875_);
  and _59581_ (_08879_, _06436_, _04731_);
  and _59582_ (_08880_, _06401_, _04726_);
  nor _59583_ (_08881_, _08880_, _08879_);
  and _59584_ (_08882_, _08881_, _08877_);
  and _59585_ (_08883_, _06417_, _04729_);
  and _59586_ (_08884_, _06415_, _04763_);
  nor _59587_ (_08885_, _08884_, _08883_);
  and _59588_ (_08886_, _06420_, _04737_);
  and _59589_ (_08887_, _06434_, _04752_);
  nor _59590_ (_08888_, _08887_, _08886_);
  and _59591_ (_08890_, _08888_, _08885_);
  and _59592_ (_08891_, _08890_, _08882_);
  and _59593_ (_08892_, _08891_, _08874_);
  and _59594_ (_08893_, _06445_, _04793_);
  and _59595_ (_08894_, _06401_, _04772_);
  nor _59596_ (_08895_, _08894_, _08893_);
  and _59597_ (_08896_, _06440_, _04791_);
  and _59598_ (_08897_, _06431_, _04781_);
  nor _59599_ (_08898_, _08897_, _08896_);
  and _59600_ (_08899_, _08898_, _08895_);
  and _59601_ (_08901_, _06420_, _04783_);
  and _59602_ (_08902_, _06423_, _04785_);
  nor _59603_ (_08903_, _08902_, _08901_);
  and _59604_ (_08904_, _06434_, _04798_);
  and _59605_ (_08905_, _06429_, _04805_);
  nor _59606_ (_08906_, _08905_, _08904_);
  and _59607_ (_08907_, _08906_, _08903_);
  and _59608_ (_08908_, _08907_, _08899_);
  and _59609_ (_08909_, _06415_, _04809_);
  and _59610_ (_08910_, _06442_, _04770_);
  nor _59611_ (_08912_, _08910_, _08909_);
  and _59612_ (_08913_, _06436_, _04777_);
  and _59613_ (_08914_, _06398_, _04811_);
  nor _59614_ (_08915_, _08914_, _08913_);
  and _59615_ (_08916_, _08915_, _08912_);
  and _59616_ (_08917_, _06407_, _04796_);
  and _59617_ (_08918_, _06447_, _04803_);
  nor _59618_ (_08919_, _08918_, _08917_);
  and _59619_ (_08920_, _06411_, _04789_);
  and _59620_ (_08921_, _06417_, _04775_);
  nor _59621_ (_08923_, _08921_, _08920_);
  and _59622_ (_08924_, _08923_, _08919_);
  and _59623_ (_08925_, _08924_, _08916_);
  and _59624_ (_08926_, _08925_, _08908_);
  and _59625_ (_08927_, _08926_, _08892_);
  and _59626_ (_08928_, _08927_, _08858_);
  and _59627_ (_08929_, _07038_, _06872_);
  not _59628_ (_08930_, _06452_);
  and _59629_ (_08931_, _06697_, _08930_);
  and _59630_ (_08932_, _08931_, _08929_);
  and _59631_ (_08934_, _08932_, _08928_);
  and _59632_ (_08935_, _08934_, \oc8051_golden_model_1.TCON [7]);
  not _59633_ (_08936_, _07038_);
  and _59634_ (_08937_, _08936_, _06872_);
  and _59635_ (_08938_, _08937_, _08931_);
  and _59636_ (_08939_, _08938_, _08928_);
  and _59637_ (_08940_, _08939_, \oc8051_golden_model_1.TL0 [7]);
  or _59638_ (_08941_, _08940_, _08935_);
  and _59639_ (_08942_, _06697_, _06452_);
  and _59640_ (_08943_, _08942_, _08929_);
  and _59641_ (_08944_, _08943_, _08928_);
  and _59642_ (_08945_, _08944_, \oc8051_golden_model_1.P0 [7]);
  not _59643_ (_08946_, _08926_);
  and _59644_ (_08947_, _08946_, _08892_);
  nor _59645_ (_08948_, _08857_, _08608_);
  and _59646_ (_08949_, _08948_, _08943_);
  and _59647_ (_08950_, _08949_, _08947_);
  and _59648_ (_08951_, _08950_, \oc8051_golden_model_1.ACC [7]);
  or _59649_ (_08952_, _08951_, _08945_);
  or _59650_ (_08953_, _08952_, _08941_);
  not _59651_ (_08954_, _06872_);
  and _59652_ (_08955_, _07038_, _08954_);
  and _59653_ (_08956_, _08955_, _08931_);
  and _59654_ (_08957_, _08956_, _08928_);
  and _59655_ (_08958_, _08957_, \oc8051_golden_model_1.TMOD [7]);
  not _59656_ (_08959_, _08892_);
  and _59657_ (_08960_, _08926_, _08959_);
  and _59658_ (_08961_, _08960_, _08858_);
  and _59659_ (_08962_, _08961_, _08943_);
  and _59660_ (_08963_, _08962_, \oc8051_golden_model_1.P1 [7]);
  or _59661_ (_08964_, _08963_, _08958_);
  and _59662_ (_08965_, _08961_, _08932_);
  and _59663_ (_08966_, _08965_, \oc8051_golden_model_1.SCON [7]);
  nor _59664_ (_08967_, _08926_, _08892_);
  and _59665_ (_08968_, _08967_, _08949_);
  and _59666_ (_08969_, _08968_, \oc8051_golden_model_1.B [7]);
  or _59667_ (_08970_, _08969_, _08966_);
  or _59668_ (_08971_, _08970_, _08964_);
  or _59669_ (_08972_, _08971_, _08953_);
  not _59670_ (_08973_, _06697_);
  nor _59671_ (_08974_, _07038_, _06872_);
  and _59672_ (_08975_, _08974_, _08928_);
  and _59673_ (_08976_, _08975_, _06452_);
  and _59674_ (_08977_, _08976_, _08973_);
  and _59675_ (_08978_, _08977_, \oc8051_golden_model_1.PCON [7]);
  and _59676_ (_08979_, _08976_, _06697_);
  and _59677_ (_08980_, _08979_, \oc8051_golden_model_1.DPH [7]);
  or _59678_ (_08981_, _08980_, _08978_);
  or _59679_ (_08982_, _08981_, _08972_);
  and _59680_ (_08983_, _08942_, _08928_);
  and _59681_ (_08984_, _08983_, _08937_);
  and _59682_ (_08985_, _08984_, \oc8051_golden_model_1.DPL [7]);
  and _59683_ (_08986_, _08975_, _08931_);
  and _59684_ (_08987_, _08986_, \oc8051_golden_model_1.TL1 [7]);
  and _59685_ (_08988_, _08955_, _08983_);
  and _59686_ (_08989_, _08988_, \oc8051_golden_model_1.SP [7]);
  or _59687_ (_08990_, _08989_, _08987_);
  or _59688_ (_08991_, _08990_, _08985_);
  and _59689_ (_08992_, _08947_, _08858_);
  and _59690_ (_08993_, _08992_, _08932_);
  and _59691_ (_08994_, _08993_, \oc8051_golden_model_1.IE [7]);
  and _59692_ (_08995_, _08967_, _08858_);
  and _59693_ (_08996_, _08995_, _08932_);
  and _59694_ (_08997_, _08996_, \oc8051_golden_model_1.IP [7]);
  or _59695_ (_08998_, _08997_, _08994_);
  and _59696_ (_08999_, _08992_, _08943_);
  and _59697_ (_09000_, _08999_, \oc8051_golden_model_1.P2 [7]);
  and _59698_ (_09001_, _08995_, _08943_);
  and _59699_ (_09002_, _09001_, \oc8051_golden_model_1.P3 [7]);
  or _59700_ (_09003_, _09002_, _09000_);
  or _59701_ (_09004_, _09003_, _08998_);
  and _59702_ (_09005_, _08961_, _08956_);
  and _59703_ (_09006_, _09005_, \oc8051_golden_model_1.SBUF [7]);
  and _59704_ (_09007_, _08960_, _08949_);
  and _59705_ (_09008_, _09007_, \oc8051_golden_model_1.PSW [7]);
  or _59706_ (_09009_, _09008_, _09006_);
  or _59707_ (_09010_, _09009_, _09004_);
  nor _59708_ (_09011_, _06697_, _06452_);
  and _59709_ (_09012_, _09011_, _08928_);
  and _59710_ (_09013_, _09012_, _08929_);
  and _59711_ (_09014_, _09013_, \oc8051_golden_model_1.TH0 [7]);
  and _59712_ (_09015_, _09012_, _08955_);
  and _59713_ (_09016_, _09015_, \oc8051_golden_model_1.TH1 [7]);
  or _59714_ (_09017_, _09016_, _09014_);
  or _59715_ (_09018_, _09017_, _09010_);
  or _59716_ (_09019_, _09018_, _08991_);
  or _59717_ (_09020_, _09019_, _08982_);
  or _59718_ (_09021_, _09020_, _08826_);
  and _59719_ (_09022_, _09021_, _07470_);
  nor _59720_ (_09023_, _07211_, _05951_);
  not _59721_ (_09024_, _09023_);
  nor _59722_ (_09025_, _07212_, _05951_);
  not _59723_ (_09026_, _09025_);
  and _59724_ (_09027_, _07209_, _06321_);
  nor _59725_ (_09028_, _09027_, _07224_);
  and _59726_ (_09029_, _09028_, _09026_);
  and _59727_ (_09030_, _09029_, _09024_);
  not _59728_ (_09031_, _09030_);
  or _59729_ (_09032_, _09031_, _09022_);
  or _59730_ (_09033_, _09032_, _08824_);
  or _59731_ (_09034_, _09030_, _06182_);
  and _59732_ (_09035_, _09034_, _09033_);
  or _59733_ (_09036_, _09035_, _06220_);
  and _59734_ (_09037_, _09036_, _08609_);
  or _59735_ (_09038_, _09037_, _06217_);
  nor _59736_ (_09039_, _08661_, _05952_);
  nor _59737_ (_09040_, _09039_, _07238_);
  and _59738_ (_09041_, _09040_, _09038_);
  nor _59739_ (_09042_, _08608_, _08042_);
  and _59740_ (_09043_, _08608_, _08042_);
  nor _59741_ (_09044_, _09043_, _09042_);
  and _59742_ (_09045_, _09044_, _07238_);
  or _59743_ (_09046_, _09045_, _09041_);
  and _59744_ (_09047_, _09046_, _08577_);
  or _59745_ (_09048_, _09047_, _08576_);
  and _59746_ (_09049_, _09048_, _08571_);
  and _59747_ (_09050_, _09042_, _07243_);
  or _59748_ (_09051_, _09050_, _09049_);
  and _59749_ (_09052_, _09051_, _07236_);
  and _59750_ (_09053_, _08574_, _07235_);
  or _59751_ (_09054_, _09053_, _07233_);
  or _59752_ (_09055_, _09054_, _09052_);
  not _59753_ (_09056_, _06366_);
  nor _59754_ (_09057_, _09056_, _06182_);
  nor _59755_ (_09058_, _08661_, _05961_);
  nor _59756_ (_09059_, _09058_, _09057_);
  and _59757_ (_09060_, _09059_, _09055_);
  not _59758_ (_09061_, _06528_);
  nor _59759_ (_09062_, _09061_, _06182_);
  not _59760_ (_09063_, _09043_);
  and _59761_ (_09064_, _09063_, _09057_);
  or _59762_ (_09065_, _09064_, _09062_);
  or _59763_ (_09066_, _09065_, _09060_);
  nand _59764_ (_09067_, _08573_, _09062_);
  and _59765_ (_09068_, _09067_, _05959_);
  and _59766_ (_09069_, _09068_, _09066_);
  or _59767_ (_09070_, _08794_, _05959_);
  nand _59768_ (_09071_, _09070_, _08569_);
  or _59769_ (_09072_, _09071_, _09069_);
  and _59770_ (_09073_, _09072_, _08570_);
  or _59771_ (_09074_, _09073_, _07435_);
  not _59772_ (_09075_, _07261_);
  not _59773_ (_09076_, _08755_);
  nand _59774_ (_09077_, _08700_, \oc8051_golden_model_1.IRAM[0] [6]);
  or _59775_ (_09078_, _08700_, _08092_);
  and _59776_ (_09079_, _09078_, _08709_);
  nand _59777_ (_09080_, _09079_, _09077_);
  nand _59778_ (_09081_, _08700_, \oc8051_golden_model_1.IRAM[2] [6]);
  or _59779_ (_09082_, _08700_, _08096_);
  and _59780_ (_09083_, _09082_, _08708_);
  nand _59781_ (_09084_, _09083_, _09081_);
  nand _59782_ (_09085_, _09084_, _09080_);
  nand _59783_ (_09086_, _09085_, _08692_);
  nand _59784_ (_09087_, _08700_, \oc8051_golden_model_1.IRAM[4] [6]);
  or _59785_ (_09088_, _08700_, _08112_);
  and _59786_ (_09089_, _09088_, _08709_);
  nand _59787_ (_09090_, _09089_, _09087_);
  nand _59788_ (_09091_, _08700_, \oc8051_golden_model_1.IRAM[6] [6]);
  or _59789_ (_09092_, _08700_, _08104_);
  and _59790_ (_09093_, _09092_, _08708_);
  nand _59791_ (_09094_, _09093_, _09091_);
  nand _59792_ (_09095_, _09094_, _09090_);
  nand _59793_ (_09096_, _09095_, _08719_);
  and _59794_ (_09097_, _09096_, _08682_);
  and _59795_ (_09098_, _09097_, _09086_);
  not _59796_ (_09099_, _08700_);
  or _59797_ (_09100_, _09099_, \oc8051_golden_model_1.IRAM[10] [6]);
  or _59798_ (_09101_, _08700_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _59799_ (_09102_, _09101_, _09100_);
  nand _59800_ (_09103_, _09102_, _08708_);
  or _59801_ (_09104_, _09099_, \oc8051_golden_model_1.IRAM[8] [6]);
  or _59802_ (_09105_, _08700_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand _59803_ (_09106_, _09105_, _09104_);
  nand _59804_ (_09107_, _09106_, _08709_);
  nand _59805_ (_09108_, _09107_, _09103_);
  nand _59806_ (_09109_, _09108_, _08692_);
  or _59807_ (_09110_, _09099_, \oc8051_golden_model_1.IRAM[14] [6]);
  or _59808_ (_09111_, _08700_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _59809_ (_09112_, _09111_, _09110_);
  nand _59810_ (_09113_, _09112_, _08708_);
  or _59811_ (_09114_, _09099_, \oc8051_golden_model_1.IRAM[12] [6]);
  or _59812_ (_09115_, _08700_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand _59813_ (_09116_, _09115_, _09114_);
  nand _59814_ (_09117_, _09116_, _08709_);
  nand _59815_ (_09118_, _09117_, _09113_);
  nand _59816_ (_09119_, _09118_, _08719_);
  and _59817_ (_09120_, _09119_, _08732_);
  and _59818_ (_09121_, _09120_, _09109_);
  nor _59819_ (_09122_, _09121_, _09098_);
  nand _59820_ (_09123_, _08700_, \oc8051_golden_model_1.IRAM[0] [5]);
  or _59821_ (_09124_, _08700_, _08194_);
  and _59822_ (_09125_, _09124_, _08709_);
  nand _59823_ (_09126_, _09125_, _09123_);
  nand _59824_ (_09127_, _08700_, \oc8051_golden_model_1.IRAM[2] [5]);
  or _59825_ (_09128_, _08700_, _08198_);
  and _59826_ (_09129_, _09128_, _08708_);
  nand _59827_ (_09130_, _09129_, _09127_);
  nand _59828_ (_09131_, _09130_, _09126_);
  nand _59829_ (_09132_, _09131_, _08692_);
  nand _59830_ (_09133_, _08700_, \oc8051_golden_model_1.IRAM[4] [5]);
  or _59831_ (_09134_, _08700_, _08214_);
  and _59832_ (_09135_, _09134_, _08709_);
  nand _59833_ (_09136_, _09135_, _09133_);
  nand _59834_ (_09137_, _08700_, \oc8051_golden_model_1.IRAM[6] [5]);
  or _59835_ (_09138_, _08700_, _08206_);
  and _59836_ (_09139_, _09138_, _08708_);
  nand _59837_ (_09140_, _09139_, _09137_);
  nand _59838_ (_09141_, _09140_, _09136_);
  nand _59839_ (_09142_, _09141_, _08719_);
  and _59840_ (_09143_, _09142_, _08682_);
  and _59841_ (_09144_, _09143_, _09132_);
  or _59842_ (_09145_, _09099_, \oc8051_golden_model_1.IRAM[10] [5]);
  or _59843_ (_09146_, _08700_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _59844_ (_09147_, _09146_, _09145_);
  nand _59845_ (_09148_, _09147_, _08708_);
  or _59846_ (_09149_, _09099_, \oc8051_golden_model_1.IRAM[8] [5]);
  or _59847_ (_09150_, _08700_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand _59848_ (_09151_, _09150_, _09149_);
  nand _59849_ (_09152_, _09151_, _08709_);
  nand _59850_ (_09153_, _09152_, _09148_);
  nand _59851_ (_09154_, _09153_, _08692_);
  or _59852_ (_09155_, _09099_, \oc8051_golden_model_1.IRAM[14] [5]);
  or _59853_ (_09156_, _08700_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _59854_ (_09157_, _09156_, _09155_);
  nand _59855_ (_09158_, _09157_, _08708_);
  or _59856_ (_09159_, _09099_, \oc8051_golden_model_1.IRAM[12] [5]);
  or _59857_ (_09160_, _08700_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand _59858_ (_09161_, _09160_, _09159_);
  nand _59859_ (_09162_, _09161_, _08709_);
  nand _59860_ (_09163_, _09162_, _09158_);
  nand _59861_ (_09164_, _09163_, _08719_);
  and _59862_ (_09165_, _09164_, _08732_);
  and _59863_ (_09166_, _09165_, _09154_);
  nor _59864_ (_09167_, _09166_, _09144_);
  nand _59865_ (_09168_, _08700_, \oc8051_golden_model_1.IRAM[0] [4]);
  or _59866_ (_09169_, _08700_, _08491_);
  and _59867_ (_09170_, _09169_, _08709_);
  nand _59868_ (_09171_, _09170_, _09168_);
  nand _59869_ (_09172_, _08700_, \oc8051_golden_model_1.IRAM[2] [4]);
  or _59870_ (_09173_, _08700_, _08495_);
  and _59871_ (_09174_, _09173_, _08708_);
  nand _59872_ (_09175_, _09174_, _09172_);
  nand _59873_ (_09176_, _09175_, _09171_);
  nand _59874_ (_09177_, _09176_, _08692_);
  nand _59875_ (_09178_, _08700_, \oc8051_golden_model_1.IRAM[4] [4]);
  or _59876_ (_09179_, _08700_, _08511_);
  and _59877_ (_09180_, _09179_, _08709_);
  nand _59878_ (_09181_, _09180_, _09178_);
  nand _59879_ (_09182_, _08700_, \oc8051_golden_model_1.IRAM[6] [4]);
  or _59880_ (_09183_, _08700_, _08503_);
  and _59881_ (_09184_, _09183_, _08708_);
  nand _59882_ (_09185_, _09184_, _09182_);
  nand _59883_ (_09186_, _09185_, _09181_);
  nand _59884_ (_09187_, _09186_, _08719_);
  and _59885_ (_09188_, _09187_, _08682_);
  and _59886_ (_09189_, _09188_, _09177_);
  or _59887_ (_09190_, _09099_, \oc8051_golden_model_1.IRAM[10] [4]);
  or _59888_ (_09191_, _08700_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _59889_ (_09192_, _09191_, _09190_);
  nand _59890_ (_09193_, _09192_, _08708_);
  or _59891_ (_09194_, _09099_, \oc8051_golden_model_1.IRAM[8] [4]);
  or _59892_ (_09195_, _08700_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand _59893_ (_09196_, _09195_, _09194_);
  nand _59894_ (_09197_, _09196_, _08709_);
  nand _59895_ (_09198_, _09197_, _09193_);
  nand _59896_ (_09199_, _09198_, _08692_);
  or _59897_ (_09200_, _09099_, \oc8051_golden_model_1.IRAM[14] [4]);
  or _59898_ (_09201_, _08700_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _59899_ (_09202_, _09201_, _09200_);
  nand _59900_ (_09203_, _09202_, _08708_);
  or _59901_ (_09204_, _09099_, \oc8051_golden_model_1.IRAM[12] [4]);
  or _59902_ (_09205_, _08700_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand _59903_ (_09206_, _09205_, _09204_);
  nand _59904_ (_09207_, _09206_, _08709_);
  nand _59905_ (_09208_, _09207_, _09203_);
  nand _59906_ (_09209_, _09208_, _08719_);
  and _59907_ (_09210_, _09209_, _08732_);
  and _59908_ (_09211_, _09210_, _09199_);
  nor _59909_ (_09212_, _09211_, _09189_);
  nand _59910_ (_09213_, _08700_, \oc8051_golden_model_1.IRAM[0] [3]);
  or _59911_ (_09214_, _08700_, _07544_);
  and _59912_ (_09215_, _09214_, _08709_);
  nand _59913_ (_09216_, _09215_, _09213_);
  nand _59914_ (_09217_, _08700_, \oc8051_golden_model_1.IRAM[2] [3]);
  or _59915_ (_09218_, _08700_, _07548_);
  and _59916_ (_09219_, _09218_, _08708_);
  nand _59917_ (_09220_, _09219_, _09217_);
  nand _59918_ (_09221_, _09220_, _09216_);
  nand _59919_ (_09222_, _09221_, _08692_);
  nand _59920_ (_09223_, _08700_, \oc8051_golden_model_1.IRAM[4] [3]);
  or _59921_ (_09224_, _08700_, _07564_);
  and _59922_ (_09225_, _09224_, _08709_);
  nand _59923_ (_09226_, _09225_, _09223_);
  nand _59924_ (_09227_, _08700_, \oc8051_golden_model_1.IRAM[6] [3]);
  or _59925_ (_09228_, _08700_, _07556_);
  and _59926_ (_09229_, _09228_, _08708_);
  nand _59927_ (_09230_, _09229_, _09227_);
  nand _59928_ (_09231_, _09230_, _09226_);
  nand _59929_ (_09232_, _09231_, _08719_);
  and _59930_ (_09233_, _09232_, _08682_);
  and _59931_ (_09234_, _09233_, _09222_);
  or _59932_ (_09235_, _09099_, \oc8051_golden_model_1.IRAM[10] [3]);
  or _59933_ (_09236_, _08700_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _59934_ (_09237_, _09236_, _09235_);
  nand _59935_ (_09238_, _09237_, _08708_);
  or _59936_ (_09239_, _09099_, \oc8051_golden_model_1.IRAM[8] [3]);
  or _59937_ (_09240_, _08700_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand _59938_ (_09241_, _09240_, _09239_);
  nand _59939_ (_09242_, _09241_, _08709_);
  nand _59940_ (_09243_, _09242_, _09238_);
  nand _59941_ (_09244_, _09243_, _08692_);
  or _59942_ (_09245_, _09099_, \oc8051_golden_model_1.IRAM[14] [3]);
  or _59943_ (_09246_, _08700_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _59944_ (_09247_, _09246_, _09245_);
  nand _59945_ (_09248_, _09247_, _08708_);
  or _59946_ (_09249_, _09099_, \oc8051_golden_model_1.IRAM[12] [3]);
  or _59947_ (_09250_, _08700_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand _59948_ (_09251_, _09250_, _09249_);
  nand _59949_ (_09252_, _09251_, _08709_);
  nand _59950_ (_09253_, _09252_, _09248_);
  nand _59951_ (_09254_, _09253_, _08719_);
  and _59952_ (_09255_, _09254_, _08732_);
  and _59953_ (_09256_, _09255_, _09244_);
  nor _59954_ (_09257_, _09256_, _09234_);
  nand _59955_ (_09258_, _08700_, \oc8051_golden_model_1.IRAM[0] [2]);
  or _59956_ (_09259_, _08700_, _07724_);
  and _59957_ (_09260_, _09259_, _08709_);
  nand _59958_ (_09261_, _09260_, _09258_);
  nand _59959_ (_09262_, _08700_, \oc8051_golden_model_1.IRAM[2] [2]);
  or _59960_ (_09263_, _08700_, _07728_);
  and _59961_ (_09264_, _09263_, _08708_);
  nand _59962_ (_09265_, _09264_, _09262_);
  nand _59963_ (_09266_, _09265_, _09261_);
  nand _59964_ (_09267_, _09266_, _08692_);
  nand _59965_ (_09268_, _08700_, \oc8051_golden_model_1.IRAM[4] [2]);
  or _59966_ (_09269_, _08700_, _07744_);
  and _59967_ (_09270_, _09269_, _08709_);
  nand _59968_ (_09271_, _09270_, _09268_);
  nand _59969_ (_09272_, _08700_, \oc8051_golden_model_1.IRAM[6] [2]);
  or _59970_ (_09273_, _08700_, _07736_);
  and _59971_ (_09274_, _09273_, _08708_);
  nand _59972_ (_09275_, _09274_, _09272_);
  nand _59973_ (_09276_, _09275_, _09271_);
  nand _59974_ (_09277_, _09276_, _08719_);
  and _59975_ (_09278_, _09277_, _08682_);
  and _59976_ (_09279_, _09278_, _09267_);
  or _59977_ (_09280_, _09099_, \oc8051_golden_model_1.IRAM[10] [2]);
  or _59978_ (_09281_, _08700_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _59979_ (_09282_, _09281_, _09280_);
  nand _59980_ (_09283_, _09282_, _08708_);
  or _59981_ (_09284_, _09099_, \oc8051_golden_model_1.IRAM[8] [2]);
  or _59982_ (_09285_, _08700_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand _59983_ (_09286_, _09285_, _09284_);
  nand _59984_ (_09287_, _09286_, _08709_);
  nand _59985_ (_09288_, _09287_, _09283_);
  nand _59986_ (_09289_, _09288_, _08692_);
  nand _59987_ (_09290_, _08700_, _07764_);
  or _59988_ (_09291_, _08700_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _59989_ (_09292_, _09291_, _09290_);
  nand _59990_ (_09293_, _09292_, _08708_);
  or _59991_ (_09294_, _09099_, \oc8051_golden_model_1.IRAM[12] [2]);
  or _59992_ (_09295_, _08700_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand _59993_ (_09296_, _09295_, _09294_);
  nand _59994_ (_09297_, _09296_, _08709_);
  nand _59995_ (_09298_, _09297_, _09293_);
  nand _59996_ (_09299_, _09298_, _08719_);
  and _59997_ (_09300_, _09299_, _08732_);
  and _59998_ (_09301_, _09300_, _09289_);
  nor _59999_ (_09302_, _09301_, _09279_);
  nand _60000_ (_09303_, _08700_, \oc8051_golden_model_1.IRAM[0] [1]);
  or _60001_ (_09304_, _08700_, _07307_);
  and _60002_ (_09305_, _09304_, _08709_);
  nand _60003_ (_09306_, _09305_, _09303_);
  nand _60004_ (_09307_, _08700_, \oc8051_golden_model_1.IRAM[2] [1]);
  or _60005_ (_09308_, _08700_, _07311_);
  and _60006_ (_09309_, _09308_, _08708_);
  nand _60007_ (_09310_, _09309_, _09307_);
  nand _60008_ (_09311_, _09310_, _09306_);
  nand _60009_ (_09312_, _09311_, _08692_);
  nand _60010_ (_09313_, _08700_, \oc8051_golden_model_1.IRAM[4] [1]);
  or _60011_ (_09314_, _08700_, _07327_);
  and _60012_ (_09315_, _09314_, _08709_);
  nand _60013_ (_09316_, _09315_, _09313_);
  nand _60014_ (_09317_, _08700_, \oc8051_golden_model_1.IRAM[6] [1]);
  or _60015_ (_09318_, _08700_, _07319_);
  and _60016_ (_09319_, _09318_, _08708_);
  nand _60017_ (_09320_, _09319_, _09317_);
  nand _60018_ (_09321_, _09320_, _09316_);
  nand _60019_ (_09322_, _09321_, _08719_);
  and _60020_ (_09323_, _09322_, _08682_);
  and _60021_ (_09324_, _09323_, _09312_);
  or _60022_ (_09325_, _09099_, \oc8051_golden_model_1.IRAM[10] [1]);
  or _60023_ (_09326_, _08700_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _60024_ (_09327_, _09326_, _09325_);
  nand _60025_ (_09328_, _09327_, _08708_);
  or _60026_ (_09329_, _09099_, \oc8051_golden_model_1.IRAM[8] [1]);
  or _60027_ (_09330_, _08700_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand _60028_ (_09331_, _09330_, _09329_);
  nand _60029_ (_09332_, _09331_, _08709_);
  nand _60030_ (_09333_, _09332_, _09328_);
  nand _60031_ (_09334_, _09333_, _08692_);
  or _60032_ (_09335_, _09099_, \oc8051_golden_model_1.IRAM[14] [1]);
  or _60033_ (_09336_, _08700_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _60034_ (_09337_, _09336_, _09335_);
  nand _60035_ (_09338_, _09337_, _08708_);
  or _60036_ (_09339_, _09099_, \oc8051_golden_model_1.IRAM[12] [1]);
  or _60037_ (_09340_, _08700_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand _60038_ (_09341_, _09340_, _09339_);
  nand _60039_ (_09342_, _09341_, _08709_);
  nand _60040_ (_09343_, _09342_, _09338_);
  nand _60041_ (_09344_, _09343_, _08719_);
  and _60042_ (_09345_, _09344_, _08732_);
  and _60043_ (_09346_, _09345_, _09334_);
  nor _60044_ (_09347_, _09346_, _09324_);
  nand _60045_ (_09348_, _08700_, \oc8051_golden_model_1.IRAM[0] [0]);
  or _60046_ (_09349_, _08700_, _07077_);
  and _60047_ (_09350_, _09349_, _08709_);
  nand _60048_ (_09351_, _09350_, _09348_);
  nand _60049_ (_09352_, _08700_, \oc8051_golden_model_1.IRAM[2] [0]);
  or _60050_ (_09353_, _08700_, _07082_);
  and _60051_ (_09354_, _09353_, _08708_);
  nand _60052_ (_09355_, _09354_, _09352_);
  nand _60053_ (_09356_, _09355_, _09351_);
  nand _60054_ (_09357_, _09356_, _08692_);
  nand _60055_ (_09358_, _08700_, \oc8051_golden_model_1.IRAM[4] [0]);
  or _60056_ (_09359_, _08700_, _07100_);
  and _60057_ (_09360_, _09359_, _08709_);
  nand _60058_ (_09361_, _09360_, _09358_);
  nand _60059_ (_09362_, _08700_, \oc8051_golden_model_1.IRAM[6] [0]);
  or _60060_ (_09363_, _08700_, _07092_);
  and _60061_ (_09364_, _09363_, _08708_);
  nand _60062_ (_09365_, _09364_, _09362_);
  nand _60063_ (_09366_, _09365_, _09361_);
  nand _60064_ (_09367_, _09366_, _08719_);
  and _60065_ (_09368_, _09367_, _08682_);
  and _60066_ (_09369_, _09368_, _09357_);
  or _60067_ (_09370_, _09099_, \oc8051_golden_model_1.IRAM[10] [0]);
  or _60068_ (_09371_, _08700_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _60069_ (_09372_, _09371_, _09370_);
  nand _60070_ (_09373_, _09372_, _08708_);
  or _60071_ (_09374_, _09099_, \oc8051_golden_model_1.IRAM[8] [0]);
  or _60072_ (_09375_, _08700_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand _60073_ (_09376_, _09375_, _09374_);
  nand _60074_ (_09377_, _09376_, _08709_);
  nand _60075_ (_09378_, _09377_, _09373_);
  nand _60076_ (_09379_, _09378_, _08692_);
  nand _60077_ (_09380_, _08700_, \oc8051_golden_model_1.IRAM[14] [0]);
  or _60078_ (_09381_, _08700_, _07119_);
  and _60079_ (_09382_, _09381_, _09380_);
  nand _60080_ (_09383_, _09382_, _08708_);
  nand _60081_ (_09384_, _08700_, _07124_);
  or _60082_ (_09385_, _08700_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand _60083_ (_09386_, _09385_, _09384_);
  nand _60084_ (_09387_, _09386_, _08709_);
  nand _60085_ (_09388_, _09387_, _09383_);
  nand _60086_ (_09389_, _09388_, _08719_);
  and _60087_ (_09390_, _09389_, _08732_);
  and _60088_ (_09391_, _09390_, _09379_);
  or _60089_ (_09392_, _09391_, _09369_);
  not _60090_ (_09393_, _09392_);
  and _60091_ (_09394_, _09393_, _09347_);
  and _60092_ (_09395_, _09394_, _09302_);
  and _60093_ (_09396_, _09395_, _09257_);
  and _60094_ (_09397_, _09396_, _09212_);
  and _60095_ (_09398_, _09397_, _09167_);
  and _60096_ (_09399_, _09398_, _09122_);
  nor _60097_ (_09400_, _09399_, _09076_);
  and _60098_ (_09401_, _09399_, _09076_);
  or _60099_ (_09402_, _09401_, _09400_);
  or _60100_ (_09403_, _09402_, _07541_);
  and _60101_ (_09404_, _09403_, _09075_);
  and _60102_ (_09405_, _09404_, _09074_);
  and _60103_ (_09406_, _08768_, _07261_);
  or _60104_ (_09407_, _09406_, _06361_);
  or _60105_ (_09408_, _09407_, _09405_);
  and _60106_ (_09409_, _08657_, \oc8051_golden_model_1.PC [7]);
  and _60107_ (_09410_, _05634_, \oc8051_golden_model_1.PC [2]);
  and _60108_ (_09411_, _09410_, \oc8051_golden_model_1.PC [3]);
  and _60109_ (_09412_, _09411_, _09409_);
  and _60110_ (_09413_, _09411_, _08657_);
  nor _60111_ (_09414_, _09413_, \oc8051_golden_model_1.PC [7]);
  nor _60112_ (_09415_, _09414_, _09412_);
  not _60113_ (_09416_, _09415_);
  nand _60114_ (_09417_, _09416_, _06361_);
  and _60115_ (_09418_, _09417_, _09408_);
  or _60116_ (_09419_, _09418_, _05940_);
  and _60117_ (_09420_, _08794_, _05940_);
  nor _60118_ (_09421_, _09420_, _07270_);
  and _60119_ (_09422_, _09421_, _09419_);
  and _60120_ (_09423_, _08649_, _07270_);
  and _60121_ (_09424_, _05938_, _05923_);
  or _60122_ (_09425_, _09424_, _09423_);
  or _60123_ (_09426_, _09425_, _09422_);
  not _60124_ (_09427_, _09424_);
  not _60125_ (_09428_, _08142_);
  not _60126_ (_09429_, _08244_);
  not _60127_ (_09430_, _08541_);
  not _60128_ (_09431_, _07776_);
  not _60129_ (_09432_, _07357_);
  and _60130_ (_09433_, _09432_, _07133_);
  and _60131_ (_09434_, _09433_, _09431_);
  and _60132_ (_09435_, _09434_, _07595_);
  and _60133_ (_09436_, _09435_, _09430_);
  and _60134_ (_09437_, _09436_, _09429_);
  and _60135_ (_09438_, _09437_, _09428_);
  nand _60136_ (_09439_, _09438_, _08552_);
  or _60137_ (_09440_, _09438_, _08552_);
  and _60138_ (_09441_, _09440_, _09439_);
  or _60139_ (_09442_, _09441_, _09427_);
  and _60140_ (_09443_, _09442_, _09426_);
  or _60141_ (_09444_, _09443_, _07281_);
  not _60142_ (_09445_, _07286_);
  or _60143_ (_09446_, _09121_, _09098_);
  or _60144_ (_09447_, _09166_, _09144_);
  or _60145_ (_09448_, _09211_, _09189_);
  or _60146_ (_09449_, _09256_, _09234_);
  or _60147_ (_09450_, _09301_, _09279_);
  or _60148_ (_09451_, _09346_, _09324_);
  and _60149_ (_09452_, _09392_, _09451_);
  and _60150_ (_09453_, _09452_, _09450_);
  and _60151_ (_09454_, _09453_, _09449_);
  and _60152_ (_09455_, _09454_, _09448_);
  and _60153_ (_09456_, _09455_, _09447_);
  and _60154_ (_09457_, _09456_, _09446_);
  nor _60155_ (_09458_, _09457_, _09076_);
  and _60156_ (_09459_, _09457_, _09076_);
  or _60157_ (_09460_, _09459_, _09458_);
  or _60158_ (_09461_, _09460_, _07282_);
  and _60159_ (_09462_, _09461_, _09445_);
  and _60160_ (_09463_, _09462_, _09444_);
  or _60161_ (_09464_, _09463_, _08551_);
  and _60162_ (_09465_, _09464_, _07535_);
  or _60163_ (_09466_, _09465_, _07878_);
  and _60164_ (_09467_, _09466_, _07877_);
  not _60165_ (_09468_, \oc8051_golden_model_1.PC [15]);
  and _60166_ (_09469_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and _60167_ (_09470_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and _60168_ (_09471_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and _60169_ (_09472_, _09471_, _09470_);
  and _60170_ (_09473_, _09472_, _09412_);
  and _60171_ (_09474_, _09473_, _09469_);
  and _60172_ (_09475_, _09474_, \oc8051_golden_model_1.PC [14]);
  and _60173_ (_09476_, _09475_, _09468_);
  nor _60174_ (_09477_, _09475_, _09468_);
  or _60175_ (_09478_, _09477_, _09476_);
  not _60176_ (_09479_, _09478_);
  nand _60177_ (_09480_, _09479_, _06361_);
  and _60178_ (_09481_, _09472_, _08659_);
  and _60179_ (_09482_, _09481_, _09469_);
  and _60180_ (_09483_, _09482_, \oc8051_golden_model_1.PC [14]);
  and _60181_ (_09485_, _09483_, _09468_);
  nor _60182_ (_09486_, _09483_, _09468_);
  or _60183_ (_09487_, _09486_, _09485_);
  or _60184_ (_09488_, _09487_, _06361_);
  and _60185_ (_09489_, _09488_, _09480_);
  and _60186_ (_09490_, _09489_, _07872_);
  and _60187_ (_09491_, _09490_, _07875_);
  or _60188_ (_40572_, _09491_, _09467_);
  not _60189_ (_09492_, \oc8051_golden_model_1.B [7]);
  nor _60190_ (_09493_, _01347_, _09492_);
  nor _60191_ (_09494_, _07942_, _09492_);
  and _60192_ (_09495_, _08575_, _07942_);
  or _60193_ (_09496_, _09495_, _09494_);
  and _60194_ (_09497_, _09496_, _06536_);
  not _60195_ (_09498_, _07942_);
  nor _60196_ (_09499_, _08040_, _09498_);
  or _60197_ (_09500_, _09499_, _09494_);
  or _60198_ (_09501_, _09500_, _07215_);
  nor _60199_ (_09502_, _08634_, _09492_);
  and _60200_ (_09503_, _08649_, _08634_);
  or _60201_ (_09505_, _09503_, _09502_);
  and _60202_ (_09506_, _09505_, _06268_);
  and _60203_ (_09507_, _08768_, _07942_);
  or _60204_ (_09508_, _09507_, _09494_);
  or _60205_ (_09509_, _09508_, _07151_);
  and _60206_ (_09510_, _07942_, \oc8051_golden_model_1.ACC [7]);
  or _60207_ (_09511_, _09510_, _09494_);
  and _60208_ (_09512_, _09511_, _07141_);
  nor _60209_ (_09513_, _07141_, _09492_);
  or _60210_ (_09514_, _09513_, _06341_);
  or _60211_ (_09515_, _09514_, _09512_);
  and _60212_ (_09516_, _09515_, _06273_);
  and _60213_ (_09517_, _09516_, _09509_);
  and _60214_ (_09518_, _08773_, _08634_);
  or _60215_ (_09519_, _09518_, _09502_);
  and _60216_ (_09520_, _09519_, _06272_);
  or _60217_ (_09521_, _09520_, _06461_);
  or _60218_ (_09522_, _09521_, _09517_);
  or _60219_ (_09523_, _09500_, _07166_);
  and _60220_ (_09524_, _09523_, _09522_);
  or _60221_ (_09525_, _09524_, _06464_);
  or _60222_ (_09526_, _09511_, _06465_);
  and _60223_ (_09527_, _09526_, _06269_);
  and _60224_ (_09528_, _09527_, _09525_);
  or _60225_ (_09529_, _09528_, _09506_);
  and _60226_ (_09530_, _09529_, _06262_);
  and _60227_ (_09531_, _06370_, _06491_);
  or _60228_ (_09532_, _09502_, _08789_);
  and _60229_ (_09533_, _09532_, _06261_);
  and _60230_ (_09534_, _09533_, _09519_);
  or _60231_ (_09535_, _09534_, _09531_);
  or _60232_ (_09536_, _09535_, _09530_);
  not _60233_ (_09537_, _09531_);
  and _60234_ (_09538_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and _60235_ (_09539_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and _60236_ (_09540_, _09539_, _09538_);
  and _60237_ (_09541_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and _60238_ (_09542_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor _60239_ (_09543_, _09542_, _09541_);
  nor _60240_ (_09544_, _09543_, _09540_);
  and _60241_ (_09545_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and _60242_ (_09546_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and _60243_ (_09547_, _09546_, _09545_);
  and _60244_ (_09548_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and _60245_ (_09549_, _09548_, _09539_);
  and _60246_ (_09550_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  nor _60247_ (_09551_, _09548_, _09539_);
  nor _60248_ (_09552_, _09551_, _09549_);
  and _60249_ (_09553_, _09552_, _09550_);
  nor _60250_ (_09554_, _09553_, _09549_);
  and _60251_ (_09555_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and _60252_ (_09556_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and _60253_ (_09557_, _09556_, _09555_);
  nor _60254_ (_09558_, _09556_, _09555_);
  nor _60255_ (_09559_, _09558_, _09557_);
  not _60256_ (_09560_, _09559_);
  nor _60257_ (_09561_, _09560_, _09554_);
  and _60258_ (_09562_, _09560_, _09554_);
  nor _60259_ (_09563_, _09562_, _09561_);
  and _60260_ (_09564_, _09563_, _09547_);
  nor _60261_ (_09565_, _09563_, _09547_);
  nor _60262_ (_09566_, _09565_, _09564_);
  and _60263_ (_09567_, _09566_, _09544_);
  and _60264_ (_09568_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and _60265_ (_09569_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and _60266_ (_09570_, _09569_, _09568_);
  nor _60267_ (_09571_, _09569_, _09568_);
  nor _60268_ (_09572_, _09571_, _09570_);
  and _60269_ (_09573_, _09572_, _09540_);
  nor _60270_ (_09574_, _09572_, _09540_);
  nor _60271_ (_09575_, _09574_, _09573_);
  and _60272_ (_09576_, _09575_, _09557_);
  nor _60273_ (_09577_, _09575_, _09557_);
  nor _60274_ (_09578_, _09577_, _09576_);
  and _60275_ (_09579_, _09578_, _09538_);
  nor _60276_ (_09580_, _09578_, _09538_);
  nor _60277_ (_09581_, _09580_, _09579_);
  and _60278_ (_09582_, _09581_, _09567_);
  nor _60279_ (_09583_, _09564_, _09561_);
  not _60280_ (_09584_, _09583_);
  nor _60281_ (_09585_, _09581_, _09567_);
  nor _60282_ (_09586_, _09585_, _09582_);
  and _60283_ (_09587_, _09586_, _09584_);
  nor _60284_ (_09588_, _09587_, _09582_);
  nor _60285_ (_09589_, _09576_, _09573_);
  not _60286_ (_09590_, _09589_);
  and _60287_ (_09591_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and _60288_ (_09592_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and _60289_ (_09593_, _09592_, _09591_);
  nor _60290_ (_09594_, _09592_, _09591_);
  nor _60291_ (_09595_, _09594_, _09593_);
  and _60292_ (_09596_, _09595_, _09570_);
  nor _60293_ (_09597_, _09595_, _09570_);
  nor _60294_ (_09598_, _09597_, _09596_);
  and _60295_ (_09599_, _09598_, _09579_);
  nor _60296_ (_09600_, _09598_, _09579_);
  nor _60297_ (_09601_, _09600_, _09599_);
  and _60298_ (_09602_, _09601_, _09590_);
  nor _60299_ (_09603_, _09601_, _09590_);
  nor _60300_ (_09604_, _09603_, _09602_);
  not _60301_ (_09605_, _09604_);
  nor _60302_ (_09606_, _09605_, _09588_);
  and _60303_ (_09607_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not _60304_ (_09608_, _09607_);
  nor _60305_ (_09609_, _09608_, _09569_);
  nor _60306_ (_09610_, _09609_, _09596_);
  nor _60307_ (_09611_, _09602_, _09599_);
  nor _60308_ (_09612_, _09611_, _09610_);
  and _60309_ (_09613_, _09611_, _09610_);
  nor _60310_ (_09614_, _09613_, _09612_);
  and _60311_ (_09615_, _09614_, _09606_);
  or _60312_ (_09616_, _09612_, _09593_);
  or _60313_ (_09617_, _09616_, _09615_);
  and _60314_ (_09618_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and _60315_ (_09619_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and _60316_ (_09620_, _09619_, _09618_);
  not _60317_ (_09621_, _09618_);
  and _60318_ (_09622_, _09619_, _09621_);
  and _60319_ (_09623_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and _60320_ (_09624_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and _60321_ (_09625_, _09624_, _09539_);
  and _60322_ (_09626_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  and _60323_ (_09627_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  nor _60324_ (_09628_, _09627_, _09626_);
  nor _60325_ (_09629_, _09628_, _09625_);
  and _60326_ (_09630_, _09629_, _09623_);
  nor _60327_ (_09631_, _09629_, _09623_);
  nor _60328_ (_09632_, _09631_, _09630_);
  and _60329_ (_09633_, _09632_, _09622_);
  nor _60330_ (_09634_, _09633_, _09620_);
  nor _60331_ (_09635_, _09552_, _09550_);
  nor _60332_ (_09636_, _09635_, _09553_);
  not _60333_ (_09637_, _09636_);
  nor _60334_ (_09638_, _09637_, _09634_);
  and _60335_ (_09639_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and _60336_ (_09640_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and _60337_ (_09641_, _09640_, _09639_);
  nor _60338_ (_09642_, _09630_, _09625_);
  nor _60339_ (_09643_, _09546_, _09545_);
  nor _60340_ (_09644_, _09643_, _09547_);
  not _60341_ (_09645_, _09644_);
  nor _60342_ (_09646_, _09645_, _09642_);
  and _60343_ (_09647_, _09645_, _09642_);
  nor _60344_ (_09648_, _09647_, _09646_);
  and _60345_ (_09649_, _09648_, _09641_);
  nor _60346_ (_09650_, _09648_, _09641_);
  nor _60347_ (_09651_, _09650_, _09649_);
  and _60348_ (_09652_, _09637_, _09634_);
  nor _60349_ (_09653_, _09652_, _09638_);
  and _60350_ (_09654_, _09653_, _09651_);
  nor _60351_ (_09655_, _09654_, _09638_);
  not _60352_ (_09656_, _09655_);
  nor _60353_ (_09657_, _09566_, _09544_);
  nor _60354_ (_09658_, _09657_, _09567_);
  and _60355_ (_09660_, _09658_, _09656_);
  nor _60356_ (_09661_, _09649_, _09646_);
  not _60357_ (_09663_, _09661_);
  nor _60358_ (_09664_, _09658_, _09656_);
  nor _60359_ (_09666_, _09664_, _09660_);
  and _60360_ (_09667_, _09666_, _09663_);
  nor _60361_ (_09669_, _09667_, _09660_);
  nor _60362_ (_09670_, _09586_, _09584_);
  nor _60363_ (_09672_, _09670_, _09587_);
  not _60364_ (_09673_, _09672_);
  nor _60365_ (_09675_, _09673_, _09669_);
  and _60366_ (_09676_, _09605_, _09588_);
  nor _60367_ (_09678_, _09676_, _09606_);
  and _60368_ (_09679_, _09678_, _09675_);
  and _60369_ (_09681_, _09679_, _09614_);
  and _60370_ (_09682_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and _60371_ (_09684_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and _60372_ (_09685_, _09684_, _09682_);
  and _60373_ (_09687_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and _60374_ (_09688_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor _60375_ (_09690_, _09688_, _09618_);
  nor _60376_ (_09691_, _09690_, _09685_);
  and _60377_ (_09693_, _09691_, _09687_);
  nor _60378_ (_09694_, _09693_, _09685_);
  and _60379_ (_09696_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor _60380_ (_09697_, _09696_, _09682_);
  nor _60381_ (_09698_, _09697_, _09620_);
  not _60382_ (_09699_, _09698_);
  nor _60383_ (_09700_, _09699_, _09694_);
  and _60384_ (_09701_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and _60385_ (_09702_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and _60386_ (_09703_, _09702_, _09624_);
  nor _60387_ (_09704_, _09702_, _09624_);
  nor _60388_ (_09705_, _09704_, _09703_);
  and _60389_ (_09706_, _09705_, _09701_);
  nor _60390_ (_09707_, _09705_, _09701_);
  nor _60391_ (_09708_, _09707_, _09706_);
  and _60392_ (_09709_, _09699_, _09694_);
  nor _60393_ (_09710_, _09709_, _09700_);
  and _60394_ (_09711_, _09710_, _09708_);
  nor _60395_ (_09712_, _09711_, _09700_);
  nor _60396_ (_09713_, _09632_, _09622_);
  nor _60397_ (_09714_, _09713_, _09633_);
  not _60398_ (_09715_, _09714_);
  nor _60399_ (_09716_, _09715_, _09712_);
  and _60400_ (_09717_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and _60401_ (_09718_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and _60402_ (_09719_, _09718_, _09717_);
  nor _60403_ (_09720_, _09706_, _09703_);
  nor _60404_ (_09721_, _09640_, _09639_);
  nor _60405_ (_09722_, _09721_, _09641_);
  not _60406_ (_09723_, _09722_);
  nor _60407_ (_09724_, _09723_, _09720_);
  and _60408_ (_09725_, _09723_, _09720_);
  nor _60409_ (_09726_, _09725_, _09724_);
  and _60410_ (_09727_, _09726_, _09719_);
  nor _60411_ (_09728_, _09726_, _09719_);
  nor _60412_ (_09729_, _09728_, _09727_);
  and _60413_ (_09730_, _09715_, _09712_);
  nor _60414_ (_09731_, _09730_, _09716_);
  and _60415_ (_09732_, _09731_, _09729_);
  nor _60416_ (_09733_, _09732_, _09716_);
  nor _60417_ (_09734_, _09653_, _09651_);
  nor _60418_ (_09735_, _09734_, _09654_);
  not _60419_ (_09736_, _09735_);
  nor _60420_ (_09737_, _09736_, _09733_);
  nor _60421_ (_09738_, _09727_, _09724_);
  not _60422_ (_09739_, _09738_);
  and _60423_ (_09740_, _09736_, _09733_);
  nor _60424_ (_09741_, _09740_, _09737_);
  and _60425_ (_09742_, _09741_, _09739_);
  nor _60426_ (_09743_, _09742_, _09737_);
  nor _60427_ (_09744_, _09666_, _09663_);
  nor _60428_ (_09745_, _09744_, _09667_);
  not _60429_ (_09746_, _09745_);
  nor _60430_ (_09747_, _09746_, _09743_);
  and _60431_ (_09748_, _09673_, _09669_);
  nor _60432_ (_09749_, _09748_, _09675_);
  and _60433_ (_09750_, _09749_, _09747_);
  nor _60434_ (_09751_, _09678_, _09675_);
  nor _60435_ (_09752_, _09751_, _09679_);
  and _60436_ (_09753_, _09752_, _09750_);
  nor _60437_ (_09755_, _09752_, _09750_);
  nor _60438_ (_09757_, _09755_, _09753_);
  and _60439_ (_09758_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and _60440_ (_09760_, _09758_, _09618_);
  and _60441_ (_09761_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and _60442_ (_09763_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor _60443_ (_09764_, _09763_, _09684_);
  nor _60444_ (_09766_, _09764_, _09760_);
  and _60445_ (_09767_, _09766_, _09761_);
  nor _60446_ (_09769_, _09767_, _09760_);
  not _60447_ (_09770_, _09769_);
  nor _60448_ (_09772_, _09691_, _09687_);
  nor _60449_ (_09773_, _09772_, _09693_);
  and _60450_ (_09775_, _09773_, _09770_);
  and _60451_ (_09776_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and _60452_ (_09778_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and _60453_ (_09779_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and _60454_ (_09781_, _09779_, _09778_);
  nor _60455_ (_09782_, _09779_, _09778_);
  nor _60456_ (_09784_, _09782_, _09781_);
  and _60457_ (_09785_, _09784_, _09776_);
  nor _60458_ (_09787_, _09784_, _09776_);
  nor _60459_ (_09788_, _09787_, _09785_);
  nor _60460_ (_09790_, _09773_, _09770_);
  nor _60461_ (_09791_, _09790_, _09775_);
  and _60462_ (_09792_, _09791_, _09788_);
  nor _60463_ (_09793_, _09792_, _09775_);
  nor _60464_ (_09794_, _09710_, _09708_);
  nor _60465_ (_09795_, _09794_, _09711_);
  not _60466_ (_09796_, _09795_);
  nor _60467_ (_09797_, _09796_, _09793_);
  and _60468_ (_09798_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and _60469_ (_09799_, _09798_, _09718_);
  nor _60470_ (_09800_, _09785_, _09781_);
  nor _60471_ (_09801_, _09718_, _09717_);
  nor _60472_ (_09802_, _09801_, _09719_);
  not _60473_ (_09803_, _09802_);
  nor _60474_ (_09804_, _09803_, _09800_);
  and _60475_ (_09805_, _09803_, _09800_);
  nor _60476_ (_09806_, _09805_, _09804_);
  and _60477_ (_09807_, _09806_, _09799_);
  nor _60478_ (_09808_, _09806_, _09799_);
  nor _60479_ (_09809_, _09808_, _09807_);
  and _60480_ (_09810_, _09796_, _09793_);
  nor _60481_ (_09811_, _09810_, _09797_);
  and _60482_ (_09812_, _09811_, _09809_);
  nor _60483_ (_09813_, _09812_, _09797_);
  nor _60484_ (_09814_, _09731_, _09729_);
  nor _60485_ (_09815_, _09814_, _09732_);
  not _60486_ (_09816_, _09815_);
  nor _60487_ (_09817_, _09816_, _09813_);
  nor _60488_ (_09818_, _09807_, _09804_);
  not _60489_ (_09819_, _09818_);
  and _60490_ (_09820_, _09816_, _09813_);
  nor _60491_ (_09821_, _09820_, _09817_);
  and _60492_ (_09822_, _09821_, _09819_);
  nor _60493_ (_09823_, _09822_, _09817_);
  nor _60494_ (_09824_, _09741_, _09739_);
  nor _60495_ (_09825_, _09824_, _09742_);
  not _60496_ (_09826_, _09825_);
  nor _60497_ (_09827_, _09826_, _09823_);
  and _60498_ (_09828_, _09746_, _09743_);
  nor _60499_ (_09829_, _09828_, _09747_);
  and _60500_ (_09830_, _09829_, _09827_);
  nor _60501_ (_09831_, _09749_, _09747_);
  nor _60502_ (_09832_, _09831_, _09750_);
  nand _60503_ (_09833_, _09832_, _09830_);
  and _60504_ (_09834_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and _60505_ (_09835_, _09834_, _09758_);
  and _60506_ (_09836_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor _60507_ (_09837_, _09834_, _09758_);
  nor _60508_ (_09838_, _09837_, _09835_);
  and _60509_ (_09839_, _09838_, _09836_);
  nor _60510_ (_09840_, _09839_, _09835_);
  not _60511_ (_09841_, _09840_);
  nor _60512_ (_09842_, _09766_, _09761_);
  nor _60513_ (_09843_, _09842_, _09767_);
  and _60514_ (_09844_, _09843_, _09841_);
  and _60515_ (_09845_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and _60516_ (_09846_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and _60517_ (_09847_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and _60518_ (_09848_, _09847_, _09846_);
  nor _60519_ (_09849_, _09847_, _09846_);
  nor _60520_ (_09850_, _09849_, _09848_);
  and _60521_ (_09851_, _09850_, _09845_);
  nor _60522_ (_09852_, _09850_, _09845_);
  nor _60523_ (_09853_, _09852_, _09851_);
  nor _60524_ (_09854_, _09843_, _09841_);
  nor _60525_ (_09855_, _09854_, _09844_);
  and _60526_ (_09856_, _09855_, _09853_);
  nor _60527_ (_09857_, _09856_, _09844_);
  not _60528_ (_09858_, _09857_);
  nor _60529_ (_09859_, _09791_, _09788_);
  nor _60530_ (_09860_, _09859_, _09792_);
  and _60531_ (_09861_, _09860_, _09858_);
  nor _60532_ (_09862_, _09851_, _09848_);
  and _60533_ (_09863_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and _60534_ (_09864_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor _60535_ (_09865_, _09864_, _09863_);
  nor _60536_ (_09866_, _09865_, _09799_);
  not _60537_ (_09867_, _09866_);
  nor _60538_ (_09868_, _09867_, _09862_);
  and _60539_ (_09869_, _09867_, _09862_);
  nor _60540_ (_09870_, _09869_, _09868_);
  nor _60541_ (_09871_, _09860_, _09858_);
  nor _60542_ (_09872_, _09871_, _09861_);
  and _60543_ (_09873_, _09872_, _09870_);
  nor _60544_ (_09874_, _09873_, _09861_);
  nor _60545_ (_09875_, _09811_, _09809_);
  nor _60546_ (_09876_, _09875_, _09812_);
  not _60547_ (_09877_, _09876_);
  nor _60548_ (_09878_, _09877_, _09874_);
  and _60549_ (_09879_, _09877_, _09874_);
  nor _60550_ (_09880_, _09879_, _09878_);
  and _60551_ (_09881_, _09880_, _09868_);
  nor _60552_ (_09882_, _09881_, _09878_);
  nor _60553_ (_09883_, _09821_, _09819_);
  nor _60554_ (_09884_, _09883_, _09822_);
  not _60555_ (_09885_, _09884_);
  nor _60556_ (_09886_, _09885_, _09882_);
  and _60557_ (_09887_, _09826_, _09823_);
  nor _60558_ (_09888_, _09887_, _09827_);
  and _60559_ (_09889_, _09888_, _09886_);
  nor _60560_ (_09890_, _09829_, _09827_);
  nor _60561_ (_09891_, _09890_, _09830_);
  and _60562_ (_09892_, _09891_, _09889_);
  nor _60563_ (_09893_, _09891_, _09889_);
  nor _60564_ (_09894_, _09893_, _09892_);
  and _60565_ (_09895_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and _60566_ (_09896_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and _60567_ (_09897_, _09896_, _09895_);
  and _60568_ (_09898_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor _60569_ (_09899_, _09896_, _09895_);
  nor _60570_ (_09900_, _09899_, _09897_);
  and _60571_ (_09901_, _09900_, _09898_);
  nor _60572_ (_09902_, _09901_, _09897_);
  not _60573_ (_09903_, _09902_);
  nor _60574_ (_09904_, _09838_, _09836_);
  nor _60575_ (_09905_, _09904_, _09839_);
  and _60576_ (_09906_, _09905_, _09903_);
  and _60577_ (_09907_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and _60578_ (_09908_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and _60579_ (_09909_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and _60580_ (_09910_, _09909_, _09908_);
  nor _60581_ (_09911_, _09909_, _09908_);
  nor _60582_ (_09912_, _09911_, _09910_);
  and _60583_ (_09913_, _09912_, _09907_);
  nor _60584_ (_09914_, _09912_, _09907_);
  nor _60585_ (_09915_, _09914_, _09913_);
  nor _60586_ (_09916_, _09905_, _09903_);
  nor _60587_ (_09917_, _09916_, _09906_);
  and _60588_ (_09918_, _09917_, _09915_);
  nor _60589_ (_09919_, _09918_, _09906_);
  not _60590_ (_09920_, _09919_);
  nor _60591_ (_09921_, _09855_, _09853_);
  nor _60592_ (_09922_, _09921_, _09856_);
  and _60593_ (_09923_, _09922_, _09920_);
  not _60594_ (_09924_, _09798_);
  nor _60595_ (_09925_, _09913_, _09910_);
  nor _60596_ (_09926_, _09925_, _09924_);
  and _60597_ (_09927_, _09925_, _09924_);
  nor _60598_ (_09928_, _09927_, _09926_);
  nor _60599_ (_09929_, _09922_, _09920_);
  nor _60600_ (_09930_, _09929_, _09923_);
  and _60601_ (_09931_, _09930_, _09928_);
  nor _60602_ (_09932_, _09931_, _09923_);
  not _60603_ (_09933_, _09932_);
  nor _60604_ (_09934_, _09872_, _09870_);
  nor _60605_ (_09935_, _09934_, _09873_);
  and _60606_ (_09936_, _09935_, _09933_);
  nor _60607_ (_09937_, _09935_, _09933_);
  nor _60608_ (_09938_, _09937_, _09936_);
  and _60609_ (_09939_, _09938_, _09926_);
  nor _60610_ (_09940_, _09939_, _09936_);
  nor _60611_ (_09941_, _09880_, _09868_);
  nor _60612_ (_09942_, _09941_, _09881_);
  not _60613_ (_09943_, _09942_);
  nor _60614_ (_09944_, _09943_, _09940_);
  and _60615_ (_09945_, _09885_, _09882_);
  nor _60616_ (_09946_, _09945_, _09886_);
  and _60617_ (_09947_, _09946_, _09944_);
  nor _60618_ (_09948_, _09888_, _09886_);
  nor _60619_ (_09949_, _09948_, _09889_);
  nand _60620_ (_09950_, _09949_, _09947_);
  or _60621_ (_09951_, _09949_, _09947_);
  and _60622_ (_09952_, _09951_, _09950_);
  and _60623_ (_09953_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and _60624_ (_09954_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and _60625_ (_09955_, _09954_, _09953_);
  and _60626_ (_09956_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor _60627_ (_09957_, _09954_, _09953_);
  nor _60628_ (_09958_, _09957_, _09955_);
  and _60629_ (_09959_, _09958_, _09956_);
  nor _60630_ (_09960_, _09959_, _09955_);
  not _60631_ (_09961_, _09960_);
  nor _60632_ (_09962_, _09900_, _09898_);
  nor _60633_ (_09963_, _09962_, _09901_);
  and _60634_ (_09964_, _09963_, _09961_);
  and _60635_ (_09965_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and _60636_ (_09966_, _09965_, _09909_);
  and _60637_ (_09967_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and _60638_ (_09968_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor _60639_ (_09969_, _09968_, _09967_);
  nor _60640_ (_09970_, _09969_, _09966_);
  nor _60641_ (_09971_, _09963_, _09961_);
  nor _60642_ (_09972_, _09971_, _09964_);
  and _60643_ (_09973_, _09972_, _09970_);
  nor _60644_ (_09974_, _09973_, _09964_);
  not _60645_ (_09975_, _09974_);
  nor _60646_ (_09976_, _09917_, _09915_);
  nor _60647_ (_09977_, _09976_, _09918_);
  and _60648_ (_09978_, _09977_, _09975_);
  nor _60649_ (_09979_, _09977_, _09975_);
  nor _60650_ (_09980_, _09979_, _09978_);
  and _60651_ (_09981_, _09980_, _09966_);
  nor _60652_ (_09982_, _09981_, _09978_);
  not _60653_ (_09983_, _09982_);
  nor _60654_ (_09984_, _09930_, _09928_);
  nor _60655_ (_09985_, _09984_, _09931_);
  and _60656_ (_09986_, _09985_, _09983_);
  nor _60657_ (_09987_, _09938_, _09926_);
  nor _60658_ (_09988_, _09987_, _09939_);
  and _60659_ (_09989_, _09988_, _09986_);
  and _60660_ (_09990_, _09943_, _09940_);
  nor _60661_ (_09991_, _09990_, _09944_);
  and _60662_ (_09992_, _09991_, _09989_);
  nor _60663_ (_09993_, _09946_, _09944_);
  nor _60664_ (_09994_, _09993_, _09947_);
  and _60665_ (_09995_, _09994_, _09992_);
  nor _60666_ (_09996_, _09994_, _09992_);
  nor _60667_ (_09997_, _09996_, _09995_);
  and _60668_ (_09998_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and _60669_ (_09999_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and _60670_ (_10000_, _09999_, _09998_);
  and _60671_ (_10001_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor _60672_ (_10002_, _09999_, _09998_);
  nor _60673_ (_10003_, _10002_, _10000_);
  and _60674_ (_10004_, _10003_, _10001_);
  nor _60675_ (_10005_, _10004_, _10000_);
  not _60676_ (_10006_, _10005_);
  nor _60677_ (_10007_, _09958_, _09956_);
  nor _60678_ (_10008_, _10007_, _09959_);
  and _60679_ (_10009_, _10008_, _10006_);
  nor _60680_ (_10010_, _10008_, _10006_);
  nor _60681_ (_10011_, _10010_, _10009_);
  and _60682_ (_10012_, _10011_, _09965_);
  nor _60683_ (_10013_, _10012_, _10009_);
  not _60684_ (_10014_, _10013_);
  nor _60685_ (_10015_, _09972_, _09970_);
  nor _60686_ (_10016_, _10015_, _09973_);
  and _60687_ (_10017_, _10016_, _10014_);
  nor _60688_ (_10018_, _09980_, _09966_);
  nor _60689_ (_10019_, _10018_, _09981_);
  and _60690_ (_10020_, _10019_, _10017_);
  nor _60691_ (_10021_, _09985_, _09983_);
  nor _60692_ (_10022_, _10021_, _09986_);
  and _60693_ (_10023_, _10022_, _10020_);
  nor _60694_ (_10024_, _09988_, _09986_);
  nor _60695_ (_10025_, _10024_, _09989_);
  and _60696_ (_10026_, _10025_, _10023_);
  nor _60697_ (_10027_, _09991_, _09989_);
  nor _60698_ (_10028_, _10027_, _09992_);
  and _60699_ (_10029_, _10028_, _10026_);
  and _60700_ (_10030_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and _60701_ (_10031_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and _60702_ (_10032_, _10031_, _10030_);
  nor _60703_ (_10033_, _10003_, _10001_);
  nor _60704_ (_10034_, _10033_, _10004_);
  and _60705_ (_10035_, _10034_, _10032_);
  nor _60706_ (_10036_, _10011_, _09965_);
  nor _60707_ (_10037_, _10036_, _10012_);
  and _60708_ (_10038_, _10037_, _10035_);
  nor _60709_ (_10039_, _10016_, _10014_);
  nor _60710_ (_10040_, _10039_, _10017_);
  and _60711_ (_10041_, _10040_, _10038_);
  nor _60712_ (_10042_, _10019_, _10017_);
  nor _60713_ (_10043_, _10042_, _10020_);
  and _60714_ (_10044_, _10043_, _10041_);
  nor _60715_ (_10045_, _10022_, _10020_);
  nor _60716_ (_10046_, _10045_, _10023_);
  and _60717_ (_10047_, _10046_, _10044_);
  nor _60718_ (_10048_, _10025_, _10023_);
  nor _60719_ (_10049_, _10048_, _10026_);
  and _60720_ (_10050_, _10049_, _10047_);
  nor _60721_ (_10051_, _10028_, _10026_);
  nor _60722_ (_10052_, _10051_, _10029_);
  and _60723_ (_10053_, _10052_, _10050_);
  nor _60724_ (_10054_, _10053_, _10029_);
  not _60725_ (_10055_, _10054_);
  and _60726_ (_10056_, _10055_, _09997_);
  or _60727_ (_10057_, _10056_, _09995_);
  nand _60728_ (_10058_, _10057_, _09952_);
  and _60729_ (_10059_, _10058_, _09950_);
  not _60730_ (_10060_, _10059_);
  and _60731_ (_10061_, _10060_, _09894_);
  or _60732_ (_10062_, _10061_, _09892_);
  or _60733_ (_10063_, _09832_, _09830_);
  and _60734_ (_10064_, _10063_, _09833_);
  nand _60735_ (_10065_, _10064_, _10062_);
  and _60736_ (_10066_, _10065_, _09833_);
  not _60737_ (_10067_, _10066_);
  and _60738_ (_10068_, _10067_, _09757_);
  or _60739_ (_10069_, _10068_, _09753_);
  nor _60740_ (_10070_, _09679_, _09606_);
  and _60741_ (_10071_, _10070_, _09614_);
  nor _60742_ (_10072_, _10070_, _09614_);
  or _60743_ (_10073_, _10072_, _10071_);
  and _60744_ (_10074_, _10073_, _10069_);
  or _60745_ (_10075_, _10074_, _09681_);
  or _60746_ (_10076_, _10075_, _09617_);
  or _60747_ (_10077_, _10076_, _09537_);
  and _60748_ (_10078_, _10077_, _06258_);
  and _60749_ (_10079_, _10078_, _09536_);
  not _60750_ (_10080_, _07215_);
  and _60751_ (_10081_, _08808_, _08634_);
  or _60752_ (_10082_, _10081_, _09502_);
  and _60753_ (_10083_, _10082_, _06257_);
  or _60754_ (_10084_, _10083_, _10080_);
  or _60755_ (_10085_, _10084_, _10079_);
  and _60756_ (_10086_, _10085_, _09501_);
  or _60757_ (_10087_, _10086_, _07460_);
  and _60758_ (_10088_, _08755_, _07942_);
  or _60759_ (_10089_, _09494_, _07208_);
  or _60760_ (_10090_, _10089_, _10088_);
  and _60761_ (_10091_, _10090_, _05982_);
  and _60762_ (_10092_, _10091_, _10087_);
  and _60763_ (_10093_, _06370_, _05944_);
  not _60764_ (_10094_, _05982_);
  and _60765_ (_10095_, _09021_, _07942_);
  or _60766_ (_10096_, _10095_, _09494_);
  and _60767_ (_10097_, _10096_, _10094_);
  or _60768_ (_10098_, _10097_, _10093_);
  or _60769_ (_10099_, _10098_, _10092_);
  not _60770_ (_10100_, _10093_);
  not _60771_ (_10101_, \oc8051_golden_model_1.B [1]);
  nor _60772_ (_10102_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor _60773_ (_10103_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and _60774_ (_10104_, _10103_, _10102_);
  and _60775_ (_10105_, _10104_, _10101_);
  not _60776_ (_10106_, \oc8051_golden_model_1.B [0]);
  and _60777_ (_10107_, _10106_, \oc8051_golden_model_1.ACC [7]);
  nor _60778_ (_10108_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and _60779_ (_10109_, _10108_, _10107_);
  and _60780_ (_10110_, _10109_, _10105_);
  and _60781_ (_10111_, \oc8051_golden_model_1.B [0], _08572_);
  not _60782_ (_10112_, _10111_);
  and _60783_ (_10113_, _10108_, _10105_);
  and _60784_ (_10114_, _10113_, _10112_);
  or _60785_ (_10115_, _10114_, _08572_);
  not _60786_ (_10116_, \oc8051_golden_model_1.ACC [6]);
  and _60787_ (_10117_, \oc8051_golden_model_1.B [0], _10116_);
  nor _60788_ (_10118_, _10117_, _08572_);
  nor _60789_ (_10119_, _10118_, _10101_);
  not _60790_ (_10120_, _10119_);
  and _60791_ (_10121_, _10108_, _10104_);
  and _60792_ (_10122_, _10121_, _10120_);
  nor _60793_ (_10123_, _10122_, _10115_);
  nor _60794_ (_10124_, _10123_, _10110_);
  and _60795_ (_10125_, _10122_, \oc8051_golden_model_1.B [0]);
  nor _60796_ (_10126_, _10125_, _10116_);
  and _60797_ (_10127_, _10126_, _10101_);
  nor _60798_ (_10128_, _10126_, _10101_);
  nor _60799_ (_10129_, _10128_, _10127_);
  nor _60800_ (_10130_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor _60801_ (_10131_, _10130_, _09758_);
  nor _60802_ (_10132_, _10131_, \oc8051_golden_model_1.ACC [4]);
  and _60803_ (_10133_, \oc8051_golden_model_1.ACC [4], _10106_);
  nor _60804_ (_10134_, _10133_, \oc8051_golden_model_1.ACC [5]);
  not _60805_ (_10135_, \oc8051_golden_model_1.ACC [4]);
  and _60806_ (_10136_, _10135_, \oc8051_golden_model_1.B [0]);
  nor _60807_ (_10137_, _10136_, _10134_);
  nor _60808_ (_10138_, _10137_, _10132_);
  not _60809_ (_10139_, _10138_);
  and _60810_ (_10140_, _10139_, _10129_);
  nor _60811_ (_10141_, _10124_, \oc8051_golden_model_1.B [2]);
  nor _60812_ (_10142_, _10141_, _10127_);
  not _60813_ (_10143_, _10142_);
  nor _60814_ (_10144_, _10143_, _10140_);
  not _60815_ (_10145_, \oc8051_golden_model_1.B [3]);
  nor _60816_ (_10146_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and _60817_ (_10147_, _10146_, _10102_);
  and _60818_ (_10148_, _10147_, _10145_);
  and _60819_ (_10149_, \oc8051_golden_model_1.B [2], _08572_);
  not _60820_ (_10150_, _10149_);
  and _60821_ (_10151_, _10150_, _10148_);
  not _60822_ (_10152_, _10151_);
  nor _60823_ (_10153_, _10152_, _10144_);
  nor _60824_ (_10154_, _10153_, _10124_);
  nor _60825_ (_10155_, _10154_, _10110_);
  and _60826_ (_10156_, _10147_, \oc8051_golden_model_1.ACC [7]);
  nor _60827_ (_10157_, _10156_, _10148_);
  nor _60828_ (_10158_, _10155_, \oc8051_golden_model_1.B [3]);
  not _60829_ (_10159_, \oc8051_golden_model_1.B [2]);
  nor _60830_ (_10160_, _10139_, _10129_);
  nor _60831_ (_10161_, _10160_, _10140_);
  not _60832_ (_10162_, _10161_);
  and _60833_ (_10163_, _10162_, _10153_);
  nor _60834_ (_10164_, _10153_, _10126_);
  nor _60835_ (_10165_, _10164_, _10163_);
  and _60836_ (_10166_, _10165_, _10159_);
  nor _60837_ (_10167_, _10165_, _10159_);
  nor _60838_ (_10168_, _10167_, _10166_);
  not _60839_ (_10169_, _10168_);
  not _60840_ (_10170_, \oc8051_golden_model_1.ACC [5]);
  nor _60841_ (_10171_, _10153_, _10170_);
  and _60842_ (_10172_, _10153_, _10131_);
  or _60843_ (_10173_, _10172_, _10171_);
  and _60844_ (_10174_, _10173_, _10101_);
  nor _60845_ (_10175_, _10173_, _10101_);
  nor _60846_ (_10176_, _10175_, _10136_);
  nor _60847_ (_10177_, _10176_, _10174_);
  nor _60848_ (_10178_, _10177_, _10169_);
  or _60849_ (_10179_, _10178_, _10166_);
  nor _60850_ (_10180_, _10179_, _10158_);
  nor _60851_ (_10181_, _10180_, _10157_);
  nor _60852_ (_10182_, _10181_, _10155_);
  nor _60853_ (_10183_, _10182_, _10110_);
  not _60854_ (_10184_, _10181_);
  and _60855_ (_10185_, _10177_, _10169_);
  nor _60856_ (_10186_, _10185_, _10178_);
  nor _60857_ (_10187_, _10186_, _10184_);
  nor _60858_ (_10188_, _10181_, _10165_);
  nor _60859_ (_10189_, _10188_, _10187_);
  and _60860_ (_10190_, _10189_, _10145_);
  nor _60861_ (_10191_, _10189_, _10145_);
  nor _60862_ (_10192_, _10191_, _10190_);
  not _60863_ (_10193_, _10192_);
  nor _60864_ (_10194_, _10181_, _10173_);
  nor _60865_ (_10195_, _10175_, _10174_);
  and _60866_ (_10196_, _10195_, _10136_);
  nor _60867_ (_10197_, _10195_, _10136_);
  nor _60868_ (_10198_, _10197_, _10196_);
  and _60869_ (_10199_, _10198_, _10181_);
  or _60870_ (_10200_, _10199_, _10194_);
  nor _60871_ (_10201_, _10200_, \oc8051_golden_model_1.B [2]);
  and _60872_ (_10202_, _10200_, \oc8051_golden_model_1.B [2]);
  nor _60873_ (_10203_, _10136_, _10133_);
  and _60874_ (_10204_, _10181_, _10203_);
  nor _60875_ (_10205_, _10181_, \oc8051_golden_model_1.ACC [4]);
  nor _60876_ (_10206_, _10205_, _10204_);
  and _60877_ (_10207_, _10206_, _10101_);
  nor _60878_ (_10208_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor _60879_ (_10209_, _10208_, _09953_);
  nor _60880_ (_10210_, _10209_, \oc8051_golden_model_1.ACC [2]);
  and _60881_ (_10211_, _10106_, \oc8051_golden_model_1.ACC [2]);
  nor _60882_ (_10212_, _10211_, \oc8051_golden_model_1.ACC [3]);
  not _60883_ (_10213_, \oc8051_golden_model_1.ACC [2]);
  and _60884_ (_10214_, \oc8051_golden_model_1.B [0], _10213_);
  nor _60885_ (_10215_, _10214_, _10212_);
  nor _60886_ (_10216_, _10215_, _10210_);
  not _60887_ (_10217_, _10216_);
  nor _60888_ (_10218_, _10206_, _10101_);
  nor _60889_ (_10219_, _10218_, _10207_);
  and _60890_ (_10220_, _10219_, _10217_);
  nor _60891_ (_10221_, _10220_, _10207_);
  nor _60892_ (_10222_, _10221_, _10202_);
  nor _60893_ (_10223_, _10222_, _10201_);
  nor _60894_ (_10224_, _10223_, _10193_);
  nor _60895_ (_10225_, _10183_, \oc8051_golden_model_1.B [4]);
  nor _60896_ (_10226_, _10225_, _10190_);
  not _60897_ (_10227_, _10226_);
  nor _60898_ (_10228_, _10227_, _10224_);
  not _60899_ (_10229_, \oc8051_golden_model_1.B [5]);
  and _60900_ (_10230_, _10146_, _10229_);
  not _60901_ (_10231_, _10230_);
  and _60902_ (_10232_, \oc8051_golden_model_1.B [4], _08572_);
  nor _60903_ (_10233_, _10232_, _10231_);
  not _60904_ (_10234_, _10233_);
  nor _60905_ (_10235_, _10234_, _10228_);
  nor _60906_ (_10236_, _10235_, _10183_);
  nor _60907_ (_10237_, _10236_, _10110_);
  and _60908_ (_10238_, _10146_, \oc8051_golden_model_1.ACC [7]);
  nor _60909_ (_10239_, _10238_, _10230_);
  nor _60910_ (_10240_, _10237_, \oc8051_golden_model_1.B [5]);
  not _60911_ (_10241_, \oc8051_golden_model_1.B [4]);
  and _60912_ (_10242_, _10223_, _10193_);
  nor _60913_ (_10243_, _10242_, _10224_);
  not _60914_ (_10244_, _10243_);
  and _60915_ (_10245_, _10244_, _10235_);
  nor _60916_ (_10246_, _10235_, _10189_);
  nor _60917_ (_10247_, _10246_, _10245_);
  and _60918_ (_10248_, _10247_, _10241_);
  nor _60919_ (_10249_, _10247_, _10241_);
  nor _60920_ (_10250_, _10249_, _10248_);
  not _60921_ (_10251_, _10250_);
  nor _60922_ (_10252_, _10235_, _10200_);
  nor _60923_ (_10253_, _10202_, _10201_);
  and _60924_ (_10254_, _10253_, _10221_);
  nor _60925_ (_10255_, _10253_, _10221_);
  nor _60926_ (_10256_, _10255_, _10254_);
  not _60927_ (_10257_, _10256_);
  and _60928_ (_10258_, _10257_, _10235_);
  nor _60929_ (_10259_, _10258_, _10252_);
  nor _60930_ (_10260_, _10259_, \oc8051_golden_model_1.B [3]);
  and _60931_ (_10261_, _10259_, \oc8051_golden_model_1.B [3]);
  nor _60932_ (_10262_, _10219_, _10217_);
  nor _60933_ (_10263_, _10262_, _10220_);
  not _60934_ (_10264_, _10263_);
  and _60935_ (_10265_, _10264_, _10235_);
  nor _60936_ (_10266_, _10235_, _10206_);
  nor _60937_ (_10267_, _10266_, _10265_);
  and _60938_ (_10268_, _10267_, _10159_);
  nor _60939_ (_10269_, _10235_, _06055_);
  and _60940_ (_10270_, _10235_, _10209_);
  or _60941_ (_10271_, _10270_, _10269_);
  and _60942_ (_10272_, _10271_, _10101_);
  nor _60943_ (_10273_, _10271_, _10101_);
  nor _60944_ (_10274_, _10273_, _10214_);
  nor _60945_ (_10275_, _10274_, _10272_);
  nor _60946_ (_10276_, _10267_, _10159_);
  nor _60947_ (_10277_, _10276_, _10268_);
  not _60948_ (_10278_, _10277_);
  nor _60949_ (_10279_, _10278_, _10275_);
  nor _60950_ (_10280_, _10279_, _10268_);
  nor _60951_ (_10281_, _10280_, _10261_);
  nor _60952_ (_10282_, _10281_, _10260_);
  nor _60953_ (_10283_, _10282_, _10251_);
  or _60954_ (_10284_, _10283_, _10248_);
  nor _60955_ (_10285_, _10284_, _10240_);
  nor _60956_ (_10286_, _10285_, _10239_);
  nor _60957_ (_10287_, _10286_, _10237_);
  not _60958_ (_10288_, _10286_);
  and _60959_ (_10289_, _10282_, _10251_);
  nor _60960_ (_10290_, _10289_, _10283_);
  nor _60961_ (_10291_, _10290_, _10288_);
  nor _60962_ (_10292_, _10286_, _10247_);
  nor _60963_ (_10293_, _10292_, _10291_);
  and _60964_ (_10294_, _10293_, _10229_);
  nor _60965_ (_10295_, _10293_, _10229_);
  nor _60966_ (_10296_, _10295_, _10294_);
  not _60967_ (_10297_, _10296_);
  nor _60968_ (_10298_, _10286_, _10259_);
  nor _60969_ (_10299_, _10261_, _10260_);
  nor _60970_ (_10300_, _10299_, _10280_);
  and _60971_ (_10301_, _10299_, _10280_);
  or _60972_ (_10302_, _10301_, _10300_);
  and _60973_ (_10303_, _10302_, _10286_);
  or _60974_ (_10304_, _10303_, _10298_);
  and _60975_ (_10305_, _10304_, _10241_);
  nor _60976_ (_10306_, _10304_, _10241_);
  and _60977_ (_10307_, _10278_, _10275_);
  nor _60978_ (_10308_, _10307_, _10279_);
  nor _60979_ (_10309_, _10308_, _10288_);
  nor _60980_ (_10310_, _10286_, _10267_);
  nor _60981_ (_10311_, _10310_, _10309_);
  and _60982_ (_10312_, _10311_, _10145_);
  nor _60983_ (_10313_, _10273_, _10272_);
  nor _60984_ (_10314_, _10313_, _10214_);
  and _60985_ (_10315_, _10313_, _10214_);
  or _60986_ (_10316_, _10315_, _10314_);
  nor _60987_ (_10317_, _10316_, _10288_);
  nor _60988_ (_10318_, _10286_, _10271_);
  nor _60989_ (_10319_, _10318_, _10317_);
  and _60990_ (_10320_, _10319_, _10159_);
  nor _60991_ (_10321_, _10319_, _10159_);
  nor _60992_ (_10322_, _10214_, _10211_);
  and _60993_ (_10323_, _10286_, _10322_);
  nor _60994_ (_10324_, _10286_, \oc8051_golden_model_1.ACC [2]);
  nor _60995_ (_10325_, _10324_, _10323_);
  and _60996_ (_10326_, _10325_, _10101_);
  and _60997_ (_10327_, _06042_, \oc8051_golden_model_1.B [0]);
  not _60998_ (_10328_, _10327_);
  nor _60999_ (_10329_, _10325_, _10101_);
  nor _61000_ (_10330_, _10329_, _10326_);
  and _61001_ (_10331_, _10330_, _10328_);
  nor _61002_ (_10332_, _10331_, _10326_);
  nor _61003_ (_10333_, _10332_, _10321_);
  nor _61004_ (_10334_, _10333_, _10320_);
  nor _61005_ (_10335_, _10311_, _10145_);
  nor _61006_ (_10336_, _10335_, _10312_);
  not _61007_ (_10337_, _10336_);
  nor _61008_ (_10338_, _10337_, _10334_);
  nor _61009_ (_10339_, _10338_, _10312_);
  nor _61010_ (_10340_, _10339_, _10306_);
  nor _61011_ (_10341_, _10340_, _10305_);
  nor _61012_ (_10342_, _10341_, _10297_);
  nor _61013_ (_10343_, _10342_, _10294_);
  and _61014_ (_10344_, \oc8051_golden_model_1.ACC [7], _09492_);
  nor _61015_ (_10345_, _10344_, _10146_);
  nor _61016_ (_10346_, _10345_, _10343_);
  not _61017_ (_10347_, _10146_);
  nor _61018_ (_10348_, _10287_, _10110_);
  nor _61019_ (_10349_, _10348_, _10347_);
  nor _61020_ (_10350_, _10349_, _10346_);
  and _61021_ (_10351_, _10350_, _10287_);
  or _61022_ (_10352_, _10351_, _10110_);
  nor _61023_ (_10353_, _10352_, _09492_);
  nor _61024_ (_10354_, _10352_, \oc8051_golden_model_1.B [7]);
  nor _61025_ (_10355_, _10354_, _09607_);
  not _61026_ (_10356_, _10355_);
  not _61027_ (_10357_, \oc8051_golden_model_1.B [6]);
  and _61028_ (_10358_, _10341_, _10297_);
  nor _61029_ (_10359_, _10358_, _10342_);
  nor _61030_ (_10360_, _10359_, _10350_);
  not _61031_ (_10361_, _10350_);
  nor _61032_ (_10362_, _10361_, _10293_);
  nor _61033_ (_10363_, _10362_, _10360_);
  nor _61034_ (_10364_, _10363_, _10357_);
  and _61035_ (_10365_, _10363_, _10357_);
  nor _61036_ (_10366_, _10306_, _10305_);
  nor _61037_ (_10367_, _10366_, _10339_);
  and _61038_ (_10368_, _10366_, _10339_);
  or _61039_ (_10369_, _10368_, _10367_);
  nor _61040_ (_10370_, _10369_, _10350_);
  nor _61041_ (_10371_, _10361_, _10304_);
  nor _61042_ (_10372_, _10371_, _10370_);
  nor _61043_ (_10373_, _10372_, _10229_);
  and _61044_ (_10374_, _10372_, _10229_);
  not _61045_ (_10375_, _10374_);
  and _61046_ (_10376_, _10337_, _10334_);
  nor _61047_ (_10377_, _10376_, _10338_);
  nor _61048_ (_10378_, _10377_, _10350_);
  nor _61049_ (_10379_, _10361_, _10311_);
  nor _61050_ (_10380_, _10379_, _10378_);
  nor _61051_ (_10381_, _10380_, _10241_);
  and _61052_ (_10382_, _10350_, _10319_);
  nor _61053_ (_10383_, _10321_, _10320_);
  and _61054_ (_10384_, _10383_, _10332_);
  nor _61055_ (_10385_, _10383_, _10332_);
  nor _61056_ (_10386_, _10385_, _10384_);
  nor _61057_ (_10387_, _10386_, _10350_);
  or _61058_ (_10388_, _10387_, _10382_);
  and _61059_ (_10389_, _10388_, _10145_);
  nor _61060_ (_10390_, _10388_, _10145_);
  nor _61061_ (_10391_, _10390_, _10389_);
  nor _61062_ (_10392_, _10330_, _10328_);
  nor _61063_ (_10393_, _10392_, _10331_);
  nor _61064_ (_10394_, _10393_, _10350_);
  nor _61065_ (_10395_, _10361_, _10325_);
  nor _61066_ (_10396_, _10395_, _10394_);
  nor _61067_ (_10397_, _10396_, _10159_);
  and _61068_ (_10398_, _10396_, _10159_);
  nor _61069_ (_10399_, _10398_, _10397_);
  and _61070_ (_10400_, _10399_, _10391_);
  and _61071_ (_10401_, _10350_, _06042_);
  nor _61072_ (_10402_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  nor _61073_ (_10403_, _10402_, _10030_);
  nor _61074_ (_10404_, _10350_, _10403_);
  nor _61075_ (_10405_, _10404_, _10401_);
  and _61076_ (_10406_, _10405_, _10101_);
  nor _61077_ (_10407_, _10405_, _10101_);
  and _61078_ (_10408_, _10106_, \oc8051_golden_model_1.ACC [0]);
  not _61079_ (_10409_, _10408_);
  nor _61080_ (_10410_, _10409_, _10407_);
  nor _61081_ (_10411_, _10410_, _10406_);
  and _61082_ (_10412_, _10411_, _10400_);
  and _61083_ (_10413_, _10397_, _10391_);
  nor _61084_ (_10414_, _10413_, _10390_);
  not _61085_ (_10415_, _10414_);
  nor _61086_ (_10416_, _10415_, _10412_);
  and _61087_ (_10417_, _10380_, _10241_);
  nor _61088_ (_10418_, _10417_, _10416_);
  or _61089_ (_10419_, _10418_, _10381_);
  and _61090_ (_10420_, _10419_, _10375_);
  nor _61091_ (_10421_, _10420_, _10373_);
  nor _61092_ (_10422_, _10421_, _10365_);
  or _61093_ (_10423_, _10422_, _10364_);
  and _61094_ (_10424_, _10423_, _10356_);
  nor _61095_ (_10425_, _10424_, _10353_);
  nor _61096_ (_10426_, _10417_, _10381_);
  nor _61097_ (_10427_, _10374_, _10373_);
  and _61098_ (_10428_, _10427_, _10426_);
  nor _61099_ (_10429_, _10365_, _10364_);
  and _61100_ (_10430_, _10429_, _10356_);
  and _61101_ (_10431_, _10430_, _10428_);
  nor _61102_ (_10432_, _10407_, _10406_);
  and _61103_ (_10433_, \oc8051_golden_model_1.B [0], _06097_);
  not _61104_ (_10434_, _10433_);
  and _61105_ (_10435_, _10434_, _10432_);
  and _61106_ (_10436_, _10435_, _10409_);
  and _61107_ (_10437_, _10436_, _10400_);
  and _61108_ (_10438_, _10437_, _10431_);
  nor _61109_ (_10439_, _10438_, _10425_);
  or _61110_ (_10440_, _10439_, _10110_);
  and _61111_ (_10441_, _10440_, _10352_);
  or _61112_ (_10442_, _10441_, _10100_);
  and _61113_ (_10443_, _10442_, _10099_);
  and _61114_ (_10444_, _10443_, _06219_);
  and _61115_ (_10445_, _08825_, _07942_);
  or _61116_ (_10446_, _10445_, _09494_);
  and _61117_ (_10447_, _10446_, _06218_);
  or _61118_ (_10448_, _10447_, _06369_);
  or _61119_ (_10449_, _10448_, _10444_);
  and _61120_ (_10450_, _09044_, _07942_);
  or _61121_ (_10451_, _10450_, _09494_);
  or _61122_ (_10452_, _10451_, _07237_);
  and _61123_ (_10453_, _10452_, _07240_);
  and _61124_ (_10454_, _10453_, _10449_);
  or _61125_ (_10455_, _10454_, _09497_);
  and _61126_ (_10456_, _10455_, _07242_);
  or _61127_ (_10457_, _09494_, _08043_);
  and _61128_ (_10458_, _10446_, _06375_);
  and _61129_ (_10459_, _10458_, _10457_);
  or _61130_ (_10460_, _10459_, _10456_);
  and _61131_ (_10461_, _10460_, _07234_);
  and _61132_ (_10462_, _09511_, _06545_);
  and _61133_ (_10463_, _10462_, _10457_);
  or _61134_ (_10464_, _10463_, _06366_);
  or _61135_ (_10465_, _10464_, _10461_);
  nor _61136_ (_10466_, _09043_, _09498_);
  or _61137_ (_10467_, _09494_, _09056_);
  or _61138_ (_10468_, _10467_, _10466_);
  and _61139_ (_10469_, _10468_, _09061_);
  and _61140_ (_10470_, _10469_, _10465_);
  nor _61141_ (_10471_, _08573_, _09498_);
  or _61142_ (_10472_, _10471_, _09494_);
  and _61143_ (_10473_, _10472_, _06528_);
  or _61144_ (_10474_, _10473_, _06568_);
  or _61145_ (_10475_, _10474_, _10470_);
  or _61146_ (_10476_, _09508_, _06926_);
  and _61147_ (_10477_, _10476_, _05928_);
  and _61148_ (_10478_, _10477_, _10475_);
  and _61149_ (_10479_, _09505_, _05927_);
  or _61150_ (_10480_, _10479_, _06278_);
  or _61151_ (_10481_, _10480_, _10478_);
  and _61152_ (_10482_, _08550_, _07942_);
  or _61153_ (_10483_, _09494_, _06279_);
  or _61154_ (_10484_, _10483_, _10482_);
  and _61155_ (_10485_, _10484_, _01347_);
  and _61156_ (_10486_, _10485_, _10481_);
  or _61157_ (_10487_, _10486_, _09493_);
  and _61158_ (_40573_, _10487_, _42618_);
  nor _61159_ (_10488_, _01347_, _08572_);
  nor _61160_ (_10489_, _07939_, _08572_);
  not _61161_ (_10490_, _07939_);
  nor _61162_ (_10491_, _09043_, _10490_);
  or _61163_ (_10492_, _10491_, _10489_);
  and _61164_ (_10493_, _10492_, _06366_);
  and _61165_ (_10494_, _08040_, _08572_);
  nor _61166_ (_10495_, _10494_, _07043_);
  and _61167_ (_10496_, _06370_, _06544_);
  not _61168_ (_10497_, _10496_);
  nor _61169_ (_10498_, _08755_, \oc8051_golden_model_1.ACC [7]);
  and _61170_ (_10499_, _08755_, \oc8051_golden_model_1.ACC [7]);
  nor _61171_ (_10500_, _10499_, _10498_);
  and _61172_ (_10501_, _06345_, _06535_);
  nor _61173_ (_10502_, _10501_, _06884_);
  or _61174_ (_10503_, _10502_, _10500_);
  nor _61175_ (_10504_, _08040_, _08572_);
  nor _61176_ (_10505_, _10504_, _10494_);
  and _61177_ (_10506_, _07041_, _06535_);
  or _61178_ (_10507_, _10506_, _06703_);
  nor _61179_ (_10508_, _10507_, _06887_);
  not _61180_ (_10509_, _10508_);
  and _61181_ (_10510_, _10509_, _10505_);
  or _61182_ (_10511_, _06182_, _05975_);
  nor _61183_ (_10512_, _08040_, _10490_);
  or _61184_ (_10513_, _10512_, _10489_);
  or _61185_ (_10514_, _10513_, _07215_);
  not _61186_ (_10515_, _05984_);
  and _61187_ (_10516_, _06370_, _05976_);
  not _61188_ (_10517_, _10516_);
  and _61189_ (_10518_, _07949_, \oc8051_golden_model_1.PSW [7]);
  and _61190_ (_10519_, _10518_, _07908_);
  and _61191_ (_10520_, _10519_, _07892_);
  and _61192_ (_10521_, _10520_, _07607_);
  and _61193_ (_10522_, _10521_, _06286_);
  nor _61194_ (_10523_, _10521_, _06286_);
  or _61195_ (_10524_, _10523_, _10522_);
  nor _61196_ (_10525_, _10524_, _08572_);
  and _61197_ (_10526_, _10524_, _08572_);
  nor _61198_ (_10527_, _10526_, _10525_);
  not _61199_ (_10528_, _10527_);
  nor _61200_ (_10529_, _10520_, _07607_);
  nor _61201_ (_10530_, _10529_, _10521_);
  nor _61202_ (_10531_, _10530_, _10116_);
  and _61203_ (_10532_, _10519_, _07883_);
  nor _61204_ (_10533_, _10532_, _07896_);
  nor _61205_ (_10534_, _10533_, _10520_);
  and _61206_ (_10535_, _10534_, _10170_);
  nor _61207_ (_10536_, _10534_, _10170_);
  nor _61208_ (_10537_, _10519_, _07883_);
  nor _61209_ (_10538_, _10537_, _10532_);
  nor _61210_ (_10539_, _10538_, _10135_);
  nor _61211_ (_10540_, _10539_, _10536_);
  nor _61212_ (_10541_, _10540_, _10535_);
  nor _61213_ (_10542_, _10536_, _10535_);
  not _61214_ (_10543_, _10542_);
  and _61215_ (_10544_, _10538_, _10135_);
  or _61216_ (_10545_, _10544_, _10539_);
  or _61217_ (_10546_, _10545_, _10543_);
  nor _61218_ (_10547_, _08807_, _06473_);
  nor _61219_ (_10548_, _10547_, _10519_);
  nor _61220_ (_10549_, _10548_, _06055_);
  and _61221_ (_10550_, _10548_, _06055_);
  nor _61222_ (_10551_, _10550_, _10549_);
  nor _61223_ (_10552_, _10518_, _06657_);
  nor _61224_ (_10553_, _10552_, _08807_);
  nor _61225_ (_10554_, _10553_, _10213_);
  and _61226_ (_10555_, _10553_, _10213_);
  nor _61227_ (_10556_, _10555_, _10554_);
  and _61228_ (_10557_, _10556_, _10551_);
  not _61229_ (_10558_, \oc8051_golden_model_1.PSW [7]);
  nor _61230_ (_10559_, _06251_, _10558_);
  nor _61231_ (_10560_, _10559_, _07005_);
  nor _61232_ (_10561_, _10560_, _10518_);
  nor _61233_ (_10562_, _10561_, _06042_);
  and _61234_ (_10563_, _06251_, _10558_);
  nor _61235_ (_10564_, _10563_, _10559_);
  and _61236_ (_10565_, _10564_, _06097_);
  and _61237_ (_10566_, _10561_, _06042_);
  nor _61238_ (_10567_, _10562_, _10566_);
  not _61239_ (_10568_, _10567_);
  nor _61240_ (_10569_, _10568_, _10565_);
  or _61241_ (_10570_, _10569_, _10562_);
  and _61242_ (_10571_, _10570_, _10557_);
  and _61243_ (_10572_, _10554_, _10551_);
  or _61244_ (_10573_, _10572_, _10549_);
  nor _61245_ (_10574_, _10573_, _10571_);
  nor _61246_ (_10575_, _10574_, _10546_);
  nor _61247_ (_10576_, _10575_, _10541_);
  and _61248_ (_10577_, _10530_, _10116_);
  nor _61249_ (_10578_, _10531_, _10577_);
  not _61250_ (_10579_, _10578_);
  nor _61251_ (_10580_, _10579_, _10576_);
  or _61252_ (_10581_, _10580_, _10531_);
  and _61253_ (_10582_, _10581_, _10528_);
  nor _61254_ (_10583_, _10581_, _10528_);
  or _61255_ (_10584_, _10583_, _10582_);
  or _61256_ (_10585_, _10584_, _10517_);
  and _61257_ (_10586_, _06343_, _05976_);
  and _61258_ (_10587_, _06345_, _05976_);
  nor _61259_ (_10588_, _10587_, _10586_);
  and _61260_ (_10589_, _09392_, \oc8051_golden_model_1.PSW [7]);
  and _61261_ (_10590_, _10589_, _09451_);
  and _61262_ (_10591_, _10590_, _09450_);
  and _61263_ (_10592_, _10591_, _09449_);
  and _61264_ (_10593_, _10592_, _09448_);
  and _61265_ (_10594_, _10593_, _09447_);
  and _61266_ (_10595_, _10594_, _09446_);
  nor _61267_ (_10596_, _10595_, _09076_);
  and _61268_ (_10597_, _10595_, _09076_);
  nor _61269_ (_10598_, _10597_, _10596_);
  and _61270_ (_10599_, _10598_, \oc8051_golden_model_1.ACC [7]);
  nor _61271_ (_10600_, _10598_, \oc8051_golden_model_1.ACC [7]);
  nor _61272_ (_10601_, _10600_, _10599_);
  not _61273_ (_10602_, _10601_);
  nor _61274_ (_10603_, _10594_, _09446_);
  nor _61275_ (_10604_, _10603_, _10595_);
  nor _61276_ (_10605_, _10604_, _10116_);
  nor _61277_ (_10606_, _10593_, _09447_);
  nor _61278_ (_10607_, _10606_, _10594_);
  and _61279_ (_10608_, _10607_, _10170_);
  nor _61280_ (_10609_, _10607_, _10170_);
  nor _61281_ (_10610_, _10609_, _10608_);
  not _61282_ (_10611_, _10610_);
  nor _61283_ (_10612_, _10592_, _09448_);
  nor _61284_ (_10613_, _10612_, _10593_);
  nor _61285_ (_10614_, _10613_, _10135_);
  and _61286_ (_10615_, _10613_, _10135_);
  or _61287_ (_10616_, _10615_, _10614_);
  or _61288_ (_10617_, _10616_, _10611_);
  nor _61289_ (_10618_, _10591_, _09449_);
  nor _61290_ (_10619_, _10618_, _10592_);
  nor _61291_ (_10620_, _10619_, _06055_);
  and _61292_ (_10621_, _10619_, _06055_);
  nor _61293_ (_10622_, _10621_, _10620_);
  nor _61294_ (_10623_, _10590_, _09450_);
  nor _61295_ (_10624_, _10623_, _10591_);
  nor _61296_ (_10625_, _10624_, _10213_);
  and _61297_ (_10626_, _10624_, _10213_);
  nor _61298_ (_10627_, _10626_, _10625_);
  and _61299_ (_10628_, _10627_, _10622_);
  nor _61300_ (_10629_, _10589_, _09451_);
  nor _61301_ (_10630_, _10629_, _10590_);
  nor _61302_ (_10631_, _10630_, _06042_);
  and _61303_ (_10632_, _10630_, _06042_);
  nor _61304_ (_10633_, _09392_, \oc8051_golden_model_1.PSW [7]);
  nor _61305_ (_10634_, _10633_, _10589_);
  and _61306_ (_10635_, _10634_, _06097_);
  nor _61307_ (_10636_, _10635_, _10632_);
  or _61308_ (_10637_, _10636_, _10631_);
  and _61309_ (_10638_, _10637_, _10628_);
  and _61310_ (_10639_, _10625_, _10622_);
  or _61311_ (_10640_, _10639_, _10620_);
  nor _61312_ (_10641_, _10640_, _10638_);
  nor _61313_ (_10642_, _10641_, _10617_);
  and _61314_ (_10643_, _10614_, _10610_);
  nor _61315_ (_10644_, _10643_, _10609_);
  not _61316_ (_10645_, _10644_);
  nor _61317_ (_10646_, _10645_, _10642_);
  and _61318_ (_10647_, _10604_, _10116_);
  nor _61319_ (_10648_, _10605_, _10647_);
  not _61320_ (_10649_, _10648_);
  nor _61321_ (_10650_, _10649_, _10646_);
  or _61322_ (_10651_, _10650_, _10605_);
  and _61323_ (_10652_, _10651_, _10602_);
  nor _61324_ (_10653_, _10651_, _10602_);
  or _61325_ (_10654_, _10653_, _10652_);
  or _61326_ (_10655_, _10654_, _10588_);
  not _61327_ (_10656_, _10588_);
  and _61328_ (_10657_, _07133_, \oc8051_golden_model_1.PSW [7]);
  and _61329_ (_10658_, _10657_, _09432_);
  and _61330_ (_10659_, _10658_, _09431_);
  and _61331_ (_10661_, _10659_, _07595_);
  and _61332_ (_10662_, _10661_, _09430_);
  and _61333_ (_10663_, _10662_, _09429_);
  and _61334_ (_10664_, _10663_, _09428_);
  and _61335_ (_10665_, _10664_, _08040_);
  nor _61336_ (_10666_, _10664_, _08040_);
  or _61337_ (_10667_, _10666_, _10665_);
  nor _61338_ (_10668_, _10667_, _08572_);
  and _61339_ (_10669_, _10667_, _08572_);
  nor _61340_ (_10670_, _10669_, _10668_);
  not _61341_ (_10672_, _10670_);
  nor _61342_ (_10673_, _10663_, _09428_);
  nor _61343_ (_10674_, _10673_, _10664_);
  nor _61344_ (_10675_, _10674_, _10116_);
  nor _61345_ (_10676_, _10662_, _09429_);
  nor _61346_ (_10677_, _10676_, _10663_);
  and _61347_ (_10678_, _10677_, _10170_);
  nor _61348_ (_10679_, _10677_, _10170_);
  nor _61349_ (_10680_, _10661_, _09430_);
  nor _61350_ (_10681_, _10680_, _10662_);
  nor _61351_ (_10683_, _10681_, _10135_);
  nor _61352_ (_10684_, _10683_, _10679_);
  nor _61353_ (_10685_, _10684_, _10678_);
  nor _61354_ (_10686_, _10679_, _10678_);
  not _61355_ (_10687_, _10686_);
  and _61356_ (_10688_, _10681_, _10135_);
  or _61357_ (_10689_, _10688_, _10683_);
  or _61358_ (_10690_, _10689_, _10687_);
  nor _61359_ (_10691_, _10659_, _07595_);
  nor _61360_ (_10692_, _10691_, _10661_);
  nor _61361_ (_10694_, _10692_, _06055_);
  and _61362_ (_10695_, _10692_, _06055_);
  nor _61363_ (_10696_, _10695_, _10694_);
  nor _61364_ (_10697_, _10658_, _09431_);
  nor _61365_ (_10698_, _10697_, _10659_);
  nor _61366_ (_10699_, _10698_, _10213_);
  and _61367_ (_10700_, _10698_, _10213_);
  nor _61368_ (_10701_, _10700_, _10699_);
  and _61369_ (_10702_, _10701_, _10696_);
  nor _61370_ (_10703_, _10657_, _09432_);
  nor _61371_ (_10705_, _10703_, _10658_);
  nor _61372_ (_10706_, _10705_, _06042_);
  and _61373_ (_10707_, _10705_, _06042_);
  nor _61374_ (_10708_, _07133_, \oc8051_golden_model_1.PSW [7]);
  nor _61375_ (_10709_, _10708_, _10657_);
  and _61376_ (_10710_, _10709_, _06097_);
  nor _61377_ (_10711_, _10710_, _10707_);
  or _61378_ (_10712_, _10711_, _10706_);
  nand _61379_ (_10713_, _10712_, _10702_);
  and _61380_ (_10714_, _10699_, _10696_);
  nor _61381_ (_10716_, _10714_, _10694_);
  and _61382_ (_10717_, _10716_, _10713_);
  nor _61383_ (_10718_, _10717_, _10690_);
  nor _61384_ (_10719_, _10718_, _10685_);
  and _61385_ (_10720_, _10674_, _10116_);
  nor _61386_ (_10721_, _10675_, _10720_);
  not _61387_ (_10722_, _10721_);
  nor _61388_ (_10723_, _10722_, _10719_);
  or _61389_ (_10724_, _10723_, _10675_);
  and _61390_ (_10725_, _10724_, _10672_);
  nor _61391_ (_10727_, _10724_, _10672_);
  or _61392_ (_10728_, _10727_, _10725_);
  and _61393_ (_10729_, _07041_, _05976_);
  and _61394_ (_10730_, _06327_, _05976_);
  nor _61395_ (_10731_, _10730_, _10729_);
  and _61396_ (_10732_, _06336_, _05972_);
  and _61397_ (_10733_, _10732_, _05976_);
  not _61398_ (_10734_, _10733_);
  and _61399_ (_10735_, _10734_, _10731_);
  or _61400_ (_10736_, _10735_, _10728_);
  not _61401_ (_10737_, _10735_);
  nor _61402_ (_10738_, _10049_, _10047_);
  nor _61403_ (_10739_, _10738_, _10050_);
  or _61404_ (_10740_, _10739_, _09537_);
  not _61405_ (_10741_, _06700_);
  nor _61406_ (_10742_, _07794_, _06741_);
  and _61407_ (_10743_, _10742_, _10741_);
  not _61408_ (_10744_, _10743_);
  nand _61409_ (_10745_, _10744_, _08040_);
  nor _61410_ (_10746_, _08636_, _08572_);
  and _61411_ (_10747_, _08773_, _08636_);
  or _61412_ (_10748_, _10747_, _10746_);
  or _61413_ (_10749_, _10748_, _06273_);
  and _61414_ (_10750_, _10749_, _07166_);
  not _61415_ (_10751_, _06784_);
  nor _61416_ (_10752_, _06345_, _07209_);
  and _61417_ (_10753_, _10752_, _07212_);
  nor _61418_ (_10754_, _10753_, _06014_);
  nor _61419_ (_10755_, _10754_, _10751_);
  not _61420_ (_10756_, _10755_);
  nand _61421_ (_10757_, _10756_, _08040_);
  and _61422_ (_10758_, _06370_, _06706_);
  not _61423_ (_10759_, _10758_);
  nor _61424_ (_10760_, _06781_, _08572_);
  and _61425_ (_10761_, _06781_, _08572_);
  nor _61426_ (_10762_, _10761_, _10760_);
  nand _61427_ (_10763_, _10762_, _10755_);
  and _61428_ (_10764_, _10763_, _10759_);
  and _61429_ (_10765_, _10764_, _10757_);
  and _61430_ (_10766_, _10758_, _08755_);
  or _61431_ (_10767_, _10766_, _10765_);
  not _61432_ (_10768_, _06015_);
  nor _61433_ (_10769_, _06341_, _10768_);
  and _61434_ (_10770_, _10769_, _10767_);
  and _61435_ (_10771_, _08768_, _07939_);
  or _61436_ (_10772_, _10771_, _10489_);
  and _61437_ (_10773_, _10772_, _06341_);
  or _61438_ (_10774_, _10773_, _10770_);
  and _61439_ (_10775_, _06370_, _06271_);
  not _61440_ (_10776_, _10775_);
  and _61441_ (_10777_, _10776_, _10774_);
  nor _61442_ (_10778_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor _61443_ (_10779_, _10778_, _06055_);
  and _61444_ (_10780_, _10779_, \oc8051_golden_model_1.ACC [4]);
  and _61445_ (_10781_, _10780_, \oc8051_golden_model_1.ACC [5]);
  and _61446_ (_10782_, _10781_, \oc8051_golden_model_1.ACC [6]);
  and _61447_ (_10783_, _10782_, \oc8051_golden_model_1.ACC [7]);
  nor _61448_ (_10784_, _10782_, \oc8051_golden_model_1.ACC [7]);
  nor _61449_ (_10785_, _10784_, _10783_);
  nor _61450_ (_10786_, _10780_, \oc8051_golden_model_1.ACC [5]);
  nor _61451_ (_10787_, _10786_, _10781_);
  nor _61452_ (_10788_, _10781_, \oc8051_golden_model_1.ACC [6]);
  nor _61453_ (_10789_, _10788_, _10782_);
  nor _61454_ (_10790_, _10789_, _10787_);
  not _61455_ (_10791_, _10790_);
  and _61456_ (_10792_, _10791_, _10785_);
  not _61457_ (_10793_, _10792_);
  nor _61458_ (_10794_, _10783_, \oc8051_golden_model_1.PSW [7]);
  and _61459_ (_10795_, _10794_, _10793_);
  nor _61460_ (_10796_, _10795_, _10790_);
  or _61461_ (_10797_, _10796_, _10785_);
  and _61462_ (_10798_, _10793_, _10775_);
  and _61463_ (_10799_, _10798_, _10797_);
  or _61464_ (_10800_, _10799_, _06272_);
  or _61465_ (_10801_, _10800_, _10777_);
  and _61466_ (_10802_, _10801_, _10750_);
  and _61467_ (_10803_, _10513_, _06461_);
  or _61468_ (_10804_, _10803_, _10744_);
  or _61469_ (_10805_, _10804_, _10802_);
  and _61470_ (_10806_, _10805_, _10745_);
  or _61471_ (_10807_, _10806_, _07174_);
  or _61472_ (_10808_, _08755_, _07175_);
  and _61473_ (_10809_, _10808_, _06465_);
  and _61474_ (_10810_, _10809_, _10807_);
  and _61475_ (_10811_, _06370_, _06266_);
  nor _61476_ (_10812_, _08042_, _06465_);
  or _61477_ (_10813_, _10812_, _10811_);
  or _61478_ (_10814_, _10813_, _10810_);
  nand _61479_ (_10815_, _10811_, _06055_);
  and _61480_ (_10816_, _10815_, _10814_);
  or _61481_ (_10817_, _10816_, _06268_);
  and _61482_ (_10818_, _08649_, _08636_);
  or _61483_ (_10819_, _10818_, _10746_);
  or _61484_ (_10820_, _10819_, _06269_);
  and _61485_ (_10821_, _10820_, _06262_);
  and _61486_ (_10822_, _10821_, _10817_);
  or _61487_ (_10823_, _10746_, _08789_);
  and _61488_ (_10824_, _10823_, _06261_);
  and _61489_ (_10825_, _10824_, _10748_);
  or _61490_ (_10826_, _10825_, _09531_);
  or _61491_ (_10827_, _10826_, _10822_);
  and _61492_ (_10828_, _10827_, _10740_);
  or _61493_ (_10829_, _10828_, _10737_);
  and _61494_ (_10830_, _10829_, _10736_);
  or _61495_ (_10831_, _10830_, _10656_);
  and _61496_ (_10832_, _10831_, _06517_);
  and _61497_ (_10833_, _10832_, _10655_);
  and _61498_ (_10834_, _08390_, \oc8051_golden_model_1.PSW [7]);
  and _61499_ (_10835_, _10834_, _08341_);
  and _61500_ (_10836_, _10835_, _08440_);
  and _61501_ (_10837_, _10836_, _08292_);
  and _61502_ (_10838_, _10837_, _08544_);
  and _61503_ (_10839_, _10838_, _08247_);
  and _61504_ (_10840_, _10839_, _08145_);
  nor _61505_ (_10841_, _10840_, _08042_);
  and _61506_ (_10842_, _10840_, _08042_);
  nor _61507_ (_10843_, _10842_, _10841_);
  and _61508_ (_10844_, _10843_, \oc8051_golden_model_1.ACC [7]);
  nor _61509_ (_10845_, _10843_, \oc8051_golden_model_1.ACC [7]);
  nor _61510_ (_10846_, _10845_, _10844_);
  not _61511_ (_10847_, _10846_);
  nor _61512_ (_10848_, _10839_, _08145_);
  nor _61513_ (_10849_, _10848_, _10840_);
  nor _61514_ (_10850_, _10849_, _10116_);
  nor _61515_ (_10851_, _10838_, _08247_);
  nor _61516_ (_10852_, _10851_, _10839_);
  and _61517_ (_10853_, _10852_, _10170_);
  nor _61518_ (_10854_, _10852_, _10170_);
  nor _61519_ (_10855_, _10837_, _08544_);
  nor _61520_ (_10856_, _10855_, _10838_);
  nor _61521_ (_10857_, _10856_, _10135_);
  nor _61522_ (_10858_, _10857_, _10854_);
  nor _61523_ (_10859_, _10858_, _10853_);
  nor _61524_ (_10860_, _10854_, _10853_);
  not _61525_ (_10861_, _10860_);
  and _61526_ (_10862_, _10856_, _10135_);
  or _61527_ (_10863_, _10862_, _10857_);
  or _61528_ (_10864_, _10863_, _10861_);
  nor _61529_ (_10865_, _10836_, _08292_);
  nor _61530_ (_10866_, _10865_, _10837_);
  nor _61531_ (_10867_, _10866_, _06055_);
  and _61532_ (_10868_, _10866_, _06055_);
  nor _61533_ (_10869_, _10868_, _10867_);
  nor _61534_ (_10870_, _10835_, _08440_);
  nor _61535_ (_10871_, _10870_, _10836_);
  nor _61536_ (_10872_, _10871_, _10213_);
  and _61537_ (_10873_, _10871_, _10213_);
  nor _61538_ (_10874_, _10873_, _10872_);
  and _61539_ (_10875_, _10874_, _10869_);
  nor _61540_ (_10876_, _10834_, _08341_);
  nor _61541_ (_10877_, _10876_, _10835_);
  nor _61542_ (_10878_, _10877_, _06042_);
  and _61543_ (_10879_, _10877_, _06042_);
  nor _61544_ (_10880_, _08390_, \oc8051_golden_model_1.PSW [7]);
  nor _61545_ (_10881_, _10880_, _10834_);
  and _61546_ (_10882_, _10881_, _06097_);
  nor _61547_ (_10883_, _10882_, _10879_);
  or _61548_ (_10884_, _10883_, _10878_);
  nand _61549_ (_10885_, _10884_, _10875_);
  and _61550_ (_10886_, _10872_, _10869_);
  nor _61551_ (_10887_, _10886_, _10867_);
  and _61552_ (_10888_, _10887_, _10885_);
  nor _61553_ (_10889_, _10888_, _10864_);
  nor _61554_ (_10890_, _10889_, _10859_);
  and _61555_ (_10891_, _10849_, _10116_);
  nor _61556_ (_10892_, _10850_, _10891_);
  not _61557_ (_10893_, _10892_);
  nor _61558_ (_10894_, _10893_, _10890_);
  or _61559_ (_10895_, _10894_, _10850_);
  and _61560_ (_10896_, _10895_, _10847_);
  nor _61561_ (_10897_, _10895_, _10847_);
  or _61562_ (_10898_, _10897_, _10896_);
  and _61563_ (_10899_, _10898_, _06512_);
  or _61564_ (_10900_, _10899_, _10516_);
  or _61565_ (_10901_, _10900_, _10833_);
  and _61566_ (_10902_, _10901_, _10585_);
  or _61567_ (_10903_, _10902_, _10515_);
  or _61568_ (_10904_, _06182_, _05984_);
  and _61569_ (_10905_, _10904_, _06258_);
  and _61570_ (_10906_, _10905_, _10903_);
  and _61571_ (_10907_, _08808_, _08636_);
  or _61572_ (_10908_, _10907_, _10746_);
  and _61573_ (_10909_, _10908_, _06257_);
  or _61574_ (_10910_, _10909_, _10080_);
  or _61575_ (_10911_, _10910_, _10906_);
  and _61576_ (_10912_, _10911_, _10514_);
  or _61577_ (_10913_, _10912_, _07460_);
  and _61578_ (_10914_, _08755_, _07939_);
  or _61579_ (_10915_, _10489_, _07208_);
  or _61580_ (_10916_, _10915_, _10914_);
  and _61581_ (_10917_, _10916_, _05982_);
  and _61582_ (_10918_, _10917_, _10913_);
  and _61583_ (_10919_, _09021_, _07939_);
  or _61584_ (_10920_, _10919_, _10489_);
  and _61585_ (_10921_, _10920_, _10094_);
  or _61586_ (_10922_, _10921_, _10093_);
  or _61587_ (_10923_, _10922_, _10918_);
  or _61588_ (_10924_, _10114_, _10100_);
  and _61589_ (_10925_, _10924_, _10923_);
  or _61590_ (_10926_, _10925_, _05974_);
  and _61591_ (_10927_, _10926_, _10511_);
  or _61592_ (_10928_, _10927_, _06218_);
  and _61593_ (_10929_, _06370_, _06321_);
  not _61594_ (_10930_, _10929_);
  and _61595_ (_10931_, _08825_, _07939_);
  nor _61596_ (_10932_, _10931_, _10489_);
  nand _61597_ (_10933_, _10932_, _06218_);
  and _61598_ (_10934_, _10933_, _10930_);
  and _61599_ (_10935_, _10934_, _10928_);
  and _61600_ (_10936_, _10929_, _06182_);
  nor _61601_ (_10937_, _07211_, _05954_);
  or _61602_ (_10938_, _10937_, _10936_);
  or _61603_ (_10939_, _10938_, _10935_);
  not _61604_ (_10940_, _10937_);
  or _61605_ (_10941_, _10940_, _10505_);
  and _61606_ (_10942_, _10941_, _10508_);
  and _61607_ (_10943_, _10942_, _10939_);
  or _61608_ (_10944_, _10943_, _10510_);
  and _61609_ (_10945_, _07209_, _06535_);
  not _61610_ (_10946_, _10945_);
  and _61611_ (_10947_, _10946_, _10944_);
  not _61612_ (_10948_, _10502_);
  and _61613_ (_10949_, _10945_, _10505_);
  or _61614_ (_10950_, _10949_, _10948_);
  or _61615_ (_10951_, _10950_, _10947_);
  and _61616_ (_10952_, _10951_, _10503_);
  or _61617_ (_10953_, _10952_, _06533_);
  and _61618_ (_10954_, _06370_, _06535_);
  not _61619_ (_10955_, _10954_);
  or _61620_ (_10956_, _08575_, _06534_);
  and _61621_ (_10957_, _10956_, _10955_);
  nand _61622_ (_10958_, _10957_, _10953_);
  nor _61623_ (_10959_, _06182_, \oc8051_golden_model_1.ACC [7]);
  and _61624_ (_10960_, _06182_, \oc8051_golden_model_1.ACC [7]);
  nor _61625_ (_10961_, _10960_, _10959_);
  nand _61626_ (_10962_, _10954_, _10961_);
  and _61627_ (_10963_, _10962_, _07237_);
  and _61628_ (_10964_, _10963_, _10958_);
  and _61629_ (_10965_, _09044_, _07939_);
  nor _61630_ (_10966_, _10965_, _10489_);
  and _61631_ (_10967_, _10966_, _06369_);
  or _61632_ (_10968_, _10967_, _10964_);
  and _61633_ (_10969_, _10968_, _07240_);
  nor _61634_ (_10970_, _10489_, _07240_);
  nor _61635_ (_10971_, _07482_, _05960_);
  not _61636_ (_10972_, _10971_);
  and _61637_ (_10973_, _06886_, _06544_);
  and _61638_ (_10974_, _07041_, _06544_);
  nor _61639_ (_10975_, _10974_, _10973_);
  and _61640_ (_10976_, _06327_, _06544_);
  not _61641_ (_10977_, _10976_);
  and _61642_ (_10978_, _10977_, _10975_);
  and _61643_ (_10979_, _10978_, _10972_);
  not _61644_ (_10980_, _10979_);
  or _61645_ (_10981_, _10980_, _10970_);
  or _61646_ (_10982_, _10981_, _10969_);
  nor _61647_ (_10983_, _07153_, _05960_);
  nand _61648_ (_10984_, _10983_, _10499_);
  and _61649_ (_10985_, _06336_, _06544_);
  nor _61650_ (_10986_, _10985_, _10976_);
  not _61651_ (_10987_, _10986_);
  nand _61652_ (_10988_, _10987_, _10504_);
  and _61653_ (_10989_, _10988_, _06543_);
  and _61654_ (_10990_, _10989_, _10984_);
  and _61655_ (_10991_, _10990_, _10982_);
  nor _61656_ (_10992_, _08574_, _06543_);
  or _61657_ (_10993_, _10992_, _10991_);
  and _61658_ (_10994_, _10993_, _10497_);
  nor _61659_ (_10995_, _10960_, _10497_);
  or _61660_ (_10996_, _10995_, _06375_);
  nor _61661_ (_10997_, _10996_, _10994_);
  nor _61662_ (_10998_, _06755_, _06711_);
  not _61663_ (_10999_, _10998_);
  or _61664_ (_11000_, _10932_, _07242_);
  nor _61665_ (_11001_, _11000_, _08573_);
  or _61666_ (_11002_, _11001_, _10999_);
  or _61667_ (_11003_, _11002_, _10997_);
  nand _61668_ (_11004_, _10999_, _10494_);
  and _61669_ (_11005_, _11004_, _07043_);
  and _61670_ (_11006_, _11005_, _11003_);
  or _61671_ (_11007_, _11006_, _10495_);
  and _61672_ (_11008_, _07209_, _06527_);
  not _61673_ (_11009_, _11008_);
  and _61674_ (_11010_, _11009_, _11007_);
  and _61675_ (_11011_, _06343_, _06527_);
  and _61676_ (_11012_, _06345_, _06527_);
  nor _61677_ (_11013_, _11012_, _11011_);
  not _61678_ (_11014_, _11013_);
  nor _61679_ (_11015_, _11009_, _10494_);
  or _61680_ (_11016_, _11015_, _11014_);
  or _61681_ (_11017_, _11016_, _11010_);
  nand _61682_ (_11018_, _11014_, _10498_);
  and _61683_ (_11019_, _11018_, _06531_);
  and _61684_ (_11020_, _11019_, _11017_);
  and _61685_ (_11021_, _06370_, _06527_);
  nor _61686_ (_11022_, _11021_, _06530_);
  not _61687_ (_11023_, _11022_);
  not _61688_ (_11024_, _11021_);
  nand _61689_ (_11025_, _11024_, _08573_);
  and _61690_ (_11026_, _11025_, _11023_);
  or _61691_ (_11027_, _11026_, _11020_);
  nand _61692_ (_11028_, _11021_, _10959_);
  and _61693_ (_11029_, _11028_, _09056_);
  and _61694_ (_11030_, _11029_, _11027_);
  or _61695_ (_11031_, _11030_, _10493_);
  nor _61696_ (_11032_, _07041_, _06353_);
  nor _61697_ (_11033_, _11032_, _05958_);
  nor _61698_ (_11034_, _07211_, _05958_);
  or _61699_ (_11035_, _11034_, _11033_);
  and _61700_ (_11036_, _10732_, _06364_);
  nor _61701_ (_11037_, _11036_, _11035_);
  and _61702_ (_11038_, _11037_, _11031_);
  and _61703_ (_11039_, _06343_, _06364_);
  and _61704_ (_11040_, _06345_, _06364_);
  or _61705_ (_11041_, _11040_, _11039_);
  and _61706_ (_11042_, _10674_, \oc8051_golden_model_1.ACC [6]);
  and _61707_ (_11043_, _10677_, \oc8051_golden_model_1.ACC [5]);
  nand _61708_ (_11044_, _10681_, \oc8051_golden_model_1.ACC [4]);
  and _61709_ (_11045_, _10692_, \oc8051_golden_model_1.ACC [3]);
  and _61710_ (_11046_, _10698_, \oc8051_golden_model_1.ACC [2]);
  and _61711_ (_11047_, _10705_, \oc8051_golden_model_1.ACC [1]);
  nor _61712_ (_11048_, _10707_, _10706_);
  not _61713_ (_11049_, _11048_);
  and _61714_ (_11050_, _10709_, \oc8051_golden_model_1.ACC [0]);
  and _61715_ (_11051_, _11050_, _11049_);
  nor _61716_ (_11052_, _11051_, _11047_);
  nor _61717_ (_11053_, _11052_, _10701_);
  nor _61718_ (_11054_, _11053_, _11046_);
  nor _61719_ (_11055_, _11054_, _10696_);
  or _61720_ (_11056_, _11055_, _11045_);
  nand _61721_ (_11057_, _11056_, _10689_);
  and _61722_ (_11058_, _11057_, _11044_);
  nor _61723_ (_11059_, _11058_, _10686_);
  or _61724_ (_11060_, _11059_, _11043_);
  and _61725_ (_11061_, _11060_, _10722_);
  nor _61726_ (_11062_, _11061_, _11042_);
  and _61727_ (_11063_, _11062_, _10670_);
  nor _61728_ (_11064_, _11062_, _10670_);
  or _61729_ (_11065_, _11064_, _11037_);
  nor _61730_ (_11066_, _11065_, _11063_);
  or _61731_ (_11067_, _11066_, _11041_);
  or _61732_ (_11068_, _11067_, _11038_);
  not _61733_ (_11069_, _11041_);
  nand _61734_ (_11070_, _10604_, \oc8051_golden_model_1.ACC [6]);
  and _61735_ (_11071_, _10607_, \oc8051_golden_model_1.ACC [5]);
  nand _61736_ (_11072_, _10613_, \oc8051_golden_model_1.ACC [4]);
  and _61737_ (_11073_, _10619_, \oc8051_golden_model_1.ACC [3]);
  and _61738_ (_11074_, _10624_, \oc8051_golden_model_1.ACC [2]);
  and _61739_ (_11075_, _10630_, \oc8051_golden_model_1.ACC [1]);
  nor _61740_ (_11076_, _10632_, _10631_);
  not _61741_ (_11077_, _11076_);
  and _61742_ (_11078_, _10634_, \oc8051_golden_model_1.ACC [0]);
  and _61743_ (_11079_, _11078_, _11077_);
  nor _61744_ (_11080_, _11079_, _11075_);
  nor _61745_ (_11081_, _11080_, _10627_);
  nor _61746_ (_11082_, _11081_, _11074_);
  nor _61747_ (_11083_, _11082_, _10622_);
  or _61748_ (_11084_, _11083_, _11073_);
  nand _61749_ (_11085_, _11084_, _10616_);
  and _61750_ (_11086_, _11085_, _11072_);
  nor _61751_ (_11087_, _11086_, _10610_);
  or _61752_ (_11088_, _11087_, _11071_);
  nand _61753_ (_11089_, _11088_, _10649_);
  and _61754_ (_11090_, _11089_, _11070_);
  nor _61755_ (_11091_, _11090_, _10601_);
  and _61756_ (_11092_, _11090_, _10601_);
  nor _61757_ (_11093_, _11092_, _11091_);
  or _61758_ (_11094_, _11093_, _11069_);
  and _61759_ (_11095_, _11094_, _06541_);
  and _61760_ (_11096_, _11095_, _11068_);
  and _61761_ (_11097_, _06370_, _06364_);
  nand _61762_ (_11098_, _10849_, \oc8051_golden_model_1.ACC [6]);
  and _61763_ (_11099_, _10852_, \oc8051_golden_model_1.ACC [5]);
  nand _61764_ (_11100_, _10856_, \oc8051_golden_model_1.ACC [4]);
  and _61765_ (_11101_, _10866_, \oc8051_golden_model_1.ACC [3]);
  and _61766_ (_11102_, _10871_, \oc8051_golden_model_1.ACC [2]);
  and _61767_ (_11103_, _10877_, \oc8051_golden_model_1.ACC [1]);
  nor _61768_ (_11104_, _10879_, _10878_);
  not _61769_ (_11105_, _11104_);
  and _61770_ (_11106_, _10881_, \oc8051_golden_model_1.ACC [0]);
  and _61771_ (_11107_, _11106_, _11105_);
  nor _61772_ (_11108_, _11107_, _11103_);
  nor _61773_ (_11109_, _11108_, _10874_);
  nor _61774_ (_11110_, _11109_, _11102_);
  nor _61775_ (_11111_, _11110_, _10869_);
  or _61776_ (_11112_, _11111_, _11101_);
  nand _61777_ (_11113_, _11112_, _10863_);
  and _61778_ (_11114_, _11113_, _11100_);
  nor _61779_ (_11115_, _11114_, _10860_);
  or _61780_ (_11116_, _11115_, _11099_);
  nand _61781_ (_11117_, _11116_, _10893_);
  and _61782_ (_11118_, _11117_, _11098_);
  nor _61783_ (_11119_, _11118_, _10846_);
  and _61784_ (_11120_, _11118_, _10846_);
  nor _61785_ (_11121_, _11120_, _11119_);
  and _61786_ (_11122_, _11121_, _06540_);
  or _61787_ (_11123_, _11122_, _11097_);
  or _61788_ (_11124_, _11123_, _11096_);
  nor _61789_ (_11125_, _05973_, _05958_);
  not _61790_ (_11126_, _11125_);
  not _61791_ (_11127_, _11097_);
  and _61792_ (_11128_, _10530_, \oc8051_golden_model_1.ACC [6]);
  and _61793_ (_11129_, _10534_, \oc8051_golden_model_1.ACC [5]);
  nand _61794_ (_11130_, _10538_, \oc8051_golden_model_1.ACC [4]);
  and _61795_ (_11131_, _10548_, \oc8051_golden_model_1.ACC [3]);
  and _61796_ (_11132_, _10553_, \oc8051_golden_model_1.ACC [2]);
  and _61797_ (_11133_, _10561_, \oc8051_golden_model_1.ACC [1]);
  and _61798_ (_11134_, _10564_, \oc8051_golden_model_1.ACC [0]);
  and _61799_ (_11135_, _11134_, _10568_);
  nor _61800_ (_11136_, _11135_, _11133_);
  nor _61801_ (_11137_, _11136_, _10556_);
  nor _61802_ (_11138_, _11137_, _11132_);
  nor _61803_ (_11139_, _11138_, _10551_);
  or _61804_ (_11140_, _11139_, _11131_);
  nand _61805_ (_11141_, _11140_, _10545_);
  and _61806_ (_11142_, _11141_, _11130_);
  nor _61807_ (_11143_, _11142_, _10542_);
  or _61808_ (_11144_, _11143_, _11129_);
  and _61809_ (_11145_, _11144_, _10579_);
  nor _61810_ (_11146_, _11145_, _11128_);
  nor _61811_ (_11147_, _11146_, _10527_);
  and _61812_ (_11148_, _11146_, _10527_);
  nor _61813_ (_11149_, _11148_, _11147_);
  or _61814_ (_11150_, _11149_, _11127_);
  and _61815_ (_11151_, _11150_, _11126_);
  and _61816_ (_11152_, _11151_, _11124_);
  nand _61817_ (_11153_, _11125_, \oc8051_golden_model_1.ACC [6]);
  and _61818_ (_11154_, _07209_, _06280_);
  and _61819_ (_11155_, _06327_, _06280_);
  or _61820_ (_11156_, _11155_, _07045_);
  nor _61821_ (_11157_, _11156_, _11154_);
  nand _61822_ (_11158_, _11157_, _11153_);
  or _61823_ (_11159_, _11158_, _11152_);
  nor _61824_ (_11160_, _08142_, _10116_);
  not _61825_ (_11161_, _11160_);
  nand _61826_ (_11162_, _08142_, _10116_);
  and _61827_ (_11163_, _11162_, _11161_);
  nor _61828_ (_11164_, _08244_, _10170_);
  and _61829_ (_11165_, _08244_, _10170_);
  nor _61830_ (_11166_, _11165_, _11164_);
  nor _61831_ (_11167_, _08541_, _10135_);
  not _61832_ (_11168_, _11167_);
  nand _61833_ (_11169_, _08541_, _10135_);
  and _61834_ (_11170_, _11169_, _11168_);
  nor _61835_ (_11171_, _07594_, _06055_);
  and _61836_ (_11172_, _07594_, _06055_);
  nor _61837_ (_11173_, _07776_, _10213_);
  and _61838_ (_11174_, _07776_, _10213_);
  nor _61839_ (_11175_, _11174_, _11173_);
  nor _61840_ (_11176_, _07357_, _06042_);
  and _61841_ (_11177_, _07357_, _06042_);
  nor _61842_ (_11178_, _11177_, _11176_);
  and _61843_ (_11179_, _07133_, \oc8051_golden_model_1.ACC [0]);
  and _61844_ (_11180_, _11179_, _11178_);
  nor _61845_ (_11181_, _11180_, _11176_);
  not _61846_ (_11182_, _11181_);
  and _61847_ (_11183_, _11182_, _11175_);
  nor _61848_ (_11184_, _11183_, _11173_);
  nor _61849_ (_11185_, _11184_, _11172_);
  or _61850_ (_11186_, _11185_, _11171_);
  and _61851_ (_11187_, _11186_, _11170_);
  nor _61852_ (_11188_, _11187_, _11167_);
  not _61853_ (_11189_, _11188_);
  and _61854_ (_11190_, _11189_, _11166_);
  or _61855_ (_11191_, _11190_, _11164_);
  and _61856_ (_11192_, _11191_, _11163_);
  nor _61857_ (_11193_, _11192_, _11160_);
  and _61858_ (_11194_, _11193_, _10505_);
  nor _61859_ (_11195_, _11193_, _10505_);
  or _61860_ (_11196_, _11195_, _11194_);
  or _61861_ (_11197_, _11196_, _11157_);
  and _61862_ (_11198_, _11197_, _11159_);
  and _61863_ (_11199_, _06343_, _06280_);
  and _61864_ (_11200_, _06345_, _06280_);
  or _61865_ (_11201_, _11200_, _11199_);
  or _61866_ (_11202_, _11201_, _11198_);
  not _61867_ (_11203_, _11201_);
  and _61868_ (_11204_, _09446_, \oc8051_golden_model_1.ACC [6]);
  or _61869_ (_11205_, _09446_, \oc8051_golden_model_1.ACC [6]);
  not _61870_ (_11206_, _11204_);
  and _61871_ (_11207_, _11206_, _11205_);
  and _61872_ (_11208_, _09447_, \oc8051_golden_model_1.ACC [5]);
  and _61873_ (_11209_, _09167_, _10170_);
  or _61874_ (_11210_, _11209_, _11208_);
  and _61875_ (_11211_, _09448_, \oc8051_golden_model_1.ACC [4]);
  not _61876_ (_11212_, _11211_);
  or _61877_ (_11213_, _09448_, \oc8051_golden_model_1.ACC [4]);
  and _61878_ (_11214_, _11212_, _11213_);
  and _61879_ (_11215_, _09449_, \oc8051_golden_model_1.ACC [3]);
  and _61880_ (_11216_, _09257_, _06055_);
  and _61881_ (_11217_, _09450_, \oc8051_golden_model_1.ACC [2]);
  and _61882_ (_11218_, _09302_, _10213_);
  nor _61883_ (_11219_, _11217_, _11218_);
  and _61884_ (_11220_, _09451_, \oc8051_golden_model_1.ACC [1]);
  and _61885_ (_11221_, _09347_, _06042_);
  nor _61886_ (_11222_, _11220_, _11221_);
  and _61887_ (_11223_, _09392_, \oc8051_golden_model_1.ACC [0]);
  and _61888_ (_11224_, _11223_, _11222_);
  nor _61889_ (_11225_, _11224_, _11220_);
  not _61890_ (_11226_, _11225_);
  and _61891_ (_11227_, _11226_, _11219_);
  nor _61892_ (_11228_, _11227_, _11217_);
  nor _61893_ (_11229_, _11228_, _11216_);
  or _61894_ (_11230_, _11229_, _11215_);
  nand _61895_ (_11231_, _11230_, _11214_);
  and _61896_ (_11232_, _11231_, _11212_);
  nor _61897_ (_11233_, _11232_, _11210_);
  or _61898_ (_11234_, _11233_, _11208_);
  and _61899_ (_11235_, _11234_, _11207_);
  nor _61900_ (_11236_, _11235_, _11204_);
  and _61901_ (_11237_, _11236_, _10500_);
  nor _61902_ (_11238_, _11236_, _10500_);
  or _61903_ (_11239_, _11238_, _11237_);
  or _61904_ (_11240_, _11239_, _11203_);
  and _61905_ (_11241_, _11240_, _06285_);
  and _61906_ (_11242_, _11241_, _11202_);
  and _61907_ (_11243_, _06370_, _06280_);
  nor _61908_ (_11244_, _08144_, _10116_);
  not _61909_ (_11245_, _11244_);
  and _61910_ (_11246_, _08144_, _10116_);
  nor _61911_ (_11247_, _11246_, _11244_);
  nor _61912_ (_11248_, _08246_, _10170_);
  and _61913_ (_11249_, _08246_, _10170_);
  nor _61914_ (_11250_, _11249_, _11248_);
  nor _61915_ (_11251_, _08543_, _10135_);
  not _61916_ (_11252_, _11251_);
  and _61917_ (_11253_, _08543_, _10135_);
  nor _61918_ (_11254_, _11253_, _11251_);
  nor _61919_ (_11255_, _08291_, _06055_);
  and _61920_ (_11256_, _08291_, _06055_);
  nor _61921_ (_11257_, _08439_, _10213_);
  and _61922_ (_11258_, _08439_, _10213_);
  nor _61923_ (_11259_, _11258_, _11257_);
  nor _61924_ (_11260_, _08340_, _06042_);
  and _61925_ (_11261_, _08340_, _06042_);
  nor _61926_ (_11262_, _11261_, _11260_);
  and _61927_ (_11263_, _08390_, \oc8051_golden_model_1.ACC [0]);
  and _61928_ (_11264_, _11263_, _11262_);
  nor _61929_ (_11265_, _11264_, _11260_);
  not _61930_ (_11266_, _11265_);
  and _61931_ (_11267_, _11266_, _11259_);
  nor _61932_ (_11268_, _11267_, _11257_);
  nor _61933_ (_11269_, _11268_, _11256_);
  or _61934_ (_11270_, _11269_, _11255_);
  nand _61935_ (_11271_, _11270_, _11254_);
  and _61936_ (_11272_, _11271_, _11252_);
  not _61937_ (_11273_, _11272_);
  and _61938_ (_11274_, _11273_, _11250_);
  or _61939_ (_11275_, _11274_, _11248_);
  nand _61940_ (_11276_, _11275_, _11247_);
  and _61941_ (_11277_, _11276_, _11245_);
  nor _61942_ (_11278_, _11277_, _08575_);
  and _61943_ (_11279_, _11277_, _08575_);
  or _61944_ (_11280_, _11279_, _11278_);
  and _61945_ (_11281_, _11280_, _06283_);
  or _61946_ (_11282_, _11281_, _11243_);
  or _61947_ (_11283_, _11282_, _11242_);
  nor _61948_ (_11284_, _05973_, _05963_);
  not _61949_ (_11285_, _11284_);
  nor _61950_ (_11286_, _06317_, _10116_);
  not _61951_ (_11287_, _11286_);
  and _61952_ (_11288_, _06317_, _10116_);
  nor _61953_ (_11289_, _11286_, _11288_);
  nor _61954_ (_11290_, _06611_, _10170_);
  and _61955_ (_11291_, _06611_, _10170_);
  nor _61956_ (_11292_, _06968_, _10135_);
  not _61957_ (_11293_, _11292_);
  and _61958_ (_11294_, _06968_, _10135_);
  nor _61959_ (_11295_, _11292_, _11294_);
  nor _61960_ (_11296_, _06213_, _06055_);
  and _61961_ (_11297_, _06213_, _06055_);
  nor _61962_ (_11298_, _06656_, _10213_);
  and _61963_ (_11299_, _06656_, _10213_);
  nor _61964_ (_11300_, _11298_, _11299_);
  nor _61965_ (_11301_, _07004_, _06042_);
  nor _61966_ (_11302_, _06251_, _06097_);
  and _61967_ (_11303_, _07004_, \oc8051_golden_model_1.ACC [1]);
  nor _61968_ (_11304_, _07004_, \oc8051_golden_model_1.ACC [1]);
  nor _61969_ (_11305_, _11304_, _11303_);
  not _61970_ (_11306_, _11305_);
  and _61971_ (_11307_, _11306_, _11302_);
  nor _61972_ (_11308_, _11307_, _11301_);
  not _61973_ (_11309_, _11308_);
  and _61974_ (_11310_, _11309_, _11300_);
  nor _61975_ (_11311_, _11310_, _11298_);
  nor _61976_ (_11312_, _11311_, _11297_);
  or _61977_ (_11313_, _11312_, _11296_);
  nand _61978_ (_11314_, _11313_, _11295_);
  and _61979_ (_11315_, _11314_, _11293_);
  nor _61980_ (_11316_, _11315_, _11291_);
  or _61981_ (_11317_, _11316_, _11290_);
  nand _61982_ (_11318_, _11317_, _11289_);
  and _61983_ (_11319_, _11318_, _11287_);
  and _61984_ (_11320_, _11319_, _10961_);
  not _61985_ (_11321_, _11243_);
  nor _61986_ (_11322_, _11319_, _10961_);
  or _61987_ (_11323_, _11322_, _11321_);
  or _61988_ (_11324_, _11323_, _11320_);
  and _61989_ (_11325_, _11324_, _11285_);
  and _61990_ (_11326_, _11325_, _11283_);
  and _61991_ (_11327_, _11284_, \oc8051_golden_model_1.ACC [6]);
  or _61992_ (_11328_, _11327_, _06568_);
  or _61993_ (_11329_, _11328_, _11326_);
  and _61994_ (_11330_, _06370_, _05779_);
  not _61995_ (_11331_, _11330_);
  or _61996_ (_11332_, _10772_, _06926_);
  and _61997_ (_11333_, _11332_, _11331_);
  and _61998_ (_11334_, _11333_, _11329_);
  nor _61999_ (_11335_, _05973_, _06567_);
  and _62000_ (_11336_, _10778_, _06097_);
  and _62001_ (_11337_, _11336_, _06055_);
  and _62002_ (_11338_, _11337_, _10135_);
  and _62003_ (_11339_, _11338_, _10170_);
  and _62004_ (_11340_, _11339_, _10116_);
  nor _62005_ (_11341_, _11340_, _08572_);
  and _62006_ (_11342_, _11340_, _08572_);
  or _62007_ (_11343_, _11342_, _11341_);
  and _62008_ (_11344_, _11343_, _11330_);
  or _62009_ (_11345_, _11344_, _11335_);
  or _62010_ (_11346_, _11345_, _11334_);
  nand _62011_ (_11347_, _11335_, _10558_);
  and _62012_ (_11348_, _11347_, _05928_);
  and _62013_ (_11349_, _11348_, _11346_);
  and _62014_ (_11350_, _10819_, _05927_);
  or _62015_ (_11351_, _11350_, _06278_);
  or _62016_ (_11352_, _11351_, _11349_);
  and _62017_ (_11353_, _06370_, _05938_);
  not _62018_ (_11354_, _11353_);
  and _62019_ (_11355_, _08550_, _07939_);
  or _62020_ (_11356_, _11355_, _10489_);
  or _62021_ (_11357_, _11356_, _06279_);
  and _62022_ (_11358_, _11357_, _11354_);
  and _62023_ (_11359_, _11358_, _11352_);
  nor _62024_ (_11360_, _05973_, _06277_);
  and _62025_ (_11361_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and _62026_ (_11362_, _11361_, \oc8051_golden_model_1.ACC [2]);
  and _62027_ (_11363_, _11362_, \oc8051_golden_model_1.ACC [3]);
  and _62028_ (_11364_, _11363_, \oc8051_golden_model_1.ACC [4]);
  and _62029_ (_11365_, _11364_, \oc8051_golden_model_1.ACC [5]);
  and _62030_ (_11366_, _11365_, \oc8051_golden_model_1.ACC [6]);
  nor _62031_ (_11367_, _11366_, _08572_);
  and _62032_ (_11368_, _11366_, _08572_);
  or _62033_ (_11369_, _11368_, _11367_);
  and _62034_ (_11370_, _11369_, _11353_);
  or _62035_ (_11371_, _11370_, _11360_);
  or _62036_ (_11372_, _11371_, _11359_);
  nand _62037_ (_11373_, _11360_, _06097_);
  and _62038_ (_11374_, _11373_, _01347_);
  and _62039_ (_11375_, _11374_, _11372_);
  or _62040_ (_11376_, _11375_, _10488_);
  and _62041_ (_40574_, _11376_, _42618_);
  not _62042_ (_11377_, \oc8051_golden_model_1.PCON [7]);
  nor _62043_ (_11378_, _01347_, _11377_);
  nor _62044_ (_11379_, _07951_, _11377_);
  not _62045_ (_11380_, _07951_);
  nor _62046_ (_11381_, _08573_, _11380_);
  or _62047_ (_11382_, _11381_, _11379_);
  and _62048_ (_11383_, _11382_, _06528_);
  and _62049_ (_11384_, _08575_, _07951_);
  or _62050_ (_11385_, _11384_, _11379_);
  and _62051_ (_11386_, _11385_, _06536_);
  and _62052_ (_11387_, _08768_, _07951_);
  or _62053_ (_11388_, _11387_, _11379_);
  or _62054_ (_11389_, _11388_, _07151_);
  and _62055_ (_11390_, _07951_, \oc8051_golden_model_1.ACC [7]);
  or _62056_ (_11391_, _11390_, _11379_);
  and _62057_ (_11392_, _11391_, _07141_);
  nor _62058_ (_11393_, _07141_, _11377_);
  or _62059_ (_11394_, _11393_, _06341_);
  or _62060_ (_11395_, _11394_, _11392_);
  and _62061_ (_11396_, _11395_, _07166_);
  and _62062_ (_11397_, _11396_, _11389_);
  nor _62063_ (_11398_, _08040_, _11380_);
  or _62064_ (_11399_, _11398_, _11379_);
  and _62065_ (_11400_, _11399_, _06461_);
  or _62066_ (_11401_, _11400_, _11397_);
  and _62067_ (_11402_, _11401_, _06465_);
  and _62068_ (_11403_, _11391_, _06464_);
  or _62069_ (_11404_, _11403_, _10080_);
  or _62070_ (_11405_, _11404_, _11402_);
  or _62071_ (_11406_, _11399_, _07215_);
  and _62072_ (_11407_, _11406_, _11405_);
  or _62073_ (_11408_, _11407_, _07460_);
  and _62074_ (_11409_, _08755_, _07951_);
  or _62075_ (_11410_, _11379_, _07208_);
  or _62076_ (_11411_, _11410_, _11409_);
  and _62077_ (_11412_, _11411_, _05982_);
  and _62078_ (_11413_, _11412_, _11408_);
  and _62079_ (_11414_, _09021_, _07951_);
  or _62080_ (_11415_, _11414_, _11379_);
  and _62081_ (_11416_, _11415_, _10094_);
  or _62082_ (_11417_, _11416_, _06218_);
  or _62083_ (_11418_, _11417_, _11413_);
  and _62084_ (_11419_, _08825_, _07951_);
  or _62085_ (_11420_, _11419_, _11379_);
  or _62086_ (_11421_, _11420_, _06219_);
  and _62087_ (_11422_, _11421_, _11418_);
  or _62088_ (_11423_, _11422_, _06369_);
  and _62089_ (_11424_, _09044_, _07951_);
  or _62090_ (_11425_, _11424_, _11379_);
  or _62091_ (_11426_, _11425_, _07237_);
  and _62092_ (_11427_, _11426_, _07240_);
  and _62093_ (_11428_, _11427_, _11423_);
  or _62094_ (_11429_, _11428_, _11386_);
  and _62095_ (_11430_, _11429_, _07242_);
  or _62096_ (_11431_, _11379_, _08043_);
  and _62097_ (_11432_, _11420_, _06375_);
  and _62098_ (_11433_, _11432_, _11431_);
  or _62099_ (_11434_, _11433_, _11430_);
  and _62100_ (_11435_, _11434_, _07234_);
  and _62101_ (_11436_, _11391_, _06545_);
  and _62102_ (_11437_, _11436_, _11431_);
  or _62103_ (_11438_, _11437_, _06366_);
  or _62104_ (_11439_, _11438_, _11435_);
  nor _62105_ (_11440_, _09043_, _11380_);
  or _62106_ (_11441_, _11379_, _09056_);
  or _62107_ (_11442_, _11441_, _11440_);
  and _62108_ (_11443_, _11442_, _09061_);
  and _62109_ (_11444_, _11443_, _11439_);
  or _62110_ (_11445_, _11444_, _11383_);
  and _62111_ (_11446_, _11445_, _06926_);
  and _62112_ (_11447_, _11388_, _06568_);
  or _62113_ (_11448_, _11447_, _06278_);
  or _62114_ (_11449_, _11448_, _11446_);
  and _62115_ (_11450_, _08550_, _07951_);
  or _62116_ (_11451_, _11379_, _06279_);
  or _62117_ (_11452_, _11451_, _11450_);
  and _62118_ (_11453_, _11452_, _01347_);
  and _62119_ (_11454_, _11453_, _11449_);
  or _62120_ (_11455_, _11454_, _11378_);
  and _62121_ (_40575_, _11455_, _42618_);
  and _62122_ (_11456_, _01351_, \oc8051_golden_model_1.TMOD [7]);
  not _62123_ (_11457_, _07914_);
  and _62124_ (_11458_, _11457_, \oc8051_golden_model_1.TMOD [7]);
  nor _62125_ (_11459_, _08573_, _11457_);
  or _62126_ (_11460_, _11459_, _11458_);
  and _62127_ (_11461_, _11460_, _06528_);
  and _62128_ (_11462_, _08575_, _07914_);
  or _62129_ (_11463_, _11462_, _11458_);
  and _62130_ (_11464_, _11463_, _06536_);
  and _62131_ (_11465_, _08768_, _07914_);
  or _62132_ (_11466_, _11465_, _11458_);
  or _62133_ (_11467_, _11466_, _07151_);
  and _62134_ (_11468_, _07914_, \oc8051_golden_model_1.ACC [7]);
  or _62135_ (_11469_, _11468_, _11458_);
  and _62136_ (_11470_, _11469_, _07141_);
  and _62137_ (_11471_, _07142_, \oc8051_golden_model_1.TMOD [7]);
  or _62138_ (_11472_, _11471_, _06341_);
  or _62139_ (_11473_, _11472_, _11470_);
  and _62140_ (_11474_, _11473_, _07166_);
  and _62141_ (_11475_, _11474_, _11467_);
  nor _62142_ (_11476_, _08040_, _11457_);
  or _62143_ (_11477_, _11476_, _11458_);
  and _62144_ (_11478_, _11477_, _06461_);
  or _62145_ (_11479_, _11478_, _11475_);
  and _62146_ (_11480_, _11479_, _06465_);
  and _62147_ (_11481_, _11469_, _06464_);
  or _62148_ (_11482_, _11481_, _10080_);
  or _62149_ (_11483_, _11482_, _11480_);
  or _62150_ (_11484_, _11477_, _07215_);
  and _62151_ (_11485_, _11484_, _11483_);
  or _62152_ (_11486_, _11485_, _07460_);
  and _62153_ (_11487_, _08755_, _07914_);
  or _62154_ (_11488_, _11458_, _07208_);
  or _62155_ (_11489_, _11488_, _11487_);
  and _62156_ (_11490_, _11489_, _05982_);
  and _62157_ (_11491_, _11490_, _11486_);
  and _62158_ (_11492_, _09021_, _07914_);
  or _62159_ (_11493_, _11492_, _11458_);
  and _62160_ (_11494_, _11493_, _10094_);
  or _62161_ (_11495_, _11494_, _06218_);
  or _62162_ (_11496_, _11495_, _11491_);
  and _62163_ (_11497_, _08825_, _07914_);
  or _62164_ (_11498_, _11497_, _11458_);
  or _62165_ (_11499_, _11498_, _06219_);
  and _62166_ (_11500_, _11499_, _11496_);
  or _62167_ (_11501_, _11500_, _06369_);
  and _62168_ (_11502_, _09044_, _07914_);
  or _62169_ (_11503_, _11502_, _11458_);
  or _62170_ (_11504_, _11503_, _07237_);
  and _62171_ (_11505_, _11504_, _07240_);
  and _62172_ (_11506_, _11505_, _11501_);
  or _62173_ (_11507_, _11506_, _11464_);
  and _62174_ (_11508_, _11507_, _07242_);
  or _62175_ (_11509_, _11458_, _08043_);
  and _62176_ (_11510_, _11498_, _06375_);
  and _62177_ (_11511_, _11510_, _11509_);
  or _62178_ (_11512_, _11511_, _11508_);
  and _62179_ (_11513_, _11512_, _07234_);
  and _62180_ (_11514_, _11469_, _06545_);
  and _62181_ (_11515_, _11514_, _11509_);
  or _62182_ (_11516_, _11515_, _06366_);
  or _62183_ (_11517_, _11516_, _11513_);
  nor _62184_ (_11518_, _09043_, _11457_);
  or _62185_ (_11519_, _11458_, _09056_);
  or _62186_ (_11520_, _11519_, _11518_);
  and _62187_ (_11521_, _11520_, _09061_);
  and _62188_ (_11522_, _11521_, _11517_);
  or _62189_ (_11523_, _11522_, _11461_);
  and _62190_ (_11524_, _11523_, _06926_);
  and _62191_ (_11525_, _11466_, _06568_);
  or _62192_ (_11526_, _11525_, _06278_);
  or _62193_ (_11527_, _11526_, _11524_);
  and _62194_ (_11528_, _08550_, _07914_);
  or _62195_ (_11529_, _11458_, _06279_);
  or _62196_ (_11530_, _11529_, _11528_);
  and _62197_ (_11531_, _11530_, _01347_);
  and _62198_ (_11532_, _11531_, _11527_);
  or _62199_ (_11533_, _11532_, _11456_);
  and _62200_ (_40576_, _11533_, _42618_);
  not _62201_ (_11534_, \oc8051_golden_model_1.DPL [7]);
  nor _62202_ (_11535_, _01347_, _11534_);
  nor _62203_ (_11536_, _07960_, _11534_);
  not _62204_ (_11537_, _07960_);
  nor _62205_ (_11538_, _08573_, _11537_);
  or _62206_ (_11539_, _11538_, _11536_);
  and _62207_ (_11540_, _11539_, _06528_);
  and _62208_ (_11541_, _08575_, _07960_);
  or _62209_ (_11542_, _11541_, _11536_);
  and _62210_ (_11543_, _11542_, _06536_);
  nor _62211_ (_11544_, _08040_, _11537_);
  or _62212_ (_11545_, _11544_, _11536_);
  or _62213_ (_11546_, _11545_, _07215_);
  and _62214_ (_11547_, _08768_, _07960_);
  or _62215_ (_11548_, _11547_, _11536_);
  or _62216_ (_11549_, _11548_, _07151_);
  and _62217_ (_11550_, _07960_, \oc8051_golden_model_1.ACC [7]);
  or _62218_ (_11551_, _11550_, _11536_);
  and _62219_ (_11552_, _11551_, _07141_);
  nor _62220_ (_11553_, _07141_, _11534_);
  or _62221_ (_11554_, _11553_, _06341_);
  or _62222_ (_11555_, _11554_, _11552_);
  and _62223_ (_11556_, _11555_, _07166_);
  and _62224_ (_11557_, _11556_, _11549_);
  and _62225_ (_11558_, _11545_, _06461_);
  or _62226_ (_11559_, _11558_, _06464_);
  or _62227_ (_11560_, _11559_, _11557_);
  nor _62228_ (_11561_, _06019_, _05973_);
  not _62229_ (_11562_, _11561_);
  or _62230_ (_11563_, _11551_, _06465_);
  and _62231_ (_11564_, _11563_, _11562_);
  and _62232_ (_11565_, _11564_, _11560_);
  and _62233_ (_11566_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and _62234_ (_11567_, _11566_, \oc8051_golden_model_1.DPL [2]);
  and _62235_ (_11568_, _11567_, \oc8051_golden_model_1.DPL [3]);
  and _62236_ (_11569_, _11568_, \oc8051_golden_model_1.DPL [4]);
  and _62237_ (_11570_, _11569_, \oc8051_golden_model_1.DPL [5]);
  and _62238_ (_11571_, _11570_, \oc8051_golden_model_1.DPL [6]);
  nor _62239_ (_11572_, _11571_, \oc8051_golden_model_1.DPL [7]);
  and _62240_ (_11573_, _11571_, \oc8051_golden_model_1.DPL [7]);
  nor _62241_ (_11574_, _11573_, _11572_);
  and _62242_ (_11575_, _11574_, _11561_);
  or _62243_ (_11576_, _11575_, _11565_);
  and _62244_ (_11577_, _11576_, _06374_);
  nor _62245_ (_11578_, _08608_, _06374_);
  or _62246_ (_11579_, _11578_, _10080_);
  or _62247_ (_11580_, _11579_, _11577_);
  and _62248_ (_11581_, _11580_, _11546_);
  or _62249_ (_11582_, _11581_, _07460_);
  and _62250_ (_11583_, _08755_, _07960_);
  or _62251_ (_11584_, _11536_, _07208_);
  or _62252_ (_11585_, _11584_, _11583_);
  and _62253_ (_11586_, _11585_, _05982_);
  and _62254_ (_11587_, _11586_, _11582_);
  and _62255_ (_11588_, _09021_, _07960_);
  or _62256_ (_11589_, _11588_, _11536_);
  and _62257_ (_11590_, _11589_, _10094_);
  or _62258_ (_11591_, _11590_, _06218_);
  or _62259_ (_11592_, _11591_, _11587_);
  and _62260_ (_11593_, _08825_, _07960_);
  or _62261_ (_11594_, _11593_, _11536_);
  or _62262_ (_11595_, _11594_, _06219_);
  and _62263_ (_11596_, _11595_, _11592_);
  or _62264_ (_11597_, _11596_, _06369_);
  and _62265_ (_11598_, _09044_, _07960_);
  or _62266_ (_11599_, _11598_, _11536_);
  or _62267_ (_11600_, _11599_, _07237_);
  and _62268_ (_11601_, _11600_, _07240_);
  and _62269_ (_11602_, _11601_, _11597_);
  or _62270_ (_11603_, _11602_, _11543_);
  and _62271_ (_11604_, _11603_, _07242_);
  or _62272_ (_11605_, _11536_, _08043_);
  and _62273_ (_11606_, _11594_, _06375_);
  and _62274_ (_11607_, _11606_, _11605_);
  or _62275_ (_11608_, _11607_, _11604_);
  and _62276_ (_11609_, _11608_, _07234_);
  and _62277_ (_11610_, _11551_, _06545_);
  and _62278_ (_11611_, _11610_, _11605_);
  or _62279_ (_11612_, _11611_, _06366_);
  or _62280_ (_11613_, _11612_, _11609_);
  nor _62281_ (_11614_, _09043_, _11537_);
  or _62282_ (_11615_, _11536_, _09056_);
  or _62283_ (_11616_, _11615_, _11614_);
  and _62284_ (_11617_, _11616_, _09061_);
  and _62285_ (_11618_, _11617_, _11613_);
  or _62286_ (_11619_, _11618_, _11540_);
  and _62287_ (_11620_, _11619_, _06926_);
  and _62288_ (_11621_, _11548_, _06568_);
  or _62289_ (_11622_, _11621_, _06278_);
  or _62290_ (_11623_, _11622_, _11620_);
  and _62291_ (_11624_, _08550_, _07960_);
  or _62292_ (_11625_, _11536_, _06279_);
  or _62293_ (_11626_, _11625_, _11624_);
  and _62294_ (_11627_, _11626_, _01347_);
  and _62295_ (_11628_, _11627_, _11623_);
  or _62296_ (_11629_, _11628_, _11535_);
  and _62297_ (_40577_, _11629_, _42618_);
  not _62298_ (_11630_, \oc8051_golden_model_1.DPH [7]);
  nor _62299_ (_11631_, _01347_, _11630_);
  nor _62300_ (_11632_, _07963_, _11630_);
  not _62301_ (_11633_, _08186_);
  nor _62302_ (_11634_, _08573_, _11633_);
  or _62303_ (_11635_, _11634_, _11632_);
  and _62304_ (_11636_, _11635_, _06528_);
  and _62305_ (_11637_, _08575_, _08186_);
  or _62306_ (_11638_, _11637_, _11632_);
  and _62307_ (_11639_, _11638_, _06536_);
  nor _62308_ (_11640_, _08040_, _11633_);
  or _62309_ (_11641_, _11640_, _11632_);
  or _62310_ (_11642_, _11641_, _07215_);
  and _62311_ (_11643_, _08768_, _08186_);
  or _62312_ (_11644_, _11643_, _11632_);
  or _62313_ (_11645_, _11644_, _07151_);
  and _62314_ (_11646_, _07963_, \oc8051_golden_model_1.ACC [7]);
  or _62315_ (_11647_, _11646_, _11632_);
  and _62316_ (_11648_, _11647_, _07141_);
  nor _62317_ (_11649_, _07141_, _11630_);
  or _62318_ (_11650_, _11649_, _06341_);
  or _62319_ (_11651_, _11650_, _11648_);
  and _62320_ (_11652_, _11651_, _07166_);
  and _62321_ (_11653_, _11652_, _11645_);
  and _62322_ (_11654_, _11641_, _06461_);
  or _62323_ (_11655_, _11654_, _06464_);
  or _62324_ (_11656_, _11655_, _11653_);
  or _62325_ (_11657_, _11647_, _06465_);
  and _62326_ (_11658_, _11657_, _11562_);
  and _62327_ (_11659_, _11658_, _11656_);
  and _62328_ (_11660_, _11573_, \oc8051_golden_model_1.DPH [0]);
  and _62329_ (_11661_, _11660_, \oc8051_golden_model_1.DPH [1]);
  and _62330_ (_11662_, _11661_, \oc8051_golden_model_1.DPH [2]);
  and _62331_ (_11663_, _11662_, \oc8051_golden_model_1.DPH [3]);
  and _62332_ (_11664_, _11663_, \oc8051_golden_model_1.DPH [4]);
  and _62333_ (_11665_, _11664_, \oc8051_golden_model_1.DPH [5]);
  and _62334_ (_11666_, _11665_, \oc8051_golden_model_1.DPH [6]);
  nor _62335_ (_11667_, _11666_, _11630_);
  and _62336_ (_11668_, _11666_, _11630_);
  or _62337_ (_11669_, _11668_, _11667_);
  and _62338_ (_11670_, _11669_, _11561_);
  or _62339_ (_11671_, _11670_, _11659_);
  and _62340_ (_11672_, _11671_, _06374_);
  and _62341_ (_11673_, _06373_, _06182_);
  or _62342_ (_11674_, _11673_, _10080_);
  or _62343_ (_11675_, _11674_, _11672_);
  and _62344_ (_11676_, _11675_, _11642_);
  or _62345_ (_11677_, _11676_, _07460_);
  or _62346_ (_11678_, _11632_, _07208_);
  and _62347_ (_11679_, _08755_, _07963_);
  or _62348_ (_11680_, _11679_, _11678_);
  and _62349_ (_11681_, _11680_, _05982_);
  and _62350_ (_11682_, _11681_, _11677_);
  and _62351_ (_11683_, _09021_, _07963_);
  or _62352_ (_11684_, _11683_, _11632_);
  and _62353_ (_11685_, _11684_, _10094_);
  or _62354_ (_11686_, _11685_, _06218_);
  or _62355_ (_11687_, _11686_, _11682_);
  and _62356_ (_11688_, _08825_, _07963_);
  or _62357_ (_11689_, _11688_, _11632_);
  or _62358_ (_11690_, _11689_, _06219_);
  and _62359_ (_11691_, _11690_, _11687_);
  or _62360_ (_11692_, _11691_, _06369_);
  and _62361_ (_11693_, _09044_, _07963_);
  or _62362_ (_11694_, _11693_, _11632_);
  or _62363_ (_11695_, _11694_, _07237_);
  and _62364_ (_11696_, _11695_, _07240_);
  and _62365_ (_11697_, _11696_, _11692_);
  or _62366_ (_11698_, _11697_, _11639_);
  and _62367_ (_11699_, _11698_, _07242_);
  or _62368_ (_11700_, _11632_, _08043_);
  and _62369_ (_11701_, _11689_, _06375_);
  and _62370_ (_11702_, _11701_, _11700_);
  or _62371_ (_11703_, _11702_, _11699_);
  and _62372_ (_11704_, _11703_, _07234_);
  and _62373_ (_11705_, _11647_, _06545_);
  and _62374_ (_11706_, _11705_, _11700_);
  or _62375_ (_11707_, _11706_, _06366_);
  or _62376_ (_11708_, _11707_, _11704_);
  nor _62377_ (_11709_, _09043_, _11633_);
  or _62378_ (_11710_, _11632_, _09056_);
  or _62379_ (_11711_, _11710_, _11709_);
  and _62380_ (_11712_, _11711_, _09061_);
  and _62381_ (_11713_, _11712_, _11708_);
  or _62382_ (_11714_, _11713_, _11636_);
  and _62383_ (_11715_, _11714_, _06926_);
  and _62384_ (_11716_, _11644_, _06568_);
  or _62385_ (_11717_, _11716_, _06278_);
  or _62386_ (_11718_, _11717_, _11715_);
  and _62387_ (_11719_, _08550_, _08186_);
  or _62388_ (_11720_, _11632_, _06279_);
  or _62389_ (_11721_, _11720_, _11719_);
  and _62390_ (_11722_, _11721_, _01347_);
  and _62391_ (_11723_, _11722_, _11718_);
  or _62392_ (_11724_, _11723_, _11631_);
  and _62393_ (_40580_, _11724_, _42618_);
  and _62394_ (_11725_, _01351_, \oc8051_golden_model_1.TL1 [7]);
  not _62395_ (_11726_, _07968_);
  and _62396_ (_11727_, _11726_, \oc8051_golden_model_1.TL1 [7]);
  nor _62397_ (_11728_, _08573_, _11726_);
  or _62398_ (_11729_, _11728_, _11727_);
  and _62399_ (_11730_, _11729_, _06528_);
  and _62400_ (_11731_, _08575_, _07968_);
  or _62401_ (_11732_, _11731_, _11727_);
  and _62402_ (_11733_, _11732_, _06536_);
  and _62403_ (_11734_, _08768_, _07968_);
  or _62404_ (_11735_, _11734_, _11727_);
  or _62405_ (_11736_, _11735_, _07151_);
  and _62406_ (_11737_, _07968_, \oc8051_golden_model_1.ACC [7]);
  or _62407_ (_11738_, _11737_, _11727_);
  and _62408_ (_11739_, _11738_, _07141_);
  and _62409_ (_11740_, _07142_, \oc8051_golden_model_1.TL1 [7]);
  or _62410_ (_11741_, _11740_, _06341_);
  or _62411_ (_11742_, _11741_, _11739_);
  and _62412_ (_11743_, _11742_, _07166_);
  and _62413_ (_11744_, _11743_, _11736_);
  nor _62414_ (_11745_, _08040_, _11726_);
  or _62415_ (_11746_, _11745_, _11727_);
  and _62416_ (_11747_, _11746_, _06461_);
  or _62417_ (_11748_, _11747_, _11744_);
  and _62418_ (_11749_, _11748_, _06465_);
  and _62419_ (_11750_, _11738_, _06464_);
  or _62420_ (_11751_, _11750_, _10080_);
  or _62421_ (_11752_, _11751_, _11749_);
  or _62422_ (_11753_, _11746_, _07215_);
  and _62423_ (_11754_, _11753_, _11752_);
  or _62424_ (_11755_, _11754_, _07460_);
  and _62425_ (_11756_, _08755_, _07968_);
  or _62426_ (_11757_, _11727_, _07208_);
  or _62427_ (_11758_, _11757_, _11756_);
  and _62428_ (_11759_, _11758_, _05982_);
  and _62429_ (_11760_, _11759_, _11755_);
  and _62430_ (_11761_, _09021_, _07968_);
  or _62431_ (_11762_, _11761_, _11727_);
  and _62432_ (_11763_, _11762_, _10094_);
  or _62433_ (_11764_, _11763_, _06218_);
  or _62434_ (_11765_, _11764_, _11760_);
  and _62435_ (_11766_, _08825_, _07968_);
  or _62436_ (_11767_, _11766_, _11727_);
  or _62437_ (_11768_, _11767_, _06219_);
  and _62438_ (_11769_, _11768_, _11765_);
  or _62439_ (_11770_, _11769_, _06369_);
  and _62440_ (_11771_, _09044_, _07968_);
  or _62441_ (_11772_, _11771_, _11727_);
  or _62442_ (_11773_, _11772_, _07237_);
  and _62443_ (_11774_, _11773_, _07240_);
  and _62444_ (_11775_, _11774_, _11770_);
  or _62445_ (_11776_, _11775_, _11733_);
  and _62446_ (_11777_, _11776_, _07242_);
  or _62447_ (_11778_, _11727_, _08043_);
  and _62448_ (_11779_, _11767_, _06375_);
  and _62449_ (_11780_, _11779_, _11778_);
  or _62450_ (_11781_, _11780_, _11777_);
  and _62451_ (_11782_, _11781_, _07234_);
  and _62452_ (_11783_, _11738_, _06545_);
  and _62453_ (_11784_, _11783_, _11778_);
  or _62454_ (_11785_, _11784_, _06366_);
  or _62455_ (_11786_, _11785_, _11782_);
  nor _62456_ (_11787_, _09043_, _11726_);
  or _62457_ (_11788_, _11727_, _09056_);
  or _62458_ (_11789_, _11788_, _11787_);
  and _62459_ (_11790_, _11789_, _09061_);
  and _62460_ (_11791_, _11790_, _11786_);
  or _62461_ (_11792_, _11791_, _11730_);
  and _62462_ (_11793_, _11792_, _06926_);
  and _62463_ (_11794_, _11735_, _06568_);
  or _62464_ (_11795_, _11794_, _06278_);
  or _62465_ (_11796_, _11795_, _11793_);
  and _62466_ (_11797_, _08550_, _07968_);
  or _62467_ (_11798_, _11727_, _06279_);
  or _62468_ (_11799_, _11798_, _11797_);
  and _62469_ (_11800_, _11799_, _01347_);
  and _62470_ (_11801_, _11800_, _11796_);
  or _62471_ (_11802_, _11801_, _11725_);
  and _62472_ (_40581_, _11802_, _42618_);
  and _62473_ (_11803_, _01351_, \oc8051_golden_model_1.TL0 [7]);
  not _62474_ (_11804_, _07919_);
  and _62475_ (_11805_, _11804_, \oc8051_golden_model_1.TL0 [7]);
  nor _62476_ (_11806_, _08573_, _11804_);
  or _62477_ (_11807_, _11806_, _11805_);
  and _62478_ (_11808_, _11807_, _06528_);
  and _62479_ (_11809_, _08575_, _07919_);
  or _62480_ (_11810_, _11809_, _11805_);
  and _62481_ (_11811_, _11810_, _06536_);
  nor _62482_ (_11812_, _08040_, _11804_);
  or _62483_ (_11813_, _11812_, _11805_);
  or _62484_ (_11814_, _11813_, _07215_);
  and _62485_ (_11815_, _08768_, _07919_);
  or _62486_ (_11816_, _11815_, _11805_);
  or _62487_ (_11817_, _11816_, _07151_);
  and _62488_ (_11818_, _07919_, \oc8051_golden_model_1.ACC [7]);
  or _62489_ (_11819_, _11818_, _11805_);
  and _62490_ (_11820_, _11819_, _07141_);
  and _62491_ (_11821_, _07142_, \oc8051_golden_model_1.TL0 [7]);
  or _62492_ (_11822_, _11821_, _06341_);
  or _62493_ (_11823_, _11822_, _11820_);
  and _62494_ (_11824_, _11823_, _07166_);
  and _62495_ (_11825_, _11824_, _11817_);
  and _62496_ (_11826_, _11813_, _06461_);
  or _62497_ (_11827_, _11826_, _11825_);
  and _62498_ (_11828_, _11827_, _06465_);
  and _62499_ (_11829_, _11819_, _06464_);
  or _62500_ (_11830_, _11829_, _10080_);
  or _62501_ (_11831_, _11830_, _11828_);
  and _62502_ (_11832_, _11831_, _11814_);
  or _62503_ (_11833_, _11832_, _07460_);
  and _62504_ (_11834_, _08755_, _07919_);
  or _62505_ (_11835_, _11805_, _07208_);
  or _62506_ (_11836_, _11835_, _11834_);
  and _62507_ (_11837_, _11836_, _05982_);
  and _62508_ (_11838_, _11837_, _11833_);
  and _62509_ (_11839_, _09021_, _07919_);
  or _62510_ (_11840_, _11839_, _11805_);
  and _62511_ (_11841_, _11840_, _10094_);
  or _62512_ (_11842_, _11841_, _06218_);
  or _62513_ (_11843_, _11842_, _11838_);
  and _62514_ (_11844_, _08825_, _07919_);
  or _62515_ (_11845_, _11844_, _11805_);
  or _62516_ (_11846_, _11845_, _06219_);
  and _62517_ (_11847_, _11846_, _11843_);
  or _62518_ (_11848_, _11847_, _06369_);
  and _62519_ (_11849_, _09044_, _07919_);
  or _62520_ (_11850_, _11849_, _11805_);
  or _62521_ (_11851_, _11850_, _07237_);
  and _62522_ (_11852_, _11851_, _07240_);
  and _62523_ (_11853_, _11852_, _11848_);
  or _62524_ (_11854_, _11853_, _11811_);
  and _62525_ (_11855_, _11854_, _07242_);
  or _62526_ (_11856_, _11805_, _08043_);
  and _62527_ (_11857_, _11845_, _06375_);
  and _62528_ (_11858_, _11857_, _11856_);
  or _62529_ (_11859_, _11858_, _11855_);
  and _62530_ (_11860_, _11859_, _07234_);
  and _62531_ (_11861_, _11819_, _06545_);
  and _62532_ (_11862_, _11861_, _11856_);
  or _62533_ (_11863_, _11862_, _06366_);
  or _62534_ (_11864_, _11863_, _11860_);
  nor _62535_ (_11865_, _09043_, _11804_);
  or _62536_ (_11866_, _11805_, _09056_);
  or _62537_ (_11867_, _11866_, _11865_);
  and _62538_ (_11868_, _11867_, _09061_);
  and _62539_ (_11869_, _11868_, _11864_);
  or _62540_ (_11870_, _11869_, _11808_);
  and _62541_ (_11871_, _11870_, _06926_);
  and _62542_ (_11872_, _11816_, _06568_);
  or _62543_ (_11873_, _11872_, _06278_);
  or _62544_ (_11874_, _11873_, _11871_);
  and _62545_ (_11875_, _08550_, _07919_);
  or _62546_ (_11876_, _11805_, _06279_);
  or _62547_ (_11877_, _11876_, _11875_);
  and _62548_ (_11878_, _11877_, _01347_);
  and _62549_ (_11879_, _11878_, _11874_);
  or _62550_ (_11880_, _11879_, _11803_);
  and _62551_ (_40582_, _11880_, _42618_);
  and _62552_ (_11881_, _01351_, \oc8051_golden_model_1.TCON [7]);
  not _62553_ (_11882_, _07928_);
  and _62554_ (_11883_, _11882_, \oc8051_golden_model_1.TCON [7]);
  and _62555_ (_11884_, _08575_, _07928_);
  or _62556_ (_11885_, _11884_, _11883_);
  and _62557_ (_11886_, _11885_, _06536_);
  nor _62558_ (_11887_, _08040_, _11882_);
  or _62559_ (_11888_, _11887_, _11883_);
  or _62560_ (_11889_, _11888_, _07215_);
  not _62561_ (_11890_, _08616_);
  and _62562_ (_11891_, _11890_, \oc8051_golden_model_1.TCON [7]);
  and _62563_ (_11892_, _08649_, _08616_);
  or _62564_ (_11893_, _11892_, _11891_);
  and _62565_ (_11894_, _11893_, _06268_);
  and _62566_ (_11895_, _08768_, _07928_);
  or _62567_ (_11896_, _11895_, _11883_);
  or _62568_ (_11897_, _11896_, _07151_);
  and _62569_ (_11898_, _07928_, \oc8051_golden_model_1.ACC [7]);
  or _62570_ (_11899_, _11898_, _11883_);
  and _62571_ (_11900_, _11899_, _07141_);
  and _62572_ (_11901_, _07142_, \oc8051_golden_model_1.TCON [7]);
  or _62573_ (_11902_, _11901_, _06341_);
  or _62574_ (_11903_, _11902_, _11900_);
  and _62575_ (_11904_, _11903_, _06273_);
  and _62576_ (_11905_, _11904_, _11897_);
  and _62577_ (_11906_, _08773_, _08616_);
  or _62578_ (_11907_, _11906_, _11891_);
  and _62579_ (_11908_, _11907_, _06272_);
  or _62580_ (_11909_, _11908_, _06461_);
  or _62581_ (_11910_, _11909_, _11905_);
  or _62582_ (_11911_, _11888_, _07166_);
  and _62583_ (_11912_, _11911_, _11910_);
  or _62584_ (_11913_, _11912_, _06464_);
  or _62585_ (_11914_, _11899_, _06465_);
  and _62586_ (_11915_, _11914_, _06269_);
  and _62587_ (_11916_, _11915_, _11913_);
  or _62588_ (_11917_, _11916_, _11894_);
  and _62589_ (_11918_, _11917_, _06262_);
  and _62590_ (_11919_, _08790_, _08616_);
  or _62591_ (_11920_, _11919_, _11891_);
  and _62592_ (_11921_, _11920_, _06261_);
  or _62593_ (_11922_, _11921_, _11918_);
  and _62594_ (_11923_, _11922_, _06258_);
  and _62595_ (_11924_, _08808_, _08616_);
  or _62596_ (_11925_, _11924_, _11891_);
  and _62597_ (_11926_, _11925_, _06257_);
  or _62598_ (_11927_, _11926_, _10080_);
  or _62599_ (_11928_, _11927_, _11923_);
  and _62600_ (_11929_, _11928_, _11889_);
  or _62601_ (_11930_, _11929_, _07460_);
  and _62602_ (_11931_, _08755_, _07928_);
  or _62603_ (_11932_, _11883_, _07208_);
  or _62604_ (_11933_, _11932_, _11931_);
  and _62605_ (_11934_, _11933_, _05982_);
  and _62606_ (_11935_, _11934_, _11930_);
  and _62607_ (_11936_, _09021_, _07928_);
  or _62608_ (_11937_, _11936_, _11883_);
  and _62609_ (_11938_, _11937_, _10094_);
  or _62610_ (_11939_, _11938_, _06218_);
  or _62611_ (_11940_, _11939_, _11935_);
  and _62612_ (_11941_, _08825_, _07928_);
  or _62613_ (_11942_, _11941_, _11883_);
  or _62614_ (_11943_, _11942_, _06219_);
  and _62615_ (_11944_, _11943_, _11940_);
  or _62616_ (_11945_, _11944_, _06369_);
  and _62617_ (_11946_, _09044_, _07928_);
  or _62618_ (_11947_, _11946_, _11883_);
  or _62619_ (_11948_, _11947_, _07237_);
  and _62620_ (_11949_, _11948_, _07240_);
  and _62621_ (_11950_, _11949_, _11945_);
  or _62622_ (_11951_, _11950_, _11886_);
  and _62623_ (_11952_, _11951_, _07242_);
  or _62624_ (_11953_, _11883_, _08043_);
  and _62625_ (_11954_, _11942_, _06375_);
  and _62626_ (_11955_, _11954_, _11953_);
  or _62627_ (_11956_, _11955_, _11952_);
  and _62628_ (_11957_, _11956_, _07234_);
  and _62629_ (_11958_, _11899_, _06545_);
  and _62630_ (_11959_, _11958_, _11953_);
  or _62631_ (_11960_, _11959_, _06366_);
  or _62632_ (_11961_, _11960_, _11957_);
  nor _62633_ (_11962_, _09043_, _11882_);
  or _62634_ (_11963_, _11883_, _09056_);
  or _62635_ (_11964_, _11963_, _11962_);
  and _62636_ (_11965_, _11964_, _09061_);
  and _62637_ (_11966_, _11965_, _11961_);
  nor _62638_ (_11967_, _08573_, _11882_);
  or _62639_ (_11968_, _11967_, _11883_);
  and _62640_ (_11969_, _11968_, _06528_);
  or _62641_ (_11970_, _11969_, _06568_);
  or _62642_ (_11971_, _11970_, _11966_);
  or _62643_ (_11972_, _11896_, _06926_);
  and _62644_ (_11973_, _11972_, _05928_);
  and _62645_ (_11974_, _11973_, _11971_);
  and _62646_ (_11975_, _11893_, _05927_);
  or _62647_ (_11976_, _11975_, _06278_);
  or _62648_ (_11977_, _11976_, _11974_);
  and _62649_ (_11978_, _08550_, _07928_);
  or _62650_ (_11979_, _11883_, _06279_);
  or _62651_ (_11980_, _11979_, _11978_);
  and _62652_ (_11981_, _11980_, _01347_);
  and _62653_ (_11982_, _11981_, _11977_);
  or _62654_ (_11983_, _11982_, _11881_);
  and _62655_ (_40583_, _11983_, _42618_);
  and _62656_ (_11984_, _01351_, \oc8051_golden_model_1.TH1 [7]);
  not _62657_ (_11985_, _07910_);
  and _62658_ (_11986_, _11985_, \oc8051_golden_model_1.TH1 [7]);
  nor _62659_ (_11987_, _08573_, _11985_);
  or _62660_ (_11988_, _11987_, _11986_);
  and _62661_ (_11989_, _11988_, _06528_);
  and _62662_ (_11990_, _08575_, _07910_);
  or _62663_ (_11991_, _11990_, _11986_);
  and _62664_ (_11992_, _11991_, _06536_);
  nor _62665_ (_11993_, _08040_, _11985_);
  or _62666_ (_11994_, _11993_, _11986_);
  or _62667_ (_11995_, _11994_, _07215_);
  and _62668_ (_11996_, _08768_, _07910_);
  or _62669_ (_11997_, _11996_, _11986_);
  or _62670_ (_11998_, _11997_, _07151_);
  and _62671_ (_11999_, _07910_, \oc8051_golden_model_1.ACC [7]);
  or _62672_ (_12000_, _11999_, _11986_);
  and _62673_ (_12001_, _12000_, _07141_);
  and _62674_ (_12002_, _07142_, \oc8051_golden_model_1.TH1 [7]);
  or _62675_ (_12003_, _12002_, _06341_);
  or _62676_ (_12004_, _12003_, _12001_);
  and _62677_ (_12005_, _12004_, _07166_);
  and _62678_ (_12006_, _12005_, _11998_);
  and _62679_ (_12007_, _11994_, _06461_);
  or _62680_ (_12008_, _12007_, _12006_);
  and _62681_ (_12009_, _12008_, _06465_);
  and _62682_ (_12010_, _12000_, _06464_);
  or _62683_ (_12011_, _12010_, _10080_);
  or _62684_ (_12012_, _12011_, _12009_);
  and _62685_ (_12013_, _12012_, _11995_);
  or _62686_ (_12014_, _12013_, _07460_);
  and _62687_ (_12015_, _08755_, _07910_);
  or _62688_ (_12016_, _11986_, _07208_);
  or _62689_ (_12017_, _12016_, _12015_);
  and _62690_ (_12018_, _12017_, _05982_);
  and _62691_ (_12019_, _12018_, _12014_);
  and _62692_ (_12020_, _09021_, _07910_);
  or _62693_ (_12021_, _12020_, _11986_);
  and _62694_ (_12022_, _12021_, _10094_);
  or _62695_ (_12023_, _12022_, _06218_);
  or _62696_ (_12024_, _12023_, _12019_);
  and _62697_ (_12025_, _08825_, _07910_);
  or _62698_ (_12026_, _12025_, _11986_);
  or _62699_ (_12027_, _12026_, _06219_);
  and _62700_ (_12028_, _12027_, _12024_);
  or _62701_ (_12029_, _12028_, _06369_);
  and _62702_ (_12030_, _09044_, _07910_);
  or _62703_ (_12031_, _12030_, _11986_);
  or _62704_ (_12032_, _12031_, _07237_);
  and _62705_ (_12033_, _12032_, _07240_);
  and _62706_ (_12034_, _12033_, _12029_);
  or _62707_ (_12035_, _12034_, _11992_);
  and _62708_ (_12036_, _12035_, _07242_);
  or _62709_ (_12037_, _11986_, _08043_);
  and _62710_ (_12038_, _12026_, _06375_);
  and _62711_ (_12039_, _12038_, _12037_);
  or _62712_ (_12040_, _12039_, _12036_);
  and _62713_ (_12041_, _12040_, _07234_);
  and _62714_ (_12042_, _12000_, _06545_);
  and _62715_ (_12043_, _12042_, _12037_);
  or _62716_ (_12044_, _12043_, _06366_);
  or _62717_ (_12045_, _12044_, _12041_);
  nor _62718_ (_12046_, _09043_, _11985_);
  or _62719_ (_12047_, _11986_, _09056_);
  or _62720_ (_12048_, _12047_, _12046_);
  and _62721_ (_12049_, _12048_, _09061_);
  and _62722_ (_12050_, _12049_, _12045_);
  or _62723_ (_12051_, _12050_, _11989_);
  and _62724_ (_12052_, _12051_, _06926_);
  and _62725_ (_12053_, _11997_, _06568_);
  or _62726_ (_12054_, _12053_, _06278_);
  or _62727_ (_12055_, _12054_, _12052_);
  and _62728_ (_12056_, _08550_, _07910_);
  or _62729_ (_12057_, _11986_, _06279_);
  or _62730_ (_12058_, _12057_, _12056_);
  and _62731_ (_12059_, _12058_, _01347_);
  and _62732_ (_12060_, _12059_, _12055_);
  or _62733_ (_12061_, _12060_, _11984_);
  and _62734_ (_40584_, _12061_, _42618_);
  and _62735_ (_12062_, _01351_, \oc8051_golden_model_1.TH0 [7]);
  not _62736_ (_12063_, _07922_);
  and _62737_ (_12064_, _12063_, \oc8051_golden_model_1.TH0 [7]);
  nor _62738_ (_12065_, _08573_, _12063_);
  or _62739_ (_12066_, _12065_, _12064_);
  and _62740_ (_12067_, _12066_, _06528_);
  and _62741_ (_12068_, _08575_, _07922_);
  or _62742_ (_12069_, _12068_, _12064_);
  and _62743_ (_12070_, _12069_, _06536_);
  nor _62744_ (_12071_, _08040_, _12063_);
  or _62745_ (_12072_, _12071_, _12064_);
  or _62746_ (_12073_, _12072_, _07215_);
  and _62747_ (_12074_, _08768_, _07922_);
  or _62748_ (_12075_, _12074_, _12064_);
  or _62749_ (_12076_, _12075_, _07151_);
  and _62750_ (_12077_, _07922_, \oc8051_golden_model_1.ACC [7]);
  or _62751_ (_12078_, _12077_, _12064_);
  and _62752_ (_12079_, _12078_, _07141_);
  and _62753_ (_12080_, _07142_, \oc8051_golden_model_1.TH0 [7]);
  or _62754_ (_12081_, _12080_, _06341_);
  or _62755_ (_12082_, _12081_, _12079_);
  and _62756_ (_12083_, _12082_, _07166_);
  and _62757_ (_12084_, _12083_, _12076_);
  and _62758_ (_12085_, _12072_, _06461_);
  or _62759_ (_12086_, _12085_, _12084_);
  and _62760_ (_12087_, _12086_, _06465_);
  and _62761_ (_12088_, _12078_, _06464_);
  or _62762_ (_12089_, _12088_, _10080_);
  or _62763_ (_12090_, _12089_, _12087_);
  and _62764_ (_12091_, _12090_, _12073_);
  or _62765_ (_12092_, _12091_, _07460_);
  and _62766_ (_12093_, _08755_, _07922_);
  or _62767_ (_12094_, _12064_, _07208_);
  or _62768_ (_12095_, _12094_, _12093_);
  and _62769_ (_12096_, _12095_, _05982_);
  and _62770_ (_12097_, _12096_, _12092_);
  and _62771_ (_12098_, _09021_, _07922_);
  or _62772_ (_12099_, _12098_, _12064_);
  and _62773_ (_12100_, _12099_, _10094_);
  or _62774_ (_12101_, _12100_, _06218_);
  or _62775_ (_12102_, _12101_, _12097_);
  and _62776_ (_12103_, _08825_, _07922_);
  or _62777_ (_12104_, _12103_, _12064_);
  or _62778_ (_12105_, _12104_, _06219_);
  and _62779_ (_12106_, _12105_, _12102_);
  or _62780_ (_12107_, _12106_, _06369_);
  and _62781_ (_12108_, _09044_, _07922_);
  or _62782_ (_12109_, _12108_, _12064_);
  or _62783_ (_12110_, _12109_, _07237_);
  and _62784_ (_12111_, _12110_, _07240_);
  and _62785_ (_12112_, _12111_, _12107_);
  or _62786_ (_12113_, _12112_, _12070_);
  and _62787_ (_12114_, _12113_, _07242_);
  or _62788_ (_12115_, _12064_, _08043_);
  and _62789_ (_12116_, _12104_, _06375_);
  and _62790_ (_12117_, _12116_, _12115_);
  or _62791_ (_12118_, _12117_, _12114_);
  and _62792_ (_12119_, _12118_, _07234_);
  and _62793_ (_12120_, _12078_, _06545_);
  and _62794_ (_12121_, _12120_, _12115_);
  or _62795_ (_12122_, _12121_, _06366_);
  or _62796_ (_12123_, _12122_, _12119_);
  nor _62797_ (_12124_, _09043_, _12063_);
  or _62798_ (_12125_, _12064_, _09056_);
  or _62799_ (_12126_, _12125_, _12124_);
  and _62800_ (_12127_, _12126_, _09061_);
  and _62801_ (_12128_, _12127_, _12123_);
  or _62802_ (_12129_, _12128_, _12067_);
  and _62803_ (_12130_, _12129_, _06926_);
  and _62804_ (_12131_, _12075_, _06568_);
  or _62805_ (_12132_, _12131_, _06278_);
  or _62806_ (_12133_, _12132_, _12130_);
  and _62807_ (_12134_, _08550_, _07922_);
  or _62808_ (_12135_, _12064_, _06279_);
  or _62809_ (_12136_, _12135_, _12134_);
  and _62810_ (_12137_, _12136_, _01347_);
  and _62811_ (_12138_, _12137_, _12133_);
  or _62812_ (_12139_, _12138_, _12062_);
  and _62813_ (_40585_, _12139_, _42618_);
  not _62814_ (_12140_, _06379_);
  nor _62815_ (_12141_, _11360_, _11353_);
  not _62816_ (_12142_, _05616_);
  and _62817_ (_12143_, _09409_, _12142_);
  and _62818_ (_12144_, _12143_, _09472_);
  and _62819_ (_12145_, _12144_, _09469_);
  and _62820_ (_12146_, _12145_, \oc8051_golden_model_1.PC [14]);
  and _62821_ (_12147_, _12146_, _09468_);
  nor _62822_ (_12148_, _12146_, _09468_);
  or _62823_ (_12149_, _12148_, _12147_);
  nor _62824_ (_12150_, _12149_, _12141_);
  and _62825_ (_12151_, _11203_, _11157_);
  nor _62826_ (_12152_, _12151_, _12149_);
  nor _62827_ (_12153_, _11097_, _06540_);
  and _62828_ (_12154_, _11069_, _11037_);
  nor _62829_ (_12155_, _12154_, _12149_);
  not _62830_ (_12156_, _07042_);
  and _62831_ (_12157_, _10998_, _12156_);
  nor _62832_ (_12158_, _11008_, _07040_);
  not _62833_ (_12159_, _12158_);
  or _62834_ (_12160_, _12159_, _11012_);
  nor _62835_ (_12161_, _12160_, _11011_);
  and _62836_ (_12162_, _12161_, _12157_);
  nor _62837_ (_12163_, _12162_, _12149_);
  nor _62838_ (_12164_, _10496_, _06542_);
  nor _62839_ (_12165_, _12149_, _10979_);
  nor _62840_ (_12166_, _10954_, _06533_);
  nor _62841_ (_12167_, _07482_, _05954_);
  nor _62842_ (_12168_, _12167_, _10509_);
  and _62843_ (_12169_, _12168_, _10940_);
  nor _62844_ (_12170_, _12169_, _12149_);
  nor _62845_ (_12171_, _09487_, _09030_);
  nor _62846_ (_12172_, _10093_, _05974_);
  nor _62847_ (_12173_, _09479_, _05982_);
  nor _62848_ (_12174_, _06006_, _05973_);
  not _62849_ (_12175_, _12174_);
  not _62850_ (_12176_, _06371_);
  not _62851_ (_12177_, _06347_);
  and _62852_ (_12178_, _09412_, \oc8051_golden_model_1.PC [8]);
  and _62853_ (_12179_, _12178_, \oc8051_golden_model_1.PC [9]);
  and _62854_ (_12180_, _12179_, \oc8051_golden_model_1.PC [10]);
  and _62855_ (_12181_, _12180_, \oc8051_golden_model_1.PC [11]);
  and _62856_ (_12182_, _12181_, \oc8051_golden_model_1.PC [12]);
  and _62857_ (_12183_, _12182_, \oc8051_golden_model_1.PC [13]);
  and _62858_ (_12184_, _12183_, \oc8051_golden_model_1.PC [14]);
  nor _62859_ (_12185_, _12183_, \oc8051_golden_model_1.PC [14]);
  nor _62860_ (_12186_, _12185_, _12184_);
  not _62861_ (_12187_, _12186_);
  nor _62862_ (_12188_, _12187_, _08608_);
  and _62863_ (_12189_, _12187_, _08608_);
  nor _62864_ (_12190_, _12189_, _12188_);
  not _62865_ (_12191_, _12190_);
  nor _62866_ (_12192_, _12182_, \oc8051_golden_model_1.PC [13]);
  nor _62867_ (_12193_, _12192_, _12183_);
  not _62868_ (_12194_, _12193_);
  nor _62869_ (_12195_, _12194_, _08608_);
  and _62870_ (_12196_, _12194_, _08608_);
  nor _62871_ (_12197_, _12181_, \oc8051_golden_model_1.PC [12]);
  nor _62872_ (_12198_, _12197_, _12182_);
  not _62873_ (_12199_, _12198_);
  nor _62874_ (_12200_, _12199_, _08608_);
  nor _62875_ (_12201_, _12179_, \oc8051_golden_model_1.PC [10]);
  nor _62876_ (_12202_, _12201_, _12180_);
  not _62877_ (_12203_, _12202_);
  nor _62878_ (_12204_, _12203_, _08608_);
  not _62879_ (_12205_, _12204_);
  nor _62880_ (_12206_, _12180_, \oc8051_golden_model_1.PC [11]);
  nor _62881_ (_12207_, _12206_, _12181_);
  not _62882_ (_12208_, _12207_);
  nor _62883_ (_12209_, _12208_, _08608_);
  and _62884_ (_12210_, _12208_, _08608_);
  nor _62885_ (_12211_, _12210_, _12209_);
  and _62886_ (_12212_, _12203_, _08608_);
  nor _62887_ (_12213_, _12212_, _12204_);
  and _62888_ (_12214_, _12213_, _12211_);
  nor _62889_ (_12215_, _12178_, \oc8051_golden_model_1.PC [9]);
  nor _62890_ (_12216_, _12215_, _12179_);
  not _62891_ (_12217_, _12216_);
  nor _62892_ (_12218_, _12217_, _08608_);
  and _62893_ (_12219_, _12217_, _08608_);
  nor _62894_ (_12220_, _12219_, _12218_);
  nor _62895_ (_12221_, _09416_, _08608_);
  and _62896_ (_12222_, _09416_, _08608_);
  and _62897_ (_12223_, _09411_, _08656_);
  nor _62898_ (_12224_, _12223_, \oc8051_golden_model_1.PC [6]);
  nor _62899_ (_12225_, _12224_, _09413_);
  not _62900_ (_12226_, _12225_);
  nor _62901_ (_12227_, _12226_, _08857_);
  and _62902_ (_12228_, _12226_, _08857_);
  nor _62903_ (_12229_, _12228_, _12227_);
  not _62904_ (_12230_, _12229_);
  and _62905_ (_12231_, _09411_, \oc8051_golden_model_1.PC [4]);
  nor _62906_ (_12232_, _12231_, \oc8051_golden_model_1.PC [5]);
  nor _62907_ (_12233_, _12232_, _12223_);
  not _62908_ (_12234_, _12233_);
  nor _62909_ (_12235_, _12234_, _08926_);
  and _62910_ (_12236_, _12234_, _08926_);
  nor _62911_ (_12237_, _09411_, \oc8051_golden_model_1.PC [4]);
  nor _62912_ (_12238_, _12237_, _12231_);
  not _62913_ (_12239_, _12238_);
  nor _62914_ (_12240_, _12239_, _08892_);
  nor _62915_ (_12241_, _09410_, \oc8051_golden_model_1.PC [3]);
  nor _62916_ (_12242_, _12241_, _09411_);
  not _62917_ (_12243_, _12242_);
  nor _62918_ (_12244_, _12243_, _06452_);
  and _62919_ (_12245_, _12243_, _06452_);
  nor _62920_ (_12246_, _05634_, \oc8051_golden_model_1.PC [2]);
  nor _62921_ (_12247_, _12246_, _09410_);
  not _62922_ (_12248_, _12247_);
  nor _62923_ (_12249_, _12248_, _06697_);
  nor _62924_ (_12250_, _07038_, _06111_);
  nor _62925_ (_12251_, _06872_, \oc8051_golden_model_1.PC [0]);
  and _62926_ (_12252_, _07038_, _06111_);
  nor _62927_ (_12253_, _12252_, _12250_);
  and _62928_ (_12254_, _12253_, _12251_);
  nor _62929_ (_12255_, _12254_, _12250_);
  and _62930_ (_12256_, _12248_, _06697_);
  nor _62931_ (_12257_, _12256_, _12249_);
  not _62932_ (_12258_, _12257_);
  nor _62933_ (_12259_, _12258_, _12255_);
  nor _62934_ (_12260_, _12259_, _12249_);
  nor _62935_ (_12261_, _12260_, _12245_);
  nor _62936_ (_12262_, _12261_, _12244_);
  and _62937_ (_12263_, _12239_, _08892_);
  nor _62938_ (_12264_, _12263_, _12240_);
  not _62939_ (_12265_, _12264_);
  nor _62940_ (_12266_, _12265_, _12262_);
  nor _62941_ (_12267_, _12266_, _12240_);
  nor _62942_ (_12268_, _12267_, _12236_);
  nor _62943_ (_12269_, _12268_, _12235_);
  nor _62944_ (_12270_, _12269_, _12230_);
  nor _62945_ (_12271_, _12270_, _12227_);
  nor _62946_ (_12272_, _12271_, _12222_);
  or _62947_ (_12273_, _12272_, _12221_);
  nor _62948_ (_12274_, _09412_, \oc8051_golden_model_1.PC [8]);
  nor _62949_ (_12275_, _12274_, _12178_);
  not _62950_ (_12276_, _12275_);
  nor _62951_ (_12277_, _12276_, _08608_);
  and _62952_ (_12278_, _12276_, _08608_);
  nor _62953_ (_12279_, _12278_, _12277_);
  and _62954_ (_12280_, _12279_, _12273_);
  and _62955_ (_12281_, _12280_, _12220_);
  and _62956_ (_12282_, _12281_, _12214_);
  nor _62957_ (_12283_, _12277_, _12218_);
  not _62958_ (_12284_, _12283_);
  and _62959_ (_12285_, _12284_, _12214_);
  or _62960_ (_12286_, _12285_, _12209_);
  nor _62961_ (_12287_, _12286_, _12282_);
  and _62962_ (_12288_, _12287_, _12205_);
  and _62963_ (_12289_, _12199_, _08608_);
  nor _62964_ (_12290_, _12289_, _12200_);
  not _62965_ (_12291_, _12290_);
  nor _62966_ (_12292_, _12291_, _12288_);
  nor _62967_ (_12293_, _12292_, _12200_);
  nor _62968_ (_12294_, _12293_, _12196_);
  nor _62969_ (_12295_, _12294_, _12195_);
  nor _62970_ (_12296_, _12295_, _12191_);
  nor _62971_ (_12297_, _12296_, _12188_);
  and _62972_ (_12298_, _09479_, _08608_);
  nor _62973_ (_12299_, _09479_, _08608_);
  nor _62974_ (_12300_, _12299_, _12298_);
  and _62975_ (_12301_, _12300_, _12297_);
  nor _62976_ (_12302_, _12300_, _12297_);
  nor _62977_ (_12303_, _12302_, _12301_);
  nor _62978_ (_12304_, _08755_, _06286_);
  nor _62979_ (_12305_, _12304_, _08802_);
  or _62980_ (_12306_, _09446_, _06317_);
  or _62981_ (_12307_, _09122_, _07607_);
  and _62982_ (_12308_, _12307_, _12306_);
  and _62983_ (_12309_, _12308_, _12305_);
  or _62984_ (_12310_, _09167_, _07896_);
  or _62985_ (_12311_, _09447_, _06611_);
  and _62986_ (_12312_, _12311_, _12310_);
  or _62987_ (_12313_, _09212_, _07883_);
  or _62988_ (_12314_, _09448_, _06968_);
  and _62989_ (_12315_, _12314_, _12313_);
  and _62990_ (_12316_, _12315_, _12312_);
  and _62991_ (_12317_, _12316_, _12309_);
  or _62992_ (_12318_, _09449_, _06213_);
  or _62993_ (_12319_, _09257_, _06473_);
  and _62994_ (_12320_, _12319_, _12318_);
  or _62995_ (_12321_, _09450_, _06656_);
  or _62996_ (_12322_, _09302_, _06657_);
  and _62997_ (_12323_, _12322_, _12321_);
  and _62998_ (_12324_, _12323_, _12320_);
  or _62999_ (_12325_, _09451_, _07004_);
  or _63000_ (_12326_, _09347_, _07005_);
  and _63001_ (_12327_, _12326_, _12325_);
  or _63002_ (_12328_, _09392_, _06251_);
  nand _63003_ (_12329_, _09392_, _06251_);
  and _63004_ (_12330_, _12329_, _12328_);
  and _63005_ (_12331_, _12330_, _12327_);
  and _63006_ (_12332_, _12331_, _12324_);
  and _63007_ (_12333_, _12332_, _12317_);
  or _63008_ (_12334_, _12333_, _12303_);
  nand _63009_ (_12335_, _12332_, _12317_);
  or _63010_ (_12336_, _12335_, _09479_);
  nand _63011_ (_12337_, _12336_, _12334_);
  nor _63012_ (_12338_, _12337_, _12177_);
  not _63013_ (_12339_, _08041_);
  and _63014_ (_12340_, _08040_, _06182_);
  nor _63015_ (_12341_, _12340_, _12339_);
  nor _63016_ (_12342_, _08142_, _07607_);
  and _63017_ (_12343_, _08142_, _07607_);
  nor _63018_ (_12344_, _12343_, _12342_);
  and _63019_ (_12345_, _12344_, _12341_);
  or _63020_ (_12346_, _08244_, _07896_);
  and _63021_ (_12347_, _08244_, _07896_);
  not _63022_ (_12348_, _12347_);
  and _63023_ (_12349_, _12348_, _12346_);
  and _63024_ (_12350_, _08541_, _07883_);
  nor _63025_ (_12351_, _08541_, _07883_);
  nor _63026_ (_12352_, _12351_, _12350_);
  and _63027_ (_12353_, _12352_, _12349_);
  and _63028_ (_12354_, _12353_, _12345_);
  and _63029_ (_12355_, _07594_, _06473_);
  and _63030_ (_12356_, _07776_, _06657_);
  nor _63031_ (_12357_, _12356_, _12355_);
  or _63032_ (_12358_, _07594_, _06473_);
  or _63033_ (_12359_, _07776_, _06657_);
  and _63034_ (_12360_, _12359_, _12358_);
  and _63035_ (_12361_, _12360_, _12357_);
  or _63036_ (_12362_, _07357_, _07005_);
  and _63037_ (_12363_, _07357_, _07005_);
  not _63038_ (_12364_, _12363_);
  and _63039_ (_12365_, _12364_, _12362_);
  nand _63040_ (_12366_, _07133_, _06251_);
  or _63041_ (_12367_, _07133_, _06251_);
  and _63042_ (_12368_, _12367_, _12366_);
  and _63043_ (_12369_, _12368_, _12365_);
  and _63044_ (_12370_, _12369_, _12361_);
  and _63045_ (_12371_, _12370_, _12354_);
  nand _63046_ (_12372_, _12371_, _09479_);
  and _63047_ (_12373_, _07209_, _06260_);
  not _63048_ (_12374_, _12373_);
  not _63049_ (_12375_, _06357_);
  nor _63050_ (_12376_, _07211_, _06006_);
  nor _63051_ (_12377_, _12376_, _12375_);
  and _63052_ (_12378_, _12377_, _12374_);
  not _63053_ (_12379_, _12378_);
  not _63054_ (_12380_, _12303_);
  or _63055_ (_12381_, _12371_, _12380_);
  and _63056_ (_12382_, _12381_, _12379_);
  and _63057_ (_12383_, _12382_, _12372_);
  and _63058_ (_12384_, _09487_, _06464_);
  not _63059_ (_12385_, _12149_);
  and _63060_ (_12386_, _12385_, _07154_);
  not _63061_ (_12387_, _08654_);
  not _63062_ (_12388_, _09487_);
  and _63063_ (_12389_, _08142_, _08040_);
  and _63064_ (_12390_, _12389_, _08553_);
  and _63065_ (_12391_, _07357_, _07133_);
  and _63066_ (_12392_, _12391_, _08554_);
  nand _63067_ (_12393_, _12392_, _12390_);
  or _63068_ (_12394_, _12393_, _12388_);
  and _63069_ (_12395_, _08659_, \oc8051_golden_model_1.PC [8]);
  and _63070_ (_12396_, _12395_, \oc8051_golden_model_1.PC [9]);
  and _63071_ (_12397_, _12396_, \oc8051_golden_model_1.PC [10]);
  and _63072_ (_12398_, _12397_, \oc8051_golden_model_1.PC [11]);
  and _63073_ (_12399_, _12398_, \oc8051_golden_model_1.PC [12]);
  and _63074_ (_12400_, _12399_, \oc8051_golden_model_1.PC [13]);
  and _63075_ (_12401_, _12400_, \oc8051_golden_model_1.PC [14]);
  nor _63076_ (_12402_, _12400_, \oc8051_golden_model_1.PC [14]);
  nor _63077_ (_12403_, _12402_, _12401_);
  and _63078_ (_12404_, _12403_, _06182_);
  nor _63079_ (_12405_, _12403_, _06182_);
  nor _63080_ (_12406_, _12405_, _12404_);
  not _63081_ (_12407_, _12406_);
  nor _63082_ (_12408_, _12399_, \oc8051_golden_model_1.PC [13]);
  nor _63083_ (_12409_, _12408_, _12400_);
  nor _63084_ (_12410_, _12409_, _06182_);
  and _63085_ (_12411_, _12409_, _06182_);
  not _63086_ (_12412_, _12411_);
  nor _63087_ (_12413_, _12398_, \oc8051_golden_model_1.PC [12]);
  nor _63088_ (_12414_, _12413_, _12399_);
  and _63089_ (_12415_, _12414_, _06182_);
  nor _63090_ (_12416_, _12397_, \oc8051_golden_model_1.PC [11]);
  nor _63091_ (_12417_, _12416_, _12398_);
  and _63092_ (_12418_, _12417_, _06182_);
  nor _63093_ (_12419_, _12417_, _06182_);
  nor _63094_ (_12420_, _12396_, \oc8051_golden_model_1.PC [10]);
  nor _63095_ (_12421_, _12420_, _12397_);
  and _63096_ (_12422_, _12421_, _06182_);
  nor _63097_ (_12423_, _12421_, _06182_);
  nor _63098_ (_12424_, _12423_, _12422_);
  nor _63099_ (_12425_, _12395_, \oc8051_golden_model_1.PC [9]);
  nor _63100_ (_12426_, _12425_, _12396_);
  nor _63101_ (_12427_, _12426_, _06182_);
  and _63102_ (_12428_, _12426_, _06182_);
  not _63103_ (_12429_, _12428_);
  nor _63104_ (_12430_, _08659_, \oc8051_golden_model_1.PC [8]);
  nor _63105_ (_12431_, _12430_, _12395_);
  and _63106_ (_12432_, _12431_, _06182_);
  and _63107_ (_12433_, _08661_, _06182_);
  nor _63108_ (_12434_, _08661_, _06182_);
  nor _63109_ (_12435_, _12434_, _12433_);
  not _63110_ (_12436_, _12435_);
  and _63111_ (_12437_, _08656_, _05929_);
  nor _63112_ (_12438_, _12437_, \oc8051_golden_model_1.PC [6]);
  nor _63113_ (_12439_, _12438_, _08658_);
  not _63114_ (_12440_, _12439_);
  nor _63115_ (_12441_, _12440_, _06317_);
  and _63116_ (_12442_, _12440_, _06317_);
  nor _63117_ (_12443_, _12442_, _12441_);
  and _63118_ (_12444_, _05929_, \oc8051_golden_model_1.PC [4]);
  nor _63119_ (_12445_, _12444_, \oc8051_golden_model_1.PC [5]);
  nor _63120_ (_12446_, _12445_, _12437_);
  not _63121_ (_12447_, _12446_);
  nor _63122_ (_12448_, _12447_, _06611_);
  and _63123_ (_12449_, _12447_, _06611_);
  nor _63124_ (_12450_, _05929_, \oc8051_golden_model_1.PC [4]);
  nor _63125_ (_12451_, _12450_, _12444_);
  not _63126_ (_12452_, _12451_);
  nor _63127_ (_12453_, _12452_, _06968_);
  nor _63128_ (_12454_, _06213_, _06033_);
  and _63129_ (_12455_, _06213_, _06033_);
  nor _63130_ (_12456_, _06656_, _06085_);
  nor _63131_ (_12457_, _07004_, \oc8051_golden_model_1.PC [1]);
  nor _63132_ (_12458_, _06251_, _05630_);
  and _63133_ (_12459_, _07004_, \oc8051_golden_model_1.PC [1]);
  nor _63134_ (_12460_, _12459_, _12457_);
  and _63135_ (_12461_, _12460_, _12458_);
  nor _63136_ (_12462_, _12461_, _12457_);
  and _63137_ (_12463_, _06656_, _06085_);
  nor _63138_ (_12464_, _12463_, _12456_);
  not _63139_ (_12465_, _12464_);
  nor _63140_ (_12466_, _12465_, _12462_);
  nor _63141_ (_12467_, _12466_, _12456_);
  nor _63142_ (_12468_, _12467_, _12455_);
  nor _63143_ (_12469_, _12468_, _12454_);
  and _63144_ (_12470_, _12452_, _06968_);
  nor _63145_ (_12471_, _12470_, _12453_);
  not _63146_ (_12472_, _12471_);
  nor _63147_ (_12473_, _12472_, _12469_);
  nor _63148_ (_12474_, _12473_, _12453_);
  nor _63149_ (_12475_, _12474_, _12449_);
  or _63150_ (_12476_, _12475_, _12448_);
  and _63151_ (_12477_, _12476_, _12443_);
  nor _63152_ (_12478_, _12477_, _12441_);
  nor _63153_ (_12479_, _12478_, _12436_);
  nor _63154_ (_12480_, _12479_, _12433_);
  nor _63155_ (_12481_, _12431_, _06182_);
  nor _63156_ (_12482_, _12481_, _12432_);
  not _63157_ (_12483_, _12482_);
  nor _63158_ (_12484_, _12483_, _12480_);
  nor _63159_ (_12485_, _12484_, _12432_);
  and _63160_ (_12486_, _12485_, _12429_);
  or _63161_ (_12487_, _12486_, _12427_);
  not _63162_ (_12488_, _12487_);
  and _63163_ (_12489_, _12488_, _12424_);
  nor _63164_ (_12490_, _12489_, _12422_);
  nor _63165_ (_12491_, _12490_, _12419_);
  or _63166_ (_12492_, _12491_, _12418_);
  nor _63167_ (_12493_, _12414_, _06182_);
  nor _63168_ (_12494_, _12493_, _12415_);
  and _63169_ (_12495_, _12494_, _12492_);
  nor _63170_ (_12496_, _12495_, _12415_);
  and _63171_ (_12497_, _12496_, _12412_);
  or _63172_ (_12498_, _12497_, _12410_);
  nor _63173_ (_12499_, _12498_, _12407_);
  nor _63174_ (_12500_, _12499_, _12404_);
  nor _63175_ (_12501_, _09487_, _06182_);
  and _63176_ (_12502_, _09487_, _06182_);
  nor _63177_ (_12503_, _12502_, _12501_);
  and _63178_ (_12504_, _12503_, _12500_);
  nor _63179_ (_12505_, _12503_, _12500_);
  nor _63180_ (_12506_, _12505_, _12504_);
  and _63181_ (_12507_, _12392_, _12390_);
  or _63182_ (_12508_, _12507_, _12506_);
  nand _63183_ (_12509_, _12508_, _12394_);
  nand _63184_ (_12510_, _12509_, _12387_);
  nor _63185_ (_12511_, _10758_, _10768_);
  and _63186_ (_12512_, _12511_, _10755_);
  nor _63187_ (_12513_, _07486_, _06781_);
  and _63188_ (_12514_, _12513_, _12512_);
  or _63189_ (_12515_, _12514_, _12149_);
  not _63190_ (_12516_, _12512_);
  nor _63191_ (_12517_, _07141_, _06758_);
  or _63192_ (_12518_, _12517_, _09487_);
  nor _63193_ (_12519_, _07141_, \oc8051_golden_model_1.PC [15]);
  and _63194_ (_12520_, _12519_, _07504_);
  nand _63195_ (_12521_, _12520_, _12513_);
  and _63196_ (_12522_, _12521_, _12518_);
  or _63197_ (_12523_, _12522_, _12516_);
  and _63198_ (_12524_, _12523_, _08654_);
  and _63199_ (_12525_, _12524_, _12515_);
  nor _63200_ (_12526_, _12525_, _07154_);
  and _63201_ (_12527_, _12526_, _12510_);
  nor _63202_ (_12528_, _12527_, _12386_);
  and _63203_ (_12529_, _12528_, _07151_);
  and _63204_ (_12530_, _08390_, _08340_);
  and _63205_ (_12531_, _08762_, _12530_);
  and _63206_ (_12532_, _08144_, _08042_);
  and _63207_ (_12533_, _12532_, _08759_);
  nand _63208_ (_12534_, _12533_, _12531_);
  or _63209_ (_12535_, _12534_, _09478_);
  and _63210_ (_12536_, _12533_, _12531_);
  or _63211_ (_12537_, _12536_, _12380_);
  and _63212_ (_12538_, _12537_, _12535_);
  and _63213_ (_12539_, _12538_, _06341_);
  nor _63214_ (_12540_, _06009_, _05973_);
  nor _63215_ (_12541_, _12540_, _10775_);
  not _63216_ (_12542_, _12541_);
  or _63217_ (_12543_, _12542_, _12539_);
  or _63218_ (_12544_, _12543_, _12529_);
  and _63219_ (_12545_, _06466_, _06010_);
  not _63220_ (_12546_, _12545_);
  nor _63221_ (_12547_, _12541_, _12149_);
  nor _63222_ (_12548_, _12547_, _12546_);
  nand _63223_ (_12549_, _12548_, _12544_);
  and _63224_ (_12550_, _10743_, _07175_);
  not _63225_ (_12551_, _12550_);
  nor _63226_ (_12552_, _12545_, _12388_);
  nor _63227_ (_12553_, _12552_, _12551_);
  nand _63228_ (_12554_, _12553_, _12549_);
  nor _63229_ (_12555_, _12550_, _12149_);
  nor _63230_ (_12556_, _12555_, _06464_);
  and _63231_ (_12557_, _12556_, _12554_);
  or _63232_ (_12558_, _12557_, _12384_);
  nor _63233_ (_12559_, _06012_, _05973_);
  nor _63234_ (_12560_, _12559_, _10811_);
  nand _63235_ (_12561_, _12560_, _12558_);
  nor _63236_ (_12562_, _12560_, _12385_);
  not _63237_ (_12563_, _06013_);
  nor _63238_ (_12564_, _06267_, _12563_);
  and _63239_ (_12565_, _12564_, _06269_);
  not _63240_ (_12566_, _12565_);
  nor _63241_ (_12567_, _12566_, _12562_);
  nand _63242_ (_12568_, _12567_, _12561_);
  nor _63243_ (_12569_, _12565_, _09487_);
  not _63244_ (_12570_, _12569_);
  and _63245_ (_12571_, _12570_, _12378_);
  and _63246_ (_12572_, _12571_, _12568_);
  or _63247_ (_12573_, _12572_, _12383_);
  nor _63248_ (_12574_, _12573_, _06347_);
  or _63249_ (_12575_, _12574_, _06480_);
  nor _63250_ (_12576_, _12575_, _12338_);
  nor _63251_ (_12577_, _11256_, _11255_);
  nor _63252_ (_12578_, _12577_, _11259_);
  not _63253_ (_12579_, _11262_);
  nor _63254_ (_12580_, _08390_, \oc8051_golden_model_1.ACC [0]);
  or _63255_ (_12581_, _12580_, _11263_);
  and _63256_ (_12582_, _12581_, _12579_);
  and _63257_ (_12583_, _12582_, _12578_);
  nor _63258_ (_12584_, _11250_, _11254_);
  nor _63259_ (_12585_, _11247_, _08575_);
  and _63260_ (_12586_, _12585_, _12584_);
  and _63261_ (_12587_, _12586_, _12583_);
  nor _63262_ (_12588_, _12587_, _12303_);
  and _63263_ (_12589_, _12587_, _09478_);
  nor _63264_ (_12590_, _12589_, _12588_);
  nor _63265_ (_12591_, _12590_, _06774_);
  or _63266_ (_12592_, _12591_, _12576_);
  nand _63267_ (_12593_, _12592_, _12176_);
  nor _63268_ (_12594_, _11296_, _11297_);
  nor _63269_ (_12595_, _12594_, _11300_);
  and _63270_ (_12596_, _06251_, _06097_);
  nor _63271_ (_12597_, _12596_, _11302_);
  nor _63272_ (_12598_, _11306_, _12597_);
  and _63273_ (_12599_, _12598_, _12595_);
  nor _63274_ (_12600_, _11290_, _11291_);
  nor _63275_ (_12601_, _12600_, _11295_);
  nor _63276_ (_12602_, _11289_, _10961_);
  and _63277_ (_12603_, _12602_, _12601_);
  and _63278_ (_12604_, _12603_, _12599_);
  nand _63279_ (_12605_, _12604_, _09478_);
  or _63280_ (_12606_, _12604_, _12303_);
  and _63281_ (_12607_, _12606_, _12605_);
  or _63282_ (_12608_, _12607_, _12176_);
  nand _63283_ (_12609_, _12608_, _12593_);
  nand _63284_ (_12610_, _12609_, _12175_);
  and _63285_ (_12611_, _12174_, _12149_);
  not _63286_ (_12612_, _12611_);
  not _63287_ (_12613_, _06007_);
  nor _63288_ (_12614_, _06261_, _12613_);
  nor _63289_ (_12615_, _06355_, _06019_);
  nor _63290_ (_12616_, _07399_, _12615_);
  and _63291_ (_12617_, _12616_, _12614_);
  not _63292_ (_12618_, _06492_);
  nor _63293_ (_12619_, _06495_, _06455_);
  and _63294_ (_12620_, _12619_, _12618_);
  nor _63295_ (_12621_, _07197_, _07398_);
  and _63296_ (_12622_, _12621_, _12620_);
  and _63297_ (_12623_, _12622_, _12617_);
  and _63298_ (_12624_, _12623_, _12612_);
  nand _63299_ (_12625_, _12624_, _12610_);
  nor _63300_ (_12626_, _12623_, _09487_);
  nor _63301_ (_12627_, _06019_, _05981_);
  not _63302_ (_12628_, _12627_);
  nor _63303_ (_12629_, _11561_, _09531_);
  and _63304_ (_12630_, _12629_, _12628_);
  not _63305_ (_12631_, _12630_);
  nor _63306_ (_12632_, _12631_, _12626_);
  nand _63307_ (_12633_, _12632_, _12625_);
  nor _63308_ (_12634_, _12630_, _12385_);
  and _63309_ (_12635_, _06506_, _06020_);
  not _63310_ (_12636_, _12635_);
  nor _63311_ (_12637_, _12636_, _12634_);
  and _63312_ (_12638_, _12637_, _12633_);
  and _63313_ (_12639_, _10735_, _10588_);
  or _63314_ (_12640_, _12635_, _09487_);
  nand _63315_ (_12641_, _12640_, _12639_);
  or _63316_ (_12642_, _12641_, _12638_);
  nor _63317_ (_12643_, _10516_, _06512_);
  not _63318_ (_12644_, _12643_);
  nor _63319_ (_12645_, _12639_, _12385_);
  nor _63320_ (_12646_, _12645_, _12644_);
  nand _63321_ (_12647_, _12646_, _12642_);
  nor _63322_ (_12648_, _12643_, _09487_);
  nor _63323_ (_12649_, _12648_, _10515_);
  nand _63324_ (_12650_, _12649_, _12647_);
  nor _63325_ (_12651_, _12385_, _05984_);
  nor _63326_ (_12652_, _06257_, _06254_);
  not _63327_ (_12653_, _12652_);
  nor _63328_ (_12654_, _12653_, _12651_);
  nand _63329_ (_12655_, _12654_, _12650_);
  nor _63330_ (_12656_, _12652_, _09487_);
  nor _63331_ (_12657_, _12656_, _06373_);
  nand _63332_ (_12658_, _12657_, _12655_);
  not _63333_ (_12659_, _07216_);
  and _63334_ (_12660_, _09478_, _06373_);
  nor _63335_ (_12661_, _12660_, _12659_);
  nand _63336_ (_12662_, _12661_, _12658_);
  nor _63337_ (_12663_, _09487_, _07216_);
  nor _63338_ (_12664_, _12663_, _10094_);
  and _63339_ (_12665_, _12664_, _12662_);
  or _63340_ (_12666_, _12665_, _12173_);
  nand _63341_ (_12667_, _12666_, _12172_);
  not _63342_ (_12668_, _05946_);
  nor _63343_ (_12669_, _06323_, _12668_);
  not _63344_ (_12670_, _12669_);
  nor _63345_ (_12671_, _12172_, _12385_);
  nor _63346_ (_12672_, _12671_, _12670_);
  nand _63347_ (_12673_, _12672_, _12667_);
  and _63348_ (_12674_, _05944_, _05926_);
  nor _63349_ (_12675_, _12669_, _09487_);
  nor _63350_ (_12676_, _12675_, _12674_);
  nand _63351_ (_12678_, _12676_, _12673_);
  not _63352_ (_12679_, _12674_);
  nor _63353_ (_12680_, _12679_, _12506_);
  nor _63354_ (_12681_, _12680_, _09031_);
  and _63355_ (_12682_, _12681_, _12678_);
  or _63356_ (_12683_, _12682_, _12171_);
  nand _63357_ (_12684_, _12683_, _06219_);
  and _63358_ (_12685_, _09479_, _06218_);
  nor _63359_ (_12686_, _12685_, _10929_);
  and _63360_ (_12687_, _12686_, _12684_);
  and _63361_ (_12688_, _10929_, _09487_);
  or _63362_ (_12689_, _12688_, _12687_);
  nor _63363_ (_12690_, _05973_, _05951_);
  not _63364_ (_12691_, _12690_);
  nand _63365_ (_12692_, _12691_, _12689_);
  not _63366_ (_12693_, \oc8051_golden_model_1.DPH [0]);
  and _63367_ (_12694_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor _63368_ (_12695_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and _63369_ (_12696_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _63370_ (_12697_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _63371_ (_12699_, _12697_, _12696_);
  not _63372_ (_12700_, _12699_);
  and _63373_ (_12701_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _63374_ (_12702_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _63375_ (_12703_, _12702_, _12701_);
  not _63376_ (_12704_, _12703_);
  and _63377_ (_12705_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _63378_ (_12706_, _06001_, _05997_);
  nor _63379_ (_12707_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _63380_ (_12708_, _12707_, _12705_);
  not _63381_ (_12709_, _12708_);
  nor _63382_ (_12710_, _12709_, _12706_);
  nor _63383_ (_12711_, _12710_, _12705_);
  nor _63384_ (_12712_, _12711_, _12704_);
  nor _63385_ (_12713_, _12712_, _12701_);
  nor _63386_ (_12714_, _12713_, _12700_);
  nor _63387_ (_12715_, _12714_, _12696_);
  nor _63388_ (_12716_, _12715_, _12695_);
  nor _63389_ (_12717_, _12716_, _12694_);
  nor _63390_ (_12718_, _12717_, _12693_);
  and _63391_ (_12719_, _12718_, \oc8051_golden_model_1.DPH [1]);
  and _63392_ (_12720_, _12719_, \oc8051_golden_model_1.DPH [2]);
  and _63393_ (_12721_, _12720_, \oc8051_golden_model_1.DPH [3]);
  and _63394_ (_12722_, _12721_, \oc8051_golden_model_1.DPH [4]);
  and _63395_ (_12723_, _12722_, \oc8051_golden_model_1.DPH [5]);
  and _63396_ (_12724_, _12723_, \oc8051_golden_model_1.DPH [6]);
  and _63397_ (_12725_, _12724_, \oc8051_golden_model_1.DPH [7]);
  nor _63398_ (_12726_, _12724_, \oc8051_golden_model_1.DPH [7]);
  nor _63399_ (_12727_, _12726_, _12725_);
  and _63400_ (_12728_, _12727_, _12690_);
  nor _63401_ (_12729_, _06322_, _06217_);
  not _63402_ (_12730_, _12729_);
  nor _63403_ (_12731_, _12730_, _12728_);
  nand _63404_ (_12732_, _12731_, _12692_);
  and _63405_ (_12733_, _06321_, _05926_);
  nor _63406_ (_12734_, _12729_, _09487_);
  nor _63407_ (_12735_, _12734_, _12733_);
  nand _63408_ (_12736_, _12735_, _12732_);
  not _63409_ (_12737_, _12169_);
  and _63410_ (_12738_, _11342_, _09487_);
  nor _63411_ (_12739_, _12506_, _11342_);
  or _63412_ (_12740_, _12739_, _12738_);
  and _63413_ (_12741_, _12740_, _12733_);
  nor _63414_ (_12742_, _12741_, _12737_);
  and _63415_ (_12743_, _12742_, _12736_);
  or _63416_ (_12744_, _12743_, _12170_);
  nand _63417_ (_12745_, _12744_, _12166_);
  nor _63418_ (_12746_, _12166_, _09487_);
  nor _63419_ (_12747_, _12746_, _06369_);
  nand _63420_ (_12748_, _12747_, _12745_);
  and _63421_ (_12749_, _09478_, _06369_);
  not _63422_ (_12750_, _05955_);
  nor _63423_ (_12751_, _06536_, _12750_);
  not _63424_ (_12752_, _12751_);
  nor _63425_ (_12753_, _12752_, _12749_);
  nand _63426_ (_12754_, _12753_, _12748_);
  and _63427_ (_12755_, _06535_, _05926_);
  nor _63428_ (_12756_, _12751_, _09487_);
  nor _63429_ (_12757_, _12756_, _12755_);
  nand _63430_ (_12758_, _12757_, _12754_);
  not _63431_ (_12759_, _11342_);
  and _63432_ (_12760_, _12759_, _09487_);
  nor _63433_ (_12761_, _12506_, _12759_);
  or _63434_ (_12762_, _12761_, _12760_);
  and _63435_ (_12763_, _12762_, _12755_);
  nor _63436_ (_12764_, _12763_, _10980_);
  and _63437_ (_12765_, _12764_, _12758_);
  or _63438_ (_12766_, _12765_, _12165_);
  nand _63439_ (_12767_, _12766_, _12164_);
  nor _63440_ (_12768_, _12164_, _09487_);
  nor _63441_ (_12769_, _12768_, _06375_);
  nand _63442_ (_12770_, _12769_, _12767_);
  and _63443_ (_12771_, _09478_, _06375_);
  nor _63444_ (_12772_, _06545_, _07233_);
  not _63445_ (_12773_, _12772_);
  nor _63446_ (_12774_, _12773_, _12771_);
  nand _63447_ (_12775_, _12774_, _12770_);
  and _63448_ (_12776_, _06544_, _05926_);
  nor _63449_ (_12777_, _12772_, _09487_);
  nor _63450_ (_12778_, _12777_, _12776_);
  nand _63451_ (_12779_, _12778_, _12775_);
  not _63452_ (_12780_, _12162_);
  and _63453_ (_12781_, _12506_, _10558_);
  not _63454_ (_12782_, _12776_);
  nor _63455_ (_12783_, _09487_, _10558_);
  nor _63456_ (_12784_, _12783_, _12782_);
  not _63457_ (_12785_, _12784_);
  nor _63458_ (_12786_, _12785_, _12781_);
  nor _63459_ (_12787_, _12786_, _12780_);
  and _63460_ (_12788_, _12787_, _12779_);
  or _63461_ (_12789_, _12788_, _12163_);
  nand _63462_ (_12790_, _12789_, _11022_);
  nor _63463_ (_12791_, _11022_, _09487_);
  nor _63464_ (_12792_, _12791_, _06366_);
  nand _63465_ (_12793_, _12792_, _12790_);
  and _63466_ (_12794_, _09478_, _06366_);
  not _63467_ (_12795_, _05966_);
  nor _63468_ (_12796_, _06528_, _12795_);
  not _63469_ (_12797_, _12796_);
  nor _63470_ (_12798_, _12797_, _12794_);
  nand _63471_ (_12799_, _12798_, _12793_);
  and _63472_ (_12800_, _06527_, _05926_);
  nor _63473_ (_12801_, _12796_, _09487_);
  nor _63474_ (_12802_, _12801_, _12800_);
  nand _63475_ (_12803_, _12802_, _12799_);
  not _63476_ (_12804_, _12154_);
  and _63477_ (_12805_, _09487_, _10558_);
  nor _63478_ (_12806_, _12506_, _10558_);
  or _63479_ (_12807_, _12806_, _12805_);
  and _63480_ (_12808_, _12807_, _12800_);
  nor _63481_ (_12809_, _12808_, _12804_);
  and _63482_ (_12810_, _12809_, _12803_);
  or _63483_ (_12811_, _12810_, _12155_);
  nand _63484_ (_12812_, _12811_, _12153_);
  nor _63485_ (_12813_, _12153_, _09487_);
  nor _63486_ (_12814_, _12813_, _11125_);
  and _63487_ (_12815_, _12814_, _12812_);
  and _63488_ (_12816_, _12149_, _11125_);
  or _63489_ (_12817_, _12816_, _06551_);
  nor _63490_ (_12818_, _12817_, _12815_);
  and _63491_ (_12819_, _08040_, _06551_);
  or _63492_ (_12820_, _12819_, _12818_);
  nand _63493_ (_12821_, _12820_, _05959_);
  nor _63494_ (_12822_, _09487_, _05959_);
  nor _63495_ (_12823_, _12822_, _06365_);
  nand _63496_ (_12824_, _12823_, _12821_);
  not _63497_ (_12825_, _07959_);
  and _63498_ (_12826_, _07948_, \oc8051_golden_model_1.P0 [2]);
  and _63499_ (_12827_, _08616_, \oc8051_golden_model_1.TCON [2]);
  and _63500_ (_12828_, _08620_, \oc8051_golden_model_1.P1 [2]);
  and _63501_ (_12829_, _08622_, \oc8051_golden_model_1.SCON [2]);
  and _63502_ (_12830_, _08624_, \oc8051_golden_model_1.P2 [2]);
  and _63503_ (_12831_, _08626_, \oc8051_golden_model_1.IE [2]);
  and _63504_ (_12832_, _08628_, \oc8051_golden_model_1.P3 [2]);
  and _63505_ (_12833_, _08632_, \oc8051_golden_model_1.IP [2]);
  and _63506_ (_12834_, _08630_, \oc8051_golden_model_1.PSW [2]);
  and _63507_ (_12835_, _08636_, \oc8051_golden_model_1.ACC [2]);
  and _63508_ (_12836_, _08634_, \oc8051_golden_model_1.B [2]);
  or _63509_ (_12837_, _12836_, _12835_);
  or _63510_ (_12838_, _12837_, _12834_);
  or _63511_ (_12839_, _12838_, _12833_);
  or _63512_ (_12840_, _12839_, _12832_);
  or _63513_ (_12841_, _12840_, _12831_);
  or _63514_ (_12842_, _12841_, _12830_);
  or _63515_ (_12843_, _12842_, _12829_);
  or _63516_ (_12844_, _12843_, _12828_);
  or _63517_ (_12845_, _12844_, _12827_);
  nor _63518_ (_12846_, _12845_, _12826_);
  and _63519_ (_12847_, _12846_, _08438_);
  nor _63520_ (_12848_, _12847_, _12825_);
  not _63521_ (_12849_, _08172_);
  and _63522_ (_12850_, _07948_, \oc8051_golden_model_1.P0 [1]);
  and _63523_ (_12851_, _08616_, \oc8051_golden_model_1.TCON [1]);
  and _63524_ (_12852_, _08620_, \oc8051_golden_model_1.P1 [1]);
  and _63525_ (_12853_, _08622_, \oc8051_golden_model_1.SCON [1]);
  and _63526_ (_12854_, _08624_, \oc8051_golden_model_1.P2 [1]);
  and _63527_ (_12855_, _08626_, \oc8051_golden_model_1.IE [1]);
  and _63528_ (_12856_, _08628_, \oc8051_golden_model_1.P3 [1]);
  and _63529_ (_12857_, _08632_, \oc8051_golden_model_1.IP [1]);
  and _63530_ (_12858_, _08630_, \oc8051_golden_model_1.PSW [1]);
  and _63531_ (_12859_, _08636_, \oc8051_golden_model_1.ACC [1]);
  and _63532_ (_12860_, _08634_, \oc8051_golden_model_1.B [1]);
  or _63533_ (_12861_, _12860_, _12859_);
  or _63534_ (_12862_, _12861_, _12858_);
  or _63535_ (_12863_, _12862_, _12857_);
  or _63536_ (_12864_, _12863_, _12856_);
  or _63537_ (_12865_, _12864_, _12855_);
  or _63538_ (_12866_, _12865_, _12854_);
  or _63539_ (_12867_, _12866_, _12853_);
  or _63540_ (_12868_, _12867_, _12852_);
  or _63541_ (_12869_, _12868_, _12851_);
  nor _63542_ (_12870_, _12869_, _12850_);
  and _63543_ (_12871_, _12870_, _08339_);
  nor _63544_ (_12872_, _12871_, _12849_);
  nor _63545_ (_12873_, _12872_, _12848_);
  and _63546_ (_12874_, _08628_, \oc8051_golden_model_1.P3 [4]);
  and _63547_ (_12875_, _08626_, \oc8051_golden_model_1.IE [4]);
  nor _63548_ (_12876_, _12875_, _12874_);
  and _63549_ (_12877_, _08622_, \oc8051_golden_model_1.SCON [4]);
  and _63550_ (_12878_, _08624_, \oc8051_golden_model_1.P2 [4]);
  nor _63551_ (_12879_, _12878_, _12877_);
  and _63552_ (_12880_, _12879_, _12876_);
  and _63553_ (_12881_, _08630_, \oc8051_golden_model_1.PSW [4]);
  and _63554_ (_12882_, _08632_, \oc8051_golden_model_1.IP [4]);
  and _63555_ (_12883_, _08636_, \oc8051_golden_model_1.ACC [4]);
  and _63556_ (_12884_, _08634_, \oc8051_golden_model_1.B [4]);
  or _63557_ (_12885_, _12884_, _12883_);
  or _63558_ (_12886_, _12885_, _12882_);
  nor _63559_ (_12887_, _12886_, _12881_);
  and _63560_ (_12888_, _08616_, \oc8051_golden_model_1.TCON [4]);
  and _63561_ (_12889_, _07948_, \oc8051_golden_model_1.P0 [4]);
  and _63562_ (_12890_, _08620_, \oc8051_golden_model_1.P1 [4]);
  or _63563_ (_12891_, _12890_, _12889_);
  nor _63564_ (_12892_, _12891_, _12888_);
  and _63565_ (_12893_, _12892_, _12887_);
  and _63566_ (_12894_, _12893_, _12880_);
  and _63567_ (_12895_, _12894_, _08542_);
  and _63568_ (_12896_, _07889_, _06657_);
  not _63569_ (_12897_, _12896_);
  nor _63570_ (_12898_, _12897_, _12895_);
  nor _63571_ (_12899_, _12898_, _08788_);
  and _63572_ (_12900_, _12899_, _12873_);
  and _63573_ (_12901_, _07889_, _06656_);
  not _63574_ (_12902_, _12901_);
  and _63575_ (_12903_, _07948_, \oc8051_golden_model_1.P0 [0]);
  and _63576_ (_12904_, _08616_, \oc8051_golden_model_1.TCON [0]);
  and _63577_ (_12905_, _08620_, \oc8051_golden_model_1.P1 [0]);
  and _63578_ (_12906_, _08622_, \oc8051_golden_model_1.SCON [0]);
  and _63579_ (_12907_, _08624_, \oc8051_golden_model_1.P2 [0]);
  and _63580_ (_12908_, _08626_, \oc8051_golden_model_1.IE [0]);
  and _63581_ (_12909_, _08628_, \oc8051_golden_model_1.P3 [0]);
  and _63582_ (_12910_, _08632_, \oc8051_golden_model_1.IP [0]);
  and _63583_ (_12911_, _08630_, \oc8051_golden_model_1.PSW [0]);
  and _63584_ (_12912_, _08636_, \oc8051_golden_model_1.ACC [0]);
  and _63585_ (_12913_, _08634_, \oc8051_golden_model_1.B [0]);
  or _63586_ (_12914_, _12913_, _12912_);
  or _63587_ (_12915_, _12914_, _12911_);
  or _63588_ (_12916_, _12915_, _12910_);
  or _63589_ (_12917_, _12916_, _12909_);
  or _63590_ (_12918_, _12917_, _12908_);
  or _63591_ (_12919_, _12918_, _12907_);
  or _63592_ (_12920_, _12919_, _12906_);
  or _63593_ (_12921_, _12920_, _12905_);
  or _63594_ (_12922_, _12921_, _12904_);
  nor _63595_ (_12923_, _12922_, _12903_);
  not _63596_ (_12924_, _12923_);
  nor _63597_ (_12925_, _12924_, _08389_);
  nor _63598_ (_12926_, _12925_, _12902_);
  and _63599_ (_12927_, _08632_, \oc8051_golden_model_1.IP [6]);
  and _63600_ (_12928_, _08622_, \oc8051_golden_model_1.SCON [6]);
  nor _63601_ (_12929_, _12928_, _12927_);
  and _63602_ (_12930_, _08630_, \oc8051_golden_model_1.PSW [6]);
  and _63603_ (_12931_, _08634_, \oc8051_golden_model_1.B [6]);
  and _63604_ (_12932_, _08636_, \oc8051_golden_model_1.ACC [6]);
  or _63605_ (_12933_, _12932_, _12931_);
  nor _63606_ (_12934_, _12933_, _12930_);
  and _63607_ (_12935_, _08616_, \oc8051_golden_model_1.TCON [6]);
  and _63608_ (_12936_, _07948_, \oc8051_golden_model_1.P0 [6]);
  and _63609_ (_12937_, _08620_, \oc8051_golden_model_1.P1 [6]);
  or _63610_ (_12938_, _12937_, _12936_);
  nor _63611_ (_12939_, _12938_, _12935_);
  and _63612_ (_12940_, _08624_, \oc8051_golden_model_1.P2 [6]);
  and _63613_ (_12941_, _08628_, \oc8051_golden_model_1.P3 [6]);
  and _63614_ (_12942_, _08626_, \oc8051_golden_model_1.IE [6]);
  or _63615_ (_12943_, _12942_, _12941_);
  nor _63616_ (_12944_, _12943_, _12940_);
  and _63617_ (_12945_, _12944_, _12939_);
  and _63618_ (_12946_, _12945_, _12934_);
  and _63619_ (_12947_, _12946_, _12929_);
  and _63620_ (_12948_, _12947_, _08143_);
  and _63621_ (_12949_, _07917_, _06657_);
  not _63622_ (_12950_, _12949_);
  nor _63623_ (_12951_, _12950_, _12948_);
  nor _63624_ (_12952_, _12951_, _12926_);
  not _63625_ (_12953_, _08185_);
  and _63626_ (_12954_, _07948_, \oc8051_golden_model_1.P0 [3]);
  and _63627_ (_12955_, _08616_, \oc8051_golden_model_1.TCON [3]);
  and _63628_ (_12956_, _08620_, \oc8051_golden_model_1.P1 [3]);
  and _63629_ (_12957_, _08622_, \oc8051_golden_model_1.SCON [3]);
  and _63630_ (_12958_, _08624_, \oc8051_golden_model_1.P2 [3]);
  and _63631_ (_12959_, _08626_, \oc8051_golden_model_1.IE [3]);
  and _63632_ (_12960_, _08628_, \oc8051_golden_model_1.P3 [3]);
  and _63633_ (_12961_, _08632_, \oc8051_golden_model_1.IP [3]);
  and _63634_ (_12962_, _08630_, \oc8051_golden_model_1.PSW [3]);
  and _63635_ (_12963_, _08634_, \oc8051_golden_model_1.B [3]);
  and _63636_ (_12964_, _08636_, \oc8051_golden_model_1.ACC [3]);
  or _63637_ (_12965_, _12964_, _12963_);
  or _63638_ (_12966_, _12965_, _12962_);
  or _63639_ (_12967_, _12966_, _12961_);
  or _63640_ (_12968_, _12967_, _12960_);
  or _63641_ (_12969_, _12968_, _12959_);
  or _63642_ (_12970_, _12969_, _12958_);
  or _63643_ (_12971_, _12970_, _12957_);
  or _63644_ (_12972_, _12971_, _12956_);
  or _63645_ (_12973_, _12972_, _12955_);
  nor _63646_ (_12974_, _12973_, _12954_);
  and _63647_ (_12975_, _12974_, _08290_);
  nor _63648_ (_12976_, _12975_, _12953_);
  and _63649_ (_12977_, _07948_, \oc8051_golden_model_1.P0 [5]);
  and _63650_ (_12978_, _08616_, \oc8051_golden_model_1.TCON [5]);
  and _63651_ (_12979_, _08620_, \oc8051_golden_model_1.P1 [5]);
  and _63652_ (_12980_, _08622_, \oc8051_golden_model_1.SCON [5]);
  and _63653_ (_12981_, _08624_, \oc8051_golden_model_1.P2 [5]);
  and _63654_ (_12982_, _08626_, \oc8051_golden_model_1.IE [5]);
  and _63655_ (_12983_, _08628_, \oc8051_golden_model_1.P3 [5]);
  and _63656_ (_12984_, _08632_, \oc8051_golden_model_1.IP [5]);
  and _63657_ (_12985_, _08630_, \oc8051_golden_model_1.PSW [5]);
  and _63658_ (_12986_, _08636_, \oc8051_golden_model_1.ACC [5]);
  and _63659_ (_12987_, _08634_, \oc8051_golden_model_1.B [5]);
  or _63660_ (_12988_, _12987_, _12986_);
  or _63661_ (_12989_, _12988_, _12985_);
  or _63662_ (_12990_, _12989_, _12984_);
  or _63663_ (_12991_, _12990_, _12983_);
  or _63664_ (_12992_, _12991_, _12982_);
  or _63665_ (_12993_, _12992_, _12981_);
  or _63666_ (_12994_, _12993_, _12980_);
  or _63667_ (_12995_, _12994_, _12979_);
  or _63668_ (_12996_, _12995_, _12978_);
  nor _63669_ (_12997_, _12996_, _12977_);
  and _63670_ (_12998_, _12997_, _08245_);
  and _63671_ (_12999_, _07880_, _06657_);
  not _63672_ (_13000_, _12999_);
  nor _63673_ (_13001_, _13000_, _12998_);
  nor _63674_ (_13002_, _13001_, _12976_);
  and _63675_ (_13003_, _13002_, _12952_);
  and _63676_ (_13004_, _13003_, _12900_);
  nor _63677_ (_13005_, _09478_, _13004_);
  and _63678_ (_13006_, _12303_, _13004_);
  or _63679_ (_13007_, _13006_, _06558_);
  or _63680_ (_13008_, _13007_, _13005_);
  and _63681_ (_13009_, _13008_, _12151_);
  and _63682_ (_13010_, _13009_, _12824_);
  or _63683_ (_13011_, _13010_, _12152_);
  nor _63684_ (_13012_, _11243_, _06283_);
  nand _63685_ (_13013_, _13012_, _13011_);
  nor _63686_ (_13014_, _13012_, _09487_);
  nor _63687_ (_13015_, _13014_, _11284_);
  and _63688_ (_13016_, _13015_, _13013_);
  and _63689_ (_13017_, _12149_, _11284_);
  or _63690_ (_13018_, _13017_, _06281_);
  nor _63691_ (_13019_, _13018_, _13016_);
  and _63692_ (_13020_, _08040_, _06281_);
  or _63693_ (_13021_, _13020_, _13019_);
  nand _63694_ (_13022_, _13021_, _05964_);
  nor _63695_ (_13023_, _09487_, _05964_);
  nor _63696_ (_13024_, _13023_, _06362_);
  nand _63697_ (_13025_, _13024_, _13022_);
  nor _63698_ (_13026_, _12380_, _13004_);
  and _63699_ (_13027_, _09479_, _13004_);
  nor _63700_ (_13028_, _13027_, _13026_);
  and _63701_ (_13029_, _13028_, _06362_);
  and _63702_ (_13030_, _08569_, _07264_);
  not _63703_ (_13031_, _13030_);
  nor _63704_ (_13032_, _13031_, _13029_);
  nand _63705_ (_13033_, _13032_, _13025_);
  nor _63706_ (_13034_, _13030_, _12149_);
  nor _63707_ (_13035_, _13034_, _06568_);
  nand _63708_ (_13036_, _13035_, _13033_);
  nor _63709_ (_13037_, _11335_, _11330_);
  not _63710_ (_13038_, _13037_);
  and _63711_ (_13039_, _09487_, _06568_);
  nor _63712_ (_13040_, _13039_, _13038_);
  nand _63713_ (_13041_, _13040_, _13036_);
  nor _63714_ (_13042_, _12149_, _13037_);
  nor _63715_ (_13043_, _13042_, _06361_);
  nand _63716_ (_13044_, _13043_, _13041_);
  and _63717_ (_13045_, _06361_, _06182_);
  nor _63718_ (_13046_, _13045_, _05940_);
  nand _63719_ (_13047_, _13046_, _13044_);
  and _63720_ (_13048_, _12388_, _05940_);
  nor _63721_ (_13049_, _13048_, _05927_);
  nand _63722_ (_13050_, _13049_, _13047_);
  and _63723_ (_13051_, _13028_, _05927_);
  nor _63724_ (_13052_, _09424_, _07281_);
  not _63725_ (_13053_, _13052_);
  nor _63726_ (_13054_, _13053_, _13051_);
  nand _63727_ (_13055_, _13054_, _13050_);
  nor _63728_ (_13056_, _13052_, _12149_);
  nor _63729_ (_13057_, _13056_, _06278_);
  nand _63730_ (_13058_, _13057_, _13055_);
  not _63731_ (_13059_, _12141_);
  and _63732_ (_13060_, _09487_, _06278_);
  nor _63733_ (_13061_, _13060_, _13059_);
  and _63734_ (_13062_, _13061_, _13058_);
  or _63735_ (_13063_, _13062_, _12150_);
  nand _63736_ (_13064_, _13063_, _12140_);
  nor _63737_ (_13065_, _12140_, _06182_);
  nor _63738_ (_13066_, _13065_, _05939_);
  nand _63739_ (_13067_, _13066_, _13064_);
  and _63740_ (_13068_, _05938_, _05926_);
  and _63741_ (_13069_, _09487_, _05939_);
  nor _63742_ (_13070_, _13069_, _13068_);
  and _63743_ (_13071_, _13070_, _13067_);
  and _63744_ (_13072_, _13068_, _12385_);
  nor _63745_ (_13073_, _13072_, _13071_);
  or _63746_ (_13074_, _13073_, _01351_);
  or _63747_ (_13075_, _01347_, \oc8051_golden_model_1.PC [15]);
  and _63748_ (_13076_, _13075_, _42618_);
  and _63749_ (_40586_, _13076_, _13074_);
  not _63750_ (_13077_, _07904_);
  and _63751_ (_13078_, _13077_, \oc8051_golden_model_1.P2 [7]);
  and _63752_ (_13079_, _08575_, _07904_);
  or _63753_ (_13080_, _13079_, _13078_);
  and _63754_ (_13081_, _13080_, _06536_);
  nor _63755_ (_13082_, _08040_, _13077_);
  or _63756_ (_13083_, _13082_, _13078_);
  or _63757_ (_13084_, _13083_, _07215_);
  not _63758_ (_13085_, _08624_);
  and _63759_ (_13086_, _13085_, \oc8051_golden_model_1.P2 [7]);
  and _63760_ (_13087_, _08649_, _08624_);
  or _63761_ (_13088_, _13087_, _13086_);
  and _63762_ (_13089_, _13088_, _06268_);
  and _63763_ (_13090_, _08768_, _07904_);
  or _63764_ (_13091_, _13090_, _13078_);
  or _63765_ (_13092_, _13091_, _07151_);
  and _63766_ (_13093_, _07904_, \oc8051_golden_model_1.ACC [7]);
  or _63767_ (_13094_, _13093_, _13078_);
  and _63768_ (_13095_, _13094_, _07141_);
  and _63769_ (_13096_, _07142_, \oc8051_golden_model_1.P2 [7]);
  or _63770_ (_13097_, _13096_, _06341_);
  or _63771_ (_13098_, _13097_, _13095_);
  and _63772_ (_13099_, _13098_, _06273_);
  and _63773_ (_13100_, _13099_, _13092_);
  and _63774_ (_13101_, _08773_, _08624_);
  or _63775_ (_13102_, _13101_, _13086_);
  and _63776_ (_13103_, _13102_, _06272_);
  or _63777_ (_13104_, _13103_, _06461_);
  or _63778_ (_13105_, _13104_, _13100_);
  or _63779_ (_13106_, _13083_, _07166_);
  and _63780_ (_13107_, _13106_, _13105_);
  or _63781_ (_13108_, _13107_, _06464_);
  or _63782_ (_13109_, _13094_, _06465_);
  and _63783_ (_13110_, _13109_, _06269_);
  and _63784_ (_13111_, _13110_, _13108_);
  or _63785_ (_13112_, _13111_, _13089_);
  and _63786_ (_13113_, _13112_, _06262_);
  or _63787_ (_13114_, _13086_, _08789_);
  and _63788_ (_13115_, _13114_, _06261_);
  and _63789_ (_13116_, _13115_, _13102_);
  or _63790_ (_13117_, _13116_, _13113_);
  and _63791_ (_13118_, _13117_, _06258_);
  and _63792_ (_13119_, _08808_, _08624_);
  or _63793_ (_13120_, _13119_, _13086_);
  and _63794_ (_13121_, _13120_, _06257_);
  or _63795_ (_13122_, _13121_, _10080_);
  or _63796_ (_13123_, _13122_, _13118_);
  and _63797_ (_13124_, _13123_, _13084_);
  or _63798_ (_13125_, _13124_, _07460_);
  and _63799_ (_13126_, _08755_, _07904_);
  or _63800_ (_13127_, _13078_, _07208_);
  or _63801_ (_13128_, _13127_, _13126_);
  and _63802_ (_13129_, _13128_, _05982_);
  and _63803_ (_13130_, _13129_, _13125_);
  and _63804_ (_13131_, _09021_, _07904_);
  or _63805_ (_13132_, _13131_, _13078_);
  and _63806_ (_13133_, _13132_, _10094_);
  or _63807_ (_13134_, _13133_, _06218_);
  or _63808_ (_13135_, _13134_, _13130_);
  and _63809_ (_13136_, _08825_, _07904_);
  or _63810_ (_13137_, _13136_, _13078_);
  or _63811_ (_13138_, _13137_, _06219_);
  and _63812_ (_13139_, _13138_, _13135_);
  or _63813_ (_13140_, _13139_, _06369_);
  and _63814_ (_13141_, _09044_, _07904_);
  or _63815_ (_13142_, _13141_, _13078_);
  or _63816_ (_13143_, _13142_, _07237_);
  and _63817_ (_13144_, _13143_, _07240_);
  and _63818_ (_13145_, _13144_, _13140_);
  or _63819_ (_13146_, _13145_, _13081_);
  and _63820_ (_13147_, _13146_, _07242_);
  or _63821_ (_13148_, _13078_, _08043_);
  and _63822_ (_13149_, _13137_, _06375_);
  and _63823_ (_13150_, _13149_, _13148_);
  or _63824_ (_13151_, _13150_, _13147_);
  and _63825_ (_13152_, _13151_, _07234_);
  and _63826_ (_13153_, _13094_, _06545_);
  and _63827_ (_13154_, _13153_, _13148_);
  or _63828_ (_13155_, _13154_, _06366_);
  or _63829_ (_13156_, _13155_, _13152_);
  nor _63830_ (_13157_, _09043_, _13077_);
  or _63831_ (_13158_, _13078_, _09056_);
  or _63832_ (_13159_, _13158_, _13157_);
  and _63833_ (_13160_, _13159_, _09061_);
  and _63834_ (_13161_, _13160_, _13156_);
  nor _63835_ (_13162_, _08573_, _13077_);
  or _63836_ (_13163_, _13162_, _13078_);
  and _63837_ (_13164_, _13163_, _06528_);
  or _63838_ (_13165_, _13164_, _06568_);
  or _63839_ (_13166_, _13165_, _13161_);
  or _63840_ (_13167_, _13091_, _06926_);
  and _63841_ (_13168_, _13167_, _05928_);
  and _63842_ (_13169_, _13168_, _13166_);
  and _63843_ (_13170_, _13088_, _05927_);
  or _63844_ (_13171_, _13170_, _06278_);
  or _63845_ (_13172_, _13171_, _13169_);
  and _63846_ (_13173_, _08550_, _07904_);
  or _63847_ (_13174_, _13078_, _06279_);
  or _63848_ (_13175_, _13174_, _13173_);
  and _63849_ (_13176_, _13175_, _01347_);
  and _63850_ (_13177_, _13176_, _13172_);
  nor _63851_ (_13178_, \oc8051_golden_model_1.P2 [7], rst);
  nor _63852_ (_13179_, _13178_, _01354_);
  or _63853_ (_40587_, _13179_, _13177_);
  not _63854_ (_13180_, _07894_);
  and _63855_ (_13181_, _13180_, \oc8051_golden_model_1.P3 [7]);
  and _63856_ (_13182_, _08575_, _07894_);
  or _63857_ (_13183_, _13182_, _13181_);
  and _63858_ (_13184_, _13183_, _06536_);
  nor _63859_ (_13185_, _08040_, _13180_);
  or _63860_ (_13186_, _13185_, _13181_);
  or _63861_ (_13187_, _13186_, _07215_);
  not _63862_ (_13188_, _08628_);
  and _63863_ (_13189_, _13188_, \oc8051_golden_model_1.P3 [7]);
  and _63864_ (_13190_, _08649_, _08628_);
  or _63865_ (_13191_, _13190_, _13189_);
  and _63866_ (_13192_, _13191_, _06268_);
  and _63867_ (_13193_, _08768_, _07894_);
  or _63868_ (_13194_, _13193_, _13181_);
  or _63869_ (_13195_, _13194_, _07151_);
  and _63870_ (_13196_, _07894_, \oc8051_golden_model_1.ACC [7]);
  or _63871_ (_13197_, _13196_, _13181_);
  and _63872_ (_13198_, _13197_, _07141_);
  and _63873_ (_13199_, _07142_, \oc8051_golden_model_1.P3 [7]);
  or _63874_ (_13200_, _13199_, _06341_);
  or _63875_ (_13201_, _13200_, _13198_);
  and _63876_ (_13202_, _13201_, _06273_);
  and _63877_ (_13203_, _13202_, _13195_);
  and _63878_ (_13204_, _08773_, _08628_);
  or _63879_ (_13205_, _13204_, _13189_);
  and _63880_ (_13206_, _13205_, _06272_);
  or _63881_ (_13207_, _13206_, _06461_);
  or _63882_ (_13208_, _13207_, _13203_);
  or _63883_ (_13209_, _13186_, _07166_);
  and _63884_ (_13210_, _13209_, _13208_);
  or _63885_ (_13211_, _13210_, _06464_);
  or _63886_ (_13212_, _13197_, _06465_);
  and _63887_ (_13213_, _13212_, _06269_);
  and _63888_ (_13214_, _13213_, _13211_);
  or _63889_ (_13215_, _13214_, _13192_);
  and _63890_ (_13216_, _13215_, _06262_);
  and _63891_ (_13217_, _08790_, _08628_);
  or _63892_ (_13218_, _13217_, _13189_);
  and _63893_ (_13219_, _13218_, _06261_);
  or _63894_ (_13220_, _13219_, _13216_);
  and _63895_ (_13221_, _13220_, _06258_);
  and _63896_ (_13222_, _08808_, _08628_);
  or _63897_ (_13223_, _13222_, _13189_);
  and _63898_ (_13224_, _13223_, _06257_);
  or _63899_ (_13225_, _13224_, _10080_);
  or _63900_ (_13226_, _13225_, _13221_);
  and _63901_ (_13227_, _13226_, _13187_);
  or _63902_ (_13228_, _13227_, _07460_);
  and _63903_ (_13229_, _08755_, _07894_);
  or _63904_ (_13230_, _13181_, _07208_);
  or _63905_ (_13231_, _13230_, _13229_);
  and _63906_ (_13232_, _13231_, _05982_);
  and _63907_ (_13233_, _13232_, _13228_);
  and _63908_ (_13234_, _09021_, _07894_);
  or _63909_ (_13235_, _13234_, _13181_);
  and _63910_ (_13236_, _13235_, _10094_);
  or _63911_ (_13237_, _13236_, _06218_);
  or _63912_ (_13238_, _13237_, _13233_);
  and _63913_ (_13239_, _08825_, _07894_);
  or _63914_ (_13240_, _13239_, _13181_);
  or _63915_ (_13241_, _13240_, _06219_);
  and _63916_ (_13242_, _13241_, _13238_);
  or _63917_ (_13243_, _13242_, _06369_);
  and _63918_ (_13244_, _09044_, _07894_);
  or _63919_ (_13245_, _13244_, _13181_);
  or _63920_ (_13246_, _13245_, _07237_);
  and _63921_ (_13247_, _13246_, _07240_);
  and _63922_ (_13248_, _13247_, _13243_);
  or _63923_ (_13249_, _13248_, _13184_);
  and _63924_ (_13250_, _13249_, _07242_);
  or _63925_ (_13251_, _13181_, _08043_);
  and _63926_ (_13252_, _13240_, _06375_);
  and _63927_ (_13253_, _13252_, _13251_);
  or _63928_ (_13254_, _13253_, _13250_);
  and _63929_ (_13255_, _13254_, _07234_);
  and _63930_ (_13256_, _13197_, _06545_);
  and _63931_ (_13257_, _13256_, _13251_);
  or _63932_ (_13258_, _13257_, _06366_);
  or _63933_ (_13259_, _13258_, _13255_);
  nor _63934_ (_13260_, _09043_, _13180_);
  or _63935_ (_13261_, _13181_, _09056_);
  or _63936_ (_13262_, _13261_, _13260_);
  and _63937_ (_13263_, _13262_, _09061_);
  and _63938_ (_13264_, _13263_, _13259_);
  nor _63939_ (_13265_, _08573_, _13180_);
  or _63940_ (_13266_, _13265_, _13181_);
  and _63941_ (_13267_, _13266_, _06528_);
  or _63942_ (_13268_, _13267_, _06568_);
  or _63943_ (_13269_, _13268_, _13264_);
  or _63944_ (_13270_, _13194_, _06926_);
  and _63945_ (_13271_, _13270_, _05928_);
  and _63946_ (_13272_, _13271_, _13269_);
  and _63947_ (_13273_, _13191_, _05927_);
  or _63948_ (_13274_, _13273_, _06278_);
  or _63949_ (_13275_, _13274_, _13272_);
  and _63950_ (_13276_, _08550_, _07894_);
  or _63951_ (_13277_, _13181_, _06279_);
  or _63952_ (_13278_, _13277_, _13276_);
  and _63953_ (_13279_, _13278_, _01347_);
  and _63954_ (_13280_, _13279_, _13275_);
  nor _63955_ (_13281_, \oc8051_golden_model_1.P3 [7], rst);
  nor _63956_ (_13282_, _13281_, _01354_);
  or _63957_ (_40588_, _13282_, _13280_);
  not _63958_ (_13283_, _07926_);
  and _63959_ (_13284_, _13283_, \oc8051_golden_model_1.P0 [7]);
  and _63960_ (_13285_, _08575_, _07926_);
  or _63961_ (_13286_, _13285_, _13284_);
  and _63962_ (_13287_, _13286_, _06536_);
  nor _63963_ (_13288_, _08040_, _13283_);
  or _63964_ (_13289_, _13288_, _13284_);
  or _63965_ (_13290_, _13289_, _07215_);
  not _63966_ (_13291_, _07948_);
  and _63967_ (_13292_, _13291_, \oc8051_golden_model_1.P0 [7]);
  and _63968_ (_13293_, _08649_, _07948_);
  or _63969_ (_13294_, _13293_, _13292_);
  and _63970_ (_13295_, _13294_, _06268_);
  and _63971_ (_13296_, _08768_, _07926_);
  or _63972_ (_13297_, _13296_, _13284_);
  or _63973_ (_13298_, _13297_, _07151_);
  and _63974_ (_13299_, _07926_, \oc8051_golden_model_1.ACC [7]);
  or _63975_ (_13300_, _13299_, _13284_);
  and _63976_ (_13301_, _13300_, _07141_);
  and _63977_ (_13302_, _07142_, \oc8051_golden_model_1.P0 [7]);
  or _63978_ (_13303_, _13302_, _06341_);
  or _63979_ (_13304_, _13303_, _13301_);
  and _63980_ (_13305_, _13304_, _06273_);
  and _63981_ (_13306_, _13305_, _13298_);
  and _63982_ (_13307_, _08773_, _07948_);
  or _63983_ (_13308_, _13307_, _13292_);
  and _63984_ (_13309_, _13308_, _06272_);
  or _63985_ (_13310_, _13309_, _06461_);
  or _63986_ (_13311_, _13310_, _13306_);
  or _63987_ (_13312_, _13289_, _07166_);
  and _63988_ (_13313_, _13312_, _13311_);
  or _63989_ (_13314_, _13313_, _06464_);
  or _63990_ (_13315_, _13300_, _06465_);
  and _63991_ (_13316_, _13315_, _06269_);
  and _63992_ (_13317_, _13316_, _13314_);
  or _63993_ (_13318_, _13317_, _13295_);
  and _63994_ (_13319_, _13318_, _06262_);
  and _63995_ (_13320_, _08790_, _07948_);
  or _63996_ (_13321_, _13320_, _13292_);
  and _63997_ (_13322_, _13321_, _06261_);
  or _63998_ (_13323_, _13322_, _13319_);
  and _63999_ (_13324_, _13323_, _06258_);
  and _64000_ (_13325_, _08808_, _07948_);
  or _64001_ (_13326_, _13325_, _13292_);
  and _64002_ (_13327_, _13326_, _06257_);
  or _64003_ (_13328_, _13327_, _10080_);
  or _64004_ (_13329_, _13328_, _13324_);
  and _64005_ (_13330_, _13329_, _13290_);
  or _64006_ (_13331_, _13330_, _07460_);
  and _64007_ (_13332_, _08755_, _07926_);
  or _64008_ (_13333_, _13284_, _07208_);
  or _64009_ (_13334_, _13333_, _13332_);
  and _64010_ (_13335_, _13334_, _05982_);
  and _64011_ (_13336_, _13335_, _13331_);
  and _64012_ (_13337_, _09021_, _07926_);
  or _64013_ (_13338_, _13337_, _13284_);
  and _64014_ (_13339_, _13338_, _10094_);
  or _64015_ (_13340_, _13339_, _06218_);
  or _64016_ (_13341_, _13340_, _13336_);
  and _64017_ (_13342_, _08825_, _07926_);
  or _64018_ (_13343_, _13342_, _13284_);
  or _64019_ (_13344_, _13343_, _06219_);
  and _64020_ (_13345_, _13344_, _13341_);
  or _64021_ (_13346_, _13345_, _06369_);
  and _64022_ (_13347_, _09044_, _07926_);
  or _64023_ (_13348_, _13347_, _13284_);
  or _64024_ (_13349_, _13348_, _07237_);
  and _64025_ (_13350_, _13349_, _07240_);
  and _64026_ (_13351_, _13350_, _13346_);
  or _64027_ (_13352_, _13351_, _13287_);
  and _64028_ (_13353_, _13352_, _07242_);
  or _64029_ (_13354_, _13284_, _08043_);
  and _64030_ (_13355_, _13343_, _06375_);
  and _64031_ (_13356_, _13355_, _13354_);
  or _64032_ (_13357_, _13356_, _13353_);
  and _64033_ (_13358_, _13357_, _07234_);
  and _64034_ (_13359_, _13300_, _06545_);
  and _64035_ (_13360_, _13359_, _13354_);
  or _64036_ (_13361_, _13360_, _06366_);
  or _64037_ (_13362_, _13361_, _13358_);
  nor _64038_ (_13363_, _09043_, _13283_);
  or _64039_ (_13364_, _13284_, _09056_);
  or _64040_ (_13365_, _13364_, _13363_);
  and _64041_ (_13366_, _13365_, _09061_);
  and _64042_ (_13367_, _13366_, _13362_);
  nor _64043_ (_13368_, _08573_, _13283_);
  or _64044_ (_13369_, _13368_, _13284_);
  and _64045_ (_13370_, _13369_, _06528_);
  or _64046_ (_13371_, _13370_, _06568_);
  or _64047_ (_13372_, _13371_, _13367_);
  or _64048_ (_13373_, _13297_, _06926_);
  and _64049_ (_13374_, _13373_, _05928_);
  and _64050_ (_13375_, _13374_, _13372_);
  and _64051_ (_13376_, _13294_, _05927_);
  or _64052_ (_13377_, _13376_, _06278_);
  or _64053_ (_13378_, _13377_, _13375_);
  and _64054_ (_13379_, _08550_, _07926_);
  or _64055_ (_13380_, _13284_, _06279_);
  or _64056_ (_13381_, _13380_, _13379_);
  and _64057_ (_13382_, _13381_, _01347_);
  and _64058_ (_13383_, _13382_, _13378_);
  nor _64059_ (_13384_, \oc8051_golden_model_1.P0 [7], rst);
  nor _64060_ (_13385_, _13384_, _01354_);
  or _64061_ (_40589_, _13385_, _13383_);
  nor _64062_ (_13386_, \oc8051_golden_model_1.P1 [7], rst);
  nor _64063_ (_13387_, _13386_, _01354_);
  not _64064_ (_13388_, _07971_);
  and _64065_ (_13389_, _13388_, \oc8051_golden_model_1.P1 [7]);
  and _64066_ (_13390_, _08575_, _07971_);
  or _64067_ (_13391_, _13390_, _13389_);
  and _64068_ (_13392_, _13391_, _06536_);
  nor _64069_ (_13393_, _08040_, _13388_);
  or _64070_ (_13394_, _13393_, _13389_);
  or _64071_ (_13395_, _13394_, _07215_);
  not _64072_ (_13396_, _08620_);
  and _64073_ (_13397_, _13396_, \oc8051_golden_model_1.P1 [7]);
  and _64074_ (_13398_, _08649_, _08620_);
  or _64075_ (_13399_, _13398_, _13397_);
  and _64076_ (_13400_, _13399_, _06268_);
  and _64077_ (_13401_, _08768_, _07971_);
  or _64078_ (_13402_, _13401_, _13389_);
  or _64079_ (_13403_, _13402_, _07151_);
  and _64080_ (_13404_, _07971_, \oc8051_golden_model_1.ACC [7]);
  or _64081_ (_13405_, _13404_, _13389_);
  and _64082_ (_13406_, _13405_, _07141_);
  and _64083_ (_13407_, _07142_, \oc8051_golden_model_1.P1 [7]);
  or _64084_ (_13408_, _13407_, _06341_);
  or _64085_ (_13409_, _13408_, _13406_);
  and _64086_ (_13410_, _13409_, _06273_);
  and _64087_ (_13411_, _13410_, _13403_);
  and _64088_ (_13412_, _08773_, _08620_);
  or _64089_ (_13413_, _13412_, _13397_);
  and _64090_ (_13414_, _13413_, _06272_);
  or _64091_ (_13415_, _13414_, _06461_);
  or _64092_ (_13416_, _13415_, _13411_);
  or _64093_ (_13417_, _13394_, _07166_);
  and _64094_ (_13418_, _13417_, _13416_);
  or _64095_ (_13419_, _13418_, _06464_);
  or _64096_ (_13420_, _13405_, _06465_);
  and _64097_ (_13421_, _13420_, _06269_);
  and _64098_ (_13422_, _13421_, _13419_);
  or _64099_ (_13423_, _13422_, _13400_);
  and _64100_ (_13424_, _13423_, _06262_);
  or _64101_ (_13425_, _13397_, _08789_);
  and _64102_ (_13426_, _13425_, _06261_);
  and _64103_ (_13427_, _13426_, _13413_);
  or _64104_ (_13428_, _13427_, _13424_);
  and _64105_ (_13429_, _13428_, _06258_);
  and _64106_ (_13430_, _08808_, _08620_);
  or _64107_ (_13431_, _13430_, _13397_);
  and _64108_ (_13432_, _13431_, _06257_);
  or _64109_ (_13433_, _13432_, _10080_);
  or _64110_ (_13434_, _13433_, _13429_);
  and _64111_ (_13435_, _13434_, _13395_);
  or _64112_ (_13436_, _13435_, _07460_);
  and _64113_ (_13437_, _08755_, _07971_);
  or _64114_ (_13438_, _13389_, _07208_);
  or _64115_ (_13439_, _13438_, _13437_);
  and _64116_ (_13440_, _13439_, _05982_);
  and _64117_ (_13441_, _13440_, _13436_);
  and _64118_ (_13442_, _09021_, _07971_);
  or _64119_ (_13443_, _13442_, _13389_);
  and _64120_ (_13444_, _13443_, _10094_);
  or _64121_ (_13445_, _13444_, _06218_);
  or _64122_ (_13446_, _13445_, _13441_);
  and _64123_ (_13447_, _08825_, _07971_);
  or _64124_ (_13448_, _13447_, _13389_);
  or _64125_ (_13449_, _13448_, _06219_);
  and _64126_ (_13450_, _13449_, _13446_);
  or _64127_ (_13451_, _13450_, _06369_);
  and _64128_ (_13452_, _09044_, _07971_);
  or _64129_ (_13453_, _13452_, _13389_);
  or _64130_ (_13454_, _13453_, _07237_);
  and _64131_ (_13455_, _13454_, _07240_);
  and _64132_ (_13456_, _13455_, _13451_);
  or _64133_ (_13457_, _13456_, _13392_);
  and _64134_ (_13458_, _13457_, _07242_);
  or _64135_ (_13459_, _13389_, _08043_);
  and _64136_ (_13460_, _13448_, _06375_);
  and _64137_ (_13461_, _13460_, _13459_);
  or _64138_ (_13462_, _13461_, _13458_);
  and _64139_ (_13463_, _13462_, _07234_);
  and _64140_ (_13464_, _13405_, _06545_);
  and _64141_ (_13465_, _13464_, _13459_);
  or _64142_ (_13466_, _13465_, _06366_);
  or _64143_ (_13467_, _13466_, _13463_);
  nor _64144_ (_13468_, _09043_, _13388_);
  or _64145_ (_13469_, _13389_, _09056_);
  or _64146_ (_13470_, _13469_, _13468_);
  and _64147_ (_13471_, _13470_, _09061_);
  and _64148_ (_13472_, _13471_, _13467_);
  nor _64149_ (_13473_, _08573_, _13388_);
  or _64150_ (_13474_, _13473_, _13389_);
  and _64151_ (_13475_, _13474_, _06528_);
  or _64152_ (_13476_, _13475_, _06568_);
  or _64153_ (_13477_, _13476_, _13472_);
  or _64154_ (_13478_, _13402_, _06926_);
  and _64155_ (_13479_, _13478_, _05928_);
  and _64156_ (_13480_, _13479_, _13477_);
  and _64157_ (_13481_, _13399_, _05927_);
  or _64158_ (_13482_, _13481_, _06278_);
  or _64159_ (_13483_, _13482_, _13480_);
  and _64160_ (_13484_, _08550_, _07971_);
  or _64161_ (_13485_, _13389_, _06279_);
  or _64162_ (_13486_, _13485_, _13484_);
  and _64163_ (_13487_, _13486_, _01347_);
  and _64164_ (_13488_, _13487_, _13483_);
  or _64165_ (_40591_, _13488_, _13387_);
  and _64166_ (_13489_, _01351_, \oc8051_golden_model_1.IP [7]);
  not _64167_ (_13490_, _07946_);
  and _64168_ (_13491_, _13490_, \oc8051_golden_model_1.IP [7]);
  and _64169_ (_13492_, _08575_, _07946_);
  or _64170_ (_13493_, _13492_, _13491_);
  and _64171_ (_13494_, _13493_, _06536_);
  nor _64172_ (_13495_, _08040_, _13490_);
  or _64173_ (_13496_, _13495_, _13491_);
  or _64174_ (_13497_, _13496_, _07215_);
  not _64175_ (_13498_, _08632_);
  and _64176_ (_13499_, _13498_, \oc8051_golden_model_1.IP [7]);
  and _64177_ (_13500_, _08649_, _08632_);
  or _64178_ (_13501_, _13500_, _13499_);
  and _64179_ (_13502_, _13501_, _06268_);
  and _64180_ (_13503_, _08768_, _07946_);
  or _64181_ (_13504_, _13503_, _13491_);
  or _64182_ (_13505_, _13504_, _07151_);
  and _64183_ (_13506_, _07946_, \oc8051_golden_model_1.ACC [7]);
  or _64184_ (_13507_, _13506_, _13491_);
  and _64185_ (_13508_, _13507_, _07141_);
  and _64186_ (_13509_, _07142_, \oc8051_golden_model_1.IP [7]);
  or _64187_ (_13510_, _13509_, _06341_);
  or _64188_ (_13511_, _13510_, _13508_);
  and _64189_ (_13512_, _13511_, _06273_);
  and _64190_ (_13513_, _13512_, _13505_);
  and _64191_ (_13514_, _08773_, _08632_);
  or _64192_ (_13515_, _13514_, _13499_);
  and _64193_ (_13516_, _13515_, _06272_);
  or _64194_ (_13517_, _13516_, _06461_);
  or _64195_ (_13518_, _13517_, _13513_);
  or _64196_ (_13519_, _13496_, _07166_);
  and _64197_ (_13520_, _13519_, _13518_);
  or _64198_ (_13521_, _13520_, _06464_);
  or _64199_ (_13522_, _13507_, _06465_);
  and _64200_ (_13523_, _13522_, _06269_);
  and _64201_ (_13524_, _13523_, _13521_);
  or _64202_ (_13525_, _13524_, _13502_);
  and _64203_ (_13526_, _13525_, _06262_);
  and _64204_ (_13527_, _08790_, _08632_);
  or _64205_ (_13528_, _13527_, _13499_);
  and _64206_ (_13529_, _13528_, _06261_);
  or _64207_ (_13530_, _13529_, _13526_);
  and _64208_ (_13531_, _13530_, _06258_);
  and _64209_ (_13532_, _08808_, _08632_);
  or _64210_ (_13533_, _13532_, _13499_);
  and _64211_ (_13534_, _13533_, _06257_);
  or _64212_ (_13535_, _13534_, _10080_);
  or _64213_ (_13536_, _13535_, _13531_);
  and _64214_ (_13537_, _13536_, _13497_);
  or _64215_ (_13538_, _13537_, _07460_);
  and _64216_ (_13539_, _08755_, _07946_);
  or _64217_ (_13540_, _13491_, _07208_);
  or _64218_ (_13541_, _13540_, _13539_);
  and _64219_ (_13542_, _13541_, _05982_);
  and _64220_ (_13543_, _13542_, _13538_);
  and _64221_ (_13544_, _09021_, _07946_);
  or _64222_ (_13545_, _13544_, _13491_);
  and _64223_ (_13546_, _13545_, _10094_);
  or _64224_ (_13547_, _13546_, _06218_);
  or _64225_ (_13548_, _13547_, _13543_);
  and _64226_ (_13549_, _08825_, _07946_);
  or _64227_ (_13550_, _13549_, _13491_);
  or _64228_ (_13551_, _13550_, _06219_);
  and _64229_ (_13552_, _13551_, _13548_);
  or _64230_ (_13553_, _13552_, _06369_);
  and _64231_ (_13554_, _09044_, _07946_);
  or _64232_ (_13555_, _13554_, _13491_);
  or _64233_ (_13556_, _13555_, _07237_);
  and _64234_ (_13557_, _13556_, _07240_);
  and _64235_ (_13558_, _13557_, _13553_);
  or _64236_ (_13559_, _13558_, _13494_);
  and _64237_ (_13560_, _13559_, _07242_);
  or _64238_ (_13561_, _13491_, _08043_);
  and _64239_ (_13562_, _13550_, _06375_);
  and _64240_ (_13563_, _13562_, _13561_);
  or _64241_ (_13564_, _13563_, _13560_);
  and _64242_ (_13565_, _13564_, _07234_);
  and _64243_ (_13566_, _13507_, _06545_);
  and _64244_ (_13567_, _13566_, _13561_);
  or _64245_ (_13568_, _13567_, _06366_);
  or _64246_ (_13569_, _13568_, _13565_);
  nor _64247_ (_13570_, _09043_, _13490_);
  or _64248_ (_13571_, _13491_, _09056_);
  or _64249_ (_13572_, _13571_, _13570_);
  and _64250_ (_13573_, _13572_, _09061_);
  and _64251_ (_13574_, _13573_, _13569_);
  nor _64252_ (_13575_, _08573_, _13490_);
  or _64253_ (_13576_, _13575_, _13491_);
  and _64254_ (_13577_, _13576_, _06528_);
  or _64255_ (_13578_, _13577_, _06568_);
  or _64256_ (_13579_, _13578_, _13574_);
  or _64257_ (_13580_, _13504_, _06926_);
  and _64258_ (_13581_, _13580_, _05928_);
  and _64259_ (_13582_, _13581_, _13579_);
  and _64260_ (_13583_, _13501_, _05927_);
  or _64261_ (_13584_, _13583_, _06278_);
  or _64262_ (_13585_, _13584_, _13582_);
  and _64263_ (_13586_, _08550_, _07946_);
  or _64264_ (_13587_, _13491_, _06279_);
  or _64265_ (_13588_, _13587_, _13586_);
  and _64266_ (_13589_, _13588_, _01347_);
  and _64267_ (_13590_, _13589_, _13585_);
  or _64268_ (_13591_, _13590_, _13489_);
  and _64269_ (_40592_, _13591_, _42618_);
  and _64270_ (_13592_, _01351_, \oc8051_golden_model_1.IE [7]);
  not _64271_ (_13593_, _07900_);
  and _64272_ (_13594_, _13593_, \oc8051_golden_model_1.IE [7]);
  and _64273_ (_13595_, _08575_, _07900_);
  or _64274_ (_13596_, _13595_, _13594_);
  and _64275_ (_13597_, _13596_, _06536_);
  nor _64276_ (_13598_, _08040_, _13593_);
  or _64277_ (_13599_, _13598_, _13594_);
  or _64278_ (_13600_, _13599_, _07215_);
  not _64279_ (_13601_, _08626_);
  and _64280_ (_13602_, _13601_, \oc8051_golden_model_1.IE [7]);
  and _64281_ (_13603_, _08649_, _08626_);
  or _64282_ (_13604_, _13603_, _13602_);
  and _64283_ (_13605_, _13604_, _06268_);
  and _64284_ (_13606_, _08768_, _07900_);
  or _64285_ (_13607_, _13606_, _13594_);
  or _64286_ (_13608_, _13607_, _07151_);
  and _64287_ (_13609_, _07900_, \oc8051_golden_model_1.ACC [7]);
  or _64288_ (_13610_, _13609_, _13594_);
  and _64289_ (_13611_, _13610_, _07141_);
  and _64290_ (_13612_, _07142_, \oc8051_golden_model_1.IE [7]);
  or _64291_ (_13614_, _13612_, _06341_);
  or _64292_ (_13615_, _13614_, _13611_);
  and _64293_ (_13616_, _13615_, _06273_);
  and _64294_ (_13617_, _13616_, _13608_);
  and _64295_ (_13618_, _08773_, _08626_);
  or _64296_ (_13619_, _13618_, _13602_);
  and _64297_ (_13620_, _13619_, _06272_);
  or _64298_ (_13621_, _13620_, _06461_);
  or _64299_ (_13622_, _13621_, _13617_);
  or _64300_ (_13623_, _13599_, _07166_);
  and _64301_ (_13625_, _13623_, _13622_);
  or _64302_ (_13626_, _13625_, _06464_);
  or _64303_ (_13627_, _13610_, _06465_);
  and _64304_ (_13628_, _13627_, _06269_);
  and _64305_ (_13629_, _13628_, _13626_);
  or _64306_ (_13630_, _13629_, _13605_);
  and _64307_ (_13631_, _13630_, _06262_);
  and _64308_ (_13632_, _08790_, _08626_);
  or _64309_ (_13633_, _13632_, _13602_);
  and _64310_ (_13634_, _13633_, _06261_);
  or _64311_ (_13636_, _13634_, _13631_);
  and _64312_ (_13637_, _13636_, _06258_);
  and _64313_ (_13638_, _08808_, _08626_);
  or _64314_ (_13639_, _13638_, _13602_);
  and _64315_ (_13640_, _13639_, _06257_);
  or _64316_ (_13641_, _13640_, _10080_);
  or _64317_ (_13642_, _13641_, _13637_);
  and _64318_ (_13643_, _13642_, _13600_);
  or _64319_ (_13644_, _13643_, _07460_);
  and _64320_ (_13645_, _08755_, _07900_);
  or _64321_ (_13647_, _13594_, _07208_);
  or _64322_ (_13648_, _13647_, _13645_);
  and _64323_ (_13649_, _13648_, _05982_);
  and _64324_ (_13650_, _13649_, _13644_);
  and _64325_ (_13651_, _09021_, _07900_);
  or _64326_ (_13652_, _13651_, _13594_);
  and _64327_ (_13653_, _13652_, _10094_);
  or _64328_ (_13654_, _13653_, _06218_);
  or _64329_ (_13655_, _13654_, _13650_);
  and _64330_ (_13656_, _08825_, _07900_);
  or _64331_ (_13658_, _13656_, _13594_);
  or _64332_ (_13659_, _13658_, _06219_);
  and _64333_ (_13660_, _13659_, _13655_);
  or _64334_ (_13661_, _13660_, _06369_);
  and _64335_ (_13662_, _09044_, _07900_);
  or _64336_ (_13663_, _13662_, _13594_);
  or _64337_ (_13664_, _13663_, _07237_);
  and _64338_ (_13665_, _13664_, _07240_);
  and _64339_ (_13666_, _13665_, _13661_);
  or _64340_ (_13667_, _13666_, _13597_);
  and _64341_ (_13669_, _13667_, _07242_);
  or _64342_ (_13670_, _13594_, _08043_);
  and _64343_ (_13671_, _13658_, _06375_);
  and _64344_ (_13672_, _13671_, _13670_);
  or _64345_ (_13673_, _13672_, _13669_);
  and _64346_ (_13674_, _13673_, _07234_);
  and _64347_ (_13675_, _13610_, _06545_);
  and _64348_ (_13676_, _13675_, _13670_);
  or _64349_ (_13677_, _13676_, _06366_);
  or _64350_ (_13678_, _13677_, _13674_);
  nor _64351_ (_13680_, _09043_, _13593_);
  or _64352_ (_13681_, _13594_, _09056_);
  or _64353_ (_13682_, _13681_, _13680_);
  and _64354_ (_13683_, _13682_, _09061_);
  and _64355_ (_13684_, _13683_, _13678_);
  nor _64356_ (_13685_, _08573_, _13593_);
  or _64357_ (_13686_, _13685_, _13594_);
  and _64358_ (_13687_, _13686_, _06528_);
  or _64359_ (_13688_, _13687_, _06568_);
  or _64360_ (_13689_, _13688_, _13684_);
  or _64361_ (_13691_, _13607_, _06926_);
  and _64362_ (_13692_, _13691_, _05928_);
  and _64363_ (_13693_, _13692_, _13689_);
  and _64364_ (_13694_, _13604_, _05927_);
  or _64365_ (_13695_, _13694_, _06278_);
  or _64366_ (_13696_, _13695_, _13693_);
  and _64367_ (_13697_, _08550_, _07900_);
  or _64368_ (_13698_, _13594_, _06279_);
  or _64369_ (_13699_, _13698_, _13697_);
  and _64370_ (_13700_, _13699_, _01347_);
  and _64371_ (_13702_, _13700_, _13696_);
  or _64372_ (_13703_, _13702_, _13592_);
  and _64373_ (_40593_, _13703_, _42618_);
  and _64374_ (_13704_, _01351_, \oc8051_golden_model_1.SCON [7]);
  not _64375_ (_13705_, _07973_);
  and _64376_ (_13706_, _13705_, \oc8051_golden_model_1.SCON [7]);
  and _64377_ (_13707_, _08575_, _07973_);
  or _64378_ (_13708_, _13707_, _13706_);
  and _64379_ (_13709_, _13708_, _06536_);
  nor _64380_ (_13710_, _08040_, _13705_);
  or _64381_ (_13712_, _13710_, _13706_);
  or _64382_ (_13713_, _13712_, _07215_);
  not _64383_ (_13714_, _08622_);
  and _64384_ (_13715_, _13714_, \oc8051_golden_model_1.SCON [7]);
  and _64385_ (_13716_, _08649_, _08622_);
  or _64386_ (_13717_, _13716_, _13715_);
  and _64387_ (_13718_, _13717_, _06268_);
  and _64388_ (_13719_, _08768_, _07973_);
  or _64389_ (_13720_, _13719_, _13706_);
  or _64390_ (_13721_, _13720_, _07151_);
  and _64391_ (_13723_, _07973_, \oc8051_golden_model_1.ACC [7]);
  or _64392_ (_13724_, _13723_, _13706_);
  and _64393_ (_13725_, _13724_, _07141_);
  and _64394_ (_13726_, _07142_, \oc8051_golden_model_1.SCON [7]);
  or _64395_ (_13727_, _13726_, _06341_);
  or _64396_ (_13728_, _13727_, _13725_);
  and _64397_ (_13729_, _13728_, _06273_);
  and _64398_ (_13730_, _13729_, _13721_);
  and _64399_ (_13731_, _08773_, _08622_);
  or _64400_ (_13732_, _13731_, _13715_);
  and _64401_ (_13734_, _13732_, _06272_);
  or _64402_ (_13735_, _13734_, _06461_);
  or _64403_ (_13736_, _13735_, _13730_);
  or _64404_ (_13737_, _13712_, _07166_);
  and _64405_ (_13738_, _13737_, _13736_);
  or _64406_ (_13739_, _13738_, _06464_);
  or _64407_ (_13740_, _13724_, _06465_);
  and _64408_ (_13741_, _13740_, _06269_);
  and _64409_ (_13742_, _13741_, _13739_);
  or _64410_ (_13743_, _13742_, _13718_);
  and _64411_ (_13745_, _13743_, _06262_);
  and _64412_ (_13746_, _08790_, _08622_);
  or _64413_ (_13747_, _13746_, _13715_);
  and _64414_ (_13748_, _13747_, _06261_);
  or _64415_ (_13749_, _13748_, _13745_);
  and _64416_ (_13750_, _13749_, _06258_);
  and _64417_ (_13751_, _08808_, _08622_);
  or _64418_ (_13752_, _13751_, _13715_);
  and _64419_ (_13753_, _13752_, _06257_);
  or _64420_ (_13754_, _13753_, _10080_);
  or _64421_ (_13756_, _13754_, _13750_);
  and _64422_ (_13757_, _13756_, _13713_);
  or _64423_ (_13758_, _13757_, _07460_);
  and _64424_ (_13759_, _08755_, _07973_);
  or _64425_ (_13760_, _13706_, _07208_);
  or _64426_ (_13761_, _13760_, _13759_);
  and _64427_ (_13762_, _13761_, _05982_);
  and _64428_ (_13763_, _13762_, _13758_);
  and _64429_ (_13764_, _09021_, _07973_);
  or _64430_ (_13765_, _13764_, _13706_);
  and _64431_ (_13766_, _13765_, _10094_);
  or _64432_ (_13767_, _13766_, _06218_);
  or _64433_ (_13768_, _13767_, _13763_);
  and _64434_ (_13769_, _08825_, _07973_);
  or _64435_ (_13770_, _13769_, _13706_);
  or _64436_ (_13771_, _13770_, _06219_);
  and _64437_ (_13772_, _13771_, _13768_);
  or _64438_ (_13773_, _13772_, _06369_);
  and _64439_ (_13774_, _09044_, _07973_);
  or _64440_ (_13775_, _13774_, _13706_);
  or _64441_ (_13776_, _13775_, _07237_);
  and _64442_ (_13777_, _13776_, _07240_);
  and _64443_ (_13778_, _13777_, _13773_);
  or _64444_ (_13779_, _13778_, _13709_);
  and _64445_ (_13780_, _13779_, _07242_);
  or _64446_ (_13781_, _13706_, _08043_);
  and _64447_ (_13782_, _13770_, _06375_);
  and _64448_ (_13783_, _13782_, _13781_);
  or _64449_ (_13784_, _13783_, _13780_);
  and _64450_ (_13785_, _13784_, _07234_);
  and _64451_ (_13786_, _13724_, _06545_);
  and _64452_ (_13787_, _13786_, _13781_);
  or _64453_ (_13788_, _13787_, _06366_);
  or _64454_ (_13789_, _13788_, _13785_);
  nor _64455_ (_13790_, _09043_, _13705_);
  or _64456_ (_13791_, _13706_, _09056_);
  or _64457_ (_13792_, _13791_, _13790_);
  and _64458_ (_13793_, _13792_, _09061_);
  and _64459_ (_13794_, _13793_, _13789_);
  nor _64460_ (_13795_, _08573_, _13705_);
  or _64461_ (_13796_, _13795_, _13706_);
  and _64462_ (_13797_, _13796_, _06528_);
  or _64463_ (_13798_, _13797_, _06568_);
  or _64464_ (_13799_, _13798_, _13794_);
  or _64465_ (_13800_, _13720_, _06926_);
  and _64466_ (_13801_, _13800_, _05928_);
  and _64467_ (_13802_, _13801_, _13799_);
  and _64468_ (_13803_, _13717_, _05927_);
  or _64469_ (_13804_, _13803_, _06278_);
  or _64470_ (_13805_, _13804_, _13802_);
  and _64471_ (_13806_, _08550_, _07973_);
  or _64472_ (_13807_, _13706_, _06279_);
  or _64473_ (_13808_, _13807_, _13806_);
  and _64474_ (_13809_, _13808_, _01347_);
  and _64475_ (_13810_, _13809_, _13805_);
  or _64476_ (_13811_, _13810_, _13704_);
  and _64477_ (_40594_, _13811_, _42618_);
  not _64478_ (_13812_, \oc8051_golden_model_1.SP [7]);
  nor _64479_ (_13813_, _01347_, _13812_);
  and _64480_ (_13814_, _07602_, \oc8051_golden_model_1.SP [4]);
  and _64481_ (_13815_, _13814_, \oc8051_golden_model_1.SP [5]);
  and _64482_ (_13816_, _13815_, \oc8051_golden_model_1.SP [6]);
  or _64483_ (_13817_, _13816_, \oc8051_golden_model_1.SP [7]);
  nand _64484_ (_13818_, _13816_, \oc8051_golden_model_1.SP [7]);
  and _64485_ (_13819_, _13818_, _13817_);
  or _64486_ (_13820_, _13819_, _07271_);
  nor _64487_ (_13821_, _07956_, _13812_);
  and _64488_ (_13822_, _08575_, _08173_);
  or _64489_ (_13823_, _13822_, _13821_);
  and _64490_ (_13824_, _13823_, _06536_);
  or _64491_ (_13825_, _13819_, _07494_);
  and _64492_ (_13826_, _08768_, _08173_);
  or _64493_ (_13827_, _13826_, _13821_);
  or _64494_ (_13828_, _13827_, _07151_);
  and _64495_ (_13829_, _07956_, \oc8051_golden_model_1.ACC [7]);
  or _64496_ (_13830_, _13829_, _13821_);
  or _64497_ (_13831_, _13830_, _07142_);
  or _64498_ (_13832_, _07141_, \oc8051_golden_model_1.SP [7]);
  and _64499_ (_13833_, _13832_, _07504_);
  and _64500_ (_13834_, _13833_, _13831_);
  and _64501_ (_13835_, _13819_, _06758_);
  or _64502_ (_13836_, _13835_, _06341_);
  or _64503_ (_13837_, _13836_, _13834_);
  and _64504_ (_13838_, _13837_, _06010_);
  and _64505_ (_13839_, _13838_, _13828_);
  and _64506_ (_13840_, _13819_, _07611_);
  or _64507_ (_13841_, _13840_, _06461_);
  or _64508_ (_13842_, _13841_, _13839_);
  not _64509_ (_13843_, \oc8051_golden_model_1.SP [6]);
  not _64510_ (_13844_, \oc8051_golden_model_1.SP [5]);
  not _64511_ (_13845_, \oc8051_golden_model_1.SP [4]);
  and _64512_ (_13846_, _08672_, _13845_);
  and _64513_ (_13847_, _13846_, _13844_);
  and _64514_ (_13848_, _13847_, _13843_);
  and _64515_ (_13849_, _13848_, _06800_);
  nor _64516_ (_13850_, _13849_, _13812_);
  and _64517_ (_13851_, _13849_, _13812_);
  nor _64518_ (_13852_, _13851_, _13850_);
  nand _64519_ (_13853_, _13852_, _06461_);
  and _64520_ (_13854_, _13853_, _13842_);
  or _64521_ (_13855_, _13854_, _06464_);
  or _64522_ (_13856_, _13830_, _06465_);
  and _64523_ (_13857_, _13856_, _07303_);
  and _64524_ (_13858_, _13857_, _13855_);
  and _64525_ (_13859_, _13815_, \oc8051_golden_model_1.SP [0]);
  and _64526_ (_13860_, _13859_, \oc8051_golden_model_1.SP [6]);
  nor _64527_ (_13861_, _13860_, _13812_);
  and _64528_ (_13862_, _13860_, _13812_);
  or _64529_ (_13863_, _13862_, _13861_);
  nand _64530_ (_13864_, _13863_, _06267_);
  nand _64531_ (_13865_, _13864_, _07494_);
  or _64532_ (_13866_, _13865_, _13858_);
  nand _64533_ (_13867_, _13866_, _13825_);
  and _64534_ (_13868_, _06350_, _05944_);
  nor _64535_ (_13869_, _13868_, _07214_);
  nand _64536_ (_13870_, _13869_, _13867_);
  and _64537_ (_13871_, _06337_, _05944_);
  not _64538_ (_13872_, _08173_);
  nor _64539_ (_13873_, _08040_, _13872_);
  or _64540_ (_13874_, _13873_, _13821_);
  nor _64541_ (_13875_, _13874_, _13869_);
  nor _64542_ (_13876_, _13875_, _13871_);
  and _64543_ (_13877_, _13876_, _13870_);
  and _64544_ (_13878_, _13874_, _13871_);
  or _64545_ (_13879_, _13878_, _07460_);
  or _64546_ (_13880_, _13879_, _13877_);
  or _64547_ (_13881_, _13821_, _07208_);
  and _64548_ (_13882_, _08755_, _07956_);
  or _64549_ (_13883_, _13882_, _13881_);
  and _64550_ (_13884_, _13883_, _05982_);
  and _64551_ (_13885_, _13884_, _13880_);
  and _64552_ (_13886_, _09021_, _08173_);
  or _64553_ (_13887_, _13886_, _13821_);
  and _64554_ (_13888_, _13887_, _10094_);
  or _64555_ (_13889_, _13888_, _06218_);
  or _64556_ (_13890_, _13889_, _13885_);
  and _64557_ (_13891_, _08825_, _07956_);
  or _64558_ (_13892_, _13891_, _13821_);
  or _64559_ (_13893_, _13892_, _06219_);
  and _64560_ (_13894_, _13893_, _13890_);
  or _64561_ (_13895_, _13894_, _06217_);
  or _64562_ (_13896_, _13819_, _05952_);
  and _64563_ (_13897_, _13896_, _13895_);
  or _64564_ (_13898_, _13897_, _06369_);
  and _64565_ (_13899_, _09044_, _07956_);
  or _64566_ (_13900_, _13899_, _13821_);
  or _64567_ (_13901_, _13900_, _07237_);
  and _64568_ (_13902_, _13901_, _07240_);
  and _64569_ (_13903_, _13902_, _13898_);
  or _64570_ (_13904_, _13903_, _13824_);
  and _64571_ (_13905_, _13904_, _07242_);
  or _64572_ (_13906_, _13821_, _08043_);
  and _64573_ (_13907_, _13892_, _06375_);
  and _64574_ (_13908_, _13907_, _13906_);
  or _64575_ (_13909_, _13908_, _13905_);
  and _64576_ (_13910_, _13909_, _12772_);
  and _64577_ (_13911_, _13830_, _06545_);
  and _64578_ (_13912_, _13911_, _13906_);
  and _64579_ (_13913_, _13819_, _07233_);
  or _64580_ (_13914_, _13913_, _06366_);
  or _64581_ (_13915_, _13914_, _13912_);
  or _64582_ (_13916_, _13915_, _13910_);
  and _64583_ (_13917_, _09063_, _07956_);
  or _64584_ (_13918_, _13917_, _13821_);
  or _64585_ (_13919_, _13918_, _09056_);
  and _64586_ (_13920_, _13919_, _13916_);
  or _64587_ (_13921_, _13920_, _06528_);
  nor _64588_ (_13922_, _08573_, _13872_);
  or _64589_ (_13923_, _13821_, _09061_);
  or _64590_ (_13924_, _13923_, _13922_);
  and _64591_ (_13925_, _13924_, _06716_);
  and _64592_ (_13926_, _13925_, _13921_);
  or _64593_ (_13927_, _13848_, \oc8051_golden_model_1.SP [7]);
  nand _64594_ (_13928_, _13848_, \oc8051_golden_model_1.SP [7]);
  and _64595_ (_13929_, _13928_, _13927_);
  and _64596_ (_13930_, _13929_, _06551_);
  or _64597_ (_13931_, _13930_, _07253_);
  or _64598_ (_13932_, _13931_, _13926_);
  or _64599_ (_13933_, _13819_, _05959_);
  and _64600_ (_13934_, _13933_, _13932_);
  or _64601_ (_13935_, _13934_, _06281_);
  or _64602_ (_13936_, _13929_, _06282_);
  and _64603_ (_13937_, _13936_, _06926_);
  and _64604_ (_13938_, _13937_, _13935_);
  and _64605_ (_13939_, _13827_, _06568_);
  or _64606_ (_13940_, _13939_, _07695_);
  or _64607_ (_13941_, _13940_, _13938_);
  and _64608_ (_13942_, _13941_, _13820_);
  or _64609_ (_13943_, _13942_, _06278_);
  and _64610_ (_13944_, _08550_, _08173_);
  or _64611_ (_13945_, _13821_, _06279_);
  or _64612_ (_13946_, _13945_, _13944_);
  and _64613_ (_13947_, _13946_, _01347_);
  and _64614_ (_13948_, _13947_, _13943_);
  or _64615_ (_13949_, _13948_, _13813_);
  and _64616_ (_40595_, _13949_, _42618_);
  and _64617_ (_13950_, _01351_, \oc8051_golden_model_1.SBUF [7]);
  not _64618_ (_13951_, _07886_);
  and _64619_ (_13952_, _13951_, \oc8051_golden_model_1.SBUF [7]);
  nor _64620_ (_13953_, _08573_, _13951_);
  or _64621_ (_13954_, _13953_, _13952_);
  and _64622_ (_13955_, _13954_, _06528_);
  and _64623_ (_13956_, _08575_, _07886_);
  or _64624_ (_13957_, _13956_, _13952_);
  and _64625_ (_13958_, _13957_, _06536_);
  nor _64626_ (_13959_, _08040_, _13951_);
  or _64627_ (_13960_, _13959_, _13952_);
  or _64628_ (_13961_, _13960_, _07215_);
  and _64629_ (_13962_, _08768_, _07886_);
  or _64630_ (_13963_, _13962_, _13952_);
  or _64631_ (_13964_, _13963_, _07151_);
  and _64632_ (_13965_, _07886_, \oc8051_golden_model_1.ACC [7]);
  or _64633_ (_13966_, _13965_, _13952_);
  and _64634_ (_13967_, _13966_, _07141_);
  and _64635_ (_13968_, _07142_, \oc8051_golden_model_1.SBUF [7]);
  or _64636_ (_13969_, _13968_, _06341_);
  or _64637_ (_13970_, _13969_, _13967_);
  and _64638_ (_13971_, _13970_, _07166_);
  and _64639_ (_13972_, _13971_, _13964_);
  and _64640_ (_13973_, _13960_, _06461_);
  or _64641_ (_13974_, _13973_, _13972_);
  and _64642_ (_13975_, _13974_, _06465_);
  and _64643_ (_13976_, _13966_, _06464_);
  or _64644_ (_13977_, _13976_, _10080_);
  or _64645_ (_13978_, _13977_, _13975_);
  and _64646_ (_13979_, _13978_, _13961_);
  or _64647_ (_13980_, _13979_, _07460_);
  and _64648_ (_13981_, _08755_, _07886_);
  or _64649_ (_13982_, _13952_, _07208_);
  or _64650_ (_13983_, _13982_, _13981_);
  and _64651_ (_13984_, _13983_, _05982_);
  and _64652_ (_13985_, _13984_, _13980_);
  and _64653_ (_13986_, _09021_, _07886_);
  or _64654_ (_13987_, _13986_, _13952_);
  and _64655_ (_13988_, _13987_, _10094_);
  or _64656_ (_13989_, _13988_, _06218_);
  or _64657_ (_13990_, _13989_, _13985_);
  and _64658_ (_13991_, _08825_, _07886_);
  or _64659_ (_13992_, _13991_, _13952_);
  or _64660_ (_13993_, _13992_, _06219_);
  and _64661_ (_13994_, _13993_, _13990_);
  or _64662_ (_13995_, _13994_, _06369_);
  and _64663_ (_13996_, _09044_, _07886_);
  or _64664_ (_13997_, _13996_, _13952_);
  or _64665_ (_13998_, _13997_, _07237_);
  and _64666_ (_13999_, _13998_, _07240_);
  and _64667_ (_14000_, _13999_, _13995_);
  or _64668_ (_14001_, _14000_, _13958_);
  and _64669_ (_14002_, _14001_, _07242_);
  or _64670_ (_14003_, _13952_, _08043_);
  and _64671_ (_14004_, _13992_, _06375_);
  and _64672_ (_14005_, _14004_, _14003_);
  or _64673_ (_14006_, _14005_, _14002_);
  and _64674_ (_14007_, _14006_, _07234_);
  and _64675_ (_14008_, _13966_, _06545_);
  and _64676_ (_14009_, _14008_, _14003_);
  or _64677_ (_14010_, _14009_, _06366_);
  or _64678_ (_14011_, _14010_, _14007_);
  nor _64679_ (_14012_, _09043_, _13951_);
  or _64680_ (_14013_, _13952_, _09056_);
  or _64681_ (_14014_, _14013_, _14012_);
  and _64682_ (_14015_, _14014_, _09061_);
  and _64683_ (_14016_, _14015_, _14011_);
  or _64684_ (_14017_, _14016_, _13955_);
  and _64685_ (_14018_, _14017_, _06926_);
  and _64686_ (_14019_, _13963_, _06568_);
  or _64687_ (_14020_, _14019_, _06278_);
  or _64688_ (_14021_, _14020_, _14018_);
  and _64689_ (_14022_, _08550_, _07886_);
  or _64690_ (_14023_, _13952_, _06279_);
  or _64691_ (_14024_, _14023_, _14022_);
  and _64692_ (_14025_, _14024_, _01347_);
  and _64693_ (_14026_, _14025_, _14021_);
  or _64694_ (_14027_, _14026_, _13950_);
  and _64695_ (_40597_, _14027_, _42618_);
  nor _64696_ (_14028_, _01347_, _10558_);
  nor _64697_ (_14029_, _08630_, _10558_);
  and _64698_ (_14030_, _08649_, _08630_);
  or _64699_ (_14031_, _14030_, _14029_);
  or _64700_ (_14032_, _14031_, _05928_);
  and _64701_ (_14033_, _10664_, _08552_);
  and _64702_ (_14034_, _10667_, \oc8051_golden_model_1.ACC [7]);
  or _64703_ (_14035_, _14034_, _11064_);
  or _64704_ (_14036_, _14035_, _14033_);
  or _64705_ (_14037_, _14036_, _11037_);
  nor _64706_ (_14038_, _07935_, _10558_);
  and _64707_ (_14039_, _08575_, _07935_);
  or _64708_ (_14040_, _14039_, _14038_);
  and _64709_ (_14041_, _14040_, _06536_);
  and _64710_ (_14042_, _09021_, _07935_);
  or _64711_ (_14043_, _14042_, _14038_);
  and _64712_ (_14044_, _14043_, _10094_);
  not _64713_ (_14045_, _07935_);
  nor _64714_ (_14046_, _08040_, _14045_);
  or _64715_ (_14047_, _14046_, _14038_);
  or _64716_ (_14048_, _14047_, _07215_);
  and _64717_ (_14049_, _10605_, _10601_);
  nor _64718_ (_14050_, _14049_, _10599_);
  nand _64719_ (_14051_, _10648_, _10601_);
  or _64720_ (_14052_, _14051_, _10646_);
  and _64721_ (_14053_, _14052_, _14050_);
  and _64722_ (_14054_, _10595_, _08755_);
  or _64723_ (_14055_, _14054_, _10588_);
  or _64724_ (_14056_, _14055_, _14053_);
  not _64725_ (_14057_, _06504_);
  not _64726_ (_14058_, _06505_);
  nor _64727_ (_14059_, _13004_, _14058_);
  and _64728_ (_14060_, _08773_, _08630_);
  or _64729_ (_14061_, _14060_, _14029_);
  or _64730_ (_14062_, _14029_, _08789_);
  and _64731_ (_14063_, _14062_, _06261_);
  and _64732_ (_14064_, _14063_, _14061_);
  and _64733_ (_14065_, _12366_, _12362_);
  or _64734_ (_14066_, _12363_, _14065_);
  and _64735_ (_14067_, _14066_, _12361_);
  and _64736_ (_14068_, _12358_, _12356_);
  or _64737_ (_14069_, _14068_, _12355_);
  or _64738_ (_14070_, _14069_, _14067_);
  and _64739_ (_14071_, _14070_, _12354_);
  or _64740_ (_14072_, _12350_, _12347_);
  and _64741_ (_14073_, _12345_, _14072_);
  and _64742_ (_14074_, _14073_, _12346_);
  and _64743_ (_14075_, _12343_, _08041_);
  or _64744_ (_14076_, _14075_, _12340_);
  or _64745_ (_14077_, _14076_, _14074_);
  or _64746_ (_14078_, _14077_, _14071_);
  nor _64747_ (_14079_, _12378_, _12371_);
  and _64748_ (_14080_, _14079_, _14078_);
  and _64749_ (_14081_, _08768_, _07935_);
  or _64750_ (_14082_, _14081_, _14038_);
  or _64751_ (_14083_, _14082_, _07151_);
  and _64752_ (_14084_, _07935_, \oc8051_golden_model_1.ACC [7]);
  or _64753_ (_14085_, _14084_, _14038_);
  and _64754_ (_14086_, _14085_, _07141_);
  nor _64755_ (_14087_, _07141_, _10558_);
  or _64756_ (_14088_, _14087_, _06341_);
  or _64757_ (_14089_, _14088_, _14086_);
  and _64758_ (_14090_, _14089_, _10776_);
  and _64759_ (_14091_, _14090_, _14083_);
  nor _64760_ (_14092_, _10795_, _10776_);
  or _64761_ (_14093_, _12540_, _06467_);
  or _64762_ (_14094_, _14093_, _14092_);
  or _64763_ (_14095_, _14094_, _14091_);
  or _64764_ (_14096_, _14061_, _06273_);
  or _64765_ (_14097_, _14047_, _07166_);
  and _64766_ (_14098_, _14097_, _14096_);
  and _64767_ (_14099_, _14098_, _14095_);
  or _64768_ (_14100_, _14099_, _06464_);
  or _64769_ (_14101_, _14085_, _06465_);
  nor _64770_ (_14102_, _12559_, _06268_);
  and _64771_ (_14103_, _14102_, _14101_);
  and _64772_ (_14104_, _14103_, _14100_);
  and _64773_ (_14105_, _14031_, _06268_);
  or _64774_ (_14106_, _14105_, _14104_);
  and _64775_ (_14107_, _14106_, _12378_);
  or _64776_ (_14108_, _14107_, _14080_);
  and _64777_ (_14109_, _14108_, _12177_);
  nand _64778_ (_14110_, _12329_, _12326_);
  nand _64779_ (_14111_, _14110_, _12325_);
  and _64780_ (_14112_, _14111_, _12324_);
  nand _64781_ (_14113_, _12321_, _12318_);
  and _64782_ (_14114_, _12319_, _14113_);
  or _64783_ (_14115_, _14114_, _14112_);
  and _64784_ (_14116_, _14115_, _12317_);
  nor _64785_ (_14117_, _12306_, _08802_);
  or _64786_ (_14118_, _14117_, _12304_);
  nand _64787_ (_14119_, _12314_, _12311_);
  and _64788_ (_14120_, _12309_, _14119_);
  and _64789_ (_14121_, _14120_, _12310_);
  or _64790_ (_14122_, _14121_, _14118_);
  or _64791_ (_14123_, _14122_, _14116_);
  and _64792_ (_14124_, _12335_, _06347_);
  and _64793_ (_14125_, _14124_, _14123_);
  or _64794_ (_14126_, _14125_, _14109_);
  and _64795_ (_14127_, _14126_, _06774_);
  nand _64796_ (_14128_, _08246_, \oc8051_golden_model_1.ACC [5]);
  nor _64797_ (_14129_, _08246_, \oc8051_golden_model_1.ACC [5]);
  nor _64798_ (_14130_, _08543_, \oc8051_golden_model_1.ACC [4]);
  or _64799_ (_14131_, _14130_, _14129_);
  and _64800_ (_14132_, _14131_, _14128_);
  and _64801_ (_14133_, _14132_, _12585_);
  nor _64802_ (_14134_, _08042_, \oc8051_golden_model_1.ACC [7]);
  or _64803_ (_14135_, _08144_, \oc8051_golden_model_1.ACC [6]);
  nor _64804_ (_14136_, _14135_, _08575_);
  or _64805_ (_14137_, _14136_, _14134_);
  or _64806_ (_14138_, _14137_, _14133_);
  nand _64807_ (_14139_, _08291_, \oc8051_golden_model_1.ACC [3]);
  nor _64808_ (_14140_, _08291_, \oc8051_golden_model_1.ACC [3]);
  nor _64809_ (_14141_, _08439_, \oc8051_golden_model_1.ACC [2]);
  or _64810_ (_14142_, _14141_, _14140_);
  and _64811_ (_14143_, _14142_, _14139_);
  nor _64812_ (_14144_, _08340_, \oc8051_golden_model_1.ACC [1]);
  nor _64813_ (_14145_, _08390_, _06097_);
  nor _64814_ (_14146_, _14145_, _11262_);
  or _64815_ (_14147_, _14146_, _14144_);
  and _64816_ (_14148_, _14147_, _12578_);
  or _64817_ (_14149_, _14148_, _14143_);
  and _64818_ (_14150_, _14149_, _12586_);
  or _64819_ (_14151_, _14150_, _14138_);
  nor _64820_ (_14152_, _12587_, _06774_);
  and _64821_ (_14153_, _14152_, _14151_);
  or _64822_ (_14154_, _14153_, _14127_);
  and _64823_ (_14155_, _14154_, _12176_);
  and _64824_ (_14156_, _06251_, \oc8051_golden_model_1.ACC [0]);
  nor _64825_ (_14157_, _14156_, _11303_);
  or _64826_ (_14158_, _14157_, _11304_);
  and _64827_ (_14159_, _14158_, _12595_);
  nand _64828_ (_14160_, _06213_, \oc8051_golden_model_1.ACC [3]);
  nor _64829_ (_14161_, _06213_, \oc8051_golden_model_1.ACC [3]);
  nor _64830_ (_14162_, _06656_, \oc8051_golden_model_1.ACC [2]);
  or _64831_ (_14163_, _14162_, _14161_);
  and _64832_ (_14164_, _14163_, _14160_);
  or _64833_ (_14165_, _14164_, _14159_);
  and _64834_ (_14166_, _14165_, _12603_);
  nand _64835_ (_14167_, _06611_, \oc8051_golden_model_1.ACC [5]);
  nor _64836_ (_14168_, _06611_, \oc8051_golden_model_1.ACC [5]);
  nor _64837_ (_14169_, _06968_, \oc8051_golden_model_1.ACC [4]);
  or _64838_ (_14170_, _14169_, _14168_);
  and _64839_ (_14171_, _14170_, _14167_);
  and _64840_ (_14172_, _14171_, _12602_);
  and _64841_ (_14173_, _06182_, _08572_);
  or _64842_ (_14174_, _06317_, \oc8051_golden_model_1.ACC [6]);
  nor _64843_ (_14175_, _14174_, _10961_);
  or _64844_ (_14176_, _14175_, _14173_);
  or _64845_ (_14177_, _14176_, _14172_);
  or _64846_ (_14178_, _14177_, _14166_);
  nor _64847_ (_14179_, _12604_, _12176_);
  and _64848_ (_14180_, _14179_, _14178_);
  or _64849_ (_14181_, _14180_, _12174_);
  or _64850_ (_14182_, _14181_, _14155_);
  nand _64851_ (_14183_, _12174_, \oc8051_golden_model_1.PSW [7]);
  and _64852_ (_14184_, _14183_, _06262_);
  and _64853_ (_14185_, _14184_, _14182_);
  nor _64854_ (_14186_, _14185_, _14064_);
  nor _64855_ (_14187_, _14186_, _06455_);
  and _64856_ (_14188_, _06455_, \oc8051_golden_model_1.PSW [7]);
  and _64857_ (_14189_, _14188_, _13004_);
  or _64858_ (_14190_, _14189_, _14187_);
  nor _64859_ (_14191_, _09531_, _06505_);
  and _64860_ (_14192_, _14191_, _14190_);
  or _64861_ (_14193_, _14192_, _14059_);
  and _64862_ (_14194_, _14193_, _14057_);
  and _64863_ (_14195_, _06886_, _05976_);
  and _64864_ (_14196_, _06350_, _05976_);
  nor _64865_ (_14197_, _14196_, _14195_);
  nand _64866_ (_14198_, _14197_, _10731_);
  or _64867_ (_14199_, _13004_, \oc8051_golden_model_1.PSW [7]);
  and _64868_ (_14200_, _14199_, _06504_);
  or _64869_ (_14201_, _14200_, _14198_);
  or _64870_ (_14202_, _14201_, _14194_);
  and _64871_ (_14203_, _06337_, _05976_);
  not _64872_ (_14204_, _14203_);
  and _64873_ (_14205_, _10675_, _10670_);
  nor _64874_ (_14206_, _14205_, _10668_);
  nand _64875_ (_14207_, _10721_, _10670_);
  or _64876_ (_14208_, _14207_, _10719_);
  and _64877_ (_14209_, _14208_, _14206_);
  or _64878_ (_14210_, _14209_, _14033_);
  and _64879_ (_14211_, _14210_, _14204_);
  or _64880_ (_14212_, _14211_, _10735_);
  and _64881_ (_14213_, _14212_, _14202_);
  and _64882_ (_14214_, _14210_, _14203_);
  or _64883_ (_14215_, _14214_, _10656_);
  or _64884_ (_14216_, _14215_, _14213_);
  and _64885_ (_14217_, _14216_, _14056_);
  or _64886_ (_14218_, _14217_, _06512_);
  and _64887_ (_14219_, _10850_, _10846_);
  nor _64888_ (_14220_, _14219_, _10844_);
  nand _64889_ (_14221_, _10892_, _10846_);
  or _64890_ (_14222_, _14221_, _10890_);
  and _64891_ (_14223_, _14222_, _14220_);
  and _64892_ (_14224_, _10840_, _08043_);
  or _64893_ (_14225_, _14224_, _06517_);
  or _64894_ (_14226_, _14225_, _14223_);
  and _64895_ (_14227_, _14226_, _10517_);
  and _64896_ (_14228_, _14227_, _14218_);
  and _64897_ (_14229_, _10519_, _07941_);
  and _64898_ (_14230_, _10531_, _10527_);
  nor _64899_ (_14231_, _14230_, _10525_);
  nand _64900_ (_14232_, _10578_, _10527_);
  or _64901_ (_14233_, _14232_, _10576_);
  and _64902_ (_14234_, _14233_, _14231_);
  or _64903_ (_14235_, _14234_, _14229_);
  and _64904_ (_14236_, _14235_, _10516_);
  or _64905_ (_14237_, _14236_, _10080_);
  or _64906_ (_14238_, _14237_, _14228_);
  and _64907_ (_14239_, _14238_, _14048_);
  or _64908_ (_14240_, _14239_, _07460_);
  and _64909_ (_14241_, _08755_, _07935_);
  or _64910_ (_14242_, _14038_, _07208_);
  or _64911_ (_14243_, _14242_, _14241_);
  and _64912_ (_14244_, _14243_, _05982_);
  and _64913_ (_14245_, _14244_, _14240_);
  or _64914_ (_14246_, _14245_, _14044_);
  nor _64915_ (_14247_, _10093_, _06323_);
  and _64916_ (_14248_, _14247_, _14246_);
  nor _64917_ (_14249_, _13004_, _10558_);
  and _64918_ (_14250_, _14249_, _06323_);
  or _64919_ (_14251_, _14250_, _06218_);
  or _64920_ (_14252_, _14251_, _14248_);
  and _64921_ (_14253_, _08825_, _07935_);
  or _64922_ (_14254_, _14253_, _14038_);
  or _64923_ (_14255_, _14254_, _06219_);
  and _64924_ (_14256_, _14255_, _14252_);
  or _64925_ (_14257_, _14256_, _06322_);
  nand _64926_ (_14258_, _13004_, _10558_);
  or _64927_ (_14259_, _14258_, _06881_);
  and _64928_ (_14260_, _14259_, _14257_);
  or _64929_ (_14261_, _14260_, _06369_);
  and _64930_ (_14262_, _09044_, _07935_);
  or _64931_ (_14263_, _14262_, _14038_);
  or _64932_ (_14264_, _14263_, _07237_);
  and _64933_ (_14265_, _14264_, _07240_);
  and _64934_ (_14266_, _14265_, _14261_);
  or _64935_ (_14267_, _14266_, _14041_);
  and _64936_ (_14268_, _14267_, _07242_);
  or _64937_ (_14269_, _14038_, _08043_);
  and _64938_ (_14270_, _14254_, _06375_);
  and _64939_ (_14271_, _14270_, _14269_);
  or _64940_ (_14272_, _14271_, _14268_);
  and _64941_ (_14273_, _14272_, _07234_);
  and _64942_ (_14274_, _14085_, _06545_);
  and _64943_ (_14275_, _14274_, _14269_);
  or _64944_ (_14276_, _14275_, _06366_);
  or _64945_ (_14277_, _14276_, _14273_);
  nor _64946_ (_14278_, _09043_, _14045_);
  or _64947_ (_14279_, _14038_, _09056_);
  or _64948_ (_14280_, _14279_, _14278_);
  and _64949_ (_14281_, _14280_, _09061_);
  and _64950_ (_14282_, _14281_, _14277_);
  not _64951_ (_14283_, _11037_);
  nor _64952_ (_14284_, _08573_, _14045_);
  or _64953_ (_14285_, _14284_, _14038_);
  and _64954_ (_14286_, _14285_, _06528_);
  or _64955_ (_14287_, _14286_, _14283_);
  or _64956_ (_14288_, _14287_, _14282_);
  and _64957_ (_14289_, _14288_, _14037_);
  or _64958_ (_14290_, _14289_, _11041_);
  or _64959_ (_14291_, _11069_, _14054_);
  nor _64960_ (_14292_, _10598_, _08572_);
  or _64961_ (_14293_, _14292_, _11091_);
  or _64962_ (_14294_, _14293_, _14291_);
  and _64963_ (_14295_, _14294_, _06541_);
  and _64964_ (_14296_, _14295_, _14290_);
  not _64965_ (_14297_, _12153_);
  nor _64966_ (_14298_, _10843_, _08572_);
  or _64967_ (_14299_, _14298_, _11119_);
  or _64968_ (_14300_, _11097_, _14224_);
  or _64969_ (_14301_, _14300_, _14299_);
  and _64970_ (_14302_, _14301_, _14297_);
  or _64971_ (_14303_, _14302_, _14296_);
  and _64972_ (_14304_, _10524_, \oc8051_golden_model_1.ACC [7]);
  or _64973_ (_14305_, _14304_, _11147_);
  or _64974_ (_14306_, _11127_, _14229_);
  or _64975_ (_14307_, _14306_, _14305_);
  and _64976_ (_14308_, _14307_, _11126_);
  and _64977_ (_14309_, _14308_, _14303_);
  nand _64978_ (_14310_, _11125_, \oc8051_golden_model_1.ACC [7]);
  nand _64979_ (_14311_, _14310_, _11157_);
  or _64980_ (_14312_, _14311_, _14309_);
  and _64981_ (_14313_, _11192_, _10505_);
  not _64982_ (_14314_, _10494_);
  or _64983_ (_14315_, _11160_, _10504_);
  and _64984_ (_14316_, _14315_, _14314_);
  or _64985_ (_14317_, _14316_, _11157_);
  or _64986_ (_14318_, _14317_, _14313_);
  and _64987_ (_14319_, _14318_, _14312_);
  or _64988_ (_14320_, _14319_, _11201_);
  and _64989_ (_14321_, _11235_, _10500_);
  nor _64990_ (_14322_, _11204_, _10499_);
  nor _64991_ (_14323_, _14322_, _10498_);
  or _64992_ (_14324_, _14323_, _11203_);
  or _64993_ (_14325_, _14324_, _14321_);
  and _64994_ (_14326_, _14325_, _06285_);
  and _64995_ (_14327_, _14326_, _14320_);
  not _64996_ (_14328_, _08573_);
  not _64997_ (_14329_, _08574_);
  nand _64998_ (_14330_, _11277_, _14329_);
  and _64999_ (_14331_, _14330_, _06283_);
  and _65000_ (_14332_, _14331_, _14328_);
  or _65001_ (_14333_, _14332_, _11243_);
  or _65002_ (_14334_, _14333_, _14327_);
  nor _65003_ (_14335_, _11319_, _10959_);
  or _65004_ (_14336_, _14335_, _11321_);
  or _65005_ (_14337_, _14336_, _10960_);
  and _65006_ (_14338_, _14337_, _14334_);
  or _65007_ (_14339_, _14338_, _06568_);
  nor _65008_ (_14340_, _14082_, _06926_);
  nor _65009_ (_14341_, _14340_, _11335_);
  and _65010_ (_14342_, _14341_, _14339_);
  and _65011_ (_14343_, _11335_, \oc8051_golden_model_1.ACC [0]);
  or _65012_ (_14344_, _14343_, _05927_);
  or _65013_ (_14345_, _14344_, _14342_);
  and _65014_ (_14346_, _14345_, _14032_);
  or _65015_ (_14347_, _14346_, _06278_);
  and _65016_ (_14348_, _08550_, _07935_);
  or _65017_ (_14349_, _14038_, _06279_);
  or _65018_ (_14350_, _14349_, _14348_);
  and _65019_ (_14351_, _14350_, _01347_);
  and _65020_ (_14352_, _14351_, _14347_);
  or _65021_ (_14353_, _14352_, _14028_);
  and _65022_ (_40598_, _14353_, _42618_);
  and _65023_ (_14354_, _07535_, _07289_);
  nor _65024_ (_14355_, _14354_, _07537_);
  nor _65025_ (_14356_, _07711_, _07536_);
  nor _65026_ (_14357_, _14356_, _07859_);
  and _65027_ (_14358_, _14357_, _07535_);
  and _65028_ (_14359_, _14358_, _14355_);
  not _65029_ (_14360_, _14359_);
  nand _65030_ (_14361_, _05940_, _05630_);
  nand _65031_ (_14362_, _12580_, _09062_);
  or _65032_ (_14363_, _08390_, _08954_);
  and _65033_ (_14364_, _08390_, _08954_);
  not _65034_ (_14365_, _14364_);
  and _65035_ (_14366_, _14365_, _14363_);
  and _65036_ (_14367_, _14366_, _07238_);
  nor _65037_ (_14368_, _05978_, _05630_);
  or _65038_ (_14369_, _08390_, _06501_);
  nor _65039_ (_14370_, _12925_, _12901_);
  or _65040_ (_14371_, _14370_, _08610_);
  nor _65041_ (_14372_, _08390_, _08652_);
  nand _65042_ (_14373_, _12387_, _07133_);
  nand _65043_ (_14374_, _06758_, _05630_);
  or _65044_ (_14375_, _06758_, \oc8051_golden_model_1.ACC [0]);
  nand _65045_ (_14376_, _14375_, _14374_);
  and _65046_ (_14377_, _14376_, _08654_);
  nor _65047_ (_14378_, _14377_, _07152_);
  and _65048_ (_14379_, _14378_, _14373_);
  or _65049_ (_14380_, _14379_, _14372_);
  and _65050_ (_14381_, _14380_, _08651_);
  nand _65051_ (_14382_, _12925_, _12902_);
  and _65052_ (_14383_, _14382_, _06275_);
  or _65053_ (_14384_, _14383_, _07611_);
  or _65054_ (_14385_, _14384_, _14381_);
  nor _65055_ (_14386_, _06010_, \oc8051_golden_model_1.PC [0]);
  nor _65056_ (_14387_, _14386_, _07167_);
  and _65057_ (_14388_, _14387_, _14385_);
  and _65058_ (_14389_, _07167_, _07133_);
  or _65059_ (_14390_, _14389_, _07179_);
  or _65060_ (_14391_, _14390_, _14388_);
  and _65061_ (_14392_, _14391_, _14371_);
  or _65062_ (_14393_, _14392_, _06267_);
  or _65063_ (_14394_, _08390_, _07303_);
  and _65064_ (_14395_, _14394_, _06265_);
  and _65065_ (_14396_, _14395_, _14393_);
  nand _65066_ (_14397_, _14382_, _06264_);
  nor _65067_ (_14398_, _14397_, _12926_);
  or _65068_ (_14399_, _14398_, _14396_);
  and _65069_ (_14400_, _14399_, _06007_);
  or _65070_ (_14401_, _06007_, _05630_);
  nand _65071_ (_14402_, _06501_, _14401_);
  or _65072_ (_14403_, _14402_, _14400_);
  and _65073_ (_14404_, _14403_, _14369_);
  or _65074_ (_14405_, _14404_, _07197_);
  and _65075_ (_14406_, _09392_, _06286_);
  nand _65076_ (_14407_, _08387_, _07197_);
  or _65077_ (_14408_, _14407_, _14406_);
  and _65078_ (_14409_, _14408_, _14405_);
  or _65079_ (_14410_, _14409_, _07196_);
  and _65080_ (_14411_, _07889_, \oc8051_golden_model_1.PSW [7]);
  and _65081_ (_14412_, _14411_, _06656_);
  or _65082_ (_14413_, _14412_, _14370_);
  or _65083_ (_14414_, _14413_, _08801_);
  and _65084_ (_14415_, _14414_, _05978_);
  and _65085_ (_14416_, _14415_, _14410_);
  or _65086_ (_14417_, _14416_, _14368_);
  and _65087_ (_14418_, _14417_, _08817_);
  and _65088_ (_14419_, _08812_, _07133_);
  or _65089_ (_14420_, _14419_, _08816_);
  or _65090_ (_14421_, _14420_, _14418_);
  or _65091_ (_14422_, _09392_, _08821_);
  and _65092_ (_14423_, _14422_, _07471_);
  and _65093_ (_14424_, _14423_, _14421_);
  and _65094_ (_14425_, _08608_, _07133_);
  and _65095_ (_14426_, _08957_, \oc8051_golden_model_1.TMOD [0]);
  and _65096_ (_14427_, _08968_, \oc8051_golden_model_1.B [0]);
  or _65097_ (_14428_, _14427_, _14426_);
  and _65098_ (_14429_, _08944_, \oc8051_golden_model_1.P0 [0]);
  and _65099_ (_14430_, _08950_, \oc8051_golden_model_1.ACC [0]);
  or _65100_ (_14431_, _14430_, _14429_);
  or _65101_ (_14432_, _14431_, _14428_);
  and _65102_ (_14433_, _08934_, \oc8051_golden_model_1.TCON [0]);
  and _65103_ (_14434_, _08965_, \oc8051_golden_model_1.SCON [0]);
  or _65104_ (_14435_, _14434_, _14433_);
  and _65105_ (_14436_, _08939_, \oc8051_golden_model_1.TL0 [0]);
  and _65106_ (_14437_, _09007_, \oc8051_golden_model_1.PSW [0]);
  or _65107_ (_14438_, _14437_, _14436_);
  or _65108_ (_14439_, _14438_, _14435_);
  or _65109_ (_14440_, _14439_, _14432_);
  and _65110_ (_14441_, _08977_, \oc8051_golden_model_1.PCON [0]);
  and _65111_ (_14442_, _08979_, \oc8051_golden_model_1.DPH [0]);
  or _65112_ (_14443_, _14442_, _14441_);
  or _65113_ (_14444_, _14443_, _14440_);
  and _65114_ (_14445_, _09013_, \oc8051_golden_model_1.TH0 [0]);
  and _65115_ (_14446_, _09015_, \oc8051_golden_model_1.TH1 [0]);
  and _65116_ (_14447_, _08988_, \oc8051_golden_model_1.SP [0]);
  or _65117_ (_14448_, _14447_, _14446_);
  or _65118_ (_14449_, _14448_, _14445_);
  and _65119_ (_14450_, _08999_, \oc8051_golden_model_1.P2 [0]);
  and _65120_ (_14451_, _08993_, \oc8051_golden_model_1.IE [0]);
  or _65121_ (_14452_, _14451_, _14450_);
  and _65122_ (_14453_, _09001_, \oc8051_golden_model_1.P3 [0]);
  and _65123_ (_14454_, _08996_, \oc8051_golden_model_1.IP [0]);
  or _65124_ (_14455_, _14454_, _14453_);
  or _65125_ (_14456_, _14455_, _14452_);
  and _65126_ (_14457_, _08962_, \oc8051_golden_model_1.P1 [0]);
  and _65127_ (_14458_, _09005_, \oc8051_golden_model_1.SBUF [0]);
  or _65128_ (_14459_, _14458_, _14457_);
  or _65129_ (_14460_, _14459_, _14456_);
  and _65130_ (_14461_, _08984_, \oc8051_golden_model_1.DPL [0]);
  and _65131_ (_14462_, _08986_, \oc8051_golden_model_1.TL1 [0]);
  or _65132_ (_14463_, _14462_, _14461_);
  or _65133_ (_14464_, _14463_, _14460_);
  or _65134_ (_14465_, _14464_, _14449_);
  or _65135_ (_14466_, _14465_, _14444_);
  or _65136_ (_14467_, _14466_, _14425_);
  and _65137_ (_14468_, _14467_, _07470_);
  or _65138_ (_14469_, _14468_, _09031_);
  or _65139_ (_14470_, _14469_, _14424_);
  and _65140_ (_14471_, _09031_, _06251_);
  nor _65141_ (_14472_, _14471_, _06220_);
  and _65142_ (_14473_, _14472_, _14470_);
  and _65143_ (_14474_, _08954_, _06220_);
  or _65144_ (_14475_, _14474_, _06217_);
  or _65145_ (_14476_, _14475_, _14473_);
  nor _65146_ (_14477_, _05952_, \oc8051_golden_model_1.PC [0]);
  nor _65147_ (_14478_, _14477_, _07238_);
  and _65148_ (_14479_, _14478_, _14476_);
  or _65149_ (_14480_, _14479_, _14367_);
  and _65150_ (_14481_, _14480_, _08577_);
  nor _65151_ (_14482_, _12581_, _08577_);
  or _65152_ (_14483_, _14482_, _14481_);
  and _65153_ (_14484_, _14483_, _08571_);
  and _65154_ (_14485_, _14364_, _07243_);
  or _65155_ (_14486_, _14485_, _14484_);
  and _65156_ (_14487_, _14486_, _07236_);
  and _65157_ (_14488_, _11263_, _07235_);
  or _65158_ (_14489_, _14488_, _07233_);
  or _65159_ (_14490_, _14489_, _14487_);
  nor _65160_ (_14491_, _05961_, \oc8051_golden_model_1.PC [0]);
  nor _65161_ (_14492_, _14491_, _09057_);
  and _65162_ (_14493_, _14492_, _14490_);
  and _65163_ (_14494_, _14363_, _09057_);
  or _65164_ (_14495_, _14494_, _09062_);
  or _65165_ (_14496_, _14495_, _14493_);
  and _65166_ (_14497_, _14496_, _14362_);
  or _65167_ (_14498_, _14497_, _07253_);
  or _65168_ (_14499_, _05959_, \oc8051_golden_model_1.PC [0]);
  and _65169_ (_14500_, _14499_, _08569_);
  and _65170_ (_14501_, _14500_, _14498_);
  or _65171_ (_14502_, _08569_, _07133_);
  nand _65172_ (_14503_, _14502_, _07264_);
  or _65173_ (_14504_, _14503_, _14501_);
  nand _65174_ (_14505_, _09392_, _07435_);
  and _65175_ (_14506_, _14505_, _14504_);
  or _65176_ (_14507_, _14506_, _07261_);
  not _65177_ (_14508_, _06361_);
  nand _65178_ (_14509_, _08390_, _07261_);
  and _65179_ (_14510_, _14509_, _14508_);
  and _65180_ (_14511_, _14510_, _14507_);
  and _65181_ (_14512_, _06361_, _05630_);
  or _65182_ (_14513_, _14512_, _05940_);
  or _65183_ (_14514_, _14513_, _14511_);
  and _65184_ (_14515_, _14514_, _14361_);
  or _65185_ (_14516_, _14515_, _07270_);
  or _65186_ (_14517_, _14370_, _07539_);
  and _65187_ (_14518_, _14517_, _09427_);
  and _65188_ (_14519_, _14518_, _14516_);
  nor _65189_ (_14520_, _09427_, _07133_);
  or _65190_ (_14521_, _14520_, _14519_);
  and _65191_ (_14522_, _14521_, _07282_);
  nor _65192_ (_14523_, _09392_, _07282_);
  or _65193_ (_14524_, _14523_, _07286_);
  or _65194_ (_14525_, _14524_, _14522_);
  nand _65195_ (_14526_, _08390_, _07286_);
  and _65196_ (_14527_, _14526_, _07535_);
  and _65197_ (_14528_, _14527_, _14525_);
  or _65198_ (_14529_, _14528_, _14360_);
  or _65199_ (_14530_, _14359_, \oc8051_golden_model_1.IRAM[0] [0]);
  not _65200_ (_14531_, _07872_);
  and _65201_ (_14532_, _07872_, _07866_);
  nor _65202_ (_14533_, _07873_, _14532_);
  nand _65203_ (_14534_, _14533_, _07296_);
  or _65204_ (_14535_, _14534_, _14531_);
  and _65205_ (_14536_, _14535_, _14530_);
  and _65206_ (_14537_, _14536_, _14529_);
  and _65207_ (_14538_, _07872_, _07296_);
  and _65208_ (_14539_, _14538_, _14533_);
  nand _65209_ (_14540_, _12276_, _06361_);
  or _65210_ (_14541_, _12431_, _06361_);
  and _65211_ (_14542_, _14541_, _14540_);
  and _65212_ (_14543_, _14542_, _07872_);
  and _65213_ (_14544_, _14543_, _14539_);
  or _65214_ (_40612_, _14544_, _14537_);
  nor _65215_ (_14545_, _09452_, _09394_);
  or _65216_ (_14546_, _14545_, _07282_);
  not _65217_ (_14547_, _08565_);
  or _65218_ (_14548_, _09433_, _08556_);
  and _65219_ (_14549_, _14548_, _07061_);
  or _65220_ (_14550_, _14549_, _14547_);
  nor _65221_ (_14551_, _05959_, \oc8051_golden_model_1.PC [1]);
  or _65222_ (_14552_, _05952_, _05597_);
  or _65223_ (_14553_, _09347_, _06182_);
  nand _65224_ (_14554_, _14553_, _08338_);
  and _65225_ (_14555_, _14554_, _07197_);
  not _65226_ (_14556_, _12872_);
  nand _65227_ (_14557_, _12871_, _12849_);
  and _65228_ (_14558_, _14557_, _06264_);
  and _65229_ (_14559_, _14558_, _14556_);
  nor _65230_ (_14560_, _12871_, _08172_);
  or _65231_ (_14561_, _14560_, _08610_);
  nor _65232_ (_14562_, _08761_, _08391_);
  nand _65233_ (_14563_, _14562_, _07152_);
  and _65234_ (_14564_, _14548_, _12387_);
  nor _65235_ (_14565_, _06758_, _06042_);
  and _65236_ (_14566_, _06758_, _05597_);
  or _65237_ (_14567_, _14566_, _14565_);
  and _65238_ (_14568_, _14567_, _08654_);
  or _65239_ (_14569_, _14568_, _07152_);
  or _65240_ (_14570_, _14569_, _14564_);
  and _65241_ (_14571_, _14570_, _14563_);
  or _65242_ (_14572_, _14571_, _06275_);
  or _65243_ (_14573_, _14557_, _08651_);
  and _65244_ (_14574_, _14573_, _14572_);
  or _65245_ (_14575_, _14574_, _07611_);
  nor _65246_ (_14576_, _06010_, _05597_);
  nor _65247_ (_14577_, _14576_, _07167_);
  and _65248_ (_14578_, _14577_, _14575_);
  and _65249_ (_14579_, _09432_, _07167_);
  or _65250_ (_14580_, _14579_, _07179_);
  or _65251_ (_14581_, _14580_, _14578_);
  and _65252_ (_14582_, _14581_, _14561_);
  or _65253_ (_14583_, _14582_, _06267_);
  nand _65254_ (_14584_, _08340_, _06267_);
  and _65255_ (_14585_, _14584_, _06265_);
  and _65256_ (_14586_, _14585_, _14583_);
  or _65257_ (_14587_, _14586_, _14559_);
  and _65258_ (_14588_, _14587_, _06007_);
  or _65259_ (_14589_, _06007_, \oc8051_golden_model_1.PC [1]);
  nand _65260_ (_14590_, _06501_, _14589_);
  or _65261_ (_14591_, _14590_, _14588_);
  nand _65262_ (_14592_, _08340_, _06502_);
  and _65263_ (_14593_, _14592_, _07198_);
  and _65264_ (_14594_, _14593_, _14591_);
  or _65265_ (_14595_, _14594_, _14555_);
  and _65266_ (_14596_, _14595_, _08801_);
  nand _65267_ (_14597_, _08172_, _10558_);
  and _65268_ (_14598_, _14597_, _07196_);
  and _65269_ (_14599_, _14598_, _14557_);
  or _65270_ (_14600_, _14599_, _06254_);
  or _65271_ (_14601_, _14600_, _14596_);
  nor _65272_ (_14602_, _05978_, _05597_);
  nor _65273_ (_14603_, _14602_, _08812_);
  and _65274_ (_14604_, _14603_, _14601_);
  nor _65275_ (_14605_, _07357_, _08817_);
  or _65276_ (_14606_, _14605_, _08816_);
  or _65277_ (_14607_, _14606_, _14604_);
  or _65278_ (_14608_, _09451_, _08821_);
  and _65279_ (_14609_, _14608_, _07471_);
  and _65280_ (_14610_, _14609_, _14607_);
  nor _65281_ (_14611_, _08825_, _07357_);
  and _65282_ (_14612_, _08977_, \oc8051_golden_model_1.PCON [1]);
  and _65283_ (_14613_, _08979_, \oc8051_golden_model_1.DPH [1]);
  or _65284_ (_14614_, _14613_, _14612_);
  and _65285_ (_14615_, _08934_, \oc8051_golden_model_1.TCON [1]);
  and _65286_ (_14616_, _08957_, \oc8051_golden_model_1.TMOD [1]);
  or _65287_ (_14617_, _14616_, _14615_);
  and _65288_ (_14618_, _08939_, \oc8051_golden_model_1.TL0 [1]);
  and _65289_ (_14619_, _08962_, \oc8051_golden_model_1.P1 [1]);
  or _65290_ (_14620_, _14619_, _14618_);
  or _65291_ (_14621_, _14620_, _14617_);
  and _65292_ (_14622_, _08944_, \oc8051_golden_model_1.P0 [1]);
  and _65293_ (_14623_, _08950_, \oc8051_golden_model_1.ACC [1]);
  or _65294_ (_14624_, _14623_, _14622_);
  and _65295_ (_14625_, _08968_, \oc8051_golden_model_1.B [1]);
  and _65296_ (_14626_, _09007_, \oc8051_golden_model_1.PSW [1]);
  or _65297_ (_14627_, _14626_, _14625_);
  or _65298_ (_14628_, _14627_, _14624_);
  or _65299_ (_14629_, _14628_, _14621_);
  or _65300_ (_14630_, _14629_, _14614_);
  and _65301_ (_14631_, _08986_, \oc8051_golden_model_1.TL1 [1]);
  and _65302_ (_14632_, _09015_, \oc8051_golden_model_1.TH1 [1]);
  and _65303_ (_14633_, _08988_, \oc8051_golden_model_1.SP [1]);
  or _65304_ (_14634_, _14633_, _14632_);
  or _65305_ (_14635_, _14634_, _14631_);
  and _65306_ (_14636_, _09001_, \oc8051_golden_model_1.P3 [1]);
  and _65307_ (_14637_, _08996_, \oc8051_golden_model_1.IP [1]);
  or _65308_ (_14638_, _14637_, _14636_);
  and _65309_ (_14639_, _08999_, \oc8051_golden_model_1.P2 [1]);
  and _65310_ (_14640_, _08993_, \oc8051_golden_model_1.IE [1]);
  or _65311_ (_14641_, _14640_, _14639_);
  or _65312_ (_14642_, _14641_, _14638_);
  and _65313_ (_14643_, _08965_, \oc8051_golden_model_1.SCON [1]);
  and _65314_ (_14644_, _09005_, \oc8051_golden_model_1.SBUF [1]);
  or _65315_ (_14645_, _14644_, _14643_);
  or _65316_ (_14646_, _14645_, _14642_);
  and _65317_ (_14647_, _08984_, \oc8051_golden_model_1.DPL [1]);
  and _65318_ (_14648_, _09013_, \oc8051_golden_model_1.TH0 [1]);
  or _65319_ (_14649_, _14648_, _14647_);
  or _65320_ (_14650_, _14649_, _14646_);
  or _65321_ (_14651_, _14650_, _14635_);
  or _65322_ (_14652_, _14651_, _14630_);
  or _65323_ (_14653_, _14652_, _14611_);
  and _65324_ (_14654_, _14653_, _07470_);
  or _65325_ (_14655_, _14654_, _09031_);
  or _65326_ (_14656_, _14655_, _14610_);
  and _65327_ (_14657_, _09031_, _07004_);
  nor _65328_ (_14658_, _14657_, _06220_);
  and _65329_ (_14659_, _14658_, _14656_);
  and _65330_ (_14660_, _08936_, _06220_);
  or _65331_ (_14661_, _14660_, _06217_);
  or _65332_ (_14662_, _14661_, _14659_);
  and _65333_ (_14663_, _14662_, _14552_);
  or _65334_ (_14664_, _14663_, _07238_);
  nand _65335_ (_14665_, _08340_, _07038_);
  nor _65336_ (_14666_, _08340_, _07038_);
  not _65337_ (_14667_, _14666_);
  and _65338_ (_14668_, _14667_, _14665_);
  or _65339_ (_14669_, _14668_, _07239_);
  and _65340_ (_14670_, _14669_, _08577_);
  and _65341_ (_14671_, _14670_, _14664_);
  and _65342_ (_14672_, _11262_, _07241_);
  or _65343_ (_14673_, _14672_, _07243_);
  or _65344_ (_14674_, _14673_, _14671_);
  or _65345_ (_14675_, _14666_, _08571_);
  and _65346_ (_14676_, _14675_, _07236_);
  and _65347_ (_14677_, _14676_, _14674_);
  and _65348_ (_14678_, _11260_, _07235_);
  or _65349_ (_14679_, _14678_, _07233_);
  or _65350_ (_14680_, _14679_, _14677_);
  nor _65351_ (_14681_, _05961_, _05597_);
  nor _65352_ (_14682_, _14681_, _09057_);
  and _65353_ (_14683_, _14682_, _14680_);
  and _65354_ (_14684_, _14665_, _09057_);
  or _65355_ (_14685_, _14684_, _09062_);
  or _65356_ (_14686_, _14685_, _14683_);
  nand _65357_ (_14687_, _11261_, _09062_);
  and _65358_ (_14688_, _14687_, _05959_);
  and _65359_ (_14689_, _14688_, _14686_);
  nor _65360_ (_14690_, _14689_, _14551_);
  nor _65361_ (_14691_, _14690_, _06701_);
  and _65362_ (_14692_, _14548_, _06701_);
  or _65363_ (_14693_, _14692_, _06754_);
  or _65364_ (_14694_, _14693_, _14691_);
  not _65365_ (_14695_, _06754_);
  or _65366_ (_14696_, _14548_, _14695_);
  and _65367_ (_14697_, _14696_, _07062_);
  and _65368_ (_14698_, _14697_, _14694_);
  or _65369_ (_14699_, _14698_, _14550_);
  not _65370_ (_14700_, _07292_);
  or _65371_ (_14701_, _14548_, _14700_);
  and _65372_ (_14702_, _14701_, _07264_);
  and _65373_ (_14703_, _14702_, _14699_);
  nor _65374_ (_14704_, _14545_, _07264_);
  or _65375_ (_14705_, _14704_, _14703_);
  and _65376_ (_14706_, _14705_, _09075_);
  nor _65377_ (_14707_, _14562_, _09075_);
  or _65378_ (_14708_, _14707_, _06361_);
  or _65379_ (_14709_, _14708_, _14706_);
  not _65380_ (_14710_, _05940_);
  nand _65381_ (_14711_, _06361_, _06111_);
  and _65382_ (_14712_, _14711_, _14710_);
  and _65383_ (_14713_, _14712_, _14709_);
  and _65384_ (_14714_, _05940_, _05597_);
  or _65385_ (_14715_, _07270_, _14714_);
  or _65386_ (_14716_, _14715_, _14713_);
  or _65387_ (_14717_, _14560_, _07539_);
  and _65388_ (_14718_, _14717_, _09427_);
  and _65389_ (_14719_, _14718_, _14716_);
  nor _65390_ (_14720_, _14548_, _09427_);
  or _65391_ (_14721_, _14720_, _07281_);
  or _65392_ (_14722_, _14721_, _14719_);
  and _65393_ (_14723_, _14722_, _14546_);
  or _65394_ (_14724_, _14723_, _07286_);
  or _65395_ (_14725_, _14562_, _09445_);
  and _65396_ (_14726_, _14725_, _07535_);
  and _65397_ (_14727_, _14726_, _14724_);
  or _65398_ (_14728_, _14727_, _14360_);
  or _65399_ (_14729_, _14359_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _65400_ (_14730_, _14729_, _14535_);
  and _65401_ (_14731_, _14730_, _14728_);
  nand _65402_ (_14732_, _12217_, _06361_);
  or _65403_ (_14733_, _12426_, _06361_);
  and _65404_ (_14734_, _14733_, _14732_);
  and _65405_ (_14735_, _14734_, _07872_);
  and _65406_ (_14736_, _14735_, _14539_);
  or _65407_ (_40613_, _14736_, _14731_);
  not _65408_ (_14737_, _07279_);
  nor _65409_ (_14738_, _09452_, _09450_);
  nor _65410_ (_14739_, _14738_, _09453_);
  and _65411_ (_14740_, _14739_, _07280_);
  not _65412_ (_14741_, _07280_);
  nor _65413_ (_14742_, _09433_, _09431_);
  nor _65414_ (_14743_, _14742_, _09434_);
  and _65415_ (_14744_, _14743_, _09424_);
  not _65416_ (_14745_, _07262_);
  not _65417_ (_14746_, _07263_);
  nor _65418_ (_14747_, _06085_, _05959_);
  nand _65419_ (_14748_, _08439_, _06697_);
  nor _65420_ (_14749_, _08439_, _06697_);
  not _65421_ (_14750_, _14749_);
  and _65422_ (_14751_, _14750_, _14748_);
  and _65423_ (_14752_, _14751_, _07238_);
  or _65424_ (_14753_, _09302_, _06182_);
  nand _65425_ (_14754_, _14753_, _08437_);
  and _65426_ (_14755_, _14754_, _07197_);
  nor _65427_ (_14756_, _12847_, _07959_);
  or _65428_ (_14757_, _14756_, _08610_);
  and _65429_ (_14758_, _08556_, _07776_);
  nor _65430_ (_14759_, _08556_, _07776_);
  or _65431_ (_14760_, _14759_, _14758_);
  or _65432_ (_14761_, _14760_, _08654_);
  nor _65433_ (_14762_, _06758_, _10213_);
  and _65434_ (_14763_, _06758_, _06079_);
  nor _65435_ (_14764_, _14763_, _14762_);
  nand _65436_ (_14765_, _14764_, _08654_);
  and _65437_ (_14766_, _14765_, _14761_);
  and _65438_ (_14767_, _14766_, _08652_);
  and _65439_ (_14768_, _08761_, _08439_);
  nor _65440_ (_14769_, _08761_, _08439_);
  or _65441_ (_14770_, _14769_, _14768_);
  and _65442_ (_14771_, _14770_, _07152_);
  or _65443_ (_14772_, _14771_, _14767_);
  and _65444_ (_14773_, _14772_, _08651_);
  nand _65445_ (_14774_, _12847_, _12825_);
  and _65446_ (_14775_, _14774_, _06275_);
  or _65447_ (_14776_, _14775_, _07611_);
  or _65448_ (_14777_, _14776_, _14773_);
  nor _65449_ (_14778_, _06079_, _06010_);
  nor _65450_ (_14779_, _14778_, _07167_);
  and _65451_ (_14780_, _14779_, _14777_);
  and _65452_ (_14781_, _09431_, _07167_);
  or _65453_ (_14782_, _14781_, _07179_);
  or _65454_ (_14783_, _14782_, _14780_);
  and _65455_ (_14784_, _14783_, _14757_);
  or _65456_ (_14785_, _14784_, _06267_);
  nand _65457_ (_14786_, _08439_, _06267_);
  and _65458_ (_14787_, _14786_, _06265_);
  and _65459_ (_14788_, _14787_, _14785_);
  not _65460_ (_14789_, _12848_);
  and _65461_ (_14790_, _14774_, _14789_);
  and _65462_ (_14791_, _14790_, _06264_);
  or _65463_ (_14792_, _14791_, _14788_);
  and _65464_ (_14793_, _14792_, _06007_);
  or _65465_ (_14794_, _06085_, _06007_);
  nand _65466_ (_14795_, _06501_, _14794_);
  or _65467_ (_14796_, _14795_, _14793_);
  nand _65468_ (_14797_, _08439_, _06502_);
  and _65469_ (_14798_, _14797_, _07198_);
  and _65470_ (_14799_, _14798_, _14796_);
  or _65471_ (_14800_, _14799_, _14755_);
  and _65472_ (_14801_, _14800_, _08801_);
  and _65473_ (_14802_, _07917_, \oc8051_golden_model_1.PSW [7]);
  and _65474_ (_14803_, _14802_, _06656_);
  or _65475_ (_14804_, _14803_, _14756_);
  and _65476_ (_14805_, _14804_, _07196_);
  or _65477_ (_14806_, _14805_, _06254_);
  or _65478_ (_14807_, _14806_, _14801_);
  nor _65479_ (_14808_, _06079_, _05978_);
  nor _65480_ (_14809_, _14808_, _08812_);
  and _65481_ (_14810_, _14809_, _14807_);
  nor _65482_ (_14811_, _07776_, _08817_);
  or _65483_ (_14812_, _14811_, _08816_);
  or _65484_ (_14813_, _14812_, _14810_);
  or _65485_ (_14814_, _09450_, _08821_);
  and _65486_ (_14815_, _14814_, _07471_);
  and _65487_ (_14816_, _14815_, _14813_);
  nor _65488_ (_14817_, _08825_, _07776_);
  and _65489_ (_14818_, _08962_, \oc8051_golden_model_1.P1 [2]);
  and _65490_ (_14819_, _08965_, \oc8051_golden_model_1.SCON [2]);
  or _65491_ (_14820_, _14819_, _14818_);
  and _65492_ (_14821_, _08957_, \oc8051_golden_model_1.TMOD [2]);
  and _65493_ (_14822_, _08939_, \oc8051_golden_model_1.TL0 [2]);
  or _65494_ (_14823_, _14822_, _14821_);
  or _65495_ (_14824_, _14823_, _14820_);
  and _65496_ (_14825_, _08934_, \oc8051_golden_model_1.TCON [2]);
  and _65497_ (_14826_, _09007_, \oc8051_golden_model_1.PSW [2]);
  or _65498_ (_14827_, _14826_, _14825_);
  and _65499_ (_14828_, _09005_, \oc8051_golden_model_1.SBUF [2]);
  and _65500_ (_14829_, _08968_, \oc8051_golden_model_1.B [2]);
  or _65501_ (_14830_, _14829_, _14828_);
  or _65502_ (_14831_, _14830_, _14827_);
  or _65503_ (_14832_, _14831_, _14824_);
  and _65504_ (_14833_, _08977_, \oc8051_golden_model_1.PCON [2]);
  and _65505_ (_14834_, _08979_, \oc8051_golden_model_1.DPH [2]);
  or _65506_ (_14835_, _14834_, _14833_);
  or _65507_ (_14836_, _14835_, _14832_);
  and _65508_ (_14837_, _08986_, \oc8051_golden_model_1.TL1 [2]);
  and _65509_ (_14838_, _09015_, \oc8051_golden_model_1.TH1 [2]);
  or _65510_ (_14839_, _14838_, _14837_);
  and _65511_ (_14840_, _08988_, \oc8051_golden_model_1.SP [2]);
  or _65512_ (_14841_, _14840_, _14839_);
  and _65513_ (_14842_, _08993_, \oc8051_golden_model_1.IE [2]);
  and _65514_ (_14843_, _08996_, \oc8051_golden_model_1.IP [2]);
  or _65515_ (_14844_, _14843_, _14842_);
  and _65516_ (_14845_, _08999_, \oc8051_golden_model_1.P2 [2]);
  and _65517_ (_14846_, _09001_, \oc8051_golden_model_1.P3 [2]);
  or _65518_ (_14847_, _14846_, _14845_);
  or _65519_ (_14848_, _14847_, _14844_);
  and _65520_ (_14849_, _08944_, \oc8051_golden_model_1.P0 [2]);
  and _65521_ (_14850_, _08950_, \oc8051_golden_model_1.ACC [2]);
  or _65522_ (_14851_, _14850_, _14849_);
  or _65523_ (_14852_, _14851_, _14848_);
  and _65524_ (_14853_, _08984_, \oc8051_golden_model_1.DPL [2]);
  and _65525_ (_14854_, _09013_, \oc8051_golden_model_1.TH0 [2]);
  or _65526_ (_14855_, _14854_, _14853_);
  or _65527_ (_14856_, _14855_, _14852_);
  or _65528_ (_14857_, _14856_, _14841_);
  or _65529_ (_14858_, _14857_, _14836_);
  or _65530_ (_14859_, _14858_, _14817_);
  and _65531_ (_14860_, _14859_, _07470_);
  or _65532_ (_14861_, _14860_, _09031_);
  or _65533_ (_14862_, _14861_, _14816_);
  and _65534_ (_14863_, _09031_, _06656_);
  nor _65535_ (_14864_, _14863_, _06220_);
  and _65536_ (_14865_, _14864_, _14862_);
  and _65537_ (_14866_, _08973_, _06220_);
  or _65538_ (_14867_, _14866_, _06217_);
  or _65539_ (_14868_, _14867_, _14865_);
  nor _65540_ (_14869_, _06079_, _05952_);
  nor _65541_ (_14870_, _14869_, _07238_);
  and _65542_ (_14871_, _14870_, _14868_);
  or _65543_ (_14872_, _14871_, _14752_);
  and _65544_ (_14873_, _14872_, _08577_);
  and _65545_ (_14874_, _11259_, _07241_);
  or _65546_ (_14875_, _14874_, _14873_);
  and _65547_ (_14876_, _14875_, _08571_);
  and _65548_ (_14877_, _14749_, _07243_);
  or _65549_ (_14878_, _14877_, _14876_);
  and _65550_ (_14879_, _14878_, _07236_);
  and _65551_ (_14880_, _11257_, _07235_);
  or _65552_ (_14881_, _14880_, _07233_);
  or _65553_ (_14882_, _14881_, _14879_);
  nor _65554_ (_14883_, _06079_, _05961_);
  nor _65555_ (_14884_, _14883_, _09057_);
  and _65556_ (_14885_, _14884_, _14882_);
  and _65557_ (_14886_, _14748_, _09057_);
  or _65558_ (_14887_, _14886_, _09062_);
  or _65559_ (_14888_, _14887_, _14885_);
  nand _65560_ (_14889_, _11258_, _09062_);
  and _65561_ (_14890_, _14889_, _05959_);
  and _65562_ (_14891_, _14890_, _14888_);
  or _65563_ (_14892_, _14891_, _14747_);
  and _65564_ (_14893_, _14892_, _08569_);
  not _65565_ (_14894_, _08569_);
  and _65566_ (_14895_, _14760_, _14894_);
  or _65567_ (_14896_, _14895_, _14893_);
  and _65568_ (_14897_, _14896_, _14746_);
  nor _65569_ (_14898_, _09394_, _09302_);
  or _65570_ (_14899_, _14898_, _09395_);
  and _65571_ (_14900_, _14899_, _07263_);
  or _65572_ (_14901_, _14900_, _14897_);
  and _65573_ (_14902_, _14901_, _14745_);
  and _65574_ (_14903_, _14899_, _07262_);
  or _65575_ (_14904_, _14903_, _14902_);
  and _65576_ (_14905_, _14904_, _09075_);
  and _65577_ (_14906_, _14770_, _07261_);
  or _65578_ (_14907_, _14906_, _06361_);
  or _65579_ (_14908_, _14907_, _14905_);
  nand _65580_ (_14909_, _12248_, _06361_);
  and _65581_ (_14910_, _14909_, _14710_);
  and _65582_ (_14911_, _14910_, _14908_);
  and _65583_ (_14912_, _06079_, _05940_);
  or _65584_ (_14913_, _07270_, _14912_);
  or _65585_ (_14914_, _14913_, _14911_);
  or _65586_ (_14915_, _14756_, _07539_);
  and _65587_ (_14916_, _14915_, _09427_);
  and _65588_ (_14917_, _14916_, _14914_);
  or _65589_ (_14918_, _14917_, _14744_);
  and _65590_ (_14919_, _14918_, _14741_);
  or _65591_ (_14920_, _14919_, _14740_);
  and _65592_ (_14921_, _14920_, _14737_);
  and _65593_ (_14922_, _14739_, _07279_);
  or _65594_ (_14923_, _14922_, _07286_);
  or _65595_ (_14924_, _14923_, _14921_);
  nor _65596_ (_14925_, _08440_, _08391_);
  nor _65597_ (_14926_, _14925_, _08441_);
  or _65598_ (_14927_, _14926_, _09445_);
  and _65599_ (_14928_, _14927_, _07535_);
  and _65600_ (_14929_, _14928_, _14924_);
  or _65601_ (_14930_, _14929_, _14360_);
  or _65602_ (_14931_, _14359_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _65603_ (_14932_, _14931_, _14535_);
  and _65604_ (_14933_, _14932_, _14930_);
  nand _65605_ (_14934_, _12203_, _06361_);
  or _65606_ (_14935_, _12421_, _06361_);
  and _65607_ (_14936_, _14935_, _14934_);
  and _65608_ (_14937_, _14936_, _07872_);
  and _65609_ (_14938_, _14937_, _14539_);
  or _65610_ (_40614_, _14938_, _14933_);
  nor _65611_ (_14939_, _05959_, _06033_);
  nand _65612_ (_14940_, _08291_, _06452_);
  nor _65613_ (_14941_, _08291_, _06452_);
  not _65614_ (_14942_, _14941_);
  and _65615_ (_14943_, _14942_, _14940_);
  and _65616_ (_14944_, _14943_, _07238_);
  or _65617_ (_14945_, _09257_, _06182_);
  nand _65618_ (_14946_, _14945_, _08289_);
  and _65619_ (_14947_, _14946_, _07197_);
  nor _65620_ (_14948_, _12975_, _08185_);
  or _65621_ (_14949_, _14948_, _08610_);
  nand _65622_ (_14950_, _12975_, _12953_);
  or _65623_ (_14951_, _14950_, _08651_);
  nor _65624_ (_14952_, _14768_, _08291_);
  or _65625_ (_14953_, _14952_, _08763_);
  and _65626_ (_14954_, _14953_, _07152_);
  nor _65627_ (_14955_, _14758_, _07594_);
  nor _65628_ (_14956_, _14955_, _08557_);
  nand _65629_ (_14957_, _14956_, _12387_);
  and _65630_ (_14958_, _06758_, _05932_);
  nor _65631_ (_14959_, _06758_, _06055_);
  nor _65632_ (_14960_, _14959_, _14958_);
  and _65633_ (_14961_, _14960_, _08654_);
  nor _65634_ (_14962_, _14961_, _07152_);
  and _65635_ (_14963_, _14962_, _14957_);
  or _65636_ (_14964_, _14963_, _06275_);
  or _65637_ (_14965_, _14964_, _14954_);
  and _65638_ (_14966_, _14965_, _14951_);
  or _65639_ (_14967_, _14966_, _07611_);
  nor _65640_ (_14968_, _06010_, _05932_);
  nor _65641_ (_14969_, _14968_, _07167_);
  and _65642_ (_14970_, _14969_, _14967_);
  and _65643_ (_14971_, _07595_, _07167_);
  or _65644_ (_14972_, _14971_, _07179_);
  or _65645_ (_14973_, _14972_, _14970_);
  and _65646_ (_14974_, _14973_, _14949_);
  or _65647_ (_14975_, _14974_, _06267_);
  nand _65648_ (_14976_, _08291_, _06267_);
  and _65649_ (_14977_, _14976_, _06265_);
  and _65650_ (_14978_, _14977_, _14975_);
  not _65651_ (_14979_, _12976_);
  and _65652_ (_14980_, _14950_, _14979_);
  and _65653_ (_14981_, _14980_, _06264_);
  or _65654_ (_14982_, _14981_, _14978_);
  and _65655_ (_14983_, _14982_, _06007_);
  or _65656_ (_14984_, _06007_, _06033_);
  nand _65657_ (_14985_, _06501_, _14984_);
  or _65658_ (_14986_, _14985_, _14983_);
  nand _65659_ (_14987_, _08291_, _06502_);
  and _65660_ (_14988_, _14987_, _07198_);
  and _65661_ (_14989_, _14988_, _14986_);
  or _65662_ (_14990_, _14989_, _14947_);
  and _65663_ (_14991_, _14990_, _08801_);
  nand _65664_ (_14992_, _08185_, _10558_);
  and _65665_ (_14993_, _14992_, _07196_);
  and _65666_ (_14994_, _14993_, _14950_);
  or _65667_ (_14995_, _14994_, _06254_);
  or _65668_ (_14996_, _14995_, _14991_);
  nor _65669_ (_14997_, _05978_, _05932_);
  nor _65670_ (_14998_, _14997_, _08812_);
  and _65671_ (_14999_, _14998_, _14996_);
  nor _65672_ (_15000_, _07594_, _08817_);
  or _65673_ (_15001_, _15000_, _08816_);
  or _65674_ (_15002_, _15001_, _14999_);
  or _65675_ (_15003_, _09449_, _08821_);
  and _65676_ (_15004_, _15003_, _07471_);
  and _65677_ (_15005_, _15004_, _15002_);
  nor _65678_ (_15006_, _08825_, _07594_);
  and _65679_ (_15007_, _08944_, \oc8051_golden_model_1.P0 [3]);
  and _65680_ (_15008_, _08962_, \oc8051_golden_model_1.P1 [3]);
  or _65681_ (_15009_, _15008_, _15007_);
  and _65682_ (_15010_, _08939_, \oc8051_golden_model_1.TL0 [3]);
  and _65683_ (_15011_, _08950_, \oc8051_golden_model_1.ACC [3]);
  or _65684_ (_15012_, _15011_, _15010_);
  or _65685_ (_15013_, _15012_, _15009_);
  and _65686_ (_15014_, _08934_, \oc8051_golden_model_1.TCON [3]);
  and _65687_ (_15015_, _08957_, \oc8051_golden_model_1.TMOD [3]);
  or _65688_ (_15016_, _15015_, _15014_);
  and _65689_ (_15017_, _08965_, \oc8051_golden_model_1.SCON [3]);
  and _65690_ (_15018_, _09005_, \oc8051_golden_model_1.SBUF [3]);
  or _65691_ (_15019_, _15018_, _15017_);
  or _65692_ (_15020_, _15019_, _15016_);
  or _65693_ (_15021_, _15020_, _15013_);
  and _65694_ (_15022_, _08977_, \oc8051_golden_model_1.PCON [3]);
  and _65695_ (_15023_, _08979_, \oc8051_golden_model_1.DPH [3]);
  or _65696_ (_15024_, _15023_, _15022_);
  or _65697_ (_15025_, _15024_, _15021_);
  and _65698_ (_15026_, _09015_, \oc8051_golden_model_1.TH1 [3]);
  and _65699_ (_15027_, _08984_, \oc8051_golden_model_1.DPL [3]);
  and _65700_ (_15028_, _08986_, \oc8051_golden_model_1.TL1 [3]);
  or _65701_ (_15029_, _15028_, _15027_);
  or _65702_ (_15030_, _15029_, _15026_);
  and _65703_ (_15031_, _08999_, \oc8051_golden_model_1.P2 [3]);
  and _65704_ (_15032_, _08996_, \oc8051_golden_model_1.IP [3]);
  or _65705_ (_15033_, _15032_, _15031_);
  and _65706_ (_15034_, _08993_, \oc8051_golden_model_1.IE [3]);
  and _65707_ (_15035_, _09001_, \oc8051_golden_model_1.P3 [3]);
  or _65708_ (_15036_, _15035_, _15034_);
  or _65709_ (_15037_, _15036_, _15033_);
  and _65710_ (_15038_, _08968_, \oc8051_golden_model_1.B [3]);
  and _65711_ (_15039_, _09007_, \oc8051_golden_model_1.PSW [3]);
  or _65712_ (_15040_, _15039_, _15038_);
  or _65713_ (_15041_, _15040_, _15037_);
  and _65714_ (_15042_, _09013_, \oc8051_golden_model_1.TH0 [3]);
  and _65715_ (_15043_, _08988_, \oc8051_golden_model_1.SP [3]);
  or _65716_ (_15044_, _15043_, _15042_);
  or _65717_ (_15045_, _15044_, _15041_);
  or _65718_ (_15046_, _15045_, _15030_);
  or _65719_ (_15047_, _15046_, _15025_);
  or _65720_ (_15048_, _15047_, _15006_);
  and _65721_ (_15049_, _15048_, _07470_);
  or _65722_ (_15050_, _15049_, _09031_);
  or _65723_ (_15051_, _15050_, _15005_);
  and _65724_ (_15052_, _09031_, _06213_);
  nor _65725_ (_15053_, _15052_, _06220_);
  and _65726_ (_15054_, _15053_, _15051_);
  and _65727_ (_15055_, _08930_, _06220_);
  or _65728_ (_15056_, _15055_, _06217_);
  or _65729_ (_15057_, _15056_, _15054_);
  nor _65730_ (_15058_, _05952_, _05932_);
  nor _65731_ (_15059_, _15058_, _07238_);
  and _65732_ (_15060_, _15059_, _15057_);
  or _65733_ (_15061_, _15060_, _14944_);
  and _65734_ (_15062_, _15061_, _08577_);
  and _65735_ (_15063_, _12577_, _07241_);
  or _65736_ (_15064_, _15063_, _15062_);
  and _65737_ (_15065_, _15064_, _08571_);
  and _65738_ (_15066_, _14941_, _07243_);
  or _65739_ (_15067_, _15066_, _15065_);
  and _65740_ (_15068_, _15067_, _07236_);
  and _65741_ (_15069_, _11255_, _07235_);
  or _65742_ (_15070_, _15069_, _07233_);
  or _65743_ (_15071_, _15070_, _15068_);
  nor _65744_ (_15072_, _05961_, _05932_);
  nor _65745_ (_15073_, _15072_, _09057_);
  and _65746_ (_15074_, _15073_, _15071_);
  and _65747_ (_15075_, _14940_, _09057_);
  or _65748_ (_15076_, _15075_, _09062_);
  or _65749_ (_15077_, _15076_, _15074_);
  nand _65750_ (_15078_, _11256_, _09062_);
  and _65751_ (_15079_, _15078_, _05959_);
  and _65752_ (_15080_, _15079_, _15077_);
  or _65753_ (_15081_, _15080_, _14939_);
  and _65754_ (_15082_, _15081_, _08568_);
  nor _65755_ (_15083_, _14956_, _08568_);
  or _65756_ (_15084_, _15083_, _07292_);
  or _65757_ (_15085_, _15084_, _15082_);
  nand _65758_ (_15086_, _14956_, _14547_);
  and _65759_ (_15087_, _15086_, _14746_);
  and _65760_ (_15088_, _15087_, _15085_);
  nor _65761_ (_15089_, _09395_, _09257_);
  or _65762_ (_15090_, _15089_, _09396_);
  or _65763_ (_15091_, _15090_, _07262_);
  and _65764_ (_15092_, _15091_, _07435_);
  or _65765_ (_15093_, _15092_, _15088_);
  or _65766_ (_15094_, _15090_, _14745_);
  and _65767_ (_15095_, _15094_, _09075_);
  and _65768_ (_15096_, _15095_, _15093_);
  and _65769_ (_15097_, _14953_, _07261_);
  or _65770_ (_15098_, _15097_, _06361_);
  or _65771_ (_15099_, _15098_, _15096_);
  nand _65772_ (_15100_, _12243_, _06361_);
  and _65773_ (_15101_, _15100_, _14710_);
  and _65774_ (_15102_, _15101_, _15099_);
  and _65775_ (_15103_, _05940_, _05932_);
  or _65776_ (_15104_, _07270_, _15103_);
  or _65777_ (_15105_, _15104_, _15102_);
  and _65778_ (_15106_, _07041_, _05938_);
  nor _65779_ (_15107_, _15106_, _07510_);
  or _65780_ (_15108_, _14948_, _07539_);
  and _65781_ (_15109_, _15108_, _15107_);
  and _65782_ (_15110_, _15109_, _15105_);
  not _65783_ (_15111_, _15107_);
  nor _65784_ (_15112_, _09434_, _07595_);
  nor _65785_ (_15113_, _15112_, _09435_);
  and _65786_ (_15114_, _15113_, _15111_);
  and _65787_ (_15115_, _10732_, _05938_);
  or _65788_ (_15116_, _15115_, _15114_);
  or _65789_ (_15117_, _15116_, _15110_);
  not _65790_ (_15118_, _15115_);
  or _65791_ (_15119_, _15118_, _15113_);
  and _65792_ (_15120_, _15119_, _07282_);
  and _65793_ (_15121_, _15120_, _15117_);
  or _65794_ (_15122_, _09453_, _09449_);
  nor _65795_ (_15123_, _09454_, _07282_);
  and _65796_ (_15124_, _15123_, _15122_);
  or _65797_ (_15125_, _15124_, _07286_);
  or _65798_ (_15126_, _15125_, _15121_);
  nor _65799_ (_15127_, _08441_, _08292_);
  nor _65800_ (_15128_, _15127_, _08442_);
  or _65801_ (_15129_, _15128_, _09445_);
  and _65802_ (_15130_, _15129_, _07535_);
  and _65803_ (_15131_, _15130_, _15126_);
  or _65804_ (_15132_, _15131_, _14360_);
  or _65805_ (_15133_, _14359_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _65806_ (_15134_, _15133_, _14535_);
  and _65807_ (_15135_, _15134_, _15132_);
  nand _65808_ (_15136_, _12208_, _06361_);
  or _65809_ (_15137_, _12417_, _06361_);
  and _65810_ (_15138_, _15137_, _15136_);
  and _65811_ (_15139_, _15138_, _07872_);
  and _65812_ (_15140_, _15139_, _14539_);
  or _65813_ (_40615_, _15140_, _15135_);
  nor _65814_ (_15141_, _09396_, _09212_);
  or _65815_ (_15142_, _15141_, _09397_);
  and _65816_ (_15143_, _15142_, _07263_);
  or _65817_ (_15144_, _12451_, _05952_);
  nor _65818_ (_15145_, _12452_, _05978_);
  and _65819_ (_15146_, _12451_, _06758_);
  nor _65820_ (_15147_, _06758_, _10135_);
  or _65821_ (_15148_, _15147_, _15146_);
  and _65822_ (_15149_, _15148_, _08654_);
  and _65823_ (_15150_, _08557_, _08541_);
  nor _65824_ (_15151_, _08557_, _08541_);
  or _65825_ (_15152_, _15151_, _15150_);
  and _65826_ (_15153_, _15152_, _12387_);
  or _65827_ (_15154_, _15153_, _15149_);
  and _65828_ (_15155_, _15154_, _07155_);
  and _65829_ (_15156_, _09448_, _07154_);
  or _65830_ (_15157_, _15156_, _15155_);
  and _65831_ (_15159_, _15157_, _08652_);
  and _65832_ (_15160_, _08763_, _08543_);
  nor _65833_ (_15161_, _08763_, _08543_);
  or _65834_ (_15162_, _15161_, _15160_);
  and _65835_ (_15163_, _15162_, _07152_);
  or _65836_ (_15164_, _15163_, _15159_);
  and _65837_ (_15165_, _15164_, _08651_);
  nand _65838_ (_15166_, _12897_, _12895_);
  and _65839_ (_15167_, _15166_, _06275_);
  or _65840_ (_15168_, _15167_, _07611_);
  or _65841_ (_15169_, _15168_, _15165_);
  nor _65842_ (_15170_, _12451_, _06010_);
  nor _65843_ (_15171_, _15170_, _07167_);
  and _65844_ (_15172_, _15171_, _15169_);
  and _65845_ (_15173_, _09430_, _07167_);
  or _65846_ (_15174_, _15173_, _07179_);
  or _65847_ (_15175_, _15174_, _15172_);
  nor _65848_ (_15176_, _12896_, _12895_);
  or _65849_ (_15177_, _15176_, _08610_);
  and _65850_ (_15178_, _15177_, _15175_);
  or _65851_ (_15179_, _15178_, _06267_);
  nand _65852_ (_15180_, _08543_, _06267_);
  and _65853_ (_15181_, _15180_, _06265_);
  and _65854_ (_15182_, _15181_, _15179_);
  not _65855_ (_15183_, _12898_);
  and _65856_ (_15184_, _15166_, _15183_);
  and _65857_ (_15185_, _15184_, _06264_);
  or _65858_ (_15186_, _15185_, _15182_);
  and _65859_ (_15187_, _15186_, _06007_);
  or _65860_ (_15188_, _12452_, _06007_);
  nand _65861_ (_15189_, _15188_, _06501_);
  or _65862_ (_15190_, _15189_, _15187_);
  nand _65863_ (_15191_, _08543_, _06502_);
  and _65864_ (_15192_, _15191_, _15190_);
  or _65865_ (_15193_, _15192_, _07197_);
  and _65866_ (_15194_, _09448_, _06286_);
  nand _65867_ (_15195_, _08488_, _07197_);
  or _65868_ (_15196_, _15195_, _15194_);
  and _65869_ (_15197_, _15196_, _15193_);
  or _65870_ (_15198_, _15197_, _07196_);
  and _65871_ (_15199_, _14411_, _06657_);
  or _65872_ (_15200_, _15199_, _15176_);
  or _65873_ (_15201_, _15200_, _08801_);
  and _65874_ (_15202_, _15201_, _05978_);
  and _65875_ (_15203_, _15202_, _15198_);
  or _65876_ (_15204_, _15203_, _15145_);
  and _65877_ (_15205_, _15204_, _08817_);
  nor _65878_ (_15206_, _08541_, _08817_);
  or _65879_ (_15207_, _15206_, _08816_);
  or _65880_ (_15208_, _15207_, _15205_);
  or _65881_ (_15209_, _09448_, _08821_);
  and _65882_ (_15210_, _15209_, _07471_);
  and _65883_ (_15211_, _15210_, _15208_);
  nor _65884_ (_15212_, _08825_, _08541_);
  and _65885_ (_15213_, _08962_, \oc8051_golden_model_1.P1 [4]);
  and _65886_ (_15214_, _08965_, \oc8051_golden_model_1.SCON [4]);
  or _65887_ (_15215_, _15214_, _15213_);
  and _65888_ (_15216_, _08944_, \oc8051_golden_model_1.P0 [4]);
  and _65889_ (_15217_, _08939_, \oc8051_golden_model_1.TL0 [4]);
  or _65890_ (_15218_, _15217_, _15216_);
  or _65891_ (_15219_, _15218_, _15215_);
  and _65892_ (_15220_, _08934_, \oc8051_golden_model_1.TCON [4]);
  and _65893_ (_15221_, _08957_, \oc8051_golden_model_1.TMOD [4]);
  or _65894_ (_15222_, _15221_, _15220_);
  and _65895_ (_15223_, _09005_, \oc8051_golden_model_1.SBUF [4]);
  and _65896_ (_15224_, _09007_, \oc8051_golden_model_1.PSW [4]);
  or _65897_ (_15225_, _15224_, _15223_);
  or _65898_ (_15226_, _15225_, _15222_);
  or _65899_ (_15227_, _15226_, _15219_);
  and _65900_ (_15228_, _08977_, \oc8051_golden_model_1.PCON [4]);
  and _65901_ (_15229_, _08979_, \oc8051_golden_model_1.DPH [4]);
  or _65902_ (_15230_, _15229_, _15228_);
  or _65903_ (_15231_, _15230_, _15227_);
  and _65904_ (_15232_, _09015_, \oc8051_golden_model_1.TH1 [4]);
  and _65905_ (_15233_, _08986_, \oc8051_golden_model_1.TL1 [4]);
  and _65906_ (_15234_, _08988_, \oc8051_golden_model_1.SP [4]);
  or _65907_ (_15235_, _15234_, _15233_);
  or _65908_ (_15236_, _15235_, _15232_);
  and _65909_ (_15237_, _08950_, \oc8051_golden_model_1.ACC [4]);
  and _65910_ (_15238_, _08968_, \oc8051_golden_model_1.B [4]);
  or _65911_ (_15239_, _15238_, _15237_);
  and _65912_ (_15240_, _08993_, \oc8051_golden_model_1.IE [4]);
  and _65913_ (_15241_, _08996_, \oc8051_golden_model_1.IP [4]);
  or _65914_ (_15242_, _15241_, _15240_);
  and _65915_ (_15243_, _08999_, \oc8051_golden_model_1.P2 [4]);
  and _65916_ (_15244_, _09001_, \oc8051_golden_model_1.P3 [4]);
  or _65917_ (_15245_, _15244_, _15243_);
  or _65918_ (_15246_, _15245_, _15242_);
  or _65919_ (_15247_, _15246_, _15239_);
  and _65920_ (_15248_, _08984_, \oc8051_golden_model_1.DPL [4]);
  and _65921_ (_15249_, _09013_, \oc8051_golden_model_1.TH0 [4]);
  or _65922_ (_15250_, _15249_, _15248_);
  or _65923_ (_15251_, _15250_, _15247_);
  or _65924_ (_15252_, _15251_, _15236_);
  or _65925_ (_15253_, _15252_, _15231_);
  or _65926_ (_15254_, _15253_, _15212_);
  and _65927_ (_15255_, _15254_, _07470_);
  or _65928_ (_15256_, _15255_, _09031_);
  or _65929_ (_15257_, _15256_, _15211_);
  and _65930_ (_15258_, _09031_, _06968_);
  nor _65931_ (_15259_, _15258_, _06220_);
  and _65932_ (_15260_, _15259_, _15257_);
  and _65933_ (_15261_, _08959_, _06220_);
  or _65934_ (_15262_, _15261_, _06217_);
  or _65935_ (_15263_, _15262_, _15260_);
  and _65936_ (_15264_, _15263_, _15144_);
  or _65937_ (_15265_, _15264_, _07238_);
  nand _65938_ (_15266_, _08892_, _08543_);
  nor _65939_ (_15267_, _08892_, _08543_);
  not _65940_ (_15268_, _15267_);
  and _65941_ (_15269_, _15268_, _15266_);
  or _65942_ (_15270_, _15269_, _07239_);
  and _65943_ (_15271_, _15270_, _08577_);
  and _65944_ (_15272_, _15271_, _15265_);
  and _65945_ (_15273_, _11254_, _07241_);
  or _65946_ (_15274_, _15273_, _07243_);
  or _65947_ (_15275_, _15274_, _15272_);
  or _65948_ (_15276_, _15267_, _08571_);
  and _65949_ (_15277_, _15276_, _07236_);
  and _65950_ (_15278_, _15277_, _15275_);
  and _65951_ (_15279_, _11251_, _07235_);
  or _65952_ (_15280_, _15279_, _07233_);
  or _65953_ (_15281_, _15280_, _15278_);
  nor _65954_ (_15282_, _12451_, _05961_);
  nor _65955_ (_15283_, _15282_, _09057_);
  and _65956_ (_15284_, _15283_, _15281_);
  and _65957_ (_15285_, _15266_, _09057_);
  or _65958_ (_15286_, _15285_, _09062_);
  or _65959_ (_15287_, _15286_, _15284_);
  nand _65960_ (_15288_, _11253_, _09062_);
  and _65961_ (_15289_, _15288_, _05959_);
  and _65962_ (_15290_, _15289_, _15287_);
  nor _65963_ (_15291_, _12452_, _05959_);
  nor _65964_ (_15292_, _15291_, _07292_);
  nand _65965_ (_15293_, _15292_, _08568_);
  or _65966_ (_15294_, _15293_, _15290_);
  or _65967_ (_15295_, _15152_, _08569_);
  and _65968_ (_15296_, _15295_, _14746_);
  and _65969_ (_15297_, _15296_, _15294_);
  or _65970_ (_15298_, _15297_, _15143_);
  and _65971_ (_15299_, _15298_, _14745_);
  and _65972_ (_15300_, _15142_, _07262_);
  or _65973_ (_15301_, _15300_, _15299_);
  and _65974_ (_15302_, _15301_, _09075_);
  and _65975_ (_15303_, _15162_, _07261_);
  or _65976_ (_15304_, _15303_, _06361_);
  or _65977_ (_15305_, _15304_, _15302_);
  nand _65978_ (_15306_, _12239_, _06361_);
  and _65979_ (_15307_, _15306_, _14710_);
  and _65980_ (_15308_, _15307_, _15305_);
  and _65981_ (_15309_, _12451_, _05940_);
  or _65982_ (_15310_, _15309_, _07270_);
  or _65983_ (_15311_, _15310_, _15308_);
  or _65984_ (_15312_, _15176_, _07539_);
  and _65985_ (_15313_, _15312_, _09427_);
  and _65986_ (_15314_, _15313_, _15311_);
  or _65987_ (_15315_, _09435_, _09430_);
  nor _65988_ (_15316_, _09436_, _09427_);
  and _65989_ (_15317_, _15316_, _15315_);
  or _65990_ (_15318_, _15317_, _07280_);
  or _65991_ (_15319_, _15318_, _15314_);
  nor _65992_ (_15320_, _09454_, _09448_);
  nor _65993_ (_15321_, _15320_, _09455_);
  or _65994_ (_15322_, _15321_, _14741_);
  and _65995_ (_15323_, _15322_, _14737_);
  and _65996_ (_15324_, _15323_, _15319_);
  and _65997_ (_15325_, _15321_, _07279_);
  or _65998_ (_15326_, _15325_, _07286_);
  or _65999_ (_15327_, _15326_, _15324_);
  nor _66000_ (_15328_, _08544_, _08442_);
  nor _66001_ (_15329_, _15328_, _08545_);
  or _66002_ (_15330_, _15329_, _09445_);
  and _66003_ (_15331_, _15330_, _07535_);
  and _66004_ (_15332_, _15331_, _15327_);
  or _66005_ (_15333_, _15332_, _14360_);
  or _66006_ (_15334_, _14359_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _66007_ (_15335_, _15334_, _14535_);
  and _66008_ (_15336_, _15335_, _15333_);
  nand _66009_ (_15337_, _12199_, _06361_);
  or _66010_ (_15338_, _12414_, _06361_);
  and _66011_ (_15339_, _15338_, _15337_);
  and _66012_ (_15340_, _15339_, _07872_);
  and _66013_ (_15341_, _15340_, _14539_);
  or _66014_ (_40616_, _15341_, _15336_);
  nor _66015_ (_15342_, _09397_, _09167_);
  or _66016_ (_15343_, _15342_, _09398_);
  and _66017_ (_15344_, _15343_, _07262_);
  not _66018_ (_15345_, _08563_);
  nor _66019_ (_15346_, _15150_, _08244_);
  or _66020_ (_15347_, _15346_, _08558_);
  and _66021_ (_15348_, _15347_, _15345_);
  or _66022_ (_15349_, _15348_, _08569_);
  nand _66023_ (_15350_, _08926_, _08246_);
  nor _66024_ (_15351_, _08926_, _08246_);
  not _66025_ (_15352_, _15351_);
  and _66026_ (_15353_, _15352_, _15350_);
  and _66027_ (_15354_, _15353_, _07238_);
  nor _66028_ (_15355_, _12999_, _12998_);
  or _66029_ (_15356_, _15355_, _08610_);
  nor _66030_ (_15357_, _15160_, _08246_);
  or _66031_ (_15358_, _15357_, _08764_);
  and _66032_ (_15359_, _15358_, _07152_);
  or _66033_ (_15360_, _09447_, _07155_);
  and _66034_ (_15361_, _15347_, _12387_);
  nand _66035_ (_15362_, _12447_, _06758_);
  or _66036_ (_15363_, _06758_, \oc8051_golden_model_1.ACC [5]);
  and _66037_ (_15364_, _15363_, _15362_);
  and _66038_ (_15365_, _15364_, _08654_);
  or _66039_ (_15366_, _15365_, _07154_);
  or _66040_ (_15367_, _15366_, _15361_);
  and _66041_ (_15368_, _15367_, _08652_);
  and _66042_ (_15369_, _15368_, _15360_);
  or _66043_ (_15370_, _15369_, _15359_);
  and _66044_ (_15371_, _15370_, _08651_);
  nand _66045_ (_15372_, _13000_, _12998_);
  and _66046_ (_15373_, _15372_, _06275_);
  or _66047_ (_15374_, _15373_, _07611_);
  or _66048_ (_15375_, _15374_, _15371_);
  nor _66049_ (_15376_, _12446_, _06010_);
  nor _66050_ (_15377_, _15376_, _07167_);
  and _66051_ (_15378_, _15377_, _15375_);
  and _66052_ (_15379_, _09429_, _07167_);
  or _66053_ (_15380_, _15379_, _07179_);
  or _66054_ (_15381_, _15380_, _15378_);
  and _66055_ (_15382_, _15381_, _15356_);
  or _66056_ (_15383_, _15382_, _06267_);
  nand _66057_ (_15384_, _08246_, _06267_);
  and _66058_ (_15385_, _15384_, _06265_);
  and _66059_ (_15386_, _15385_, _15383_);
  not _66060_ (_15387_, _13001_);
  and _66061_ (_15388_, _15372_, _06264_);
  and _66062_ (_15389_, _15388_, _15387_);
  or _66063_ (_15390_, _15389_, _15386_);
  and _66064_ (_15391_, _15390_, _06007_);
  or _66065_ (_15392_, _12447_, _06007_);
  nand _66066_ (_15393_, _15392_, _06501_);
  or _66067_ (_15394_, _15393_, _15391_);
  nand _66068_ (_15395_, _08246_, _06502_);
  and _66069_ (_15396_, _15395_, _15394_);
  or _66070_ (_15397_, _15396_, _07197_);
  and _66071_ (_15398_, _09447_, _06286_);
  nand _66072_ (_15399_, _08191_, _07197_);
  or _66073_ (_15400_, _15399_, _15398_);
  and _66074_ (_15401_, _15400_, _08801_);
  and _66075_ (_15402_, _15401_, _15397_);
  nand _66076_ (_15403_, _12999_, _10558_);
  and _66077_ (_15404_, _15403_, _07196_);
  and _66078_ (_15405_, _15404_, _15372_);
  or _66079_ (_15406_, _15405_, _06254_);
  or _66080_ (_15407_, _15406_, _15402_);
  nor _66081_ (_15408_, _12446_, _05978_);
  nor _66082_ (_15409_, _15408_, _08812_);
  and _66083_ (_15410_, _15409_, _15407_);
  nor _66084_ (_15411_, _08244_, _08817_);
  or _66085_ (_15412_, _15411_, _08816_);
  or _66086_ (_15413_, _15412_, _15410_);
  or _66087_ (_15414_, _09447_, _08821_);
  and _66088_ (_15415_, _15414_, _07471_);
  and _66089_ (_15416_, _15415_, _15413_);
  nor _66090_ (_15417_, _08825_, _08244_);
  and _66091_ (_15418_, _09005_, \oc8051_golden_model_1.SBUF [5]);
  and _66092_ (_15419_, _08968_, \oc8051_golden_model_1.B [5]);
  or _66093_ (_15420_, _15419_, _15418_);
  and _66094_ (_15421_, _08934_, \oc8051_golden_model_1.TCON [5]);
  and _66095_ (_15422_, _09007_, \oc8051_golden_model_1.PSW [5]);
  or _66096_ (_15423_, _15422_, _15421_);
  or _66097_ (_15424_, _15423_, _15420_);
  and _66098_ (_15425_, _08944_, \oc8051_golden_model_1.P0 [5]);
  and _66099_ (_15426_, _08965_, \oc8051_golden_model_1.SCON [5]);
  or _66100_ (_15427_, _15426_, _15425_);
  and _66101_ (_15428_, _08957_, \oc8051_golden_model_1.TMOD [5]);
  and _66102_ (_15429_, _08962_, \oc8051_golden_model_1.P1 [5]);
  or _66103_ (_15430_, _15429_, _15428_);
  or _66104_ (_15431_, _15430_, _15427_);
  or _66105_ (_15432_, _15431_, _15424_);
  and _66106_ (_15433_, _08977_, \oc8051_golden_model_1.PCON [5]);
  and _66107_ (_15434_, _08979_, \oc8051_golden_model_1.DPH [5]);
  or _66108_ (_15435_, _15434_, _15433_);
  or _66109_ (_15436_, _15435_, _15432_);
  and _66110_ (_15437_, _09013_, \oc8051_golden_model_1.TH0 [5]);
  and _66111_ (_15438_, _08986_, \oc8051_golden_model_1.TL1 [5]);
  and _66112_ (_15439_, _08988_, \oc8051_golden_model_1.SP [5]);
  or _66113_ (_15440_, _15439_, _15438_);
  or _66114_ (_15441_, _15440_, _15437_);
  and _66115_ (_15442_, _08999_, \oc8051_golden_model_1.P2 [5]);
  and _66116_ (_15443_, _09001_, \oc8051_golden_model_1.P3 [5]);
  or _66117_ (_15444_, _15443_, _15442_);
  and _66118_ (_15445_, _08993_, \oc8051_golden_model_1.IE [5]);
  and _66119_ (_15446_, _08996_, \oc8051_golden_model_1.IP [5]);
  or _66120_ (_15447_, _15446_, _15445_);
  or _66121_ (_15448_, _15447_, _15444_);
  and _66122_ (_15449_, _08939_, \oc8051_golden_model_1.TL0 [5]);
  and _66123_ (_15450_, _08950_, \oc8051_golden_model_1.ACC [5]);
  or _66124_ (_15451_, _15450_, _15449_);
  or _66125_ (_15452_, _15451_, _15448_);
  and _66126_ (_15453_, _08984_, \oc8051_golden_model_1.DPL [5]);
  and _66127_ (_15454_, _09015_, \oc8051_golden_model_1.TH1 [5]);
  or _66128_ (_15455_, _15454_, _15453_);
  or _66129_ (_15456_, _15455_, _15452_);
  or _66130_ (_15457_, _15456_, _15441_);
  or _66131_ (_15458_, _15457_, _15436_);
  or _66132_ (_15459_, _15458_, _15417_);
  and _66133_ (_15460_, _15459_, _07470_);
  or _66134_ (_15461_, _15460_, _09031_);
  or _66135_ (_15462_, _15461_, _15416_);
  and _66136_ (_15463_, _09031_, _06611_);
  nor _66137_ (_15464_, _15463_, _06220_);
  and _66138_ (_15465_, _15464_, _15462_);
  and _66139_ (_15466_, _08946_, _06220_);
  or _66140_ (_15467_, _15466_, _06217_);
  or _66141_ (_15468_, _15467_, _15465_);
  nor _66142_ (_15469_, _12446_, _05952_);
  nor _66143_ (_15470_, _15469_, _07238_);
  and _66144_ (_15471_, _15470_, _15468_);
  or _66145_ (_15472_, _15471_, _15354_);
  and _66146_ (_15473_, _15472_, _08577_);
  and _66147_ (_15474_, _11250_, _07241_);
  or _66148_ (_15475_, _15474_, _15473_);
  and _66149_ (_15476_, _15475_, _08571_);
  and _66150_ (_15477_, _15351_, _07243_);
  or _66151_ (_15478_, _15477_, _15476_);
  and _66152_ (_15479_, _15478_, _07236_);
  and _66153_ (_15480_, _11248_, _07235_);
  or _66154_ (_15481_, _15480_, _07233_);
  or _66155_ (_15482_, _15481_, _15479_);
  nor _66156_ (_15483_, _12446_, _05961_);
  nor _66157_ (_15484_, _15483_, _09057_);
  and _66158_ (_15485_, _15484_, _15482_);
  and _66159_ (_15486_, _15350_, _09057_);
  or _66160_ (_15487_, _15486_, _09062_);
  or _66161_ (_15488_, _15487_, _15485_);
  nand _66162_ (_15489_, _11249_, _09062_);
  and _66163_ (_15490_, _15489_, _05959_);
  and _66164_ (_15491_, _15490_, _15488_);
  or _66165_ (_15492_, _08567_, _08564_);
  nor _66166_ (_15493_, _12447_, _05959_);
  or _66167_ (_15494_, _15493_, _08566_);
  or _66168_ (_15495_, _15494_, _15492_);
  or _66169_ (_15496_, _15495_, _15491_);
  and _66170_ (_15497_, _15496_, _15349_);
  and _66171_ (_15498_, _15347_, _08563_);
  or _66172_ (_15499_, _15498_, _07263_);
  or _66173_ (_15500_, _15499_, _15497_);
  or _66174_ (_15501_, _15343_, _14746_);
  and _66175_ (_15502_, _15501_, _14745_);
  and _66176_ (_15503_, _15502_, _15500_);
  or _66177_ (_15504_, _15503_, _15344_);
  and _66178_ (_15505_, _15504_, _09075_);
  and _66179_ (_15506_, _15358_, _07261_);
  or _66180_ (_15507_, _15506_, _06361_);
  or _66181_ (_15508_, _15507_, _15505_);
  nand _66182_ (_15509_, _12234_, _06361_);
  and _66183_ (_15510_, _15509_, _14710_);
  and _66184_ (_15511_, _15510_, _15508_);
  and _66185_ (_15512_, _12446_, _05940_);
  or _66186_ (_15513_, _15512_, _07270_);
  or _66187_ (_15514_, _15513_, _15511_);
  or _66188_ (_15515_, _15355_, _07539_);
  and _66189_ (_15516_, _15515_, _15107_);
  and _66190_ (_15517_, _15516_, _15514_);
  nor _66191_ (_15518_, _09436_, _09429_);
  nor _66192_ (_15519_, _15518_, _09437_);
  and _66193_ (_15520_, _15519_, _15111_);
  or _66194_ (_15521_, _15520_, _15115_);
  or _66195_ (_15522_, _15521_, _15517_);
  or _66196_ (_15523_, _15519_, _15118_);
  and _66197_ (_15524_, _15523_, _07282_);
  and _66198_ (_15525_, _15524_, _15522_);
  or _66199_ (_15526_, _09455_, _09447_);
  nor _66200_ (_15527_, _09456_, _07282_);
  and _66201_ (_15528_, _15527_, _15526_);
  or _66202_ (_15529_, _15528_, _07286_);
  or _66203_ (_15530_, _15529_, _15525_);
  nor _66204_ (_15531_, _08545_, _08247_);
  nor _66205_ (_15532_, _15531_, _08546_);
  or _66206_ (_15533_, _15532_, _09445_);
  and _66207_ (_15534_, _15533_, _07535_);
  and _66208_ (_15535_, _15534_, _15530_);
  or _66209_ (_15536_, _15535_, _14360_);
  or _66210_ (_15537_, _14359_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _66211_ (_15538_, _15537_, _14535_);
  and _66212_ (_15539_, _15538_, _15536_);
  nand _66213_ (_15540_, _12194_, _06361_);
  or _66214_ (_15541_, _12409_, _06361_);
  and _66215_ (_15542_, _15541_, _15540_);
  and _66216_ (_15543_, _15542_, _07872_);
  and _66217_ (_15544_, _15543_, _14539_);
  or _66218_ (_40618_, _15544_, _15539_);
  nor _66219_ (_15545_, _12440_, _05959_);
  nand _66220_ (_15546_, _08857_, _08144_);
  nor _66221_ (_15547_, _08857_, _08144_);
  not _66222_ (_15548_, _15547_);
  and _66223_ (_15549_, _15548_, _15546_);
  and _66224_ (_15550_, _15549_, _07238_);
  nor _66225_ (_15551_, _12949_, _12948_);
  or _66226_ (_15552_, _15551_, _08610_);
  nor _66227_ (_15553_, _08764_, _08144_);
  or _66228_ (_15554_, _15553_, _08765_);
  and _66229_ (_15555_, _15554_, _07152_);
  or _66230_ (_15556_, _09446_, _07155_);
  nor _66231_ (_15557_, _08558_, _08142_);
  or _66232_ (_15558_, _15557_, _08559_);
  and _66233_ (_15559_, _15558_, _12387_);
  nand _66234_ (_15560_, _12440_, _06758_);
  or _66235_ (_15561_, _06758_, \oc8051_golden_model_1.ACC [6]);
  and _66236_ (_15562_, _15561_, _15560_);
  and _66237_ (_15563_, _15562_, _08654_);
  or _66238_ (_15564_, _15563_, _07154_);
  or _66239_ (_15565_, _15564_, _15559_);
  and _66240_ (_15566_, _15565_, _08652_);
  and _66241_ (_15567_, _15566_, _15556_);
  or _66242_ (_15568_, _15567_, _15555_);
  and _66243_ (_15569_, _15568_, _08651_);
  nand _66244_ (_15570_, _12950_, _12948_);
  and _66245_ (_15571_, _15570_, _06275_);
  or _66246_ (_15572_, _15571_, _07611_);
  or _66247_ (_15573_, _15572_, _15569_);
  nor _66248_ (_15574_, _12439_, _06010_);
  nor _66249_ (_15575_, _15574_, _07167_);
  and _66250_ (_15576_, _15575_, _15573_);
  and _66251_ (_15577_, _09428_, _07167_);
  or _66252_ (_15578_, _15577_, _07179_);
  or _66253_ (_15579_, _15578_, _15576_);
  and _66254_ (_15580_, _15579_, _15552_);
  or _66255_ (_15581_, _15580_, _06267_);
  nand _66256_ (_15582_, _08144_, _06267_);
  and _66257_ (_15583_, _15582_, _06265_);
  and _66258_ (_15584_, _15583_, _15581_);
  not _66259_ (_15585_, _12951_);
  and _66260_ (_15586_, _15570_, _15585_);
  and _66261_ (_15587_, _15586_, _06264_);
  or _66262_ (_15588_, _15587_, _15584_);
  and _66263_ (_15589_, _15588_, _06007_);
  or _66264_ (_15590_, _12440_, _06007_);
  nand _66265_ (_15591_, _15590_, _06501_);
  or _66266_ (_15592_, _15591_, _15589_);
  nand _66267_ (_15593_, _08144_, _06502_);
  and _66268_ (_15594_, _15593_, _15592_);
  or _66269_ (_15595_, _15594_, _07197_);
  and _66270_ (_15596_, _09446_, _06286_);
  nand _66271_ (_15597_, _08089_, _07197_);
  or _66272_ (_15598_, _15597_, _15596_);
  and _66273_ (_15599_, _15598_, _08801_);
  and _66274_ (_15600_, _15599_, _15595_);
  and _66275_ (_15601_, _14802_, _06657_);
  or _66276_ (_15602_, _15601_, _15551_);
  and _66277_ (_15603_, _15602_, _07196_);
  or _66278_ (_15604_, _15603_, _06254_);
  or _66279_ (_15605_, _15604_, _15600_);
  nor _66280_ (_15606_, _12439_, _05978_);
  nor _66281_ (_15607_, _15606_, _08812_);
  and _66282_ (_15608_, _15607_, _15605_);
  nor _66283_ (_15609_, _08142_, _08817_);
  or _66284_ (_15610_, _15609_, _08816_);
  or _66285_ (_15611_, _15610_, _15608_);
  or _66286_ (_15612_, _09446_, _08821_);
  and _66287_ (_15613_, _15612_, _07471_);
  and _66288_ (_15614_, _15613_, _15611_);
  nor _66289_ (_15615_, _08825_, _08142_);
  and _66290_ (_15616_, _08962_, \oc8051_golden_model_1.P1 [6]);
  and _66291_ (_15617_, _08965_, \oc8051_golden_model_1.SCON [6]);
  or _66292_ (_15618_, _15617_, _15616_);
  and _66293_ (_15619_, _08944_, \oc8051_golden_model_1.P0 [6]);
  and _66294_ (_15620_, _09005_, \oc8051_golden_model_1.SBUF [6]);
  or _66295_ (_15621_, _15620_, _15619_);
  or _66296_ (_15622_, _15621_, _15618_);
  and _66297_ (_15623_, _08957_, \oc8051_golden_model_1.TMOD [6]);
  and _66298_ (_15624_, _09007_, \oc8051_golden_model_1.PSW [6]);
  or _66299_ (_15625_, _15624_, _15623_);
  and _66300_ (_15626_, _08934_, \oc8051_golden_model_1.TCON [6]);
  and _66301_ (_15627_, _08950_, \oc8051_golden_model_1.ACC [6]);
  or _66302_ (_15628_, _15627_, _15626_);
  or _66303_ (_15629_, _15628_, _15625_);
  or _66304_ (_15630_, _15629_, _15622_);
  and _66305_ (_15631_, _08977_, \oc8051_golden_model_1.PCON [6]);
  and _66306_ (_15632_, _08979_, \oc8051_golden_model_1.DPH [6]);
  or _66307_ (_15633_, _15632_, _15631_);
  or _66308_ (_15634_, _15633_, _15630_);
  and _66309_ (_15635_, _08986_, \oc8051_golden_model_1.TL1 [6]);
  and _66310_ (_15636_, _08984_, \oc8051_golden_model_1.DPL [6]);
  and _66311_ (_15637_, _09015_, \oc8051_golden_model_1.TH1 [6]);
  or _66312_ (_15638_, _15637_, _15636_);
  or _66313_ (_15639_, _15638_, _15635_);
  and _66314_ (_15640_, _08999_, \oc8051_golden_model_1.P2 [6]);
  and _66315_ (_15641_, _09001_, \oc8051_golden_model_1.P3 [6]);
  or _66316_ (_15642_, _15641_, _15640_);
  and _66317_ (_15643_, _08993_, \oc8051_golden_model_1.IE [6]);
  and _66318_ (_15644_, _08996_, \oc8051_golden_model_1.IP [6]);
  or _66319_ (_15645_, _15644_, _15643_);
  or _66320_ (_15646_, _15645_, _15642_);
  and _66321_ (_15647_, _08939_, \oc8051_golden_model_1.TL0 [6]);
  and _66322_ (_15648_, _08968_, \oc8051_golden_model_1.B [6]);
  or _66323_ (_15649_, _15648_, _15647_);
  or _66324_ (_15650_, _15649_, _15646_);
  and _66325_ (_15651_, _09013_, \oc8051_golden_model_1.TH0 [6]);
  and _66326_ (_15652_, _08988_, \oc8051_golden_model_1.SP [6]);
  or _66327_ (_15653_, _15652_, _15651_);
  or _66328_ (_15654_, _15653_, _15650_);
  or _66329_ (_15655_, _15654_, _15639_);
  or _66330_ (_15656_, _15655_, _15634_);
  or _66331_ (_15657_, _15656_, _15615_);
  and _66332_ (_15658_, _15657_, _07470_);
  or _66333_ (_15659_, _15658_, _09031_);
  or _66334_ (_15660_, _15659_, _15614_);
  and _66335_ (_15661_, _09031_, _06317_);
  nor _66336_ (_15662_, _15661_, _06220_);
  and _66337_ (_15663_, _15662_, _15660_);
  not _66338_ (_15664_, _08857_);
  and _66339_ (_15665_, _15664_, _06220_);
  or _66340_ (_15666_, _15665_, _06217_);
  or _66341_ (_15667_, _15666_, _15663_);
  nor _66342_ (_15668_, _12439_, _05952_);
  nor _66343_ (_15669_, _15668_, _07238_);
  and _66344_ (_15670_, _15669_, _15667_);
  or _66345_ (_15671_, _15670_, _15550_);
  and _66346_ (_15672_, _15671_, _08577_);
  and _66347_ (_15673_, _11247_, _07241_);
  or _66348_ (_15674_, _15673_, _15672_);
  and _66349_ (_15675_, _15674_, _08571_);
  and _66350_ (_15676_, _15547_, _07243_);
  or _66351_ (_15677_, _15676_, _15675_);
  and _66352_ (_15678_, _15677_, _07236_);
  and _66353_ (_15679_, _11244_, _07235_);
  or _66354_ (_15680_, _15679_, _07233_);
  or _66355_ (_15681_, _15680_, _15678_);
  nor _66356_ (_15682_, _12439_, _05961_);
  nor _66357_ (_15683_, _15682_, _09057_);
  and _66358_ (_15684_, _15683_, _15681_);
  and _66359_ (_15685_, _15546_, _09057_);
  or _66360_ (_15686_, _15685_, _09062_);
  or _66361_ (_15687_, _15686_, _15684_);
  nand _66362_ (_15688_, _11246_, _09062_);
  and _66363_ (_15689_, _15688_, _05959_);
  and _66364_ (_15690_, _15689_, _15687_);
  or _66365_ (_15691_, _15690_, _15545_);
  and _66366_ (_15692_, _15691_, _08568_);
  not _66367_ (_15693_, _08568_);
  and _66368_ (_15694_, _15558_, _15693_);
  or _66369_ (_15695_, _15694_, _07292_);
  or _66370_ (_15696_, _15695_, _15692_);
  or _66371_ (_15697_, _15558_, _08565_);
  and _66372_ (_15698_, _15697_, _14746_);
  and _66373_ (_15699_, _15698_, _15696_);
  nor _66374_ (_15700_, _09398_, _09122_);
  or _66375_ (_15701_, _15700_, _09399_);
  or _66376_ (_15702_, _15701_, _07262_);
  and _66377_ (_15703_, _15702_, _07435_);
  or _66378_ (_15704_, _15703_, _15699_);
  or _66379_ (_15705_, _15701_, _14745_);
  and _66380_ (_15706_, _15705_, _09075_);
  and _66381_ (_15707_, _15706_, _15704_);
  and _66382_ (_15708_, _15554_, _07261_);
  or _66383_ (_15709_, _15708_, _06361_);
  or _66384_ (_15710_, _15709_, _15707_);
  nand _66385_ (_15711_, _12226_, _06361_);
  and _66386_ (_15712_, _15711_, _14710_);
  and _66387_ (_15713_, _15712_, _15710_);
  and _66388_ (_15714_, _12439_, _05940_);
  or _66389_ (_15715_, _15714_, _07270_);
  or _66390_ (_15716_, _15715_, _15713_);
  or _66391_ (_15717_, _15551_, _07539_);
  and _66392_ (_15718_, _15717_, _09427_);
  and _66393_ (_15719_, _15718_, _15716_);
  nor _66394_ (_15720_, _09437_, _09428_);
  nor _66395_ (_15721_, _15720_, _09438_);
  and _66396_ (_15722_, _15721_, _09424_);
  or _66397_ (_15723_, _15722_, _07280_);
  or _66398_ (_15724_, _15723_, _15719_);
  nor _66399_ (_15725_, _09456_, _09446_);
  nor _66400_ (_15726_, _15725_, _09457_);
  or _66401_ (_15727_, _15726_, _14741_);
  and _66402_ (_15728_, _15727_, _14737_);
  and _66403_ (_15729_, _15728_, _15724_);
  and _66404_ (_15730_, _15726_, _07279_);
  or _66405_ (_15731_, _15730_, _07286_);
  or _66406_ (_15732_, _15731_, _15729_);
  nor _66407_ (_15733_, _08546_, _08145_);
  nor _66408_ (_15734_, _15733_, _08547_);
  or _66409_ (_15735_, _15734_, _09445_);
  and _66410_ (_15736_, _15735_, _07535_);
  and _66411_ (_15737_, _15736_, _15732_);
  or _66412_ (_15738_, _15737_, _14360_);
  or _66413_ (_15739_, _14359_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _66414_ (_15740_, _15739_, _14535_);
  and _66415_ (_15741_, _15740_, _15738_);
  or _66416_ (_15742_, _12186_, _14508_);
  or _66417_ (_15743_, _12403_, _06361_);
  and _66418_ (_15744_, _15743_, _15742_);
  and _66419_ (_15745_, _15744_, _07872_);
  and _66420_ (_15746_, _15745_, _14539_);
  or _66421_ (_40619_, _15746_, _15741_);
  nand _66422_ (_15747_, _14359_, _09464_);
  or _66423_ (_15748_, _14359_, _07980_);
  and _66424_ (_15749_, _15748_, _14535_);
  nand _66425_ (_15750_, _15749_, _15747_);
  or _66426_ (_15751_, _14535_, _09489_);
  and _66427_ (_40620_, _15751_, _15750_);
  and _66428_ (_15752_, _14354_, _07453_);
  and _66429_ (_15753_, _15752_, _14357_);
  not _66430_ (_15754_, _15753_);
  or _66431_ (_15755_, _15754_, _14528_);
  or _66432_ (_15756_, _15753_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand _66433_ (_15757_, _14533_, _07598_);
  or _66434_ (_15758_, _15757_, _14531_);
  and _66435_ (_15759_, _15758_, _15756_);
  and _66436_ (_15760_, _15759_, _15755_);
  and _66437_ (_15761_, _07872_, _07598_);
  and _66438_ (_15762_, _15761_, _14533_);
  and _66439_ (_15763_, _15762_, _14543_);
  or _66440_ (_40623_, _15763_, _15760_);
  or _66441_ (_15764_, _15754_, _14727_);
  or _66442_ (_15765_, _15753_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _66443_ (_15766_, _15765_, _15758_);
  and _66444_ (_15767_, _15766_, _15764_);
  and _66445_ (_15768_, _15762_, _14735_);
  or _66446_ (_40626_, _15768_, _15767_);
  or _66447_ (_15769_, _15754_, _14929_);
  or _66448_ (_15770_, _15753_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _66449_ (_15771_, _15770_, _15758_);
  and _66450_ (_15772_, _15771_, _15769_);
  and _66451_ (_15773_, _15762_, _14937_);
  or _66452_ (_40627_, _15773_, _15772_);
  or _66453_ (_15774_, _15754_, _15131_);
  or _66454_ (_15775_, _15753_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _66455_ (_15776_, _15775_, _15758_);
  and _66456_ (_15777_, _15776_, _15774_);
  and _66457_ (_15778_, _15762_, _15139_);
  or _66458_ (_40628_, _15778_, _15777_);
  or _66459_ (_15779_, _15754_, _15332_);
  or _66460_ (_15780_, _15753_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _66461_ (_15781_, _15780_, _15758_);
  and _66462_ (_15782_, _15781_, _15779_);
  and _66463_ (_15783_, _15762_, _15340_);
  or _66464_ (_40629_, _15783_, _15782_);
  or _66465_ (_15784_, _15754_, _15535_);
  or _66466_ (_15785_, _15753_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _66467_ (_15786_, _15785_, _15758_);
  and _66468_ (_15787_, _15786_, _15784_);
  and _66469_ (_15788_, _15762_, _15543_);
  or _66470_ (_40630_, _15788_, _15787_);
  or _66471_ (_15789_, _15754_, _15737_);
  or _66472_ (_15790_, _15753_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _66473_ (_15791_, _15790_, _15758_);
  and _66474_ (_15792_, _15791_, _15789_);
  and _66475_ (_15793_, _15762_, _15745_);
  or _66476_ (_40632_, _15793_, _15792_);
  or _66477_ (_15794_, _15754_, _09465_);
  or _66478_ (_15795_, _15753_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _66479_ (_15796_, _15795_, _15758_);
  and _66480_ (_15797_, _15796_, _15794_);
  and _66481_ (_15798_, _15762_, _09490_);
  or _66482_ (_40633_, _15798_, _15797_);
  not _66483_ (_15799_, _07537_);
  nor _66484_ (_15800_, _15799_, _07289_);
  and _66485_ (_15801_, _15800_, _14357_);
  not _66486_ (_15802_, _15801_);
  or _66487_ (_15803_, _15802_, _14528_);
  or _66488_ (_15804_, _15801_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand _66489_ (_15805_, _14533_, _08668_);
  or _66490_ (_15806_, _15805_, _14531_);
  and _66491_ (_15807_, _15806_, _15804_);
  and _66492_ (_15808_, _15807_, _15803_);
  and _66493_ (_15809_, _08668_, _07872_);
  and _66494_ (_15810_, _15809_, _14533_);
  and _66495_ (_15811_, _15810_, _14543_);
  or _66496_ (_40637_, _15811_, _15808_);
  or _66497_ (_15812_, _15802_, _14727_);
  or _66498_ (_15813_, _15801_, \oc8051_golden_model_1.IRAM[2] [1]);
  and _66499_ (_15814_, _15813_, _15806_);
  and _66500_ (_15815_, _15814_, _15812_);
  and _66501_ (_15816_, _15810_, _14735_);
  or _66502_ (_40638_, _15816_, _15815_);
  or _66503_ (_15817_, _15802_, _14929_);
  or _66504_ (_15818_, _15801_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _66505_ (_15819_, _15818_, _15806_);
  and _66506_ (_15820_, _15819_, _15817_);
  and _66507_ (_15821_, _15810_, _14937_);
  or _66508_ (_40640_, _15821_, _15820_);
  or _66509_ (_15822_, _15802_, _15131_);
  or _66510_ (_15823_, _15801_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _66511_ (_15824_, _15823_, _15806_);
  and _66512_ (_15825_, _15824_, _15822_);
  and _66513_ (_15826_, _15810_, _15139_);
  or _66514_ (_40641_, _15826_, _15825_);
  or _66515_ (_15827_, _15802_, _15332_);
  or _66516_ (_15828_, _15801_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _66517_ (_15829_, _15828_, _15806_);
  and _66518_ (_15830_, _15829_, _15827_);
  and _66519_ (_15831_, _15810_, _15340_);
  or _66520_ (_40642_, _15831_, _15830_);
  or _66521_ (_15832_, _15802_, _15535_);
  or _66522_ (_15833_, _15801_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _66523_ (_15834_, _15833_, _15806_);
  and _66524_ (_15835_, _15834_, _15832_);
  and _66525_ (_15836_, _15810_, _15543_);
  or _66526_ (_40643_, _15836_, _15835_);
  or _66527_ (_15837_, _15802_, _15737_);
  or _66528_ (_15838_, _15801_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _66529_ (_15839_, _15838_, _15806_);
  and _66530_ (_15840_, _15839_, _15837_);
  and _66531_ (_15841_, _15810_, _15745_);
  or _66532_ (_40644_, _15841_, _15840_);
  or _66533_ (_15842_, _15802_, _09465_);
  or _66534_ (_15843_, _15801_, \oc8051_golden_model_1.IRAM[2] [7]);
  and _66535_ (_15844_, _15843_, _15806_);
  and _66536_ (_15845_, _15844_, _15842_);
  and _66537_ (_15846_, _15810_, _09490_);
  or _66538_ (_40646_, _15846_, _15845_);
  and _66539_ (_15847_, _14357_, _07538_);
  or _66540_ (_15848_, _15847_, \oc8051_golden_model_1.IRAM[3] [0]);
  nand _66541_ (_15849_, _14533_, _07295_);
  or _66542_ (_15850_, _15849_, _14531_);
  and _66543_ (_15851_, _15850_, _15848_);
  not _66544_ (_15852_, _15847_);
  or _66545_ (_15853_, _15852_, _14528_);
  and _66546_ (_15854_, _15853_, _15851_);
  and _66547_ (_15855_, _07872_, _07295_);
  and _66548_ (_15856_, _15855_, _14533_);
  and _66549_ (_15857_, _15856_, _14543_);
  or _66550_ (_40649_, _15857_, _15854_);
  or _66551_ (_15858_, _15847_, \oc8051_golden_model_1.IRAM[3] [1]);
  and _66552_ (_15859_, _15858_, _15850_);
  or _66553_ (_15860_, _15852_, _14727_);
  and _66554_ (_15861_, _15860_, _15859_);
  and _66555_ (_15862_, _15856_, _14735_);
  or _66556_ (_40651_, _15862_, _15861_);
  nor _66557_ (_15863_, _15847_, _07728_);
  and _66558_ (_15864_, _15847_, _14929_);
  or _66559_ (_15865_, _15864_, _15863_);
  and _66560_ (_15866_, _15865_, _15850_);
  and _66561_ (_15867_, _15856_, _14937_);
  or _66562_ (_40652_, _15867_, _15866_);
  or _66563_ (_15868_, _15847_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _66564_ (_15869_, _15868_, _15850_);
  or _66565_ (_15870_, _15852_, _15131_);
  and _66566_ (_15871_, _15870_, _15869_);
  and _66567_ (_15872_, _15856_, _15139_);
  or _66568_ (_40653_, _15872_, _15871_);
  or _66569_ (_15873_, _15847_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _66570_ (_15874_, _15873_, _15850_);
  or _66571_ (_15875_, _15852_, _15332_);
  and _66572_ (_15876_, _15875_, _15874_);
  and _66573_ (_15877_, _15856_, _15340_);
  or _66574_ (_40654_, _15877_, _15876_);
  or _66575_ (_15878_, _15847_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _66576_ (_15879_, _15878_, _15850_);
  or _66577_ (_15880_, _15852_, _15535_);
  and _66578_ (_15881_, _15880_, _15879_);
  and _66579_ (_15882_, _15856_, _15543_);
  or _66580_ (_40655_, _15882_, _15881_);
  or _66581_ (_15883_, _15847_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _66582_ (_15884_, _15883_, _15850_);
  or _66583_ (_15885_, _15852_, _15737_);
  and _66584_ (_15886_, _15885_, _15884_);
  and _66585_ (_15887_, _15856_, _15745_);
  or _66586_ (_40657_, _15887_, _15886_);
  or _66587_ (_15888_, _15847_, \oc8051_golden_model_1.IRAM[3] [7]);
  and _66588_ (_15889_, _15888_, _15850_);
  or _66589_ (_15890_, _15852_, _09465_);
  and _66590_ (_15891_, _15890_, _15889_);
  and _66591_ (_15892_, _15856_, _09490_);
  or _66592_ (_40658_, _15892_, _15891_);
  and _66593_ (_15893_, _07859_, _07711_);
  and _66594_ (_15894_, _15893_, _14355_);
  not _66595_ (_15895_, _15894_);
  or _66596_ (_15896_, _15895_, _14528_);
  not _66597_ (_15897_, _07869_);
  and _66598_ (_15898_, _14532_, _15897_);
  and _66599_ (_15899_, _15898_, _07296_);
  not _66600_ (_15900_, _15899_);
  or _66601_ (_15901_, _15894_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _66602_ (_15902_, _15901_, _15900_);
  and _66603_ (_15903_, _15902_, _15896_);
  and _66604_ (_15904_, _15899_, _14543_);
  or _66605_ (_40662_, _15904_, _15903_);
  or _66606_ (_15905_, _15895_, _14727_);
  or _66607_ (_15906_, _15894_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _66608_ (_15907_, _15906_, _15900_);
  and _66609_ (_15908_, _15907_, _15905_);
  and _66610_ (_15909_, _15899_, _14735_);
  or _66611_ (_40663_, _15909_, _15908_);
  or _66612_ (_15910_, _15895_, _14929_);
  or _66613_ (_15911_, _15894_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _66614_ (_15912_, _15911_, _15900_);
  and _66615_ (_15913_, _15912_, _15910_);
  and _66616_ (_15914_, _15899_, _14937_);
  or _66617_ (_40665_, _15914_, _15913_);
  or _66618_ (_15915_, _15895_, _15131_);
  or _66619_ (_15916_, _15894_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _66620_ (_15917_, _15916_, _15900_);
  and _66621_ (_15918_, _15917_, _15915_);
  and _66622_ (_15919_, _15899_, _15139_);
  or _66623_ (_40666_, _15919_, _15918_);
  or _66624_ (_15920_, _15895_, _15332_);
  or _66625_ (_15921_, _15894_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _66626_ (_15922_, _15921_, _15900_);
  and _66627_ (_15923_, _15922_, _15920_);
  and _66628_ (_15924_, _15899_, _15340_);
  or _66629_ (_40667_, _15924_, _15923_);
  or _66630_ (_15925_, _15895_, _15535_);
  or _66631_ (_15926_, _15894_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _66632_ (_15927_, _15926_, _15900_);
  and _66633_ (_15928_, _15927_, _15925_);
  and _66634_ (_15929_, _15899_, _15543_);
  or _66635_ (_40668_, _15929_, _15928_);
  or _66636_ (_15930_, _15895_, _15737_);
  or _66637_ (_15931_, _15894_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _66638_ (_15932_, _15931_, _15900_);
  and _66639_ (_15933_, _15932_, _15930_);
  and _66640_ (_15934_, _15899_, _15745_);
  or _66641_ (_40669_, _15934_, _15933_);
  or _66642_ (_15935_, _15895_, _09465_);
  or _66643_ (_15936_, _15894_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _66644_ (_15937_, _15936_, _15900_);
  and _66645_ (_15938_, _15937_, _15935_);
  and _66646_ (_15939_, _15899_, _09490_);
  or _66647_ (_40671_, _15939_, _15938_);
  and _66648_ (_15940_, _15893_, _15752_);
  not _66649_ (_15941_, _15940_);
  or _66650_ (_15942_, _15941_, _14528_);
  and _66651_ (_15943_, _15898_, _07598_);
  not _66652_ (_15944_, _15943_);
  or _66653_ (_15945_, _15940_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _66654_ (_15946_, _15945_, _15944_);
  and _66655_ (_15947_, _15946_, _15942_);
  and _66656_ (_15948_, _15943_, _14543_);
  or _66657_ (_40673_, _15948_, _15947_);
  or _66658_ (_15949_, _15941_, _14727_);
  or _66659_ (_15950_, _15940_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _66660_ (_15951_, _15950_, _15944_);
  and _66661_ (_15952_, _15951_, _15949_);
  and _66662_ (_15953_, _15943_, _14735_);
  or _66663_ (_40674_, _15953_, _15952_);
  or _66664_ (_15954_, _15941_, _14929_);
  or _66665_ (_15955_, _15940_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _66666_ (_15956_, _15955_, _15944_);
  and _66667_ (_15957_, _15956_, _15954_);
  and _66668_ (_15958_, _15943_, _14937_);
  or _66669_ (_40677_, _15958_, _15957_);
  or _66670_ (_15959_, _15941_, _15131_);
  or _66671_ (_15960_, _15940_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _66672_ (_15961_, _15960_, _15944_);
  and _66673_ (_15962_, _15961_, _15959_);
  and _66674_ (_15963_, _15943_, _15139_);
  or _66675_ (_40678_, _15963_, _15962_);
  or _66676_ (_15964_, _15941_, _15332_);
  or _66677_ (_15965_, _15940_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _66678_ (_15966_, _15965_, _15944_);
  and _66679_ (_15967_, _15966_, _15964_);
  and _66680_ (_15968_, _15943_, _15340_);
  or _66681_ (_40679_, _15968_, _15967_);
  or _66682_ (_15969_, _15941_, _15535_);
  or _66683_ (_15970_, _15940_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _66684_ (_15971_, _15970_, _15944_);
  and _66685_ (_15972_, _15971_, _15969_);
  and _66686_ (_15973_, _15943_, _15543_);
  or _66687_ (_40680_, _15973_, _15972_);
  or _66688_ (_15974_, _15941_, _15737_);
  or _66689_ (_15975_, _15940_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _66690_ (_15976_, _15975_, _15944_);
  and _66691_ (_15977_, _15976_, _15974_);
  and _66692_ (_15978_, _15943_, _15745_);
  or _66693_ (_40681_, _15978_, _15977_);
  or _66694_ (_15979_, _15941_, _09465_);
  or _66695_ (_15980_, _15940_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _66696_ (_15981_, _15980_, _15944_);
  and _66697_ (_15982_, _15981_, _15979_);
  and _66698_ (_15983_, _15943_, _09490_);
  or _66699_ (_40683_, _15983_, _15982_);
  and _66700_ (_15984_, _15893_, _15800_);
  not _66701_ (_15985_, _15984_);
  or _66702_ (_15986_, _15985_, _14528_);
  and _66703_ (_15987_, _15898_, _08668_);
  not _66704_ (_15988_, _15987_);
  or _66705_ (_15989_, _15984_, \oc8051_golden_model_1.IRAM[6] [0]);
  and _66706_ (_15990_, _15989_, _15988_);
  and _66707_ (_15991_, _15990_, _15986_);
  and _66708_ (_15992_, _15987_, _14543_);
  or _66709_ (_40685_, _15992_, _15991_);
  or _66710_ (_15993_, _15985_, _14727_);
  or _66711_ (_15994_, _15984_, \oc8051_golden_model_1.IRAM[6] [1]);
  and _66712_ (_15995_, _15994_, _15988_);
  and _66713_ (_15996_, _15995_, _15993_);
  and _66714_ (_15997_, _15987_, _14735_);
  or _66715_ (_40688_, _15997_, _15996_);
  or _66716_ (_15998_, _15985_, _14929_);
  or _66717_ (_15999_, _15984_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _66718_ (_16000_, _15999_, _15988_);
  and _66719_ (_16001_, _16000_, _15998_);
  and _66720_ (_16002_, _15987_, _14937_);
  or _66721_ (_40689_, _16002_, _16001_);
  or _66722_ (_16003_, _15985_, _15131_);
  or _66723_ (_16004_, _15984_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _66724_ (_16005_, _16004_, _15988_);
  and _66725_ (_16006_, _16005_, _16003_);
  and _66726_ (_16007_, _15987_, _15139_);
  or _66727_ (_40690_, _16007_, _16006_);
  or _66728_ (_16008_, _15985_, _15332_);
  or _66729_ (_16009_, _15984_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _66730_ (_16010_, _16009_, _15988_);
  and _66731_ (_16011_, _16010_, _16008_);
  and _66732_ (_16012_, _15987_, _15340_);
  or _66733_ (_40691_, _16012_, _16011_);
  or _66734_ (_16013_, _15985_, _15535_);
  or _66735_ (_16014_, _15984_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _66736_ (_16015_, _16014_, _15988_);
  and _66737_ (_16016_, _16015_, _16013_);
  and _66738_ (_16017_, _15987_, _15543_);
  or _66739_ (_40692_, _16017_, _16016_);
  or _66740_ (_16018_, _15985_, _15737_);
  or _66741_ (_16019_, _15984_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _66742_ (_16020_, _16019_, _15988_);
  and _66743_ (_16021_, _16020_, _16018_);
  and _66744_ (_16022_, _15987_, _15745_);
  or _66745_ (_40694_, _16022_, _16021_);
  or _66746_ (_16023_, _15985_, _09465_);
  or _66747_ (_16024_, _15984_, \oc8051_golden_model_1.IRAM[6] [7]);
  and _66748_ (_16025_, _16024_, _15988_);
  and _66749_ (_16026_, _16025_, _16023_);
  and _66750_ (_16027_, _15987_, _09490_);
  or _66751_ (_40695_, _16027_, _16026_);
  and _66752_ (_16028_, _15898_, _07295_);
  not _66753_ (_16029_, _16028_);
  or _66754_ (_16030_, _16029_, _14543_);
  and _66755_ (_16031_, _15893_, _07538_);
  and _66756_ (_16032_, _16031_, _14528_);
  nor _66757_ (_16033_, _16031_, _07092_);
  or _66758_ (_16034_, _16033_, _16028_);
  or _66759_ (_16035_, _16034_, _16032_);
  and _66760_ (_40698_, _16035_, _16030_);
  or _66761_ (_16036_, _16031_, \oc8051_golden_model_1.IRAM[7] [1]);
  and _66762_ (_16037_, _16036_, _16029_);
  not _66763_ (_16038_, _16031_);
  or _66764_ (_16039_, _16038_, _14727_);
  and _66765_ (_16040_, _16039_, _16037_);
  and _66766_ (_16041_, _16028_, _14735_);
  or _66767_ (_40700_, _16041_, _16040_);
  nor _66768_ (_16042_, _16031_, _07736_);
  and _66769_ (_16043_, _16031_, _14929_);
  or _66770_ (_16044_, _16043_, _16042_);
  and _66771_ (_16045_, _16044_, _16029_);
  and _66772_ (_16046_, _16028_, _14937_);
  or _66773_ (_40701_, _16046_, _16045_);
  or _66774_ (_16047_, _16038_, _15131_);
  or _66775_ (_16048_, _16031_, \oc8051_golden_model_1.IRAM[7] [3]);
  and _66776_ (_16049_, _16048_, _16029_);
  and _66777_ (_16050_, _16049_, _16047_);
  and _66778_ (_16051_, _16028_, _15139_);
  or _66779_ (_40702_, _16051_, _16050_);
  or _66780_ (_16052_, _16031_, \oc8051_golden_model_1.IRAM[7] [4]);
  and _66781_ (_16053_, _16052_, _16029_);
  or _66782_ (_16054_, _16038_, _15332_);
  and _66783_ (_16055_, _16054_, _16053_);
  and _66784_ (_16056_, _16028_, _15340_);
  or _66785_ (_40703_, _16056_, _16055_);
  or _66786_ (_16057_, _16038_, _15535_);
  or _66787_ (_16058_, _16031_, \oc8051_golden_model_1.IRAM[7] [5]);
  and _66788_ (_16059_, _16058_, _16029_);
  and _66789_ (_16060_, _16059_, _16057_);
  and _66790_ (_16061_, _16028_, _15543_);
  or _66791_ (_40704_, _16061_, _16060_);
  or _66792_ (_16062_, _16031_, \oc8051_golden_model_1.IRAM[7] [6]);
  and _66793_ (_16063_, _16062_, _16029_);
  or _66794_ (_16064_, _16038_, _15737_);
  and _66795_ (_16065_, _16064_, _16063_);
  and _66796_ (_16066_, _16028_, _15745_);
  or _66797_ (_40706_, _16066_, _16065_);
  or _66798_ (_16067_, _16031_, \oc8051_golden_model_1.IRAM[7] [7]);
  and _66799_ (_16068_, _16067_, _16029_);
  or _66800_ (_16069_, _16038_, _09465_);
  and _66801_ (_16070_, _16069_, _16068_);
  and _66802_ (_16071_, _16028_, _09490_);
  or _66803_ (_40707_, _16071_, _16070_);
  and _66804_ (_16072_, _14356_, _07858_);
  and _66805_ (_16073_, _16072_, _14355_);
  not _66806_ (_16074_, _16073_);
  or _66807_ (_16075_, _16074_, _14528_);
  or _66808_ (_16076_, _16073_, \oc8051_golden_model_1.IRAM[8] [0]);
  not _66809_ (_16077_, _07873_);
  or _66810_ (_16078_, _16077_, _07864_);
  and _66811_ (_16079_, _16078_, _16076_);
  and _66812_ (_16080_, _16079_, _16075_);
  not _66813_ (_16081_, _07866_);
  and _66814_ (_16082_, _07873_, _16081_);
  and _66815_ (_16083_, _16082_, _07296_);
  and _66816_ (_16084_, _16083_, _14543_);
  or _66817_ (_40711_, _16084_, _16080_);
  or _66818_ (_16085_, _16074_, _14727_);
  or _66819_ (_16086_, _16073_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _66820_ (_16087_, _16086_, _16078_);
  and _66821_ (_16088_, _16087_, _16085_);
  and _66822_ (_16089_, _16083_, _14735_);
  or _66823_ (_40712_, _16089_, _16088_);
  or _66824_ (_16090_, _16074_, _14929_);
  or _66825_ (_16091_, _16073_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _66826_ (_16092_, _16091_, _16078_);
  and _66827_ (_16093_, _16092_, _16090_);
  and _66828_ (_16094_, _16083_, _14937_);
  or _66829_ (_40714_, _16094_, _16093_);
  or _66830_ (_16095_, _16074_, _15131_);
  or _66831_ (_16096_, _16073_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _66832_ (_16097_, _16096_, _16078_);
  and _66833_ (_16098_, _16097_, _16095_);
  and _66834_ (_16099_, _16083_, _15139_);
  or _66835_ (_40715_, _16099_, _16098_);
  or _66836_ (_16100_, _16074_, _15332_);
  or _66837_ (_16101_, _16073_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _66838_ (_16102_, _16101_, _16078_);
  and _66839_ (_16103_, _16102_, _16100_);
  and _66840_ (_16104_, _16083_, _15340_);
  or _66841_ (_40716_, _16104_, _16103_);
  or _66842_ (_16105_, _16074_, _15535_);
  or _66843_ (_16106_, _16073_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _66844_ (_16107_, _16106_, _16078_);
  and _66845_ (_16108_, _16107_, _16105_);
  and _66846_ (_16109_, _16083_, _15543_);
  or _66847_ (_40717_, _16109_, _16108_);
  or _66848_ (_16110_, _16074_, _15737_);
  or _66849_ (_16111_, _16073_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _66850_ (_16112_, _16111_, _16078_);
  and _66851_ (_16113_, _16112_, _16110_);
  and _66852_ (_16114_, _16083_, _15745_);
  or _66853_ (_40718_, _16114_, _16113_);
  or _66854_ (_16115_, _16074_, _09465_);
  or _66855_ (_16116_, _16073_, \oc8051_golden_model_1.IRAM[8] [7]);
  and _66856_ (_16117_, _16116_, _16078_);
  and _66857_ (_16118_, _16117_, _16115_);
  and _66858_ (_16119_, _16083_, _09490_);
  or _66859_ (_40720_, _16119_, _16118_);
  and _66860_ (_16120_, _16072_, _15752_);
  not _66861_ (_16121_, _16120_);
  or _66862_ (_16122_, _16121_, _14528_);
  or _66863_ (_16123_, _16120_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand _66864_ (_16124_, _07873_, _07599_);
  and _66865_ (_16125_, _16124_, _16123_);
  and _66866_ (_16126_, _16125_, _16122_);
  and _66867_ (_16127_, _16082_, _07598_);
  and _66868_ (_16128_, _16127_, _14543_);
  or _66869_ (_40723_, _16128_, _16126_);
  or _66870_ (_16129_, _16121_, _14727_);
  or _66871_ (_16130_, _16120_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _66872_ (_16131_, _16130_, _16124_);
  and _66873_ (_16132_, _16131_, _16129_);
  and _66874_ (_16133_, _16127_, _14735_);
  or _66875_ (_40724_, _16133_, _16132_);
  or _66876_ (_16134_, _16121_, _14929_);
  or _66877_ (_16135_, _16120_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _66878_ (_16136_, _16135_, _16124_);
  and _66879_ (_16137_, _16136_, _16134_);
  and _66880_ (_16138_, _16127_, _14937_);
  or _66881_ (_40726_, _16138_, _16137_);
  or _66882_ (_16139_, _16121_, _15131_);
  or _66883_ (_16140_, _16120_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _66884_ (_16141_, _16140_, _16124_);
  and _66885_ (_16142_, _16141_, _16139_);
  and _66886_ (_16143_, _16127_, _15139_);
  or _66887_ (_40727_, _16143_, _16142_);
  or _66888_ (_16144_, _16121_, _15332_);
  or _66889_ (_16145_, _16120_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _66890_ (_16146_, _16145_, _16124_);
  and _66891_ (_16147_, _16146_, _16144_);
  and _66892_ (_16148_, _16127_, _15340_);
  or _66893_ (_40728_, _16148_, _16147_);
  or _66894_ (_16149_, _16121_, _15535_);
  or _66895_ (_16150_, _16120_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _66896_ (_16151_, _16150_, _16124_);
  and _66897_ (_16152_, _16151_, _16149_);
  and _66898_ (_16153_, _16127_, _15543_);
  or _66899_ (_40729_, _16153_, _16152_);
  or _66900_ (_16154_, _16121_, _15737_);
  or _66901_ (_16155_, _16120_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _66902_ (_16156_, _16155_, _16124_);
  and _66903_ (_16157_, _16156_, _16154_);
  and _66904_ (_16158_, _16127_, _15745_);
  or _66905_ (_40730_, _16158_, _16157_);
  or _66906_ (_16159_, _16121_, _09465_);
  or _66907_ (_16160_, _16120_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _66908_ (_16161_, _16160_, _16124_);
  and _66909_ (_16162_, _16161_, _16159_);
  and _66910_ (_16163_, _16127_, _09490_);
  or _66911_ (_40732_, _16163_, _16162_);
  and _66912_ (_16164_, _16072_, _15800_);
  not _66913_ (_16165_, _16164_);
  or _66914_ (_16166_, _16165_, _14528_);
  or _66915_ (_16167_, _16164_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _66916_ (_16168_, _16082_, _08668_);
  not _66917_ (_16169_, _16168_);
  and _66918_ (_16170_, _16169_, _16167_);
  and _66919_ (_16171_, _16170_, _16166_);
  and _66920_ (_16172_, _16168_, _14543_);
  or _66921_ (_40734_, _16172_, _16171_);
  or _66922_ (_16173_, _16165_, _14727_);
  or _66923_ (_16174_, _16164_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _66924_ (_16175_, _16174_, _16169_);
  and _66925_ (_16176_, _16175_, _16173_);
  and _66926_ (_16177_, _16168_, _14735_);
  or _66927_ (_40736_, _16177_, _16176_);
  or _66928_ (_16178_, _16165_, _14929_);
  or _66929_ (_16179_, _16164_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _66930_ (_16180_, _16179_, _16169_);
  and _66931_ (_16181_, _16180_, _16178_);
  and _66932_ (_16182_, _16168_, _14937_);
  or _66933_ (_40737_, _16182_, _16181_);
  or _66934_ (_16183_, _16165_, _15131_);
  or _66935_ (_16184_, _16164_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _66936_ (_16185_, _16184_, _16169_);
  and _66937_ (_16186_, _16185_, _16183_);
  and _66938_ (_16187_, _16168_, _15139_);
  or _66939_ (_40738_, _16187_, _16186_);
  or _66940_ (_16188_, _16165_, _15332_);
  or _66941_ (_16189_, _16164_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _66942_ (_16190_, _16189_, _16169_);
  and _66943_ (_16191_, _16190_, _16188_);
  and _66944_ (_16192_, _16168_, _15340_);
  or _66945_ (_40739_, _16192_, _16191_);
  or _66946_ (_16193_, _16165_, _15535_);
  or _66947_ (_16194_, _16164_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _66948_ (_16195_, _16194_, _16169_);
  and _66949_ (_16196_, _16195_, _16193_);
  and _66950_ (_16197_, _16168_, _15543_);
  or _66951_ (_40740_, _16197_, _16196_);
  or _66952_ (_16198_, _16165_, _15737_);
  or _66953_ (_16199_, _16164_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _66954_ (_16200_, _16199_, _16169_);
  and _66955_ (_16201_, _16200_, _16198_);
  and _66956_ (_16202_, _16168_, _15745_);
  or _66957_ (_40742_, _16202_, _16201_);
  or _66958_ (_16203_, _16165_, _09465_);
  or _66959_ (_16204_, _16164_, \oc8051_golden_model_1.IRAM[10] [7]);
  and _66960_ (_16205_, _16204_, _16169_);
  and _66961_ (_16206_, _16205_, _16203_);
  and _66962_ (_16207_, _16168_, _09490_);
  or _66963_ (_40743_, _16207_, _16206_);
  not _66964_ (_16208_, _07453_);
  and _66965_ (_16209_, _14354_, _16208_);
  and _66966_ (_16210_, _16072_, _16209_);
  not _66967_ (_16211_, _16210_);
  or _66968_ (_16212_, _16211_, _14528_);
  and _66969_ (_16213_, _16082_, _07295_);
  not _66970_ (_16214_, _16213_);
  or _66971_ (_16215_, _16210_, \oc8051_golden_model_1.IRAM[11] [0]);
  and _66972_ (_16216_, _16215_, _16214_);
  and _66973_ (_16217_, _16216_, _16212_);
  and _66974_ (_16218_, _16213_, _14543_);
  or _66975_ (_40746_, _16218_, _16217_);
  and _66976_ (_16219_, _16072_, _07538_);
  or _66977_ (_16220_, _16219_, \oc8051_golden_model_1.IRAM[11] [1]);
  and _66978_ (_16221_, _16220_, _16214_);
  not _66979_ (_16222_, _16219_);
  or _66980_ (_16223_, _16222_, _14727_);
  and _66981_ (_16224_, _16223_, _16221_);
  and _66982_ (_16225_, _16213_, _14735_);
  or _66983_ (_40748_, _16225_, _16224_);
  or _66984_ (_16226_, _16211_, _14929_);
  or _66985_ (_16227_, _16210_, \oc8051_golden_model_1.IRAM[11] [2]);
  and _66986_ (_16228_, _16227_, _16214_);
  and _66987_ (_16229_, _16228_, _16226_);
  and _66988_ (_16230_, _16213_, _14937_);
  or _66989_ (_40749_, _16230_, _16229_);
  or _66990_ (_16231_, _16219_, \oc8051_golden_model_1.IRAM[11] [3]);
  and _66991_ (_16232_, _16231_, _16214_);
  or _66992_ (_16233_, _16222_, _15131_);
  and _66993_ (_16234_, _16233_, _16232_);
  and _66994_ (_16235_, _16213_, _15139_);
  or _66995_ (_40750_, _16235_, _16234_);
  or _66996_ (_16236_, _16219_, \oc8051_golden_model_1.IRAM[11] [4]);
  and _66997_ (_16237_, _16236_, _16214_);
  or _66998_ (_16238_, _16222_, _15332_);
  and _66999_ (_16239_, _16238_, _16237_);
  and _67000_ (_16240_, _16213_, _15340_);
  or _67001_ (_40751_, _16240_, _16239_);
  or _67002_ (_16241_, _16219_, \oc8051_golden_model_1.IRAM[11] [5]);
  and _67003_ (_16242_, _16241_, _16214_);
  or _67004_ (_16243_, _16222_, _15535_);
  and _67005_ (_16244_, _16243_, _16242_);
  and _67006_ (_16245_, _16213_, _15543_);
  or _67007_ (_40752_, _16245_, _16244_);
  or _67008_ (_16246_, _16219_, \oc8051_golden_model_1.IRAM[11] [6]);
  and _67009_ (_16247_, _16246_, _16214_);
  or _67010_ (_16248_, _16222_, _15737_);
  and _67011_ (_16249_, _16248_, _16247_);
  and _67012_ (_16250_, _16213_, _15745_);
  or _67013_ (_40754_, _16250_, _16249_);
  or _67014_ (_16251_, _16219_, \oc8051_golden_model_1.IRAM[11] [7]);
  and _67015_ (_16252_, _16251_, _16214_);
  or _67016_ (_16253_, _16222_, _09465_);
  and _67017_ (_16254_, _16253_, _16252_);
  and _67018_ (_16255_, _16213_, _09490_);
  or _67019_ (_40755_, _16255_, _16254_);
  not _67020_ (_16256_, _07296_);
  nand _67021_ (_16257_, _14532_, _07869_);
  or _67022_ (_16258_, _16257_, _16256_);
  nor _67023_ (_16259_, _16258_, _14543_);
  and _67024_ (_16260_, _14355_, _07861_);
  nand _67025_ (_16261_, _16260_, _14528_);
  or _67026_ (_16262_, _16260_, _07124_);
  and _67027_ (_16263_, _16262_, _16258_);
  and _67028_ (_16264_, _16263_, _16261_);
  nor _67029_ (_40759_, _16264_, _16259_);
  and _67030_ (_16265_, _07874_, _07296_);
  not _67031_ (_16266_, _16265_);
  or _67032_ (_16267_, _16260_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _67033_ (_16268_, _16267_, _16266_);
  not _67034_ (_16269_, _16260_);
  or _67035_ (_16270_, _16269_, _14727_);
  and _67036_ (_16271_, _16270_, _16268_);
  and _67037_ (_16272_, _16265_, _14735_);
  or _67038_ (_40760_, _16272_, _16271_);
  or _67039_ (_16273_, _16260_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _67040_ (_16274_, _16273_, _16266_);
  or _67041_ (_16275_, _16269_, _14929_);
  and _67042_ (_16276_, _16275_, _16274_);
  and _67043_ (_16277_, _16265_, _14937_);
  or _67044_ (_40761_, _16277_, _16276_);
  or _67045_ (_16278_, _16260_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _67046_ (_16279_, _16278_, _16266_);
  or _67047_ (_16280_, _16269_, _15131_);
  and _67048_ (_16281_, _16280_, _16279_);
  and _67049_ (_16282_, _16265_, _15139_);
  or _67050_ (_40762_, _16282_, _16281_);
  or _67051_ (_16283_, _16260_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _67052_ (_16284_, _16283_, _16266_);
  or _67053_ (_16285_, _16269_, _15332_);
  and _67054_ (_16286_, _16285_, _16284_);
  and _67055_ (_16287_, _16265_, _15340_);
  or _67056_ (_40764_, _16287_, _16286_);
  or _67057_ (_16288_, _16260_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _67058_ (_16289_, _16288_, _16266_);
  or _67059_ (_16290_, _16269_, _15535_);
  and _67060_ (_16291_, _16290_, _16289_);
  and _67061_ (_16292_, _16265_, _15543_);
  or _67062_ (_40765_, _16292_, _16291_);
  or _67063_ (_16293_, _16260_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _67064_ (_16294_, _16293_, _16266_);
  or _67065_ (_16295_, _16269_, _15737_);
  and _67066_ (_16296_, _16295_, _16294_);
  and _67067_ (_16297_, _16265_, _15745_);
  or _67068_ (_40766_, _16297_, _16296_);
  or _67069_ (_16298_, _16260_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _67070_ (_16299_, _16298_, _16266_);
  or _67071_ (_16300_, _16269_, _09465_);
  and _67072_ (_16301_, _16300_, _16299_);
  and _67073_ (_16302_, _16265_, _09490_);
  or _67074_ (_40767_, _16302_, _16301_);
  and _67075_ (_16303_, _15752_, _07861_);
  or _67076_ (_16304_, _16303_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _67077_ (_16305_, _07874_, _07598_);
  not _67078_ (_16306_, _16305_);
  and _67079_ (_16307_, _16306_, _16304_);
  not _67080_ (_16308_, _16303_);
  or _67081_ (_16309_, _16308_, _14528_);
  and _67082_ (_16310_, _16309_, _16307_);
  and _67083_ (_16311_, _16305_, _14543_);
  or _67084_ (_40771_, _16311_, _16310_);
  or _67085_ (_16312_, _16303_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _67086_ (_16313_, _16312_, _16306_);
  or _67087_ (_16314_, _16308_, _14727_);
  and _67088_ (_16315_, _16314_, _16313_);
  and _67089_ (_16316_, _16305_, _14735_);
  or _67090_ (_40772_, _16316_, _16315_);
  or _67091_ (_16317_, _16303_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _67092_ (_16318_, _16317_, _16306_);
  or _67093_ (_16319_, _16308_, _14929_);
  and _67094_ (_16320_, _16319_, _16318_);
  and _67095_ (_16321_, _16305_, _14937_);
  or _67096_ (_40773_, _16321_, _16320_);
  or _67097_ (_16322_, _16303_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _67098_ (_16323_, _16322_, _16306_);
  or _67099_ (_16324_, _16308_, _15131_);
  and _67100_ (_16325_, _16324_, _16323_);
  and _67101_ (_16326_, _16305_, _15139_);
  or _67102_ (_40774_, _16326_, _16325_);
  or _67103_ (_16327_, _16303_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _67104_ (_16328_, _16327_, _16306_);
  or _67105_ (_16329_, _16308_, _15332_);
  and _67106_ (_16330_, _16329_, _16328_);
  and _67107_ (_16331_, _16305_, _15340_);
  or _67108_ (_40776_, _16331_, _16330_);
  or _67109_ (_16332_, _16303_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _67110_ (_16333_, _16332_, _16306_);
  or _67111_ (_16334_, _16308_, _15535_);
  and _67112_ (_16335_, _16334_, _16333_);
  and _67113_ (_16336_, _16305_, _15543_);
  or _67114_ (_40777_, _16336_, _16335_);
  or _67115_ (_16337_, _16303_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _67116_ (_16338_, _16337_, _16306_);
  or _67117_ (_16339_, _16308_, _15737_);
  and _67118_ (_16340_, _16339_, _16338_);
  and _67119_ (_16341_, _16305_, _15745_);
  or _67120_ (_40778_, _16341_, _16340_);
  or _67121_ (_16342_, _16303_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _67122_ (_16343_, _16342_, _16306_);
  or _67123_ (_16344_, _16308_, _09465_);
  and _67124_ (_16345_, _16344_, _16343_);
  and _67125_ (_16346_, _16305_, _09490_);
  or _67126_ (_40779_, _16346_, _16345_);
  and _67127_ (_16347_, _15800_, _07861_);
  or _67128_ (_16348_, _16347_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _67129_ (_16349_, _08668_, _07874_);
  not _67130_ (_16350_, _16349_);
  and _67131_ (_16351_, _16350_, _16348_);
  not _67132_ (_16352_, _16347_);
  or _67133_ (_16353_, _16352_, _14528_);
  and _67134_ (_16354_, _16353_, _16351_);
  and _67135_ (_16355_, _16349_, _14543_);
  or _67136_ (_40783_, _16355_, _16354_);
  or _67137_ (_16356_, _16347_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _67138_ (_16357_, _16356_, _16350_);
  or _67139_ (_16358_, _16352_, _14727_);
  and _67140_ (_16359_, _16358_, _16357_);
  and _67141_ (_16360_, _16349_, _14735_);
  or _67142_ (_40784_, _16360_, _16359_);
  not _67143_ (_16361_, _08668_);
  or _67144_ (_16362_, _16361_, _16257_);
  nor _67145_ (_16363_, _16347_, _07764_);
  and _67146_ (_16364_, _16347_, _14929_);
  or _67147_ (_16365_, _16364_, _16363_);
  and _67148_ (_16366_, _16365_, _16362_);
  and _67149_ (_16367_, _16349_, _14937_);
  or _67150_ (_40785_, _16367_, _16366_);
  or _67151_ (_16368_, _16347_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _67152_ (_16369_, _16368_, _16350_);
  or _67153_ (_16370_, _16352_, _15131_);
  and _67154_ (_16371_, _16370_, _16369_);
  and _67155_ (_16372_, _16349_, _15139_);
  or _67156_ (_40787_, _16372_, _16371_);
  or _67157_ (_16373_, _16347_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _67158_ (_16374_, _16373_, _16350_);
  or _67159_ (_16375_, _16352_, _15332_);
  and _67160_ (_16376_, _16375_, _16374_);
  and _67161_ (_16377_, _16349_, _15340_);
  or _67162_ (_40788_, _16377_, _16376_);
  or _67163_ (_16378_, _16347_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _67164_ (_16379_, _16378_, _16350_);
  or _67165_ (_16380_, _16352_, _15535_);
  and _67166_ (_16381_, _16380_, _16379_);
  and _67167_ (_16382_, _16349_, _15543_);
  or _67168_ (_40789_, _16382_, _16381_);
  or _67169_ (_16383_, _16347_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _67170_ (_16384_, _16383_, _16350_);
  or _67171_ (_16385_, _16352_, _15737_);
  and _67172_ (_16386_, _16385_, _16384_);
  and _67173_ (_16387_, _16349_, _15745_);
  or _67174_ (_40790_, _16387_, _16386_);
  or _67175_ (_16388_, _16347_, \oc8051_golden_model_1.IRAM[14] [7]);
  and _67176_ (_16389_, _16388_, _16350_);
  or _67177_ (_16390_, _16352_, _09465_);
  and _67178_ (_16391_, _16390_, _16389_);
  and _67179_ (_16392_, _16349_, _09490_);
  or _67180_ (_40791_, _16392_, _16391_);
  not _67181_ (_16393_, _07295_);
  or _67182_ (_16394_, _16257_, _16393_);
  or _67183_ (_16395_, _14543_, _16394_);
  and _67184_ (_16396_, _14528_, _07862_);
  or _67185_ (_16397_, _07862_, _07119_);
  nand _67186_ (_16398_, _16397_, _16394_);
  or _67187_ (_16399_, _16398_, _16396_);
  and _67188_ (_40795_, _16399_, _16395_);
  or _67189_ (_16400_, _07862_, \oc8051_golden_model_1.IRAM[15] [1]);
  and _67190_ (_16401_, _16400_, _07876_);
  or _67191_ (_16402_, _14727_, _07878_);
  and _67192_ (_16403_, _16402_, _16401_);
  and _67193_ (_16404_, _14735_, _07875_);
  or _67194_ (_40796_, _16404_, _16403_);
  nor _67195_ (_16405_, _07862_, _07762_);
  and _67196_ (_16406_, _14929_, _07862_);
  or _67197_ (_16407_, _16406_, _16405_);
  and _67198_ (_16408_, _16407_, _16394_);
  and _67199_ (_16409_, _14937_, _07875_);
  or _67200_ (_40797_, _16409_, _16408_);
  or _67201_ (_16410_, _07862_, \oc8051_golden_model_1.IRAM[15] [3]);
  and _67202_ (_16411_, _16410_, _07876_);
  or _67203_ (_16412_, _15131_, _07878_);
  and _67204_ (_16413_, _16412_, _16411_);
  and _67205_ (_16414_, _15139_, _07875_);
  or _67206_ (_40799_, _16414_, _16413_);
  or _67207_ (_16415_, _15332_, _07878_);
  or _67208_ (_16416_, _07862_, \oc8051_golden_model_1.IRAM[15] [4]);
  and _67209_ (_16417_, _16416_, _07876_);
  and _67210_ (_16418_, _16417_, _16415_);
  and _67211_ (_16419_, _15340_, _07875_);
  or _67212_ (_40800_, _16419_, _16418_);
  or _67213_ (_16420_, _07862_, \oc8051_golden_model_1.IRAM[15] [5]);
  and _67214_ (_16421_, _16420_, _07876_);
  or _67215_ (_16422_, _15535_, _07878_);
  and _67216_ (_16423_, _16422_, _16421_);
  and _67217_ (_16424_, _15543_, _07875_);
  or _67218_ (_40801_, _16424_, _16423_);
  or _67219_ (_16425_, _15737_, _07878_);
  or _67220_ (_16426_, _07862_, \oc8051_golden_model_1.IRAM[15] [6]);
  and _67221_ (_16427_, _16426_, _07876_);
  and _67222_ (_16428_, _16427_, _16425_);
  and _67223_ (_16429_, _15745_, _07875_);
  or _67224_ (_40802_, _16429_, _16428_);
  nor _67225_ (_16430_, _01347_, _10106_);
  nand _67226_ (_16431_, _11263_, _07942_);
  nor _67227_ (_16432_, _07942_, _10106_);
  nor _67228_ (_16433_, _16432_, _07234_);
  nand _67229_ (_16434_, _16433_, _16431_);
  and _67230_ (_16435_, _07942_, _08954_);
  or _67231_ (_16436_, _16435_, _16432_);
  or _67232_ (_16437_, _16436_, _06219_);
  and _67233_ (_16438_, _07942_, _07133_);
  or _67234_ (_16439_, _16438_, _16432_);
  or _67235_ (_16440_, _16439_, _07215_);
  nor _67236_ (_16441_, _08390_, _09498_);
  or _67237_ (_16442_, _16441_, _16432_);
  or _67238_ (_16443_, _16442_, _07151_);
  and _67239_ (_16444_, _07942_, \oc8051_golden_model_1.ACC [0]);
  or _67240_ (_16445_, _16444_, _16432_);
  and _67241_ (_16446_, _16445_, _07141_);
  nor _67242_ (_16447_, _07141_, _10106_);
  or _67243_ (_16448_, _16447_, _06341_);
  or _67244_ (_16449_, _16448_, _16446_);
  and _67245_ (_16450_, _16449_, _06273_);
  and _67246_ (_16451_, _16450_, _16443_);
  and _67247_ (_16452_, _14382_, _08634_);
  nor _67248_ (_16453_, _08634_, _10106_);
  or _67249_ (_16454_, _16453_, _16452_);
  and _67250_ (_16455_, _16454_, _06272_);
  or _67251_ (_16456_, _16455_, _16451_);
  and _67252_ (_16457_, _16456_, _07166_);
  and _67253_ (_16458_, _16439_, _06461_);
  or _67254_ (_16459_, _16458_, _06464_);
  or _67255_ (_16460_, _16459_, _16457_);
  or _67256_ (_16461_, _16445_, _06465_);
  and _67257_ (_16462_, _16461_, _06269_);
  and _67258_ (_16463_, _16462_, _16460_);
  and _67259_ (_16464_, _16432_, _06268_);
  or _67260_ (_16465_, _16464_, _06261_);
  or _67261_ (_16466_, _16465_, _16463_);
  or _67262_ (_16467_, _16442_, _06262_);
  and _67263_ (_16468_, _16467_, _16466_);
  or _67264_ (_16469_, _16468_, _09531_);
  nor _67265_ (_16470_, _10052_, _10050_);
  nor _67266_ (_16471_, _16470_, _10053_);
  or _67267_ (_16472_, _16471_, _09537_);
  and _67268_ (_16473_, _16472_, _06258_);
  and _67269_ (_16474_, _16473_, _16469_);
  and _67270_ (_16475_, _14413_, _08634_);
  or _67271_ (_16476_, _16475_, _16453_);
  and _67272_ (_16477_, _16476_, _06257_);
  or _67273_ (_16478_, _16477_, _10080_);
  or _67274_ (_16479_, _16478_, _16474_);
  and _67275_ (_16480_, _16479_, _16440_);
  or _67276_ (_16481_, _16480_, _07460_);
  and _67277_ (_16482_, _09392_, _07942_);
  or _67278_ (_16483_, _16432_, _07208_);
  or _67279_ (_16484_, _16483_, _16482_);
  and _67280_ (_16485_, _16484_, _16481_);
  or _67281_ (_16486_, _16485_, _10094_);
  and _67282_ (_16487_, _14467_, _07942_);
  or _67283_ (_16488_, _16432_, _05982_);
  or _67284_ (_16489_, _16488_, _16487_);
  and _67285_ (_16490_, _16489_, _10100_);
  and _67286_ (_16491_, _16490_, _16486_);
  nand _67287_ (_16492_, _10439_, _06097_);
  or _67288_ (_16493_, _10433_, _10408_);
  or _67289_ (_16494_, _10439_, _16493_);
  and _67290_ (_16495_, _16494_, _10093_);
  and _67291_ (_16496_, _16495_, _16492_);
  or _67292_ (_16497_, _16496_, _06218_);
  or _67293_ (_16498_, _16497_, _16491_);
  and _67294_ (_16499_, _16498_, _16437_);
  or _67295_ (_16500_, _16499_, _06369_);
  and _67296_ (_16501_, _14366_, _07942_);
  or _67297_ (_16502_, _16501_, _16432_);
  or _67298_ (_16503_, _16502_, _07237_);
  and _67299_ (_16504_, _16503_, _07240_);
  and _67300_ (_16505_, _16504_, _16500_);
  nor _67301_ (_16506_, _12580_, _09498_);
  or _67302_ (_16507_, _16506_, _16432_);
  and _67303_ (_16508_, _16431_, _06536_);
  and _67304_ (_16509_, _16508_, _16507_);
  or _67305_ (_16510_, _16509_, _16505_);
  and _67306_ (_16511_, _16510_, _07242_);
  nand _67307_ (_16512_, _16436_, _06375_);
  nor _67308_ (_16513_, _16512_, _16441_);
  or _67309_ (_16514_, _16513_, _06545_);
  or _67310_ (_16515_, _16514_, _16511_);
  and _67311_ (_16516_, _16515_, _16434_);
  or _67312_ (_16517_, _16516_, _06366_);
  and _67313_ (_16518_, _14363_, _07942_);
  or _67314_ (_16519_, _16432_, _09056_);
  or _67315_ (_16520_, _16519_, _16518_);
  and _67316_ (_16521_, _16520_, _09061_);
  and _67317_ (_16522_, _16521_, _16517_);
  and _67318_ (_16523_, _16507_, _06528_);
  or _67319_ (_16524_, _16523_, _06568_);
  or _67320_ (_16525_, _16524_, _16522_);
  or _67321_ (_16526_, _16442_, _06926_);
  and _67322_ (_16527_, _16526_, _16525_);
  or _67323_ (_16528_, _16527_, _05927_);
  or _67324_ (_16529_, _16432_, _05928_);
  and _67325_ (_16530_, _16529_, _16528_);
  or _67326_ (_16531_, _16530_, _06278_);
  or _67327_ (_16532_, _16442_, _06279_);
  and _67328_ (_16533_, _16532_, _01347_);
  and _67329_ (_16534_, _16533_, _16531_);
  or _67330_ (_16535_, _16534_, _16430_);
  and _67331_ (_43153_, _16535_, _42618_);
  nor _67332_ (_16536_, _01347_, _10101_);
  nor _67333_ (_16537_, _07942_, _10101_);
  nor _67334_ (_16538_, _11261_, _09498_);
  or _67335_ (_16539_, _16538_, _16537_);
  or _67336_ (_16540_, _16539_, _09061_);
  or _67337_ (_16541_, _07942_, \oc8051_golden_model_1.B [1]);
  nand _67338_ (_16542_, _07942_, _07038_);
  and _67339_ (_16543_, _16542_, _06218_);
  and _67340_ (_16544_, _16543_, _16541_);
  nor _67341_ (_16545_, _08634_, _10101_);
  and _67342_ (_16546_, _14560_, _08634_);
  or _67343_ (_16547_, _16546_, _16545_);
  and _67344_ (_16548_, _16547_, _06268_);
  nor _67345_ (_16549_, _09498_, _07357_);
  or _67346_ (_16550_, _16549_, _16537_);
  or _67347_ (_16551_, _16550_, _07166_);
  and _67348_ (_16552_, _14562_, _07942_);
  not _67349_ (_16553_, _16552_);
  and _67350_ (_16554_, _16553_, _16541_);
  or _67351_ (_16555_, _16554_, _07151_);
  and _67352_ (_16556_, _07942_, \oc8051_golden_model_1.ACC [1]);
  or _67353_ (_16557_, _16556_, _16537_);
  and _67354_ (_16558_, _16557_, _07141_);
  nor _67355_ (_16559_, _07141_, _10101_);
  or _67356_ (_16560_, _16559_, _06341_);
  or _67357_ (_16561_, _16560_, _16558_);
  and _67358_ (_16562_, _16561_, _06273_);
  and _67359_ (_16563_, _16562_, _16555_);
  and _67360_ (_16564_, _14557_, _08634_);
  or _67361_ (_16565_, _16564_, _16545_);
  and _67362_ (_16566_, _16565_, _06272_);
  or _67363_ (_16567_, _16566_, _06461_);
  or _67364_ (_16568_, _16567_, _16563_);
  and _67365_ (_16569_, _16568_, _16551_);
  or _67366_ (_16570_, _16569_, _06464_);
  or _67367_ (_16571_, _16557_, _06465_);
  and _67368_ (_16572_, _16571_, _06269_);
  and _67369_ (_16573_, _16572_, _16570_);
  or _67370_ (_16574_, _16573_, _16548_);
  and _67371_ (_16575_, _16574_, _06262_);
  and _67372_ (_16576_, _16564_, _14556_);
  or _67373_ (_16577_, _16576_, _16545_);
  and _67374_ (_16578_, _16577_, _06261_);
  or _67375_ (_16579_, _16578_, _09531_);
  or _67376_ (_16580_, _16579_, _16575_);
  nor _67377_ (_16581_, _10055_, _09997_);
  nor _67378_ (_16582_, _16581_, _10056_);
  or _67379_ (_16583_, _16582_, _09537_);
  and _67380_ (_16584_, _16583_, _06258_);
  and _67381_ (_16585_, _16584_, _16580_);
  or _67382_ (_16586_, _16545_, _14597_);
  and _67383_ (_16587_, _16586_, _06257_);
  and _67384_ (_16588_, _16587_, _16565_);
  or _67385_ (_16589_, _16588_, _10080_);
  or _67386_ (_16590_, _16589_, _16585_);
  or _67387_ (_16591_, _16550_, _07215_);
  and _67388_ (_16592_, _16591_, _16590_);
  or _67389_ (_16593_, _16592_, _07460_);
  and _67390_ (_16594_, _09451_, _07942_);
  or _67391_ (_16595_, _16537_, _07208_);
  or _67392_ (_16596_, _16595_, _16594_);
  and _67393_ (_16597_, _16596_, _05982_);
  and _67394_ (_16598_, _16597_, _16593_);
  or _67395_ (_16599_, _14653_, _09498_);
  and _67396_ (_16600_, _16541_, _10094_);
  and _67397_ (_16601_, _16600_, _16599_);
  or _67398_ (_16602_, _16601_, _10093_);
  or _67399_ (_16603_, _16602_, _16598_);
  nor _67400_ (_16604_, _10434_, _10432_);
  or _67401_ (_16605_, _16604_, _10435_);
  nor _67402_ (_16606_, _16605_, _10439_);
  and _67403_ (_16607_, _10439_, _10405_);
  or _67404_ (_16608_, _16607_, _16606_);
  or _67405_ (_16609_, _16608_, _10100_);
  and _67406_ (_16610_, _16609_, _06219_);
  and _67407_ (_16611_, _16610_, _16603_);
  or _67408_ (_16612_, _16611_, _16544_);
  and _67409_ (_16613_, _16612_, _07237_);
  or _67410_ (_16614_, _14668_, _09498_);
  and _67411_ (_16615_, _16541_, _06369_);
  and _67412_ (_16616_, _16615_, _16614_);
  or _67413_ (_16617_, _16616_, _06536_);
  or _67414_ (_16618_, _16617_, _16613_);
  and _67415_ (_16619_, _11262_, _07942_);
  or _67416_ (_16620_, _16619_, _16537_);
  or _67417_ (_16621_, _16620_, _07240_);
  and _67418_ (_16622_, _16621_, _07242_);
  and _67419_ (_16623_, _16622_, _16618_);
  or _67420_ (_16624_, _14666_, _09498_);
  and _67421_ (_16625_, _16541_, _06375_);
  and _67422_ (_16626_, _16625_, _16624_);
  or _67423_ (_16627_, _16626_, _06545_);
  or _67424_ (_16628_, _16627_, _16623_);
  and _67425_ (_16629_, _16556_, _08341_);
  or _67426_ (_16630_, _16537_, _07234_);
  or _67427_ (_16631_, _16630_, _16629_);
  and _67428_ (_16632_, _16631_, _09056_);
  and _67429_ (_16633_, _16632_, _16628_);
  or _67430_ (_16634_, _16542_, _08341_);
  and _67431_ (_16635_, _16541_, _06366_);
  and _67432_ (_16636_, _16635_, _16634_);
  or _67433_ (_16637_, _16636_, _06528_);
  or _67434_ (_16638_, _16637_, _16633_);
  and _67435_ (_16639_, _16638_, _16540_);
  or _67436_ (_16640_, _16639_, _06568_);
  or _67437_ (_16641_, _16554_, _06926_);
  and _67438_ (_16642_, _16641_, _05928_);
  and _67439_ (_16643_, _16642_, _16640_);
  and _67440_ (_16644_, _16547_, _05927_);
  or _67441_ (_16645_, _16644_, _06278_);
  or _67442_ (_16646_, _16645_, _16643_);
  or _67443_ (_16647_, _16537_, _06279_);
  or _67444_ (_16648_, _16647_, _16552_);
  and _67445_ (_16649_, _16648_, _01347_);
  and _67446_ (_16650_, _16649_, _16646_);
  or _67447_ (_16651_, _16650_, _16536_);
  and _67448_ (_43154_, _16651_, _42618_);
  nor _67449_ (_16652_, _01347_, _10159_);
  nor _67450_ (_16653_, _07942_, _10159_);
  and _67451_ (_16654_, _07942_, _08973_);
  or _67452_ (_16655_, _16654_, _16653_);
  or _67453_ (_16656_, _16655_, _06219_);
  nor _67454_ (_16657_, _09498_, _07776_);
  or _67455_ (_16658_, _16657_, _16653_);
  or _67456_ (_16659_, _16658_, _07215_);
  and _67457_ (_16660_, _14774_, _08634_);
  and _67458_ (_16661_, _16660_, _14789_);
  nor _67459_ (_16662_, _08634_, _10159_);
  or _67460_ (_16663_, _16662_, _06262_);
  or _67461_ (_16664_, _16663_, _16661_);
  or _67462_ (_16665_, _16658_, _07166_);
  and _67463_ (_16666_, _14770_, _07942_);
  or _67464_ (_16667_, _16666_, _16653_);
  or _67465_ (_16668_, _16667_, _07151_);
  and _67466_ (_16669_, _07942_, \oc8051_golden_model_1.ACC [2]);
  or _67467_ (_16670_, _16669_, _16653_);
  and _67468_ (_16671_, _16670_, _07141_);
  nor _67469_ (_16672_, _07141_, _10159_);
  or _67470_ (_16673_, _16672_, _06341_);
  or _67471_ (_16674_, _16673_, _16671_);
  and _67472_ (_16675_, _16674_, _06273_);
  and _67473_ (_16676_, _16675_, _16668_);
  or _67474_ (_16677_, _16662_, _16660_);
  and _67475_ (_16678_, _16677_, _06272_);
  or _67476_ (_16679_, _16678_, _06461_);
  or _67477_ (_16680_, _16679_, _16676_);
  and _67478_ (_16681_, _16680_, _16665_);
  or _67479_ (_16682_, _16681_, _06464_);
  or _67480_ (_16683_, _16670_, _06465_);
  and _67481_ (_16684_, _16683_, _06269_);
  and _67482_ (_16685_, _16684_, _16682_);
  and _67483_ (_16686_, _14756_, _08634_);
  or _67484_ (_16687_, _16686_, _16662_);
  and _67485_ (_16688_, _16687_, _06268_);
  or _67486_ (_16689_, _16688_, _06261_);
  or _67487_ (_16690_, _16689_, _16685_);
  and _67488_ (_16691_, _16690_, _16664_);
  or _67489_ (_16692_, _16691_, _09531_);
  or _67490_ (_16693_, _10057_, _09952_);
  and _67491_ (_16694_, _16693_, _10058_);
  or _67492_ (_16695_, _16694_, _09537_);
  and _67493_ (_16696_, _16695_, _06258_);
  and _67494_ (_16697_, _16696_, _16692_);
  and _67495_ (_16698_, _14804_, _08634_);
  or _67496_ (_16699_, _16698_, _16662_);
  and _67497_ (_16700_, _16699_, _06257_);
  or _67498_ (_16701_, _16700_, _10080_);
  or _67499_ (_16702_, _16701_, _16697_);
  and _67500_ (_16703_, _16702_, _16659_);
  or _67501_ (_16704_, _16703_, _07460_);
  and _67502_ (_16705_, _09450_, _07942_);
  or _67503_ (_16706_, _16653_, _07208_);
  or _67504_ (_16707_, _16706_, _16705_);
  and _67505_ (_16708_, _16707_, _16704_);
  or _67506_ (_16709_, _16708_, _10094_);
  and _67507_ (_16710_, _14859_, _07942_);
  or _67508_ (_16711_, _16653_, _05982_);
  or _67509_ (_16712_, _16711_, _16710_);
  and _67510_ (_16713_, _16712_, _10100_);
  and _67511_ (_16714_, _16713_, _16709_);
  not _67512_ (_16715_, _10439_);
  or _67513_ (_16716_, _16715_, _10396_);
  nor _67514_ (_16717_, _10435_, _10406_);
  not _67515_ (_16718_, _16717_);
  and _67516_ (_16719_, _16718_, _10399_);
  nor _67517_ (_16720_, _16718_, _10399_);
  nor _67518_ (_16721_, _16720_, _16719_);
  or _67519_ (_16722_, _16721_, _10439_);
  and _67520_ (_16723_, _16722_, _10093_);
  and _67521_ (_16724_, _16723_, _16716_);
  or _67522_ (_16725_, _16724_, _06218_);
  or _67523_ (_16726_, _16725_, _16714_);
  and _67524_ (_16727_, _16726_, _16656_);
  or _67525_ (_16728_, _16727_, _06369_);
  and _67526_ (_16729_, _14751_, _07942_);
  or _67527_ (_16730_, _16729_, _16653_);
  or _67528_ (_16731_, _16730_, _07237_);
  and _67529_ (_16732_, _16731_, _07240_);
  and _67530_ (_16733_, _16732_, _16728_);
  and _67531_ (_16734_, _11259_, _07942_);
  or _67532_ (_16735_, _16734_, _16653_);
  and _67533_ (_16736_, _16735_, _06536_);
  or _67534_ (_16737_, _16736_, _16733_);
  and _67535_ (_16738_, _16737_, _07242_);
  or _67536_ (_16739_, _16653_, _08440_);
  and _67537_ (_16740_, _16655_, _06375_);
  and _67538_ (_16741_, _16740_, _16739_);
  or _67539_ (_16742_, _16741_, _16738_);
  and _67540_ (_16743_, _16742_, _07234_);
  and _67541_ (_16744_, _16670_, _06545_);
  and _67542_ (_16745_, _16744_, _16739_);
  or _67543_ (_16746_, _16745_, _06366_);
  or _67544_ (_16747_, _16746_, _16743_);
  and _67545_ (_16748_, _14748_, _07942_);
  or _67546_ (_16749_, _16653_, _09056_);
  or _67547_ (_16750_, _16749_, _16748_);
  and _67548_ (_16751_, _16750_, _09061_);
  and _67549_ (_16752_, _16751_, _16747_);
  nor _67550_ (_16753_, _11258_, _09498_);
  or _67551_ (_16754_, _16753_, _16653_);
  and _67552_ (_16755_, _16754_, _06528_);
  or _67553_ (_16756_, _16755_, _06568_);
  or _67554_ (_16757_, _16756_, _16752_);
  or _67555_ (_16758_, _16667_, _06926_);
  and _67556_ (_16759_, _16758_, _05928_);
  and _67557_ (_16760_, _16759_, _16757_);
  and _67558_ (_16761_, _16687_, _05927_);
  or _67559_ (_16762_, _16761_, _06278_);
  or _67560_ (_16763_, _16762_, _16760_);
  and _67561_ (_16764_, _14926_, _07942_);
  or _67562_ (_16765_, _16653_, _06279_);
  or _67563_ (_16766_, _16765_, _16764_);
  and _67564_ (_16767_, _16766_, _01347_);
  and _67565_ (_16768_, _16767_, _16763_);
  or _67566_ (_16769_, _16768_, _16652_);
  and _67567_ (_43155_, _16769_, _42618_);
  nor _67568_ (_16770_, _01347_, _10145_);
  nor _67569_ (_16771_, _07942_, _10145_);
  and _67570_ (_16772_, _07942_, _08930_);
  or _67571_ (_16773_, _16772_, _16771_);
  or _67572_ (_16774_, _16773_, _06219_);
  and _67573_ (_16775_, _15048_, _07942_);
  or _67574_ (_16776_, _16775_, _16771_);
  and _67575_ (_16777_, _16776_, _10094_);
  nor _67576_ (_16778_, _08634_, _10145_);
  and _67577_ (_16779_, _14950_, _08634_);
  or _67578_ (_16780_, _16779_, _16778_);
  or _67579_ (_16781_, _16778_, _14979_);
  and _67580_ (_16782_, _16781_, _16780_);
  or _67581_ (_16783_, _16782_, _06262_);
  and _67582_ (_16784_, _14953_, _07942_);
  or _67583_ (_16785_, _16784_, _16771_);
  or _67584_ (_16786_, _16785_, _07151_);
  and _67585_ (_16787_, _07942_, \oc8051_golden_model_1.ACC [3]);
  or _67586_ (_16788_, _16787_, _16771_);
  and _67587_ (_16789_, _16788_, _07141_);
  nor _67588_ (_16790_, _07141_, _10145_);
  or _67589_ (_16791_, _16790_, _06341_);
  or _67590_ (_16792_, _16791_, _16789_);
  and _67591_ (_16793_, _16792_, _06273_);
  and _67592_ (_16794_, _16793_, _16786_);
  and _67593_ (_16795_, _16780_, _06272_);
  or _67594_ (_16796_, _16795_, _06461_);
  or _67595_ (_16797_, _16796_, _16794_);
  nor _67596_ (_16798_, _09498_, _07594_);
  or _67597_ (_16799_, _16798_, _16771_);
  or _67598_ (_16800_, _16799_, _07166_);
  and _67599_ (_16801_, _16800_, _16797_);
  or _67600_ (_16802_, _16801_, _06464_);
  or _67601_ (_16803_, _16788_, _06465_);
  and _67602_ (_16804_, _16803_, _06269_);
  and _67603_ (_16805_, _16804_, _16802_);
  and _67604_ (_16806_, _14948_, _08634_);
  or _67605_ (_16807_, _16806_, _16778_);
  and _67606_ (_16808_, _16807_, _06268_);
  or _67607_ (_16809_, _16808_, _06261_);
  or _67608_ (_16810_, _16809_, _16805_);
  and _67609_ (_16811_, _16810_, _16783_);
  or _67610_ (_16812_, _16811_, _09531_);
  nor _67611_ (_16813_, _10060_, _09894_);
  nor _67612_ (_16814_, _16813_, _10061_);
  or _67613_ (_16815_, _16814_, _09537_);
  and _67614_ (_16816_, _16815_, _06258_);
  and _67615_ (_16817_, _16816_, _16812_);
  or _67616_ (_16818_, _16778_, _14992_);
  and _67617_ (_16819_, _16818_, _06257_);
  and _67618_ (_16820_, _16819_, _16780_);
  or _67619_ (_16821_, _16820_, _10080_);
  or _67620_ (_16822_, _16821_, _16817_);
  or _67621_ (_16823_, _16799_, _07215_);
  and _67622_ (_16824_, _16823_, _16822_);
  or _67623_ (_16825_, _16824_, _07460_);
  and _67624_ (_16826_, _09449_, _07942_);
  or _67625_ (_16827_, _16771_, _07208_);
  or _67626_ (_16828_, _16827_, _16826_);
  and _67627_ (_16829_, _16828_, _05982_);
  and _67628_ (_16830_, _16829_, _16825_);
  or _67629_ (_16831_, _16830_, _16777_);
  and _67630_ (_16832_, _16831_, _10100_);
  nor _67631_ (_16833_, _16719_, _10398_);
  nor _67632_ (_16834_, _16833_, _10391_);
  and _67633_ (_16835_, _16833_, _10391_);
  or _67634_ (_16836_, _16835_, _16834_);
  or _67635_ (_16837_, _16836_, _10439_);
  or _67636_ (_16838_, _16715_, _10388_);
  and _67637_ (_16839_, _16838_, _10093_);
  and _67638_ (_16840_, _16839_, _16837_);
  or _67639_ (_16841_, _16840_, _06218_);
  or _67640_ (_16842_, _16841_, _16832_);
  and _67641_ (_16843_, _16842_, _16774_);
  or _67642_ (_16844_, _16843_, _06369_);
  and _67643_ (_16845_, _14943_, _07942_);
  or _67644_ (_16846_, _16845_, _16771_);
  or _67645_ (_16847_, _16846_, _07237_);
  and _67646_ (_16848_, _16847_, _07240_);
  and _67647_ (_16849_, _16848_, _16844_);
  and _67648_ (_16850_, _12577_, _07942_);
  or _67649_ (_16851_, _16850_, _16771_);
  and _67650_ (_16852_, _16851_, _06536_);
  or _67651_ (_16853_, _16852_, _16849_);
  and _67652_ (_16854_, _16853_, _07242_);
  or _67653_ (_16855_, _16771_, _08292_);
  and _67654_ (_16856_, _16773_, _06375_);
  and _67655_ (_16857_, _16856_, _16855_);
  or _67656_ (_16858_, _16857_, _16854_);
  and _67657_ (_16859_, _16858_, _07234_);
  and _67658_ (_16860_, _16788_, _06545_);
  and _67659_ (_16861_, _16860_, _16855_);
  or _67660_ (_16862_, _16861_, _06366_);
  or _67661_ (_16863_, _16862_, _16859_);
  and _67662_ (_16864_, _14940_, _07942_);
  or _67663_ (_16865_, _16771_, _09056_);
  or _67664_ (_16866_, _16865_, _16864_);
  and _67665_ (_16867_, _16866_, _09061_);
  and _67666_ (_16868_, _16867_, _16863_);
  nor _67667_ (_16869_, _11256_, _09498_);
  or _67668_ (_16870_, _16869_, _16771_);
  and _67669_ (_16871_, _16870_, _06528_);
  or _67670_ (_16872_, _16871_, _06568_);
  or _67671_ (_16873_, _16872_, _16868_);
  or _67672_ (_16874_, _16785_, _06926_);
  and _67673_ (_16875_, _16874_, _05928_);
  and _67674_ (_16876_, _16875_, _16873_);
  and _67675_ (_16877_, _16807_, _05927_);
  or _67676_ (_16878_, _16877_, _06278_);
  or _67677_ (_16879_, _16878_, _16876_);
  and _67678_ (_16880_, _15128_, _07942_);
  or _67679_ (_16881_, _16771_, _06279_);
  or _67680_ (_16882_, _16881_, _16880_);
  and _67681_ (_16883_, _16882_, _01347_);
  and _67682_ (_16884_, _16883_, _16879_);
  or _67683_ (_16885_, _16884_, _16770_);
  and _67684_ (_43156_, _16885_, _42618_);
  nor _67685_ (_16886_, _01347_, _10241_);
  nor _67686_ (_16887_, _07942_, _10241_);
  and _67687_ (_16888_, _08959_, _07942_);
  or _67688_ (_16889_, _16888_, _16887_);
  or _67689_ (_16890_, _16889_, _06219_);
  and _67690_ (_16891_, _15254_, _07942_);
  or _67691_ (_16892_, _16891_, _16887_);
  and _67692_ (_16893_, _16892_, _10094_);
  nor _67693_ (_16894_, _08541_, _09498_);
  or _67694_ (_16895_, _16894_, _16887_);
  or _67695_ (_16896_, _16895_, _07215_);
  nor _67696_ (_16897_, _08634_, _10241_);
  and _67697_ (_16898_, _15176_, _08634_);
  or _67698_ (_16899_, _16898_, _16897_);
  and _67699_ (_16900_, _16899_, _06268_);
  and _67700_ (_16901_, _15162_, _07942_);
  or _67701_ (_16902_, _16901_, _16887_);
  or _67702_ (_16903_, _16902_, _07151_);
  and _67703_ (_16904_, _07942_, \oc8051_golden_model_1.ACC [4]);
  or _67704_ (_16905_, _16904_, _16887_);
  and _67705_ (_16906_, _16905_, _07141_);
  nor _67706_ (_16907_, _07141_, _10241_);
  or _67707_ (_16908_, _16907_, _06341_);
  or _67708_ (_16909_, _16908_, _16906_);
  and _67709_ (_16910_, _16909_, _06273_);
  and _67710_ (_16911_, _16910_, _16903_);
  and _67711_ (_16912_, _15166_, _08634_);
  or _67712_ (_16913_, _16912_, _16897_);
  and _67713_ (_16914_, _16913_, _06272_);
  or _67714_ (_16915_, _16914_, _06461_);
  or _67715_ (_16916_, _16915_, _16911_);
  or _67716_ (_16917_, _16895_, _07166_);
  and _67717_ (_16918_, _16917_, _16916_);
  or _67718_ (_16919_, _16918_, _06464_);
  or _67719_ (_16920_, _16905_, _06465_);
  and _67720_ (_16921_, _16920_, _06269_);
  and _67721_ (_16922_, _16921_, _16919_);
  or _67722_ (_16923_, _16922_, _16900_);
  and _67723_ (_16924_, _16923_, _06262_);
  or _67724_ (_16925_, _16897_, _15183_);
  and _67725_ (_16926_, _16925_, _06261_);
  and _67726_ (_16927_, _16926_, _16913_);
  or _67727_ (_16928_, _16927_, _09531_);
  or _67728_ (_16929_, _16928_, _16924_);
  or _67729_ (_16930_, _10064_, _10062_);
  and _67730_ (_16931_, _16930_, _10065_);
  or _67731_ (_16932_, _16931_, _09537_);
  and _67732_ (_16933_, _16932_, _06258_);
  and _67733_ (_16934_, _16933_, _16929_);
  and _67734_ (_16935_, _15200_, _08634_);
  or _67735_ (_16936_, _16935_, _16897_);
  and _67736_ (_16937_, _16936_, _06257_);
  or _67737_ (_16938_, _16937_, _10080_);
  or _67738_ (_16939_, _16938_, _16934_);
  and _67739_ (_16940_, _16939_, _16896_);
  or _67740_ (_16941_, _16940_, _07460_);
  and _67741_ (_16942_, _09448_, _07942_);
  or _67742_ (_16943_, _16887_, _07208_);
  or _67743_ (_16944_, _16943_, _16942_);
  and _67744_ (_16945_, _16944_, _05982_);
  and _67745_ (_16946_, _16945_, _16941_);
  or _67746_ (_16947_, _16946_, _16893_);
  and _67747_ (_16948_, _16947_, _10100_);
  or _67748_ (_16949_, _16715_, _10380_);
  nor _67749_ (_16950_, _16833_, _10390_);
  or _67750_ (_16951_, _16950_, _10389_);
  nand _67751_ (_16952_, _16951_, _10426_);
  or _67752_ (_16953_, _16951_, _10426_);
  and _67753_ (_16954_, _16953_, _16952_);
  or _67754_ (_16955_, _16954_, _10439_);
  and _67755_ (_16956_, _16955_, _10093_);
  and _67756_ (_16957_, _16956_, _16949_);
  or _67757_ (_16958_, _16957_, _06218_);
  or _67758_ (_16959_, _16958_, _16948_);
  and _67759_ (_16960_, _16959_, _16890_);
  or _67760_ (_16961_, _16960_, _06369_);
  and _67761_ (_16962_, _15269_, _07942_);
  or _67762_ (_16963_, _16962_, _16887_);
  or _67763_ (_16964_, _16963_, _07237_);
  and _67764_ (_16965_, _16964_, _07240_);
  and _67765_ (_16966_, _16965_, _16961_);
  and _67766_ (_16967_, _11254_, _07942_);
  or _67767_ (_16968_, _16967_, _16887_);
  and _67768_ (_16969_, _16968_, _06536_);
  or _67769_ (_16970_, _16969_, _16966_);
  and _67770_ (_16971_, _16970_, _07242_);
  or _67771_ (_16972_, _16887_, _08544_);
  and _67772_ (_16973_, _16889_, _06375_);
  and _67773_ (_16974_, _16973_, _16972_);
  or _67774_ (_16975_, _16974_, _16971_);
  and _67775_ (_16976_, _16975_, _07234_);
  and _67776_ (_16977_, _16905_, _06545_);
  and _67777_ (_16978_, _16977_, _16972_);
  or _67778_ (_16979_, _16978_, _06366_);
  or _67779_ (_16980_, _16979_, _16976_);
  and _67780_ (_16981_, _15266_, _07942_);
  or _67781_ (_16982_, _16887_, _09056_);
  or _67782_ (_16983_, _16982_, _16981_);
  and _67783_ (_16984_, _16983_, _09061_);
  and _67784_ (_16985_, _16984_, _16980_);
  nor _67785_ (_16986_, _11253_, _09498_);
  or _67786_ (_16987_, _16986_, _16887_);
  and _67787_ (_16988_, _16987_, _06528_);
  or _67788_ (_16989_, _16988_, _06568_);
  or _67789_ (_16990_, _16989_, _16985_);
  or _67790_ (_16991_, _16902_, _06926_);
  and _67791_ (_16992_, _16991_, _05928_);
  and _67792_ (_16993_, _16992_, _16990_);
  and _67793_ (_16994_, _16899_, _05927_);
  or _67794_ (_16995_, _16994_, _06278_);
  or _67795_ (_16996_, _16995_, _16993_);
  and _67796_ (_16997_, _15329_, _07942_);
  or _67797_ (_16998_, _16887_, _06279_);
  or _67798_ (_16999_, _16998_, _16997_);
  and _67799_ (_17000_, _16999_, _01347_);
  and _67800_ (_17001_, _17000_, _16996_);
  or _67801_ (_17002_, _17001_, _16886_);
  and _67802_ (_43157_, _17002_, _42618_);
  nor _67803_ (_17003_, _01347_, _10229_);
  nor _67804_ (_17004_, _07942_, _10229_);
  and _67805_ (_17005_, _15459_, _07942_);
  or _67806_ (_17006_, _17005_, _17004_);
  and _67807_ (_17007_, _17006_, _10094_);
  nor _67808_ (_17008_, _08244_, _09498_);
  or _67809_ (_17009_, _17008_, _17004_);
  or _67810_ (_17010_, _17009_, _07215_);
  nor _67811_ (_17011_, _08634_, _10229_);
  and _67812_ (_17012_, _15355_, _08634_);
  or _67813_ (_17013_, _17012_, _17011_);
  and _67814_ (_17014_, _17013_, _06268_);
  and _67815_ (_17015_, _15358_, _07942_);
  or _67816_ (_17016_, _17015_, _17004_);
  or _67817_ (_17017_, _17016_, _07151_);
  and _67818_ (_17018_, _07942_, \oc8051_golden_model_1.ACC [5]);
  or _67819_ (_17019_, _17018_, _17004_);
  and _67820_ (_17020_, _17019_, _07141_);
  nor _67821_ (_17021_, _07141_, _10229_);
  or _67822_ (_17022_, _17021_, _06341_);
  or _67823_ (_17023_, _17022_, _17020_);
  and _67824_ (_17024_, _17023_, _06273_);
  and _67825_ (_17025_, _17024_, _17017_);
  and _67826_ (_17026_, _15372_, _08634_);
  or _67827_ (_17027_, _17026_, _17011_);
  and _67828_ (_17028_, _17027_, _06272_);
  or _67829_ (_17029_, _17028_, _06461_);
  or _67830_ (_17030_, _17029_, _17025_);
  or _67831_ (_17031_, _17009_, _07166_);
  and _67832_ (_17032_, _17031_, _17030_);
  or _67833_ (_17033_, _17032_, _06464_);
  or _67834_ (_17034_, _17019_, _06465_);
  and _67835_ (_17035_, _17034_, _06269_);
  and _67836_ (_17036_, _17035_, _17033_);
  or _67837_ (_17037_, _17036_, _17014_);
  and _67838_ (_17038_, _17037_, _06262_);
  or _67839_ (_17039_, _17011_, _15387_);
  and _67840_ (_17040_, _17039_, _06261_);
  and _67841_ (_17041_, _17040_, _17027_);
  or _67842_ (_17042_, _17041_, _09531_);
  or _67843_ (_17043_, _17042_, _17038_);
  nor _67844_ (_17044_, _10067_, _09757_);
  nor _67845_ (_17045_, _17044_, _10068_);
  or _67846_ (_17046_, _17045_, _09537_);
  and _67847_ (_17047_, _17046_, _06258_);
  and _67848_ (_17048_, _17047_, _17043_);
  or _67849_ (_17049_, _17011_, _15403_);
  and _67850_ (_17050_, _17049_, _06257_);
  and _67851_ (_17051_, _17050_, _17027_);
  or _67852_ (_17052_, _17051_, _10080_);
  or _67853_ (_17053_, _17052_, _17048_);
  and _67854_ (_17054_, _17053_, _17010_);
  or _67855_ (_17055_, _17054_, _07460_);
  and _67856_ (_17056_, _09447_, _07942_);
  or _67857_ (_17057_, _17004_, _07208_);
  or _67858_ (_17058_, _17057_, _17056_);
  and _67859_ (_17059_, _17058_, _05982_);
  and _67860_ (_17060_, _17059_, _17055_);
  or _67861_ (_17061_, _17060_, _17007_);
  and _67862_ (_17062_, _17061_, _10100_);
  or _67863_ (_17063_, _16715_, _10372_);
  not _67864_ (_17064_, _10417_);
  and _67865_ (_17065_, _16952_, _17064_);
  nor _67866_ (_17066_, _17065_, _10427_);
  and _67867_ (_17067_, _17065_, _10427_);
  or _67868_ (_17068_, _17067_, _17066_);
  or _67869_ (_17069_, _17068_, _10439_);
  and _67870_ (_17070_, _17069_, _10093_);
  and _67871_ (_17071_, _17070_, _17063_);
  or _67872_ (_17072_, _17071_, _06218_);
  or _67873_ (_17073_, _17072_, _17062_);
  and _67874_ (_17074_, _08946_, _07942_);
  or _67875_ (_17075_, _17074_, _17004_);
  or _67876_ (_17076_, _17075_, _06219_);
  and _67877_ (_17077_, _17076_, _17073_);
  or _67878_ (_17078_, _17077_, _06369_);
  and _67879_ (_17079_, _15353_, _07942_);
  or _67880_ (_17080_, _17079_, _17004_);
  or _67881_ (_17081_, _17080_, _07237_);
  and _67882_ (_17082_, _17081_, _07240_);
  and _67883_ (_17083_, _17082_, _17078_);
  and _67884_ (_17084_, _11250_, _07942_);
  or _67885_ (_17085_, _17084_, _17004_);
  and _67886_ (_17086_, _17085_, _06536_);
  or _67887_ (_17087_, _17086_, _17083_);
  and _67888_ (_17088_, _17087_, _07242_);
  or _67889_ (_17089_, _17004_, _08247_);
  and _67890_ (_17090_, _17075_, _06375_);
  and _67891_ (_17091_, _17090_, _17089_);
  or _67892_ (_17092_, _17091_, _17088_);
  and _67893_ (_17093_, _17092_, _07234_);
  and _67894_ (_17094_, _17019_, _06545_);
  and _67895_ (_17095_, _17094_, _17089_);
  or _67896_ (_17096_, _17095_, _06366_);
  or _67897_ (_17097_, _17096_, _17093_);
  and _67898_ (_17098_, _15350_, _07942_);
  or _67899_ (_17099_, _17004_, _09056_);
  or _67900_ (_17100_, _17099_, _17098_);
  and _67901_ (_17101_, _17100_, _09061_);
  and _67902_ (_17102_, _17101_, _17097_);
  nor _67903_ (_17103_, _11249_, _09498_);
  or _67904_ (_17104_, _17103_, _17004_);
  and _67905_ (_17105_, _17104_, _06528_);
  or _67906_ (_17106_, _17105_, _06568_);
  or _67907_ (_17107_, _17106_, _17102_);
  or _67908_ (_17108_, _17016_, _06926_);
  and _67909_ (_17109_, _17108_, _05928_);
  and _67910_ (_17110_, _17109_, _17107_);
  and _67911_ (_17111_, _17013_, _05927_);
  or _67912_ (_17112_, _17111_, _06278_);
  or _67913_ (_17113_, _17112_, _17110_);
  and _67914_ (_17114_, _15532_, _07942_);
  or _67915_ (_17115_, _17004_, _06279_);
  or _67916_ (_17116_, _17115_, _17114_);
  and _67917_ (_17117_, _17116_, _01347_);
  and _67918_ (_17118_, _17117_, _17113_);
  or _67919_ (_17119_, _17118_, _17003_);
  and _67920_ (_43159_, _17119_, _42618_);
  nor _67921_ (_17120_, _01347_, _10357_);
  nor _67922_ (_17121_, _07942_, _10357_);
  and _67923_ (_17122_, _15664_, _07942_);
  or _67924_ (_17123_, _17122_, _17121_);
  or _67925_ (_17124_, _17123_, _06219_);
  and _67926_ (_17125_, _15657_, _07942_);
  or _67927_ (_17126_, _17125_, _17121_);
  and _67928_ (_17127_, _17126_, _10094_);
  nor _67929_ (_17128_, _08142_, _09498_);
  or _67930_ (_17129_, _17128_, _17121_);
  or _67931_ (_17130_, _17129_, _07215_);
  nor _67932_ (_17131_, _08634_, _10357_);
  and _67933_ (_17132_, _15551_, _08634_);
  or _67934_ (_17133_, _17132_, _17131_);
  and _67935_ (_17134_, _17133_, _06268_);
  and _67936_ (_17135_, _15554_, _07942_);
  or _67937_ (_17136_, _17135_, _17121_);
  or _67938_ (_17137_, _17136_, _07151_);
  and _67939_ (_17138_, _07942_, \oc8051_golden_model_1.ACC [6]);
  or _67940_ (_17139_, _17138_, _17121_);
  and _67941_ (_17140_, _17139_, _07141_);
  nor _67942_ (_17141_, _07141_, _10357_);
  or _67943_ (_17142_, _17141_, _06341_);
  or _67944_ (_17143_, _17142_, _17140_);
  and _67945_ (_17144_, _17143_, _06273_);
  and _67946_ (_17145_, _17144_, _17137_);
  and _67947_ (_17146_, _15570_, _08634_);
  or _67948_ (_17147_, _17146_, _17131_);
  and _67949_ (_17148_, _17147_, _06272_);
  or _67950_ (_17149_, _17148_, _06461_);
  or _67951_ (_17150_, _17149_, _17145_);
  or _67952_ (_17151_, _17129_, _07166_);
  and _67953_ (_17152_, _17151_, _17150_);
  or _67954_ (_17153_, _17152_, _06464_);
  or _67955_ (_17154_, _17139_, _06465_);
  and _67956_ (_17155_, _17154_, _06269_);
  and _67957_ (_17156_, _17155_, _17153_);
  or _67958_ (_17157_, _17156_, _17134_);
  and _67959_ (_17158_, _17157_, _06262_);
  or _67960_ (_17159_, _17131_, _15585_);
  and _67961_ (_17160_, _17159_, _06261_);
  and _67962_ (_17161_, _17160_, _17147_);
  or _67963_ (_17162_, _17161_, _09531_);
  or _67964_ (_17163_, _17162_, _17158_);
  nor _67965_ (_17164_, _10073_, _10069_);
  nor _67966_ (_17165_, _17164_, _10074_);
  or _67967_ (_17166_, _17165_, _09537_);
  and _67968_ (_17167_, _17166_, _06258_);
  and _67969_ (_17168_, _17167_, _17163_);
  and _67970_ (_17169_, _15602_, _08634_);
  or _67971_ (_17170_, _17169_, _17131_);
  and _67972_ (_17171_, _17170_, _06257_);
  or _67973_ (_17172_, _17171_, _10080_);
  or _67974_ (_17173_, _17172_, _17168_);
  and _67975_ (_17174_, _17173_, _17130_);
  or _67976_ (_17175_, _17174_, _07460_);
  and _67977_ (_17176_, _09446_, _07942_);
  or _67978_ (_17177_, _17121_, _07208_);
  or _67979_ (_17178_, _17177_, _17176_);
  and _67980_ (_17179_, _17178_, _05982_);
  and _67981_ (_17180_, _17179_, _17175_);
  or _67982_ (_17181_, _17180_, _17127_);
  and _67983_ (_17182_, _17181_, _10100_);
  nor _67984_ (_17183_, _17065_, _10373_);
  or _67985_ (_17184_, _17183_, _10374_);
  or _67986_ (_17185_, _17184_, _10429_);
  nand _67987_ (_17186_, _17184_, _10429_);
  and _67988_ (_17187_, _17186_, _17185_);
  or _67989_ (_17188_, _17187_, _10439_);
  nor _67990_ (_17189_, _10439_, _10100_);
  and _67991_ (_17190_, _10363_, _10093_);
  or _67992_ (_17191_, _17190_, _17189_);
  and _67993_ (_17192_, _17191_, _17188_);
  or _67994_ (_17193_, _17192_, _06218_);
  or _67995_ (_17194_, _17193_, _17182_);
  and _67996_ (_17195_, _17194_, _17124_);
  or _67997_ (_17196_, _17195_, _06369_);
  and _67998_ (_17197_, _15549_, _07942_);
  or _67999_ (_17198_, _17197_, _17121_);
  or _68000_ (_17199_, _17198_, _07237_);
  and _68001_ (_17200_, _17199_, _07240_);
  and _68002_ (_17201_, _17200_, _17196_);
  and _68003_ (_17202_, _11247_, _07942_);
  or _68004_ (_17203_, _17202_, _17121_);
  and _68005_ (_17204_, _17203_, _06536_);
  or _68006_ (_17205_, _17204_, _17201_);
  and _68007_ (_17206_, _17205_, _07242_);
  or _68008_ (_17207_, _17121_, _08145_);
  and _68009_ (_17208_, _17123_, _06375_);
  and _68010_ (_17209_, _17208_, _17207_);
  or _68011_ (_17210_, _17209_, _17206_);
  and _68012_ (_17211_, _17210_, _07234_);
  and _68013_ (_17212_, _17139_, _06545_);
  and _68014_ (_17213_, _17212_, _17207_);
  or _68015_ (_17214_, _17213_, _06366_);
  or _68016_ (_17215_, _17214_, _17211_);
  and _68017_ (_17216_, _15546_, _07942_);
  or _68018_ (_17217_, _17121_, _09056_);
  or _68019_ (_17218_, _17217_, _17216_);
  and _68020_ (_17219_, _17218_, _09061_);
  and _68021_ (_17220_, _17219_, _17215_);
  nor _68022_ (_17221_, _11246_, _09498_);
  or _68023_ (_17222_, _17221_, _17121_);
  and _68024_ (_17223_, _17222_, _06528_);
  or _68025_ (_17224_, _17223_, _06568_);
  or _68026_ (_17225_, _17224_, _17220_);
  or _68027_ (_17226_, _17136_, _06926_);
  and _68028_ (_17227_, _17226_, _05928_);
  and _68029_ (_17228_, _17227_, _17225_);
  and _68030_ (_17229_, _17133_, _05927_);
  or _68031_ (_17230_, _17229_, _06278_);
  or _68032_ (_17231_, _17230_, _17228_);
  and _68033_ (_17232_, _15734_, _07942_);
  or _68034_ (_17233_, _17121_, _06279_);
  or _68035_ (_17234_, _17233_, _17232_);
  and _68036_ (_17235_, _17234_, _01347_);
  and _68037_ (_17236_, _17235_, _17231_);
  or _68038_ (_17237_, _17236_, _17120_);
  and _68039_ (_43160_, _17237_, _42618_);
  nor _68040_ (_17238_, _01347_, _06097_);
  nand _68041_ (_17239_, _11284_, _08572_);
  nand _68042_ (_17240_, _12581_, _06283_);
  and _68043_ (_17241_, _17240_, _11321_);
  nor _68044_ (_17242_, _07133_, \oc8051_golden_model_1.ACC [0]);
  nor _68045_ (_17243_, _17242_, _11179_);
  and _68046_ (_17244_, _11154_, _17243_);
  and _68047_ (_17245_, _11156_, _17243_);
  nor _68048_ (_17246_, _10634_, _06097_);
  or _68049_ (_17247_, _17246_, _10635_);
  or _68050_ (_17248_, _11069_, _17247_);
  nand _68051_ (_17249_, _11021_, _12596_);
  nand _68052_ (_17250_, _12581_, _06533_);
  and _68053_ (_17251_, _17250_, _10955_);
  nand _68054_ (_17252_, _06251_, _05974_);
  nor _68055_ (_17253_, _07939_, _06097_);
  and _68056_ (_17254_, _14467_, _07939_);
  or _68057_ (_17255_, _17254_, _17253_);
  and _68058_ (_17256_, _17255_, _10094_);
  and _68059_ (_17257_, _07939_, _07133_);
  or _68060_ (_17258_, _17257_, _17253_);
  or _68061_ (_17259_, _17258_, _07215_);
  or _68062_ (_17260_, _17247_, _10588_);
  or _68063_ (_17261_, _10743_, _07133_);
  or _68064_ (_17262_, _10755_, _07133_);
  nor _68065_ (_17263_, _06781_, _06097_);
  and _68066_ (_17264_, _06781_, _06097_);
  nor _68067_ (_17265_, _17264_, _17263_);
  nand _68068_ (_17266_, _17265_, _10755_);
  and _68069_ (_17267_, _17266_, _10759_);
  and _68070_ (_17268_, _17267_, _17262_);
  and _68071_ (_17269_, _17268_, _07155_);
  or _68072_ (_17270_, _17269_, _09392_);
  or _68073_ (_17271_, _17268_, _10758_);
  and _68074_ (_17272_, _17271_, _06015_);
  or _68075_ (_17273_, _17272_, _07154_);
  and _68076_ (_17274_, _17273_, _07151_);
  and _68077_ (_17275_, _17274_, _17270_);
  nor _68078_ (_17276_, _08390_, _10490_);
  or _68079_ (_17277_, _17276_, _17253_);
  and _68080_ (_17278_, _17277_, _06341_);
  or _68081_ (_17279_, _17278_, _06272_);
  or _68082_ (_17280_, _17279_, _17275_);
  and _68083_ (_17281_, _14382_, _08636_);
  nor _68084_ (_17282_, _08636_, _06097_);
  or _68085_ (_17283_, _17282_, _06273_);
  or _68086_ (_17284_, _17283_, _17281_);
  and _68087_ (_17285_, _17284_, _07166_);
  and _68088_ (_17286_, _17285_, _17280_);
  and _68089_ (_17287_, _17258_, _06461_);
  or _68090_ (_17288_, _17287_, _10744_);
  or _68091_ (_17289_, _17288_, _17286_);
  and _68092_ (_17290_, _17289_, _17261_);
  or _68093_ (_17291_, _17290_, _07174_);
  or _68094_ (_17292_, _09392_, _07175_);
  and _68095_ (_17293_, _17292_, _06465_);
  and _68096_ (_17294_, _17293_, _17291_);
  and _68097_ (_17295_, _08390_, _06464_);
  or _68098_ (_17296_, _17295_, _10811_);
  or _68099_ (_17297_, _17296_, _17294_);
  nand _68100_ (_17298_, _10811_, _10135_);
  and _68101_ (_17299_, _17298_, _17297_);
  or _68102_ (_17300_, _17299_, _06268_);
  or _68103_ (_17301_, _17253_, _06269_);
  and _68104_ (_17302_, _17301_, _06262_);
  and _68105_ (_17303_, _17302_, _17300_);
  and _68106_ (_17304_, _17277_, _06261_);
  or _68107_ (_17305_, _17304_, _09531_);
  or _68108_ (_17306_, _17305_, _17303_);
  nor _68109_ (_17307_, _07211_, _05977_);
  nor _68110_ (_17308_, _17307_, _14203_);
  not _68111_ (_17309_, _14197_);
  or _68112_ (_17310_, _17309_, _10729_);
  nor _68113_ (_17311_, _17310_, _06705_);
  nand _68114_ (_17312_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nand _68115_ (_17313_, _17312_, _09531_);
  and _68116_ (_17314_, _17313_, _17311_);
  and _68117_ (_17315_, _17314_, _17308_);
  and _68118_ (_17316_, _17315_, _17306_);
  nor _68119_ (_17317_, _10709_, _06097_);
  or _68120_ (_17318_, _17317_, _10710_);
  and _68121_ (_17319_, _10737_, _17318_);
  or _68122_ (_17320_, _17319_, _10656_);
  or _68123_ (_17321_, _17320_, _17316_);
  and _68124_ (_17322_, _17321_, _17260_);
  or _68125_ (_17323_, _17322_, _06512_);
  nor _68126_ (_17324_, _10881_, _06097_);
  or _68127_ (_17325_, _17324_, _10882_);
  or _68128_ (_17326_, _17325_, _06517_);
  and _68129_ (_17327_, _17326_, _10517_);
  and _68130_ (_17328_, _17327_, _17323_);
  nor _68131_ (_17329_, _10564_, _06097_);
  or _68132_ (_17330_, _17329_, _10565_);
  and _68133_ (_17331_, _17330_, _10516_);
  or _68134_ (_17332_, _17331_, _10515_);
  or _68135_ (_17333_, _17332_, _17328_);
  nand _68136_ (_17334_, _06251_, _10515_);
  and _68137_ (_17335_, _17334_, _06258_);
  and _68138_ (_17336_, _17335_, _17333_);
  and _68139_ (_17337_, _14413_, _08636_);
  or _68140_ (_17338_, _17337_, _17282_);
  and _68141_ (_17340_, _17338_, _06257_);
  or _68142_ (_17341_, _17340_, _10080_);
  or _68143_ (_17342_, _17341_, _17336_);
  and _68144_ (_17343_, _17342_, _17259_);
  or _68145_ (_17344_, _17343_, _07460_);
  and _68146_ (_17345_, _09392_, _07939_);
  or _68147_ (_17346_, _17253_, _07208_);
  or _68148_ (_17347_, _17346_, _17345_);
  and _68149_ (_17348_, _17347_, _05982_);
  and _68150_ (_17349_, _17348_, _17344_);
  or _68151_ (_17351_, _17349_, _17256_);
  and _68152_ (_17352_, _17351_, _10100_);
  or _68153_ (_17353_, _17189_, _05974_);
  or _68154_ (_17354_, _17353_, _17352_);
  and _68155_ (_17355_, _17354_, _17252_);
  or _68156_ (_17356_, _17355_, _06218_);
  and _68157_ (_17357_, _07939_, _08954_);
  or _68158_ (_17358_, _17357_, _17253_);
  or _68159_ (_17359_, _17358_, _06219_);
  and _68160_ (_17360_, _17359_, _10930_);
  and _68161_ (_17362_, _17360_, _17356_);
  nor _68162_ (_17363_, _10930_, _06251_);
  or _68163_ (_17364_, _17363_, _10937_);
  or _68164_ (_17365_, _17364_, _17362_);
  or _68165_ (_17366_, _10940_, _17243_);
  and _68166_ (_17367_, _10946_, _10508_);
  and _68167_ (_17368_, _17367_, _17366_);
  and _68168_ (_17369_, _17368_, _17365_);
  not _68169_ (_17370_, _17367_);
  and _68170_ (_17371_, _17370_, _17243_);
  or _68171_ (_17373_, _17371_, _10501_);
  or _68172_ (_17374_, _17373_, _17369_);
  not _68173_ (_17375_, _10501_);
  nor _68174_ (_17376_, _09392_, \oc8051_golden_model_1.ACC [0]);
  nor _68175_ (_17377_, _11223_, _17376_);
  or _68176_ (_17378_, _17377_, _17375_);
  and _68177_ (_17379_, _17378_, _06885_);
  and _68178_ (_17380_, _17379_, _17374_);
  and _68179_ (_17381_, _17377_, _06884_);
  or _68180_ (_17382_, _17381_, _06533_);
  or _68181_ (_17384_, _17382_, _17380_);
  and _68182_ (_17385_, _17384_, _17251_);
  and _68183_ (_17386_, _10954_, _12597_);
  or _68184_ (_17387_, _17386_, _06369_);
  or _68185_ (_17388_, _17387_, _17385_);
  and _68186_ (_17389_, _14366_, _07939_);
  or _68187_ (_17390_, _17389_, _17253_);
  or _68188_ (_17391_, _17390_, _07237_);
  and _68189_ (_17392_, _17391_, _17388_);
  or _68190_ (_17393_, _17392_, _06536_);
  or _68191_ (_17395_, _17253_, _07240_);
  and _68192_ (_17396_, _17395_, _10977_);
  and _68193_ (_17397_, _17396_, _17393_);
  or _68194_ (_17398_, _10985_, _11179_);
  and _68195_ (_17399_, _17398_, _10987_);
  or _68196_ (_17400_, _17399_, _17397_);
  not _68197_ (_17401_, _10983_);
  not _68198_ (_17402_, _10985_);
  or _68199_ (_17403_, _17402_, _11179_);
  and _68200_ (_17404_, _17403_, _17401_);
  and _68201_ (_17405_, _17404_, _17400_);
  and _68202_ (_17406_, _10983_, _11223_);
  or _68203_ (_17407_, _17406_, _06542_);
  or _68204_ (_17408_, _17407_, _17405_);
  or _68205_ (_17409_, _11263_, _06543_);
  and _68206_ (_17410_, _17409_, _10497_);
  and _68207_ (_17411_, _17410_, _17408_);
  and _68208_ (_17412_, _11302_, _10496_);
  or _68209_ (_17413_, _17412_, _17411_);
  and _68210_ (_17414_, _17413_, _07242_);
  nand _68211_ (_17415_, _17358_, _06375_);
  nor _68212_ (_17416_, _17415_, _17276_);
  or _68213_ (_17417_, _17416_, _06711_);
  or _68214_ (_17418_, _17417_, _17414_);
  nor _68215_ (_17419_, _17242_, _06755_);
  or _68216_ (_17420_, _17419_, _10998_);
  and _68217_ (_17421_, _17420_, _17418_);
  and _68218_ (_17422_, _06350_, _06527_);
  nor _68219_ (_17423_, _17422_, _07040_);
  and _68220_ (_17424_, _17423_, _12156_);
  not _68221_ (_17425_, _17242_);
  nand _68222_ (_17426_, _17425_, _06755_);
  nand _68223_ (_17427_, _17426_, _17424_);
  or _68224_ (_17428_, _17427_, _17421_);
  and _68225_ (_17429_, _06337_, _06527_);
  not _68226_ (_17430_, _17429_);
  or _68227_ (_17431_, _17424_, _17425_);
  and _68228_ (_17432_, _17431_, _17430_);
  and _68229_ (_17433_, _17432_, _17428_);
  nor _68230_ (_17434_, _17242_, _17430_);
  or _68231_ (_17435_, _17434_, _11014_);
  or _68232_ (_17436_, _17435_, _17433_);
  nand _68233_ (_17437_, _11014_, _17376_);
  and _68234_ (_17438_, _17437_, _06531_);
  and _68235_ (_17439_, _17438_, _17436_);
  nand _68236_ (_17440_, _11024_, _12580_);
  and _68237_ (_17441_, _17440_, _11023_);
  or _68238_ (_17442_, _17441_, _17439_);
  and _68239_ (_17443_, _17442_, _17249_);
  or _68240_ (_17444_, _17443_, _06366_);
  and _68241_ (_17445_, _14363_, _07939_);
  or _68242_ (_17446_, _17253_, _09056_);
  or _68243_ (_17447_, _17446_, _17445_);
  and _68244_ (_17448_, _17447_, _11037_);
  and _68245_ (_17449_, _17448_, _17444_);
  and _68246_ (_17450_, _14283_, _17318_);
  or _68247_ (_17451_, _17450_, _11041_);
  or _68248_ (_17452_, _17451_, _17449_);
  and _68249_ (_17453_, _17452_, _17248_);
  or _68250_ (_17454_, _17453_, _06540_);
  or _68251_ (_17455_, _17325_, _06541_);
  and _68252_ (_17456_, _17455_, _11127_);
  and _68253_ (_17457_, _17456_, _17454_);
  and _68254_ (_17458_, _11097_, _17330_);
  or _68255_ (_17459_, _17458_, _11125_);
  or _68256_ (_17460_, _17459_, _17457_);
  and _68257_ (_17461_, _11125_, _10558_);
  or _68258_ (_17462_, _17461_, _07045_);
  nor _68259_ (_17463_, _17462_, _11155_);
  and _68260_ (_17464_, _17463_, _17460_);
  nor _68261_ (_17465_, _17464_, _17245_);
  nor _68262_ (_17466_, _17465_, _11154_);
  or _68263_ (_17467_, _17466_, _17244_);
  and _68264_ (_17468_, _17467_, _11203_);
  and _68265_ (_17469_, _11201_, _17377_);
  or _68266_ (_17470_, _17469_, _06283_);
  or _68267_ (_17471_, _17470_, _17468_);
  and _68268_ (_17472_, _17471_, _17241_);
  and _68269_ (_17473_, _11243_, _12597_);
  or _68270_ (_17474_, _17473_, _11284_);
  or _68271_ (_17475_, _17474_, _17472_);
  and _68272_ (_17476_, _17475_, _17239_);
  or _68273_ (_17477_, _17476_, _06568_);
  or _68274_ (_17478_, _17277_, _06926_);
  and _68275_ (_17479_, _17478_, _11331_);
  and _68276_ (_17480_, _17479_, _17477_);
  nor _68277_ (_17481_, _11335_, _06097_);
  nor _68278_ (_17482_, _17481_, _13037_);
  or _68279_ (_17483_, _17482_, _17480_);
  nand _68280_ (_17484_, _11335_, _06042_);
  and _68281_ (_17485_, _17484_, _05928_);
  and _68282_ (_17486_, _17485_, _17483_);
  and _68283_ (_17487_, _17253_, _05927_);
  or _68284_ (_17488_, _17487_, _06278_);
  or _68285_ (_17489_, _17488_, _17486_);
  or _68286_ (_17490_, _17277_, _06279_);
  and _68287_ (_17491_, _17490_, _11354_);
  and _68288_ (_17492_, _17491_, _17489_);
  nor _68289_ (_17493_, _11360_, _06097_);
  nor _68290_ (_17494_, _17493_, _12141_);
  or _68291_ (_17495_, _17494_, _17492_);
  nand _68292_ (_17496_, _11360_, _06042_);
  and _68293_ (_17497_, _17496_, _01347_);
  and _68294_ (_17498_, _17497_, _17495_);
  or _68295_ (_17499_, _17498_, _17238_);
  and _68296_ (_43161_, _17499_, _42618_);
  nor _68297_ (_17500_, _01347_, _06042_);
  or _68298_ (_17501_, _11106_, _11105_);
  nor _68299_ (_17502_, _11107_, _06541_);
  and _68300_ (_17503_, _17502_, _17501_);
  and _68301_ (_17504_, _06886_, _06364_);
  nor _68302_ (_17505_, _11035_, _17504_);
  not _68303_ (_17506_, _17423_);
  not _68304_ (_17507_, _12157_);
  nand _68305_ (_17508_, _17507_, _11177_);
  or _68306_ (_17509_, _17401_, _11220_);
  not _68307_ (_17510_, _06888_);
  and _68308_ (_17511_, _06350_, _06535_);
  not _68309_ (_17512_, _17511_);
  and _68310_ (_17513_, _17512_, _10508_);
  nor _68311_ (_17514_, _07939_, _06042_);
  nor _68312_ (_17515_, _10490_, _07357_);
  or _68313_ (_17516_, _17515_, _17514_);
  or _68314_ (_17517_, _17516_, _07215_);
  nor _68315_ (_17518_, _08636_, _06042_);
  and _68316_ (_17519_, _14557_, _08636_);
  or _68317_ (_17520_, _17519_, _17518_);
  or _68318_ (_17521_, _17518_, _14556_);
  and _68319_ (_17522_, _17521_, _06261_);
  and _68320_ (_17523_, _17522_, _17520_);
  nand _68321_ (_17524_, _10744_, _07357_);
  nand _68322_ (_17525_, _10756_, _07357_);
  nor _68323_ (_17526_, _06781_, _06042_);
  and _68324_ (_17527_, _06781_, _06042_);
  nor _68325_ (_17528_, _17527_, _17526_);
  nand _68326_ (_17529_, _17528_, _10755_);
  and _68327_ (_17530_, _17529_, _10759_);
  and _68328_ (_17531_, _17530_, _17525_);
  or _68329_ (_17532_, _17531_, _10758_);
  and _68330_ (_17533_, _17532_, _06015_);
  or _68331_ (_17534_, _17533_, _07154_);
  and _68332_ (_17535_, _17531_, _07155_);
  or _68333_ (_17536_, _17535_, _09451_);
  and _68334_ (_17537_, _17536_, _17534_);
  or _68335_ (_17538_, _17537_, _06341_);
  or _68336_ (_17539_, _07939_, \oc8051_golden_model_1.ACC [1]);
  and _68337_ (_17540_, _14562_, _07939_);
  not _68338_ (_17541_, _17540_);
  and _68339_ (_17542_, _17541_, _17539_);
  or _68340_ (_17543_, _17542_, _07151_);
  and _68341_ (_17544_, _17543_, _17538_);
  or _68342_ (_17545_, _17544_, _10775_);
  nor _68343_ (_17546_, _10779_, \oc8051_golden_model_1.PSW [6]);
  nor _68344_ (_17547_, _17546_, \oc8051_golden_model_1.ACC [1]);
  and _68345_ (_17548_, _17546_, \oc8051_golden_model_1.ACC [1]);
  nor _68346_ (_17549_, _17548_, _17547_);
  nand _68347_ (_17550_, _17549_, _10775_);
  and _68348_ (_17551_, _17550_, _06466_);
  and _68349_ (_17552_, _17551_, _17545_);
  and _68350_ (_17553_, _17520_, _06272_);
  and _68351_ (_17554_, _17516_, _06461_);
  or _68352_ (_17555_, _17554_, _10744_);
  or _68353_ (_17556_, _17555_, _17553_);
  or _68354_ (_17557_, _17556_, _17552_);
  and _68355_ (_17558_, _17557_, _17524_);
  or _68356_ (_17559_, _17558_, _07174_);
  or _68357_ (_17560_, _09451_, _07175_);
  and _68358_ (_17561_, _17560_, _06465_);
  and _68359_ (_17562_, _17561_, _17559_);
  nor _68360_ (_17563_, _08340_, _06465_);
  or _68361_ (_17564_, _17563_, _10811_);
  or _68362_ (_17565_, _17564_, _17562_);
  nand _68363_ (_17566_, _10811_, _10170_);
  and _68364_ (_17567_, _17566_, _17565_);
  or _68365_ (_17568_, _17567_, _06268_);
  and _68366_ (_17569_, _14560_, _08636_);
  or _68367_ (_17570_, _17569_, _17518_);
  or _68368_ (_17571_, _17570_, _06269_);
  and _68369_ (_17572_, _17571_, _06262_);
  and _68370_ (_17573_, _17572_, _17568_);
  or _68371_ (_17574_, _17573_, _17523_);
  and _68372_ (_17575_, _17574_, _09537_);
  nor _68373_ (_17576_, _10031_, _10030_);
  nor _68374_ (_17577_, _17576_, _10032_);
  nand _68375_ (_17578_, _17577_, _09531_);
  nand _68376_ (_17579_, _17578_, _10735_);
  or _68377_ (_17580_, _17579_, _17575_);
  nor _68378_ (_17581_, _10657_, _06097_);
  or _68379_ (_17582_, _17581_, _10708_);
  nor _68380_ (_17583_, _17582_, _11178_);
  and _68381_ (_17584_, _17582_, _11178_);
  or _68382_ (_17585_, _17584_, _10735_);
  or _68383_ (_17586_, _17585_, _17583_);
  and _68384_ (_17587_, _17586_, _10588_);
  and _68385_ (_17588_, _17587_, _17580_);
  not _68386_ (_17589_, _11222_);
  nor _68387_ (_17590_, _10589_, _06097_);
  or _68388_ (_17591_, _17590_, _10633_);
  nand _68389_ (_17592_, _17591_, _17589_);
  or _68390_ (_17593_, _17591_, _17589_);
  and _68391_ (_17594_, _17593_, _10656_);
  and _68392_ (_17595_, _17594_, _17592_);
  or _68393_ (_17596_, _17595_, _06512_);
  or _68394_ (_17597_, _17596_, _17588_);
  nor _68395_ (_17598_, _10834_, _06097_);
  or _68396_ (_17599_, _17598_, _10880_);
  nor _68397_ (_17600_, _17599_, _11262_);
  and _68398_ (_17601_, _17599_, _11262_);
  or _68399_ (_17602_, _17601_, _06517_);
  or _68400_ (_17603_, _17602_, _17600_);
  and _68401_ (_17604_, _17603_, _10517_);
  and _68402_ (_17605_, _17604_, _17597_);
  nor _68403_ (_17606_, _06251_, \oc8051_golden_model_1.ACC [0]);
  not _68404_ (_17607_, _17606_);
  and _68405_ (_17608_, _11305_, _17607_);
  nor _68406_ (_17609_, _11305_, _17607_);
  nor _68407_ (_17610_, _17609_, _17608_);
  or _68408_ (_17611_, _12597_, _10558_);
  and _68409_ (_17612_, _17611_, _17610_);
  and _68410_ (_17613_, _12598_, \oc8051_golden_model_1.PSW [7]);
  or _68411_ (_17614_, _17613_, _17612_);
  and _68412_ (_17615_, _17614_, _10516_);
  or _68413_ (_17616_, _17615_, _10515_);
  or _68414_ (_17617_, _17616_, _17605_);
  nand _68415_ (_17618_, _07004_, _10515_);
  and _68416_ (_17619_, _17618_, _06258_);
  and _68417_ (_17620_, _17619_, _17617_);
  or _68418_ (_17621_, _17518_, _14597_);
  and _68419_ (_17622_, _17621_, _06257_);
  and _68420_ (_17623_, _17622_, _17520_);
  or _68421_ (_17624_, _17623_, _10080_);
  or _68422_ (_17625_, _17624_, _17620_);
  and _68423_ (_17626_, _17625_, _17517_);
  or _68424_ (_17627_, _17626_, _07460_);
  and _68425_ (_17628_, _09451_, _07939_);
  or _68426_ (_17629_, _17514_, _07208_);
  or _68427_ (_17630_, _17629_, _17628_);
  and _68428_ (_17631_, _17630_, _05982_);
  and _68429_ (_17632_, _17631_, _17627_);
  or _68430_ (_17633_, _14653_, _10490_);
  and _68431_ (_17634_, _17539_, _10094_);
  and _68432_ (_17635_, _17634_, _17633_);
  or _68433_ (_17636_, _17635_, _10093_);
  or _68434_ (_17637_, _17636_, _17632_);
  nand _68435_ (_17638_, _10350_, _10093_);
  and _68436_ (_17639_, _17638_, _17637_);
  or _68437_ (_17640_, _17639_, _05974_);
  nand _68438_ (_17641_, _07004_, _05974_);
  and _68439_ (_17642_, _17641_, _06219_);
  and _68440_ (_17643_, _17642_, _17640_);
  nand _68441_ (_17644_, _07939_, _07038_);
  and _68442_ (_17645_, _17539_, _06218_);
  and _68443_ (_17646_, _17645_, _17644_);
  or _68444_ (_17647_, _17646_, _10929_);
  or _68445_ (_17648_, _17647_, _17643_);
  nand _68446_ (_17649_, _10929_, _07004_);
  and _68447_ (_17650_, _17649_, _10940_);
  and _68448_ (_17651_, _17650_, _17648_);
  and _68449_ (_17652_, _10937_, _11178_);
  or _68450_ (_17653_, _17652_, _17651_);
  and _68451_ (_17654_, _17653_, _17513_);
  not _68452_ (_17655_, _17513_);
  and _68453_ (_17656_, _17655_, _11178_);
  or _68454_ (_17657_, _17656_, _17654_);
  and _68455_ (_17658_, _17657_, _17510_);
  and _68456_ (_17659_, _11178_, _06888_);
  or _68457_ (_17660_, _17659_, _10948_);
  or _68458_ (_17661_, _17660_, _17658_);
  or _68459_ (_17662_, _11222_, _10502_);
  and _68460_ (_17663_, _17662_, _17661_);
  or _68461_ (_17664_, _17663_, _06533_);
  or _68462_ (_17665_, _11262_, _06534_);
  and _68463_ (_17666_, _17665_, _10955_);
  and _68464_ (_17667_, _17666_, _17664_);
  nor _68465_ (_17668_, _10955_, _11305_);
  or _68466_ (_17669_, _17668_, _17667_);
  and _68467_ (_17670_, _17669_, _07237_);
  or _68468_ (_17671_, _14668_, _10490_);
  and _68469_ (_17672_, _17539_, _06369_);
  and _68470_ (_17673_, _17672_, _17671_);
  or _68471_ (_17674_, _17673_, _06536_);
  or _68472_ (_17675_, _17674_, _17670_);
  or _68473_ (_17676_, _17514_, _07240_);
  and _68474_ (_17677_, _17676_, _10986_);
  and _68475_ (_17678_, _17677_, _17675_);
  and _68476_ (_17679_, _10987_, _11176_);
  or _68477_ (_17680_, _17679_, _10983_);
  or _68478_ (_17681_, _17680_, _17678_);
  and _68479_ (_17682_, _17681_, _17509_);
  or _68480_ (_17683_, _17682_, _06542_);
  or _68481_ (_17684_, _11260_, _06543_);
  and _68482_ (_17685_, _17684_, _10497_);
  and _68483_ (_17686_, _17685_, _17683_);
  and _68484_ (_17687_, _11301_, _10496_);
  or _68485_ (_17688_, _17687_, _17686_);
  and _68486_ (_17689_, _17688_, _07242_);
  or _68487_ (_17690_, _14666_, _10490_);
  and _68488_ (_17691_, _17539_, _06375_);
  and _68489_ (_17692_, _17691_, _17690_);
  or _68490_ (_17693_, _17692_, _17507_);
  or _68491_ (_17694_, _17693_, _17689_);
  and _68492_ (_17695_, _17694_, _17508_);
  or _68493_ (_17696_, _17695_, _17506_);
  nand _68494_ (_17697_, _17506_, _11177_);
  and _68495_ (_17698_, _17697_, _17430_);
  and _68496_ (_17699_, _17698_, _17696_);
  nor _68497_ (_17700_, _11177_, _17430_);
  or _68498_ (_17701_, _17700_, _11014_);
  or _68499_ (_17702_, _17701_, _17699_);
  nand _68500_ (_17703_, _11014_, _11221_);
  and _68501_ (_17704_, _17703_, _06531_);
  and _68502_ (_17705_, _17704_, _17702_);
  nand _68503_ (_17706_, _11024_, _11261_);
  and _68504_ (_17707_, _17706_, _11023_);
  or _68505_ (_17708_, _17707_, _17705_);
  and _68506_ (_17709_, _11021_, _06042_);
  nand _68507_ (_17710_, _17709_, _07004_);
  and _68508_ (_17711_, _17710_, _09056_);
  and _68509_ (_17712_, _17711_, _17708_);
  or _68510_ (_17713_, _17644_, _08341_);
  and _68511_ (_17714_, _17539_, _06366_);
  and _68512_ (_17715_, _17714_, _17713_);
  or _68513_ (_17716_, _17715_, _17712_);
  and _68514_ (_17717_, _17716_, _17505_);
  nor _68515_ (_17718_, _11050_, _11049_);
  nor _68516_ (_17719_, _17718_, _11051_);
  and _68517_ (_17720_, _17719_, _14283_);
  or _68518_ (_17721_, _17720_, _17717_);
  not _68519_ (_17722_, _11040_);
  and _68520_ (_17723_, _07209_, _06364_);
  not _68521_ (_17724_, _17723_);
  or _68522_ (_17725_, _17719_, _17724_);
  and _68523_ (_17726_, _17725_, _17722_);
  and _68524_ (_17727_, _17726_, _17721_);
  nor _68525_ (_17728_, _11078_, _11077_);
  nor _68526_ (_17729_, _17728_, _11079_);
  and _68527_ (_17730_, _17729_, _11040_);
  or _68528_ (_17731_, _17730_, _11039_);
  or _68529_ (_17732_, _17731_, _17727_);
  not _68530_ (_17733_, _11039_);
  or _68531_ (_17734_, _17729_, _17733_);
  and _68532_ (_17735_, _17734_, _06541_);
  and _68533_ (_17736_, _17735_, _17732_);
  or _68534_ (_17737_, _17736_, _17503_);
  and _68535_ (_17738_, _17737_, _11127_);
  or _68536_ (_17739_, _11134_, _10568_);
  nor _68537_ (_17740_, _11135_, _11127_);
  and _68538_ (_17741_, _17740_, _17739_);
  or _68539_ (_17742_, _17741_, _11125_);
  or _68540_ (_17743_, _17742_, _17738_);
  nand _68541_ (_17744_, _11125_, _06097_);
  and _68542_ (_17745_, _17744_, _11157_);
  and _68543_ (_17746_, _17745_, _17743_);
  or _68544_ (_17747_, _11179_, _11178_);
  nor _68545_ (_17748_, _11180_, _11157_);
  and _68546_ (_17749_, _17748_, _17747_);
  or _68547_ (_17750_, _17749_, _11201_);
  or _68548_ (_17751_, _17750_, _17746_);
  nor _68549_ (_17752_, _11223_, _11222_);
  nor _68550_ (_17753_, _17752_, _11224_);
  or _68551_ (_17754_, _17753_, _11203_);
  and _68552_ (_17755_, _17754_, _06285_);
  and _68553_ (_17756_, _17755_, _17751_);
  nor _68554_ (_17757_, _11263_, _11262_);
  nor _68555_ (_17758_, _17757_, _11264_);
  and _68556_ (_17759_, _17758_, _06283_);
  or _68557_ (_17760_, _17759_, _11243_);
  or _68558_ (_17761_, _17760_, _17756_);
  nor _68559_ (_17762_, _11306_, _11302_);
  nor _68560_ (_17763_, _17762_, _11307_);
  or _68561_ (_17764_, _17763_, _11321_);
  and _68562_ (_17765_, _17764_, _11285_);
  and _68563_ (_17766_, _17765_, _17761_);
  and _68564_ (_17767_, _11284_, \oc8051_golden_model_1.ACC [0]);
  or _68565_ (_17768_, _17767_, _06568_);
  or _68566_ (_17769_, _17768_, _17766_);
  or _68567_ (_17770_, _17542_, _06926_);
  and _68568_ (_17771_, _17770_, _11331_);
  and _68569_ (_17772_, _17771_, _17769_);
  nor _68570_ (_17773_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor _68571_ (_17774_, _11361_, _17773_);
  nor _68572_ (_17775_, _17774_, _11331_);
  or _68573_ (_17776_, _17775_, _11335_);
  or _68574_ (_17777_, _17776_, _17772_);
  nand _68575_ (_17778_, _11335_, _10213_);
  and _68576_ (_17779_, _17778_, _05928_);
  and _68577_ (_17780_, _17779_, _17777_);
  and _68578_ (_17781_, _17570_, _05927_);
  or _68579_ (_17782_, _17781_, _06278_);
  or _68580_ (_17783_, _17782_, _17780_);
  or _68581_ (_17784_, _17540_, _17514_);
  or _68582_ (_17785_, _17784_, _06279_);
  and _68583_ (_17786_, _17785_, _11354_);
  and _68584_ (_17787_, _17786_, _17783_);
  and _68585_ (_17788_, _17774_, _11353_);
  or _68586_ (_17789_, _17788_, _11360_);
  or _68587_ (_17790_, _17789_, _17787_);
  nand _68588_ (_17791_, _11360_, _10213_);
  and _68589_ (_17792_, _17791_, _01347_);
  and _68590_ (_17793_, _17792_, _17790_);
  or _68591_ (_17794_, _17793_, _17500_);
  and _68592_ (_43163_, _17794_, _42618_);
  nor _68593_ (_17795_, _01347_, _10213_);
  nand _68594_ (_17796_, _11284_, _06042_);
  or _68595_ (_17797_, _11266_, _11259_);
  nor _68596_ (_17798_, _11267_, _06285_);
  and _68597_ (_17799_, _17798_, _17797_);
  not _68598_ (_17800_, _11200_);
  nor _68599_ (_17801_, _11226_, _11219_);
  nor _68600_ (_17802_, _17801_, _11227_);
  or _68601_ (_17803_, _17802_, _17800_);
  and _68602_ (_17804_, _11136_, _10556_);
  nor _68603_ (_17805_, _17804_, _11137_);
  or _68604_ (_17806_, _17805_, _11127_);
  nand _68605_ (_17807_, _11014_, _11218_);
  or _68606_ (_17808_, _11219_, _10502_);
  nand _68607_ (_17809_, _06656_, _05974_);
  nor _68608_ (_17810_, _07939_, _10213_);
  nor _68609_ (_17811_, _10490_, _07776_);
  or _68610_ (_17812_, _17811_, _17810_);
  or _68611_ (_17813_, _17812_, _07215_);
  nand _68612_ (_17814_, _10744_, _07776_);
  nor _68613_ (_17815_, _10758_, _07154_);
  or _68614_ (_17816_, _17815_, _09450_);
  nor _68615_ (_17817_, _10755_, _07776_);
  or _68616_ (_17818_, _06781_, \oc8051_golden_model_1.ACC [2]);
  nand _68617_ (_17819_, _06781_, \oc8051_golden_model_1.ACC [2]);
  and _68618_ (_17820_, _17819_, _17818_);
  and _68619_ (_17821_, _17820_, _10755_);
  or _68620_ (_17822_, _17821_, _10758_);
  or _68621_ (_17823_, _17822_, _17817_);
  and _68622_ (_17824_, _17823_, _06015_);
  or _68623_ (_17825_, _17824_, _07154_);
  and _68624_ (_17826_, _17825_, _17816_);
  or _68625_ (_17827_, _17826_, _06341_);
  and _68626_ (_17828_, _14770_, _07939_);
  or _68627_ (_17829_, _17828_, _17810_);
  or _68628_ (_17830_, _17829_, _07151_);
  and _68629_ (_17831_, _17830_, _17827_);
  or _68630_ (_17832_, _17831_, _10775_);
  nor _68631_ (_17833_, _17547_, _10213_);
  and _68632_ (_17834_, _10778_, \oc8051_golden_model_1.PSW [6]);
  nor _68633_ (_17835_, _17834_, _17833_);
  nand _68634_ (_17836_, _17835_, _10775_);
  and _68635_ (_17837_, _17836_, _06466_);
  and _68636_ (_17838_, _17837_, _17832_);
  nor _68637_ (_17839_, _08636_, _10213_);
  and _68638_ (_17840_, _14774_, _08636_);
  or _68639_ (_17841_, _17840_, _17839_);
  and _68640_ (_17842_, _17841_, _06272_);
  and _68641_ (_17843_, _17812_, _06461_);
  or _68642_ (_17844_, _17843_, _10744_);
  or _68643_ (_17845_, _17844_, _17842_);
  or _68644_ (_17846_, _17845_, _17838_);
  and _68645_ (_17847_, _17846_, _17814_);
  or _68646_ (_17848_, _17847_, _07174_);
  or _68647_ (_17849_, _09450_, _07175_);
  and _68648_ (_17850_, _17849_, _06465_);
  and _68649_ (_17851_, _17850_, _17848_);
  nor _68650_ (_17852_, _08439_, _06465_);
  or _68651_ (_17853_, _17852_, _10811_);
  or _68652_ (_17854_, _17853_, _17851_);
  nand _68653_ (_17855_, _10811_, _10116_);
  and _68654_ (_17856_, _17855_, _17854_);
  or _68655_ (_17857_, _17856_, _06268_);
  and _68656_ (_17858_, _14756_, _08636_);
  or _68657_ (_17859_, _17858_, _17839_);
  or _68658_ (_17860_, _17859_, _06269_);
  and _68659_ (_17861_, _17860_, _06262_);
  and _68660_ (_17862_, _17861_, _17857_);
  or _68661_ (_17863_, _17839_, _14789_);
  and _68662_ (_17864_, _17841_, _06261_);
  and _68663_ (_17865_, _17864_, _17863_);
  or _68664_ (_17866_, _17865_, _09531_);
  or _68665_ (_17867_, _17866_, _17862_);
  nor _68666_ (_17868_, _10034_, _10032_);
  or _68667_ (_17869_, _17868_, _10035_);
  nand _68668_ (_17870_, _17869_, _09531_);
  and _68669_ (_17871_, _17870_, _10735_);
  and _68670_ (_17872_, _17871_, _17867_);
  and _68671_ (_17873_, _07357_, \oc8051_golden_model_1.ACC [1]);
  and _68672_ (_17874_, _07133_, _06097_);
  nor _68673_ (_17875_, _17874_, _11178_);
  nor _68674_ (_17876_, _17875_, _17873_);
  nor _68675_ (_17877_, _11175_, _17876_);
  and _68676_ (_17878_, _11175_, _17876_);
  nor _68677_ (_17879_, _17878_, _17877_);
  nor _68678_ (_17880_, _17243_, _11178_);
  and _68679_ (_17881_, _17880_, \oc8051_golden_model_1.PSW [7]);
  or _68680_ (_17882_, _17881_, _17879_);
  nand _68681_ (_17883_, _17881_, _17879_);
  and _68682_ (_17884_, _17883_, _10737_);
  and _68683_ (_17885_, _17884_, _17882_);
  or _68684_ (_17886_, _17885_, _17872_);
  and _68685_ (_17887_, _17886_, _10588_);
  and _68686_ (_17888_, _09347_, \oc8051_golden_model_1.ACC [1]);
  and _68687_ (_17889_, _09392_, _06097_);
  nor _68688_ (_17890_, _17889_, _11222_);
  nor _68689_ (_17891_, _17890_, _17888_);
  nor _68690_ (_17892_, _11219_, _17891_);
  and _68691_ (_17893_, _11219_, _17891_);
  nor _68692_ (_17894_, _17893_, _17892_);
  nor _68693_ (_17895_, _17377_, _11222_);
  not _68694_ (_17896_, _17895_);
  or _68695_ (_17897_, _17896_, _17894_);
  and _68696_ (_17898_, _17897_, \oc8051_golden_model_1.PSW [7]);
  nor _68697_ (_17899_, _17894_, \oc8051_golden_model_1.PSW [7]);
  nor _68698_ (_17900_, _17899_, _17898_);
  and _68699_ (_17901_, _17896_, _17894_);
  or _68700_ (_17902_, _17901_, _17900_);
  and _68701_ (_17903_, _17902_, _10656_);
  or _68702_ (_17904_, _17903_, _12644_);
  or _68703_ (_17905_, _17904_, _17887_);
  and _68704_ (_17906_, _08340_, \oc8051_golden_model_1.ACC [1]);
  and _68705_ (_17907_, _08390_, _06097_);
  nor _68706_ (_17908_, _14144_, _17907_);
  nor _68707_ (_17909_, _17908_, _17906_);
  nor _68708_ (_17910_, _11259_, _17909_);
  and _68709_ (_17911_, _11259_, _17909_);
  nor _68710_ (_17912_, _17911_, _17910_);
  and _68711_ (_17913_, _12582_, \oc8051_golden_model_1.PSW [7]);
  nand _68712_ (_17914_, _17913_, _17912_);
  or _68713_ (_17915_, _17913_, _17912_);
  and _68714_ (_17916_, _17915_, _17914_);
  or _68715_ (_17917_, _17916_, _06517_);
  nor _68716_ (_17918_, _17608_, _11303_);
  nor _68717_ (_17919_, _11300_, _17918_);
  and _68718_ (_17920_, _11300_, _17918_);
  nor _68719_ (_17921_, _17920_, _17919_);
  not _68720_ (_17922_, _17613_);
  nor _68721_ (_17923_, _17922_, _17921_);
  and _68722_ (_17924_, _17922_, _17921_);
  or _68723_ (_17925_, _17924_, _10517_);
  or _68724_ (_17926_, _17925_, _17923_);
  and _68725_ (_17927_, _17926_, _17917_);
  and _68726_ (_17928_, _17927_, _17905_);
  or _68727_ (_17929_, _17928_, _10515_);
  nand _68728_ (_17930_, _06656_, _10515_);
  and _68729_ (_17931_, _17930_, _06258_);
  and _68730_ (_17932_, _17931_, _17929_);
  and _68731_ (_17933_, _14804_, _08636_);
  or _68732_ (_17934_, _17933_, _17839_);
  and _68733_ (_17935_, _17934_, _06257_);
  or _68734_ (_17936_, _17935_, _10080_);
  or _68735_ (_17937_, _17936_, _17932_);
  and _68736_ (_17938_, _17937_, _17813_);
  or _68737_ (_17939_, _17938_, _07460_);
  and _68738_ (_17940_, _09450_, _07939_);
  or _68739_ (_17941_, _17810_, _07208_);
  or _68740_ (_17942_, _17941_, _17940_);
  and _68741_ (_17943_, _17942_, _05982_);
  and _68742_ (_17944_, _17943_, _17939_);
  and _68743_ (_17945_, _14859_, _07939_);
  or _68744_ (_17946_, _17945_, _17810_);
  and _68745_ (_17947_, _17946_, _10094_);
  or _68746_ (_17948_, _17947_, _10093_);
  or _68747_ (_17949_, _17948_, _17944_);
  or _68748_ (_17950_, _10286_, _10100_);
  and _68749_ (_17951_, _17950_, _17949_);
  or _68750_ (_17952_, _17951_, _05974_);
  and _68751_ (_17953_, _17952_, _17809_);
  or _68752_ (_17954_, _17953_, _06218_);
  and _68753_ (_17955_, _07939_, _08973_);
  or _68754_ (_17956_, _17955_, _17810_);
  or _68755_ (_17957_, _17956_, _06219_);
  and _68756_ (_17958_, _17957_, _10930_);
  and _68757_ (_17959_, _17958_, _17954_);
  nor _68758_ (_17960_, _10930_, _06656_);
  or _68759_ (_17961_, _17960_, _17959_);
  nor _68760_ (_17962_, _10937_, _06703_);
  and _68761_ (_17964_, _17962_, _17961_);
  not _68762_ (_17965_, _17962_);
  and _68763_ (_17966_, _17965_, _11175_);
  or _68764_ (_17967_, _17966_, _10506_);
  or _68765_ (_17968_, _17967_, _17964_);
  not _68766_ (_17969_, _10506_);
  or _68767_ (_17970_, _11175_, _17969_);
  and _68768_ (_17971_, _10732_, _06535_);
  not _68769_ (_17972_, _17971_);
  and _68770_ (_17973_, _17972_, _17970_);
  and _68771_ (_17974_, _17973_, _17968_);
  and _68772_ (_17975_, _17971_, _11175_);
  or _68773_ (_17976_, _17975_, _10948_);
  or _68774_ (_17977_, _17976_, _17974_);
  and _68775_ (_17978_, _17977_, _17808_);
  or _68776_ (_17979_, _17978_, _06533_);
  or _68777_ (_17980_, _11259_, _06534_);
  and _68778_ (_17981_, _17980_, _10955_);
  and _68779_ (_17982_, _17981_, _17979_);
  and _68780_ (_17983_, _10954_, _11300_);
  or _68781_ (_17984_, _17983_, _06369_);
  or _68782_ (_17985_, _17984_, _17982_);
  and _68783_ (_17986_, _14751_, _07939_);
  or _68784_ (_17987_, _17986_, _17810_);
  or _68785_ (_17988_, _17987_, _07237_);
  and _68786_ (_17989_, _17988_, _17985_);
  or _68787_ (_17990_, _17989_, _06536_);
  or _68788_ (_17991_, _17810_, _07240_);
  and _68789_ (_17992_, _17991_, _10977_);
  and _68790_ (_17993_, _17992_, _17990_);
  or _68791_ (_17994_, _10985_, _11173_);
  and _68792_ (_17995_, _17994_, _10987_);
  or _68793_ (_17996_, _17995_, _17993_);
  or _68794_ (_17997_, _17402_, _11173_);
  and _68795_ (_17998_, _17997_, _17401_);
  and _68796_ (_17999_, _17998_, _17996_);
  and _68797_ (_18000_, _10983_, _11217_);
  or _68798_ (_18001_, _18000_, _06542_);
  or _68799_ (_18002_, _18001_, _17999_);
  or _68800_ (_18003_, _11257_, _06543_);
  and _68801_ (_18004_, _18003_, _10497_);
  and _68802_ (_18005_, _18004_, _18002_);
  and _68803_ (_18006_, _11298_, _10496_);
  or _68804_ (_18007_, _18006_, _18005_);
  and _68805_ (_18008_, _18007_, _07242_);
  nand _68806_ (_18009_, _17956_, _06375_);
  nor _68807_ (_18010_, _18009_, _11258_);
  or _68808_ (_18011_, _18010_, _06711_);
  or _68809_ (_18012_, _18011_, _18008_);
  nor _68810_ (_18013_, _07042_, _06755_);
  nand _68811_ (_18014_, _11174_, _06711_);
  and _68812_ (_18015_, _18014_, _18013_);
  and _68813_ (_18016_, _18015_, _18012_);
  nor _68814_ (_18017_, _18013_, _11174_);
  or _68815_ (_18018_, _18017_, _17506_);
  or _68816_ (_18019_, _18018_, _18016_);
  nand _68817_ (_18020_, _17506_, _11174_);
  and _68818_ (_18021_, _18020_, _17430_);
  and _68819_ (_18022_, _18021_, _18019_);
  nor _68820_ (_18023_, _11174_, _17430_);
  or _68821_ (_18024_, _18023_, _11014_);
  or _68822_ (_18025_, _18024_, _18022_);
  and _68823_ (_18026_, _18025_, _17807_);
  or _68824_ (_18027_, _18026_, _06530_);
  nand _68825_ (_18028_, _11258_, _06530_);
  and _68826_ (_18029_, _18028_, _11024_);
  and _68827_ (_18030_, _18029_, _18027_);
  nor _68828_ (_18031_, _11024_, _11299_);
  or _68829_ (_18032_, _18031_, _06366_);
  or _68830_ (_18033_, _18032_, _18030_);
  and _68831_ (_18034_, _14748_, _07939_);
  or _68832_ (_18035_, _17810_, _09056_);
  or _68833_ (_18036_, _18035_, _18034_);
  and _68834_ (_18037_, _18036_, _11037_);
  and _68835_ (_18038_, _18037_, _18033_);
  and _68836_ (_18039_, _11052_, _10701_);
  nor _68837_ (_18040_, _18039_, _11053_);
  and _68838_ (_18041_, _18040_, _14283_);
  or _68839_ (_18042_, _18041_, _11041_);
  or _68840_ (_18043_, _18042_, _18038_);
  and _68841_ (_18044_, _11080_, _10627_);
  nor _68842_ (_18045_, _18044_, _11081_);
  or _68843_ (_18046_, _18045_, _11069_);
  and _68844_ (_18047_, _18046_, _06541_);
  and _68845_ (_18048_, _18047_, _18043_);
  nand _68846_ (_18049_, _11108_, _10874_);
  nor _68847_ (_18050_, _11109_, _06541_);
  and _68848_ (_18051_, _18050_, _18049_);
  or _68849_ (_18052_, _18051_, _11097_);
  or _68850_ (_18053_, _18052_, _18048_);
  and _68851_ (_18054_, _18053_, _17806_);
  or _68852_ (_18055_, _18054_, _11125_);
  nand _68853_ (_18056_, _11125_, _06042_);
  and _68854_ (_18057_, _18056_, _11157_);
  and _68855_ (_18058_, _18057_, _18055_);
  not _68856_ (_18059_, _11157_);
  nor _68857_ (_18060_, _11182_, _11175_);
  nor _68858_ (_18061_, _18060_, _11183_);
  and _68859_ (_18062_, _18061_, _18059_);
  or _68860_ (_18063_, _18062_, _11200_);
  or _68861_ (_18064_, _18063_, _18058_);
  and _68862_ (_18065_, _18064_, _17803_);
  or _68863_ (_18066_, _18065_, _11199_);
  not _68864_ (_18067_, _11199_);
  or _68865_ (_18068_, _17802_, _18067_);
  and _68866_ (_18069_, _18068_, _06285_);
  and _68867_ (_18070_, _18069_, _18066_);
  or _68868_ (_18071_, _18070_, _17799_);
  and _68869_ (_18072_, _18071_, _11321_);
  or _68870_ (_18073_, _11309_, _11300_);
  nor _68871_ (_18074_, _11310_, _11321_);
  and _68872_ (_18075_, _18074_, _18073_);
  or _68873_ (_18076_, _18075_, _11284_);
  or _68874_ (_18077_, _18076_, _18072_);
  and _68875_ (_18078_, _18077_, _17796_);
  or _68876_ (_18079_, _18078_, _06568_);
  or _68877_ (_18080_, _17829_, _06926_);
  and _68878_ (_18081_, _18080_, _11331_);
  and _68879_ (_18082_, _18081_, _18079_);
  nor _68880_ (_18083_, _17773_, _10213_);
  or _68881_ (_18084_, _18083_, _11336_);
  and _68882_ (_18085_, _18084_, _11330_);
  or _68883_ (_18086_, _18085_, _11335_);
  or _68884_ (_18087_, _18086_, _18082_);
  nand _68885_ (_18088_, _11335_, _06055_);
  and _68886_ (_18089_, _18088_, _05928_);
  and _68887_ (_18090_, _18089_, _18087_);
  and _68888_ (_18091_, _17859_, _05927_);
  or _68889_ (_18092_, _18091_, _06278_);
  or _68890_ (_18093_, _18092_, _18090_);
  and _68891_ (_18094_, _14926_, _07939_);
  or _68892_ (_18095_, _18094_, _17810_);
  or _68893_ (_18096_, _18095_, _06279_);
  and _68894_ (_18097_, _18096_, _11354_);
  and _68895_ (_18098_, _18097_, _18093_);
  nor _68896_ (_18099_, _11361_, \oc8051_golden_model_1.ACC [2]);
  nor _68897_ (_18100_, _18099_, _11362_);
  and _68898_ (_18101_, _18100_, _11353_);
  or _68899_ (_18102_, _18101_, _11360_);
  or _68900_ (_18103_, _18102_, _18098_);
  nand _68901_ (_18104_, _11360_, _06055_);
  and _68902_ (_18105_, _18104_, _01347_);
  and _68903_ (_18106_, _18105_, _18103_);
  or _68904_ (_18107_, _18106_, _17795_);
  and _68905_ (_43164_, _18107_, _42618_);
  nor _68906_ (_18108_, _01347_, _06055_);
  and _68907_ (_18109_, _11054_, _10696_);
  nor _68908_ (_18110_, _18109_, _11055_);
  and _68909_ (_18111_, _18110_, _17724_);
  or _68910_ (_18112_, _18111_, _11037_);
  nor _68911_ (_18113_, _11215_, _11216_);
  or _68912_ (_18114_, _18113_, _06885_);
  nand _68913_ (_18115_, _06213_, _05974_);
  nor _68914_ (_18116_, _07939_, _06055_);
  nor _68915_ (_18117_, _10490_, _07594_);
  or _68916_ (_18118_, _18117_, _18116_);
  or _68917_ (_18119_, _18118_, _07215_);
  and _68918_ (_18120_, _06656_, \oc8051_golden_model_1.ACC [2]);
  nor _68919_ (_18121_, _17919_, _18120_);
  nor _68920_ (_18122_, _12594_, _18121_);
  and _68921_ (_18123_, _12594_, _18121_);
  nor _68922_ (_18124_, _18123_, _18122_);
  or _68923_ (_18125_, _17923_, _18124_);
  nand _68924_ (_18126_, _17923_, _18124_);
  and _68925_ (_18127_, _18126_, _18125_);
  or _68926_ (_18128_, _18127_, _10517_);
  nor _68927_ (_18129_, _08636_, _06055_);
  and _68928_ (_18130_, _14950_, _08636_);
  or _68929_ (_18131_, _18130_, _18129_);
  or _68930_ (_18132_, _18129_, _14979_);
  and _68931_ (_18133_, _18132_, _06261_);
  and _68932_ (_18134_, _18133_, _18131_);
  nand _68933_ (_18135_, _10744_, _07594_);
  or _68934_ (_18136_, _18131_, _06273_);
  and _68935_ (_18137_, _18136_, _07166_);
  and _68936_ (_18138_, _14953_, _07939_);
  or _68937_ (_18139_, _18138_, _18116_);
  and _68938_ (_18140_, _18139_, _06341_);
  nand _68939_ (_18141_, _10756_, _07594_);
  nor _68940_ (_18142_, _06781_, _06055_);
  and _68941_ (_18143_, _06781_, _06055_);
  nor _68942_ (_18144_, _18143_, _18142_);
  nand _68943_ (_18145_, _18144_, _10755_);
  and _68944_ (_18146_, _18145_, _10759_);
  and _68945_ (_18147_, _18146_, _18141_);
  and _68946_ (_18148_, _18147_, _07155_);
  or _68947_ (_18149_, _18148_, _09449_);
  or _68948_ (_18150_, _18147_, _10758_);
  and _68949_ (_18151_, _18150_, _06015_);
  or _68950_ (_18152_, _18151_, _07154_);
  and _68951_ (_18153_, _18152_, _07151_);
  and _68952_ (_18154_, _18153_, _18149_);
  or _68953_ (_18155_, _18154_, _18140_);
  and _68954_ (_18156_, _18155_, _10776_);
  not _68955_ (_18157_, \oc8051_golden_model_1.PSW [6]);
  nor _68956_ (_18158_, _10778_, _18157_);
  nor _68957_ (_18159_, _18158_, \oc8051_golden_model_1.ACC [3]);
  nor _68958_ (_18160_, _18159_, _10779_);
  and _68959_ (_18161_, _18160_, _10775_);
  or _68960_ (_18162_, _18161_, _06272_);
  or _68961_ (_18163_, _18162_, _18156_);
  and _68962_ (_18164_, _18163_, _18137_);
  and _68963_ (_18165_, _18118_, _06461_);
  or _68964_ (_18166_, _18165_, _10744_);
  or _68965_ (_18167_, _18166_, _18164_);
  and _68966_ (_18168_, _18167_, _18135_);
  or _68967_ (_18169_, _18168_, _07174_);
  or _68968_ (_18170_, _09449_, _07175_);
  and _68969_ (_18171_, _18170_, _06465_);
  and _68970_ (_18172_, _18171_, _18169_);
  nor _68971_ (_18173_, _08291_, _06465_);
  or _68972_ (_18174_, _18173_, _10811_);
  or _68973_ (_18175_, _18174_, _18172_);
  nand _68974_ (_18176_, _10811_, _08572_);
  and _68975_ (_18177_, _18176_, _18175_);
  or _68976_ (_18178_, _18177_, _06268_);
  and _68977_ (_18179_, _14948_, _08636_);
  or _68978_ (_18180_, _18179_, _18129_);
  or _68979_ (_18181_, _18180_, _06269_);
  and _68980_ (_18182_, _18181_, _06262_);
  and _68981_ (_18183_, _18182_, _18178_);
  or _68982_ (_18184_, _18183_, _18134_);
  and _68983_ (_18185_, _18184_, _09537_);
  or _68984_ (_18186_, _10037_, _10035_);
  nor _68985_ (_18187_, _10038_, _09537_);
  nand _68986_ (_18188_, _18187_, _18186_);
  nand _68987_ (_18189_, _18188_, _10731_);
  or _68988_ (_18190_, _18189_, _18185_);
  and _68989_ (_18191_, _07776_, \oc8051_golden_model_1.ACC [2]);
  nor _68990_ (_18192_, _17877_, _18191_);
  nor _68991_ (_18193_, _11171_, _11172_);
  not _68992_ (_18194_, _18193_);
  and _68993_ (_18195_, _18194_, _18192_);
  nor _68994_ (_18196_, _18194_, _18192_);
  nor _68995_ (_18197_, _18196_, _18195_);
  nor _68996_ (_18198_, _18197_, _10558_);
  and _68997_ (_18199_, _18197_, _10558_);
  nor _68998_ (_18200_, _18199_, _18198_);
  and _68999_ (_18201_, _17879_, \oc8051_golden_model_1.PSW [7]);
  nor _69000_ (_18202_, _17880_, _10558_);
  nor _69001_ (_18203_, _18202_, _18201_);
  not _69002_ (_18204_, _18203_);
  and _69003_ (_18205_, _18204_, _18200_);
  nor _69004_ (_18206_, _18204_, _18200_);
  nor _69005_ (_18207_, _18206_, _18205_);
  and _69006_ (_18208_, _18207_, _10734_);
  or _69007_ (_18209_, _18208_, _10735_);
  and _69008_ (_18210_, _18209_, _18190_);
  and _69009_ (_18211_, _18207_, _10733_);
  or _69010_ (_18212_, _18211_, _10656_);
  or _69011_ (_18213_, _18212_, _18210_);
  and _69012_ (_18214_, _09302_, \oc8051_golden_model_1.ACC [2]);
  nor _69013_ (_18215_, _17892_, _18214_);
  nor _69014_ (_18216_, _18113_, _18215_);
  and _69015_ (_18217_, _18113_, _18215_);
  nor _69016_ (_18218_, _18217_, _18216_);
  and _69017_ (_18219_, _18218_, \oc8051_golden_model_1.PSW [7]);
  nor _69018_ (_18220_, _18218_, \oc8051_golden_model_1.PSW [7]);
  nor _69019_ (_18221_, _18220_, _18219_);
  and _69020_ (_18222_, _18221_, _17898_);
  nor _69021_ (_18223_, _18221_, _17898_);
  nor _69022_ (_18224_, _18223_, _18222_);
  or _69023_ (_18225_, _18224_, _10588_);
  and _69024_ (_18226_, _18225_, _06517_);
  and _69025_ (_18227_, _18226_, _18213_);
  and _69026_ (_18228_, _12583_, \oc8051_golden_model_1.PSW [7]);
  and _69027_ (_18229_, _08439_, \oc8051_golden_model_1.ACC [2]);
  nor _69028_ (_18230_, _17910_, _18229_);
  nor _69029_ (_18231_, _12577_, _18230_);
  and _69030_ (_18232_, _12577_, _18230_);
  nor _69031_ (_18233_, _18232_, _18231_);
  not _69032_ (_18234_, _12582_);
  or _69033_ (_18235_, _18234_, _17912_);
  or _69034_ (_18236_, _18235_, _10558_);
  and _69035_ (_18237_, _18236_, _18233_);
  or _69036_ (_18238_, _18237_, _10516_);
  or _69037_ (_18239_, _18238_, _18228_);
  and _69038_ (_18240_, _18239_, _12644_);
  or _69039_ (_18241_, _18240_, _18227_);
  and _69040_ (_18242_, _18241_, _18128_);
  or _69041_ (_18243_, _18242_, _10515_);
  nand _69042_ (_18244_, _06213_, _10515_);
  and _69043_ (_18245_, _18244_, _06258_);
  and _69044_ (_18246_, _18245_, _18243_);
  or _69045_ (_18247_, _18129_, _14992_);
  and _69046_ (_18248_, _18247_, _06257_);
  and _69047_ (_18249_, _18248_, _18131_);
  or _69048_ (_18250_, _18249_, _10080_);
  or _69049_ (_18251_, _18250_, _18246_);
  and _69050_ (_18252_, _18251_, _18119_);
  or _69051_ (_18253_, _18252_, _07460_);
  and _69052_ (_18254_, _09449_, _07939_);
  or _69053_ (_18255_, _18116_, _07208_);
  or _69054_ (_18256_, _18255_, _18254_);
  and _69055_ (_18257_, _18256_, _05982_);
  and _69056_ (_18258_, _18257_, _18253_);
  and _69057_ (_18259_, _15048_, _07939_);
  or _69058_ (_18260_, _18259_, _18116_);
  and _69059_ (_18261_, _18260_, _10094_);
  or _69060_ (_18262_, _18261_, _10093_);
  or _69061_ (_18263_, _18262_, _18258_);
  or _69062_ (_18264_, _10235_, _10100_);
  and _69063_ (_18265_, _18264_, _18263_);
  or _69064_ (_18266_, _18265_, _05974_);
  and _69065_ (_18267_, _18266_, _18115_);
  or _69066_ (_18268_, _18267_, _06218_);
  and _69067_ (_18269_, _07939_, _08930_);
  or _69068_ (_18270_, _18269_, _18116_);
  or _69069_ (_18271_, _18270_, _06219_);
  and _69070_ (_18272_, _18271_, _10930_);
  and _69071_ (_18273_, _18272_, _18268_);
  or _69072_ (_18274_, _10930_, _06213_);
  or _69073_ (_18275_, _06734_, _06328_);
  and _69074_ (_18276_, _18275_, _06535_);
  and _69075_ (_18277_, _06335_, _06535_);
  or _69076_ (_18278_, _10506_, _18277_);
  nor _69077_ (_18279_, _18278_, _18276_);
  nand _69078_ (_18280_, _18279_, _18274_);
  or _69079_ (_18281_, _18280_, _18273_);
  nor _69080_ (_18282_, _17511_, _06887_);
  or _69081_ (_18283_, _18279_, _18193_);
  and _69082_ (_18284_, _18283_, _18282_);
  and _69083_ (_18285_, _18284_, _18281_);
  not _69084_ (_18286_, _18282_);
  and _69085_ (_18287_, _18286_, _18193_);
  or _69086_ (_18288_, _18287_, _06888_);
  or _69087_ (_18289_, _18288_, _18285_);
  or _69088_ (_18290_, _18193_, _17510_);
  and _69089_ (_18291_, _18290_, _17375_);
  and _69090_ (_18292_, _18291_, _18289_);
  or _69091_ (_18293_, _18113_, _06884_);
  and _69092_ (_18294_, _18293_, _10948_);
  or _69093_ (_18295_, _18294_, _18292_);
  and _69094_ (_18296_, _18295_, _18114_);
  or _69095_ (_18297_, _18296_, _06533_);
  or _69096_ (_18298_, _12577_, _06534_);
  and _69097_ (_18299_, _18298_, _10955_);
  and _69098_ (_18300_, _18299_, _18297_);
  and _69099_ (_18301_, _10954_, _12594_);
  or _69100_ (_18302_, _18301_, _06369_);
  or _69101_ (_18303_, _18302_, _18300_);
  and _69102_ (_18304_, _14943_, _07939_);
  or _69103_ (_18305_, _18304_, _18116_);
  or _69104_ (_18306_, _18305_, _07237_);
  and _69105_ (_18307_, _18306_, _18303_);
  or _69106_ (_18308_, _18307_, _06536_);
  or _69107_ (_18309_, _18116_, _07240_);
  and _69108_ (_18310_, _18309_, _10977_);
  and _69109_ (_18311_, _18310_, _18308_);
  or _69110_ (_18312_, _10985_, _11171_);
  and _69111_ (_18313_, _18312_, _10987_);
  or _69112_ (_18314_, _18313_, _18311_);
  or _69113_ (_18315_, _17402_, _11171_);
  and _69114_ (_18316_, _18315_, _17401_);
  and _69115_ (_18317_, _18316_, _18314_);
  and _69116_ (_18318_, _10983_, _11215_);
  or _69117_ (_18319_, _18318_, _06542_);
  or _69118_ (_18320_, _18319_, _18317_);
  or _69119_ (_18321_, _11255_, _06543_);
  and _69120_ (_18322_, _18321_, _10497_);
  and _69121_ (_18323_, _18322_, _18320_);
  and _69122_ (_18324_, _11296_, _10496_);
  or _69123_ (_18325_, _18324_, _18323_);
  and _69124_ (_18326_, _18325_, _07242_);
  nand _69125_ (_18327_, _18270_, _06375_);
  nor _69126_ (_18328_, _18327_, _11256_);
  or _69127_ (_18329_, _18328_, _10999_);
  or _69128_ (_18330_, _18329_, _18326_);
  nand _69129_ (_18331_, _10999_, _11172_);
  and _69130_ (_18332_, _18331_, _07043_);
  and _69131_ (_18333_, _18332_, _11009_);
  and _69132_ (_18334_, _18333_, _18330_);
  and _69133_ (_18335_, _11009_, _07043_);
  nor _69134_ (_18336_, _18335_, _11172_);
  or _69135_ (_18337_, _18336_, _11014_);
  or _69136_ (_18338_, _18337_, _18334_);
  nand _69137_ (_18339_, _11014_, _11216_);
  and _69138_ (_18340_, _18339_, _06531_);
  and _69139_ (_18341_, _18340_, _18338_);
  nand _69140_ (_18342_, _11024_, _11256_);
  and _69141_ (_18343_, _18342_, _11023_);
  or _69142_ (_18344_, _18343_, _18341_);
  nand _69143_ (_18345_, _11021_, _11297_);
  and _69144_ (_18346_, _18345_, _09056_);
  and _69145_ (_18347_, _18346_, _18344_);
  and _69146_ (_18348_, _14940_, _07939_);
  or _69147_ (_18349_, _18348_, _18116_);
  nand _69148_ (_18350_, _18349_, _06366_);
  nand _69149_ (_18351_, _18350_, _17505_);
  or _69150_ (_18352_, _18351_, _18347_);
  and _69151_ (_18353_, _18352_, _18112_);
  and _69152_ (_18354_, _18110_, _17723_);
  or _69153_ (_18355_, _18354_, _11041_);
  or _69154_ (_18356_, _18355_, _18353_);
  and _69155_ (_18357_, _11082_, _10622_);
  nor _69156_ (_18358_, _18357_, _11083_);
  or _69157_ (_18359_, _18358_, _11069_);
  and _69158_ (_18360_, _18359_, _06541_);
  and _69159_ (_18361_, _18360_, _18356_);
  and _69160_ (_18362_, _11110_, _10869_);
  nor _69161_ (_18363_, _18362_, _11111_);
  or _69162_ (_18364_, _18363_, _11097_);
  and _69163_ (_18365_, _18364_, _14297_);
  or _69164_ (_18366_, _18365_, _18361_);
  and _69165_ (_18367_, _11138_, _10551_);
  nor _69166_ (_18368_, _18367_, _11139_);
  or _69167_ (_18369_, _18368_, _11127_);
  and _69168_ (_18370_, _18369_, _11126_);
  and _69169_ (_18371_, _18370_, _18366_);
  and _69170_ (_18372_, _11125_, \oc8051_golden_model_1.ACC [2]);
  nor _69171_ (_18373_, _18372_, _11201_);
  nand _69172_ (_18374_, _18373_, _11157_);
  or _69173_ (_18375_, _18374_, _18371_);
  nor _69174_ (_18376_, _11228_, _18113_);
  and _69175_ (_18377_, _11228_, _18113_);
  or _69176_ (_18378_, _18377_, _18376_);
  or _69177_ (_18379_, _18378_, _11203_);
  or _69178_ (_18380_, _11184_, _18194_);
  nand _69179_ (_18381_, _11184_, _18194_);
  and _69180_ (_18382_, _18381_, _18380_);
  or _69181_ (_18383_, _18382_, _11157_);
  and _69182_ (_18384_, _18383_, _06285_);
  and _69183_ (_18385_, _18384_, _18379_);
  and _69184_ (_18386_, _18385_, _18375_);
  and _69185_ (_18387_, _11268_, _12577_);
  nor _69186_ (_18388_, _11268_, _12577_);
  or _69187_ (_18389_, _18388_, _18387_);
  and _69188_ (_18390_, _18389_, _06283_);
  or _69189_ (_18391_, _18390_, _11243_);
  or _69190_ (_18392_, _18391_, _18386_);
  and _69191_ (_18393_, _11311_, _12594_);
  nor _69192_ (_18394_, _11311_, _12594_);
  or _69193_ (_18395_, _18394_, _11321_);
  or _69194_ (_18396_, _18395_, _18393_);
  and _69195_ (_18397_, _18396_, _11285_);
  and _69196_ (_18398_, _18397_, _18392_);
  and _69197_ (_18399_, _11284_, \oc8051_golden_model_1.ACC [2]);
  or _69198_ (_18400_, _18399_, _06568_);
  or _69199_ (_18401_, _18400_, _18398_);
  or _69200_ (_18402_, _18139_, _06926_);
  and _69201_ (_18403_, _18402_, _11331_);
  and _69202_ (_18404_, _18403_, _18401_);
  nor _69203_ (_18405_, _11336_, _06055_);
  or _69204_ (_18406_, _18405_, _11337_);
  and _69205_ (_18407_, _18406_, _11330_);
  or _69206_ (_18408_, _18407_, _11335_);
  or _69207_ (_18409_, _18408_, _18404_);
  nand _69208_ (_18410_, _11335_, _10135_);
  and _69209_ (_18411_, _18410_, _05928_);
  and _69210_ (_18412_, _18411_, _18409_);
  and _69211_ (_18413_, _18180_, _05927_);
  or _69212_ (_18414_, _18413_, _06278_);
  or _69213_ (_18415_, _18414_, _18412_);
  and _69214_ (_18416_, _15128_, _07939_);
  or _69215_ (_18417_, _18416_, _18116_);
  or _69216_ (_18418_, _18417_, _06279_);
  and _69217_ (_18419_, _18418_, _11354_);
  and _69218_ (_18420_, _18419_, _18415_);
  nor _69219_ (_18421_, _11362_, \oc8051_golden_model_1.ACC [3]);
  nor _69220_ (_18422_, _18421_, _11363_);
  and _69221_ (_18423_, _18422_, _11353_);
  or _69222_ (_18424_, _18423_, _11360_);
  or _69223_ (_18425_, _18424_, _18420_);
  nand _69224_ (_18426_, _11360_, _10135_);
  and _69225_ (_18427_, _18426_, _01347_);
  and _69226_ (_18428_, _18427_, _18425_);
  or _69227_ (_18429_, _18428_, _18108_);
  and _69228_ (_43165_, _18429_, _42618_);
  nor _69229_ (_18430_, _01347_, _10135_);
  or _69230_ (_18431_, _11230_, _11214_);
  and _69231_ (_18432_, _18431_, _11231_);
  or _69232_ (_18433_, _18432_, _17800_);
  or _69233_ (_18434_, _11056_, _10689_);
  and _69234_ (_18435_, _18434_, _11057_);
  and _69235_ (_18436_, _18435_, _14283_);
  nand _69236_ (_18437_, _11021_, _11294_);
  or _69237_ (_18438_, _12157_, _11169_);
  or _69238_ (_18439_, _17401_, _11211_);
  or _69239_ (_18440_, _11214_, _10502_);
  nand _69240_ (_18441_, _06968_, _05974_);
  nor _69241_ (_18442_, _07939_, _10135_);
  nor _69242_ (_18443_, _08541_, _10490_);
  or _69243_ (_18444_, _18443_, _18442_);
  or _69244_ (_18445_, _18444_, _07215_);
  nor _69245_ (_18446_, _12583_, _10558_);
  or _69246_ (_18447_, _18230_, _14140_);
  and _69247_ (_18448_, _18447_, _14139_);
  nor _69248_ (_18449_, _11254_, _18448_);
  and _69249_ (_18450_, _11254_, _18448_);
  nor _69250_ (_18451_, _18450_, _18449_);
  and _69251_ (_18452_, _18451_, \oc8051_golden_model_1.PSW [7]);
  nor _69252_ (_18453_, _18451_, \oc8051_golden_model_1.PSW [7]);
  nor _69253_ (_18454_, _18453_, _18452_);
  or _69254_ (_18455_, _18454_, _18446_);
  and _69255_ (_18456_, _18454_, _18446_);
  nor _69256_ (_18457_, _18456_, _06517_);
  and _69257_ (_18458_, _18457_, _18455_);
  or _69258_ (_18459_, _18205_, _18198_);
  nor _69259_ (_18460_, _07594_, \oc8051_golden_model_1.ACC [3]);
  nand _69260_ (_18461_, _07594_, \oc8051_golden_model_1.ACC [3]);
  and _69261_ (_18462_, _18461_, _18192_);
  or _69262_ (_18463_, _18462_, _18460_);
  nor _69263_ (_18464_, _11170_, _18463_);
  and _69264_ (_18465_, _11170_, _18463_);
  nor _69265_ (_18466_, _18465_, _18464_);
  and _69266_ (_18467_, _18466_, \oc8051_golden_model_1.PSW [7]);
  nor _69267_ (_18468_, _18466_, \oc8051_golden_model_1.PSW [7]);
  nor _69268_ (_18469_, _18468_, _18467_);
  or _69269_ (_18470_, _18469_, _18459_);
  and _69270_ (_18471_, _18469_, _18459_);
  nor _69271_ (_18472_, _10735_, _18471_);
  and _69272_ (_18473_, _18472_, _18470_);
  nand _69273_ (_18474_, _10744_, _08541_);
  nor _69274_ (_18475_, _08636_, _10135_);
  and _69275_ (_18476_, _15166_, _08636_);
  or _69276_ (_18477_, _18476_, _18475_);
  or _69277_ (_18478_, _18477_, _06273_);
  and _69278_ (_18479_, _18478_, _07166_);
  nand _69279_ (_18480_, _10756_, _08541_);
  nor _69280_ (_18481_, _06781_, _10135_);
  and _69281_ (_18482_, _06781_, _10135_);
  nor _69282_ (_18483_, _18482_, _18481_);
  nand _69283_ (_18484_, _18483_, _10755_);
  and _69284_ (_18485_, _18484_, _10759_);
  and _69285_ (_18486_, _18485_, _18480_);
  and _69286_ (_18487_, _10758_, _09448_);
  or _69287_ (_18488_, _18487_, _18486_);
  and _69288_ (_18489_, _18488_, _10769_);
  and _69289_ (_18490_, _15162_, _07939_);
  or _69290_ (_18491_, _18490_, _18442_);
  and _69291_ (_18492_, _18491_, _06341_);
  or _69292_ (_18493_, _18492_, _18489_);
  and _69293_ (_18494_, _18493_, _10776_);
  nor _69294_ (_18495_, _10779_, \oc8051_golden_model_1.ACC [4]);
  nor _69295_ (_18496_, _18495_, _10780_);
  and _69296_ (_18497_, _18496_, _10775_);
  or _69297_ (_18498_, _18497_, _06272_);
  or _69298_ (_18499_, _18498_, _18494_);
  and _69299_ (_18500_, _18499_, _18479_);
  and _69300_ (_18501_, _18444_, _06461_);
  or _69301_ (_18502_, _18501_, _10744_);
  or _69302_ (_18503_, _18502_, _18500_);
  and _69303_ (_18504_, _18503_, _18474_);
  or _69304_ (_18505_, _18504_, _07174_);
  or _69305_ (_18506_, _09448_, _07175_);
  and _69306_ (_18507_, _18506_, _06465_);
  and _69307_ (_18508_, _18507_, _18505_);
  nor _69308_ (_18509_, _08543_, _06465_);
  or _69309_ (_18510_, _18509_, _10811_);
  or _69310_ (_18511_, _18510_, _18508_);
  nand _69311_ (_18512_, _10811_, _06097_);
  and _69312_ (_18513_, _18512_, _18511_);
  or _69313_ (_18514_, _18513_, _06268_);
  and _69314_ (_18515_, _15176_, _08636_);
  or _69315_ (_18516_, _18515_, _18475_);
  or _69316_ (_18517_, _18516_, _06269_);
  and _69317_ (_18518_, _18517_, _06262_);
  and _69318_ (_18519_, _18518_, _18514_);
  or _69319_ (_18520_, _18475_, _15183_);
  and _69320_ (_18521_, _18520_, _06261_);
  and _69321_ (_18522_, _18521_, _18477_);
  or _69322_ (_18523_, _18522_, _09531_);
  or _69323_ (_18524_, _18523_, _18519_);
  nor _69324_ (_18525_, _10040_, _10038_);
  nor _69325_ (_18526_, _18525_, _10041_);
  or _69326_ (_18527_, _18526_, _09537_);
  and _69327_ (_18528_, _18527_, _10735_);
  and _69328_ (_18529_, _18528_, _18524_);
  nor _69329_ (_18530_, _18529_, _18473_);
  nor _69330_ (_18531_, _18530_, _10587_);
  or _69331_ (_18532_, _18222_, _18219_);
  and _69332_ (_18533_, _09449_, _06055_);
  or _69333_ (_18534_, _09449_, _06055_);
  and _69334_ (_18535_, _18534_, _18215_);
  or _69335_ (_18536_, _18535_, _18533_);
  nor _69336_ (_18537_, _11214_, _18536_);
  and _69337_ (_18538_, _11214_, _18536_);
  nor _69338_ (_18539_, _18538_, _18537_);
  and _69339_ (_18540_, _18539_, \oc8051_golden_model_1.PSW [7]);
  nor _69340_ (_18541_, _18539_, \oc8051_golden_model_1.PSW [7]);
  nor _69341_ (_18542_, _18541_, _18540_);
  and _69342_ (_18543_, _18542_, _18532_);
  nor _69343_ (_18544_, _18542_, _18532_);
  nor _69344_ (_18545_, _18544_, _18543_);
  and _69345_ (_18546_, _18545_, _10587_);
  or _69346_ (_18547_, _18546_, _18531_);
  or _69347_ (_18548_, _18547_, _10586_);
  not _69348_ (_18549_, _10586_);
  or _69349_ (_18550_, _18545_, _18549_);
  and _69350_ (_18551_, _18550_, _06517_);
  and _69351_ (_18552_, _18551_, _18548_);
  or _69352_ (_18553_, _18552_, _18458_);
  and _69353_ (_18554_, _18553_, _10517_);
  nor _69354_ (_18555_, _12599_, _10558_);
  or _69355_ (_18556_, _18121_, _14161_);
  and _69356_ (_18557_, _18556_, _14160_);
  nor _69357_ (_18558_, _11295_, _18557_);
  and _69358_ (_18559_, _11295_, _18557_);
  nor _69359_ (_18560_, _18559_, _18558_);
  and _69360_ (_18561_, _18560_, \oc8051_golden_model_1.PSW [7]);
  nor _69361_ (_18562_, _18560_, \oc8051_golden_model_1.PSW [7]);
  nor _69362_ (_18563_, _18562_, _18561_);
  or _69363_ (_18564_, _18563_, _18555_);
  and _69364_ (_18565_, _18563_, _18555_);
  nor _69365_ (_18566_, _18565_, _10517_);
  and _69366_ (_18567_, _18566_, _18564_);
  or _69367_ (_18568_, _18567_, _10515_);
  or _69368_ (_18569_, _18568_, _18554_);
  nand _69369_ (_18570_, _06968_, _10515_);
  and _69370_ (_18571_, _18570_, _06258_);
  and _69371_ (_18572_, _18571_, _18569_);
  and _69372_ (_18573_, _15200_, _08636_);
  or _69373_ (_18574_, _18573_, _18475_);
  and _69374_ (_18575_, _18574_, _06257_);
  or _69375_ (_18576_, _18575_, _10080_);
  or _69376_ (_18577_, _18576_, _18572_);
  and _69377_ (_18578_, _18577_, _18445_);
  or _69378_ (_18579_, _18578_, _07460_);
  and _69379_ (_18580_, _09448_, _07939_);
  or _69380_ (_18581_, _18442_, _07208_);
  or _69381_ (_18582_, _18581_, _18580_);
  and _69382_ (_18583_, _18582_, _05982_);
  and _69383_ (_18584_, _18583_, _18579_);
  and _69384_ (_18585_, _15254_, _07939_);
  or _69385_ (_18586_, _18585_, _18442_);
  and _69386_ (_18587_, _18586_, _10094_);
  or _69387_ (_18588_, _18587_, _10093_);
  or _69388_ (_18589_, _18588_, _18584_);
  or _69389_ (_18590_, _10181_, _10100_);
  and _69390_ (_18591_, _18590_, _18589_);
  or _69391_ (_18592_, _18591_, _05974_);
  and _69392_ (_18593_, _18592_, _18441_);
  or _69393_ (_18594_, _18593_, _06218_);
  and _69394_ (_18595_, _08959_, _07939_);
  or _69395_ (_18596_, _18595_, _18442_);
  or _69396_ (_18597_, _18596_, _06219_);
  and _69397_ (_18598_, _18597_, _10930_);
  and _69398_ (_18599_, _18598_, _18594_);
  nor _69399_ (_18600_, _10930_, _06968_);
  or _69400_ (_18601_, _18600_, _18277_);
  or _69401_ (_18602_, _18601_, _18599_);
  not _69402_ (_18603_, _18277_);
  or _69403_ (_18604_, _11170_, _18603_);
  and _69404_ (_18605_, _18604_, _18602_);
  or _69405_ (_18606_, _18605_, _06891_);
  not _69406_ (_18607_, _06891_);
  or _69407_ (_18608_, _11170_, _18607_);
  and _69408_ (_18609_, _18608_, _06745_);
  and _69409_ (_18610_, _18609_, _18606_);
  and _69410_ (_18611_, _11170_, _06744_);
  or _69411_ (_18612_, _18611_, _10507_);
  or _69412_ (_18613_, _18612_, _18610_);
  not _69413_ (_18614_, _10507_);
  or _69414_ (_18615_, _11170_, _18614_);
  and _69415_ (_18616_, _18615_, _17972_);
  and _69416_ (_18617_, _18616_, _18613_);
  and _69417_ (_18618_, _17971_, _11170_);
  or _69418_ (_18619_, _18618_, _10948_);
  or _69419_ (_18620_, _18619_, _18617_);
  and _69420_ (_18621_, _18620_, _18440_);
  or _69421_ (_18622_, _18621_, _06533_);
  or _69422_ (_18623_, _11254_, _06534_);
  and _69423_ (_18624_, _18623_, _10955_);
  and _69424_ (_18625_, _18624_, _18622_);
  and _69425_ (_18626_, _10954_, _11295_);
  or _69426_ (_18627_, _18626_, _06369_);
  or _69427_ (_18628_, _18627_, _18625_);
  and _69428_ (_18629_, _15269_, _07939_);
  or _69429_ (_18630_, _18629_, _18442_);
  or _69430_ (_18631_, _18630_, _07237_);
  and _69431_ (_18632_, _18631_, _18628_);
  or _69432_ (_18633_, _18632_, _06536_);
  or _69433_ (_18634_, _18442_, _07240_);
  and _69434_ (_18635_, _18634_, _10986_);
  and _69435_ (_18636_, _18635_, _18633_);
  and _69436_ (_18637_, _10987_, _11167_);
  or _69437_ (_18638_, _18637_, _10983_);
  or _69438_ (_18639_, _18638_, _18636_);
  and _69439_ (_18640_, _18639_, _18439_);
  or _69440_ (_18641_, _18640_, _06542_);
  or _69441_ (_18642_, _11251_, _06543_);
  and _69442_ (_18643_, _18642_, _10497_);
  and _69443_ (_18644_, _18643_, _18641_);
  and _69444_ (_18645_, _11292_, _10496_);
  or _69445_ (_18646_, _18645_, _18644_);
  and _69446_ (_18647_, _18646_, _07242_);
  nand _69447_ (_18648_, _18596_, _06375_);
  nor _69448_ (_18649_, _18648_, _11253_);
  or _69449_ (_18650_, _18649_, _17507_);
  or _69450_ (_18651_, _18650_, _18647_);
  and _69451_ (_18652_, _18651_, _18438_);
  or _69452_ (_18653_, _18652_, _17506_);
  or _69453_ (_18654_, _17423_, _11169_);
  and _69454_ (_18655_, _18654_, _17430_);
  and _69455_ (_18656_, _18655_, _18653_);
  and _69456_ (_18657_, _11169_, _17429_);
  or _69457_ (_18658_, _18657_, _11014_);
  or _69458_ (_18659_, _18658_, _18656_);
  or _69459_ (_18660_, _11013_, _11213_);
  and _69460_ (_18661_, _18660_, _06531_);
  and _69461_ (_18662_, _18661_, _18659_);
  nand _69462_ (_18663_, _11024_, _11253_);
  and _69463_ (_18664_, _18663_, _11023_);
  or _69464_ (_18665_, _18664_, _18662_);
  and _69465_ (_18666_, _18665_, _18437_);
  or _69466_ (_18667_, _18666_, _06366_);
  and _69467_ (_18668_, _15266_, _07939_);
  or _69468_ (_18669_, _18442_, _09056_);
  or _69469_ (_18670_, _18669_, _18668_);
  and _69470_ (_18671_, _18670_, _11037_);
  and _69471_ (_18672_, _18671_, _18667_);
  or _69472_ (_18673_, _18672_, _18436_);
  and _69473_ (_18674_, _18673_, _17722_);
  or _69474_ (_18675_, _11084_, _10616_);
  and _69475_ (_18676_, _18675_, _11085_);
  and _69476_ (_18677_, _18676_, _11040_);
  or _69477_ (_18678_, _18677_, _11039_);
  or _69478_ (_18679_, _18678_, _18674_);
  or _69479_ (_18680_, _18676_, _17733_);
  and _69480_ (_18681_, _18680_, _06541_);
  and _69481_ (_18682_, _18681_, _18679_);
  or _69482_ (_18683_, _11112_, _10863_);
  and _69483_ (_18684_, _18683_, _11113_);
  or _69484_ (_18685_, _18684_, _11097_);
  and _69485_ (_18686_, _18685_, _14297_);
  or _69486_ (_18687_, _18686_, _18682_);
  or _69487_ (_18688_, _11140_, _10545_);
  and _69488_ (_18689_, _18688_, _11141_);
  or _69489_ (_18690_, _18689_, _11127_);
  and _69490_ (_18691_, _18690_, _18687_);
  or _69491_ (_18692_, _18691_, _11125_);
  nand _69492_ (_18693_, _11125_, _06055_);
  and _69493_ (_18694_, _18693_, _11157_);
  and _69494_ (_18695_, _18694_, _18692_);
  nor _69495_ (_18696_, _11186_, _11170_);
  nor _69496_ (_18697_, _18696_, _11187_);
  and _69497_ (_18698_, _18697_, _18059_);
  or _69498_ (_18699_, _18698_, _11200_);
  or _69499_ (_18700_, _18699_, _18695_);
  and _69500_ (_18701_, _18700_, _18433_);
  or _69501_ (_18702_, _18701_, _11199_);
  or _69502_ (_18703_, _18432_, _18067_);
  and _69503_ (_18704_, _18703_, _13012_);
  and _69504_ (_18705_, _18704_, _18702_);
  or _69505_ (_18706_, _11313_, _11295_);
  and _69506_ (_18707_, _18706_, _11314_);
  and _69507_ (_18708_, _18707_, _11243_);
  or _69508_ (_18709_, _18708_, _11284_);
  or _69509_ (_18710_, _11270_, _11254_);
  and _69510_ (_18711_, _11271_, _06283_);
  and _69511_ (_18712_, _18711_, _18710_);
  or _69512_ (_18713_, _18712_, _18709_);
  or _69513_ (_18714_, _18713_, _18705_);
  nand _69514_ (_18715_, _11284_, _06055_);
  and _69515_ (_18716_, _18715_, _18714_);
  or _69516_ (_18717_, _18716_, _06568_);
  or _69517_ (_18718_, _18491_, _06926_);
  and _69518_ (_18719_, _18718_, _11331_);
  and _69519_ (_18720_, _18719_, _18717_);
  nor _69520_ (_18721_, _11337_, _10135_);
  or _69521_ (_18722_, _18721_, _11338_);
  and _69522_ (_18723_, _18722_, _11330_);
  or _69523_ (_18724_, _18723_, _11335_);
  or _69524_ (_18725_, _18724_, _18720_);
  nand _69525_ (_18726_, _11335_, _10170_);
  and _69526_ (_18727_, _18726_, _05928_);
  and _69527_ (_18728_, _18727_, _18725_);
  and _69528_ (_18729_, _18516_, _05927_);
  or _69529_ (_18730_, _18729_, _06278_);
  or _69530_ (_18731_, _18730_, _18728_);
  and _69531_ (_18732_, _15329_, _07939_);
  or _69532_ (_18733_, _18732_, _18442_);
  or _69533_ (_18734_, _18733_, _06279_);
  and _69534_ (_18735_, _18734_, _11354_);
  and _69535_ (_18736_, _18735_, _18731_);
  nor _69536_ (_18737_, _11363_, \oc8051_golden_model_1.ACC [4]);
  nor _69537_ (_18738_, _18737_, _11364_);
  and _69538_ (_18739_, _18738_, _11353_);
  or _69539_ (_18740_, _18739_, _11360_);
  or _69540_ (_18741_, _18740_, _18736_);
  nand _69541_ (_18742_, _11360_, _10170_);
  and _69542_ (_18743_, _18742_, _01347_);
  and _69543_ (_18744_, _18743_, _18741_);
  or _69544_ (_18745_, _18744_, _18430_);
  and _69545_ (_43166_, _18745_, _42618_);
  nor _69546_ (_18746_, _01347_, _10170_);
  and _69547_ (_18747_, _11058_, _10686_);
  nor _69548_ (_18748_, _18747_, _11059_);
  or _69549_ (_18749_, _18748_, _11037_);
  or _69550_ (_18750_, _11248_, _06543_);
  and _69551_ (_18752_, _18750_, _10497_);
  nand _69552_ (_18753_, _11210_, _10948_);
  or _69553_ (_18754_, _11166_, _06704_);
  and _69554_ (_18755_, _18754_, _17969_);
  and _69555_ (_18756_, _11166_, _06891_);
  nand _69556_ (_18757_, _06611_, _05974_);
  nor _69557_ (_18758_, _07939_, _10170_);
  nor _69558_ (_18759_, _08244_, _10490_);
  or _69559_ (_18760_, _18759_, _18758_);
  or _69560_ (_18761_, _18760_, _07215_);
  and _69561_ (_18762_, _06968_, \oc8051_golden_model_1.ACC [4]);
  nor _69562_ (_18763_, _18558_, _18762_);
  nor _69563_ (_18764_, _12600_, _18763_);
  and _69564_ (_18765_, _12600_, _18763_);
  nor _69565_ (_18766_, _18765_, _18764_);
  and _69566_ (_18767_, _18766_, \oc8051_golden_model_1.PSW [7]);
  nor _69567_ (_18768_, _18766_, \oc8051_golden_model_1.PSW [7]);
  nor _69568_ (_18769_, _18768_, _18767_);
  nor _69569_ (_18770_, _18565_, _18561_);
  not _69570_ (_18771_, _18770_);
  and _69571_ (_18774_, _18771_, _18769_);
  nor _69572_ (_18775_, _18771_, _18769_);
  nor _69573_ (_18776_, _18775_, _18774_);
  or _69574_ (_18777_, _18776_, _10517_);
  not _69575_ (_18778_, _10730_);
  and _69576_ (_18779_, _08541_, \oc8051_golden_model_1.ACC [4]);
  nor _69577_ (_18780_, _18464_, _18779_);
  nor _69578_ (_18781_, _11166_, _18780_);
  and _69579_ (_18782_, _11166_, _18780_);
  nor _69580_ (_18783_, _18782_, _18781_);
  and _69581_ (_18785_, _18783_, \oc8051_golden_model_1.PSW [7]);
  nor _69582_ (_18786_, _18783_, \oc8051_golden_model_1.PSW [7]);
  nor _69583_ (_18787_, _18786_, _18785_);
  nor _69584_ (_18788_, _18471_, _18467_);
  not _69585_ (_18789_, _18788_);
  and _69586_ (_18790_, _18789_, _18787_);
  nor _69587_ (_18791_, _18789_, _18787_);
  nor _69588_ (_18792_, _18791_, _18790_);
  or _69589_ (_18793_, _18792_, _18778_);
  nor _69590_ (_18794_, _08636_, _10170_);
  and _69591_ (_18796_, _15372_, _08636_);
  or _69592_ (_18797_, _18796_, _18794_);
  or _69593_ (_18798_, _18794_, _15387_);
  and _69594_ (_18799_, _18798_, _06261_);
  and _69595_ (_18800_, _18799_, _18797_);
  nand _69596_ (_18801_, _10744_, _08244_);
  nand _69597_ (_18802_, _10756_, _08244_);
  nor _69598_ (_18803_, _06781_, _10170_);
  and _69599_ (_18804_, _06781_, _10170_);
  nor _69600_ (_18805_, _18804_, _18803_);
  nand _69601_ (_18807_, _18805_, _10755_);
  and _69602_ (_18808_, _18807_, _10759_);
  and _69603_ (_18809_, _18808_, _18802_);
  and _69604_ (_18810_, _10758_, _09447_);
  or _69605_ (_18811_, _18810_, _18809_);
  and _69606_ (_18812_, _18811_, _10769_);
  and _69607_ (_18813_, _15358_, _07939_);
  or _69608_ (_18814_, _18813_, _18758_);
  and _69609_ (_18815_, _18814_, _06341_);
  or _69610_ (_18816_, _18815_, _10775_);
  or _69611_ (_18818_, _18816_, _18812_);
  nor _69612_ (_18819_, _10795_, _10787_);
  nand _69613_ (_18820_, _10795_, _10787_);
  nand _69614_ (_18821_, _18820_, _10775_);
  or _69615_ (_18822_, _18821_, _18819_);
  and _69616_ (_18823_, _18822_, _06466_);
  and _69617_ (_18824_, _18823_, _18818_);
  and _69618_ (_18825_, _18797_, _06272_);
  and _69619_ (_18826_, _18760_, _06461_);
  or _69620_ (_18827_, _18826_, _10744_);
  or _69621_ (_18829_, _18827_, _18825_);
  or _69622_ (_18830_, _18829_, _18824_);
  and _69623_ (_18831_, _18830_, _18801_);
  or _69624_ (_18832_, _18831_, _07174_);
  or _69625_ (_18833_, _09447_, _07175_);
  and _69626_ (_18834_, _18833_, _06465_);
  and _69627_ (_18835_, _18834_, _18832_);
  nor _69628_ (_18836_, _08246_, _06465_);
  or _69629_ (_18837_, _18836_, _10811_);
  or _69630_ (_18838_, _18837_, _18835_);
  nand _69631_ (_18840_, _10811_, _06042_);
  and _69632_ (_18841_, _18840_, _18838_);
  or _69633_ (_18842_, _18841_, _06268_);
  and _69634_ (_18843_, _15355_, _08636_);
  or _69635_ (_18844_, _18843_, _18794_);
  or _69636_ (_18845_, _18844_, _06269_);
  and _69637_ (_18846_, _18845_, _06262_);
  and _69638_ (_18847_, _18846_, _18842_);
  or _69639_ (_18848_, _18847_, _18800_);
  and _69640_ (_18849_, _18848_, _09537_);
  or _69641_ (_18851_, _10043_, _10041_);
  nor _69642_ (_18852_, _10044_, _09537_);
  and _69643_ (_18853_, _18852_, _18851_);
  or _69644_ (_18854_, _18853_, _10730_);
  or _69645_ (_18855_, _18854_, _18849_);
  and _69646_ (_18856_, _18855_, _18793_);
  or _69647_ (_18857_, _18856_, _17310_);
  not _69648_ (_18858_, _17310_);
  or _69649_ (_18859_, _18792_, _18858_);
  and _69650_ (_18860_, _18859_, _14204_);
  and _69651_ (_18862_, _18860_, _18857_);
  and _69652_ (_18863_, _18792_, _14203_);
  or _69653_ (_18864_, _18863_, _10656_);
  or _69654_ (_18865_, _18864_, _18862_);
  and _69655_ (_18866_, _09212_, \oc8051_golden_model_1.ACC [4]);
  nor _69656_ (_18867_, _18537_, _18866_);
  nor _69657_ (_18868_, _11210_, _18867_);
  and _69658_ (_18869_, _11210_, _18867_);
  nor _69659_ (_18870_, _18869_, _18868_);
  nor _69660_ (_18871_, _18870_, _10558_);
  and _69661_ (_18873_, _18870_, _10558_);
  nor _69662_ (_18874_, _18873_, _18871_);
  nor _69663_ (_18875_, _18543_, _18540_);
  not _69664_ (_18876_, _18875_);
  and _69665_ (_18877_, _18876_, _18874_);
  nor _69666_ (_18878_, _18876_, _18874_);
  nor _69667_ (_18879_, _18878_, _18877_);
  or _69668_ (_18880_, _18879_, _10588_);
  and _69669_ (_18881_, _18880_, _06517_);
  and _69670_ (_18882_, _18881_, _18865_);
  and _69671_ (_18884_, _08543_, \oc8051_golden_model_1.ACC [4]);
  nor _69672_ (_18885_, _18449_, _18884_);
  nor _69673_ (_18886_, _11250_, _18885_);
  and _69674_ (_18887_, _11250_, _18885_);
  nor _69675_ (_18888_, _18887_, _18886_);
  and _69676_ (_18889_, _18888_, \oc8051_golden_model_1.PSW [7]);
  nor _69677_ (_18890_, _18888_, \oc8051_golden_model_1.PSW [7]);
  nor _69678_ (_18891_, _18890_, _18889_);
  nor _69679_ (_18892_, _18456_, _18452_);
  not _69680_ (_18893_, _18892_);
  and _69681_ (_18895_, _18893_, _18891_);
  nor _69682_ (_18896_, _18893_, _18891_);
  nor _69683_ (_18897_, _18896_, _18895_);
  or _69684_ (_18898_, _18897_, _10516_);
  and _69685_ (_18899_, _18898_, _12644_);
  or _69686_ (_18900_, _18899_, _18882_);
  and _69687_ (_18901_, _18900_, _18777_);
  or _69688_ (_18902_, _18901_, _10515_);
  nand _69689_ (_18903_, _06611_, _10515_);
  and _69690_ (_18904_, _18903_, _06258_);
  and _69691_ (_18906_, _18904_, _18902_);
  or _69692_ (_18907_, _18794_, _15403_);
  and _69693_ (_18908_, _18907_, _06257_);
  and _69694_ (_18909_, _18908_, _18797_);
  or _69695_ (_18910_, _18909_, _10080_);
  or _69696_ (_18911_, _18910_, _18906_);
  and _69697_ (_18912_, _18911_, _18761_);
  or _69698_ (_18913_, _18912_, _07460_);
  and _69699_ (_18914_, _09447_, _07939_);
  or _69700_ (_18915_, _18758_, _07208_);
  or _69701_ (_18917_, _18915_, _18914_);
  and _69702_ (_18918_, _18917_, _05982_);
  and _69703_ (_18919_, _18918_, _18913_);
  and _69704_ (_18920_, _15459_, _07939_);
  or _69705_ (_18921_, _18920_, _18758_);
  and _69706_ (_18922_, _18921_, _10094_);
  or _69707_ (_18923_, _18922_, _10093_);
  or _69708_ (_18924_, _18923_, _18919_);
  or _69709_ (_18925_, _10153_, _10100_);
  and _69710_ (_18926_, _18925_, _18924_);
  or _69711_ (_18927_, _18926_, _05974_);
  and _69712_ (_18928_, _18927_, _18757_);
  or _69713_ (_18929_, _18928_, _06218_);
  and _69714_ (_18930_, _08946_, _07939_);
  or _69715_ (_18931_, _18930_, _18758_);
  or _69716_ (_18932_, _18931_, _06219_);
  and _69717_ (_18933_, _18932_, _10930_);
  and _69718_ (_18934_, _18933_, _18929_);
  nor _69719_ (_18935_, _10930_, _06611_);
  or _69720_ (_18936_, _18935_, _18277_);
  or _69721_ (_18938_, _18936_, _18934_);
  or _69722_ (_18939_, _11166_, _18603_);
  and _69723_ (_18940_, _18939_, _18607_);
  and _69724_ (_18941_, _18940_, _18938_);
  or _69725_ (_18942_, _18941_, _18756_);
  and _69726_ (_18943_, _18942_, _06745_);
  and _69727_ (_18944_, _11166_, _06744_);
  or _69728_ (_18945_, _18944_, _06703_);
  or _69729_ (_18946_, _18945_, _18943_);
  and _69730_ (_18947_, _18946_, _18755_);
  and _69731_ (_18949_, _11166_, _10506_);
  or _69732_ (_18950_, _18949_, _06887_);
  or _69733_ (_18951_, _18950_, _18947_);
  not _69734_ (_18952_, _06887_);
  or _69735_ (_18953_, _11166_, _18952_);
  and _69736_ (_18954_, _18953_, _10946_);
  and _69737_ (_18955_, _18954_, _18951_);
  and _69738_ (_18956_, _10945_, _11166_);
  or _69739_ (_18957_, _18956_, _10948_);
  or _69740_ (_18958_, _18957_, _18955_);
  and _69741_ (_18960_, _18958_, _18753_);
  or _69742_ (_18961_, _18960_, _06533_);
  or _69743_ (_18962_, _11250_, _06534_);
  and _69744_ (_18963_, _18962_, _10955_);
  and _69745_ (_18964_, _18963_, _18961_);
  and _69746_ (_18965_, _10954_, _12600_);
  or _69747_ (_18966_, _18965_, _06369_);
  or _69748_ (_18967_, _18966_, _18964_);
  and _69749_ (_18968_, _15353_, _07939_);
  or _69750_ (_18969_, _18968_, _18758_);
  or _69751_ (_18971_, _18969_, _07237_);
  and _69752_ (_18972_, _18971_, _18967_);
  or _69753_ (_18973_, _18972_, _06536_);
  and _69754_ (_18974_, _11032_, _07211_);
  or _69755_ (_18975_, _18974_, _05960_);
  or _69756_ (_18976_, _18758_, _07240_);
  and _69757_ (_18977_, _18976_, _18975_);
  and _69758_ (_18978_, _18977_, _18973_);
  and _69759_ (_18979_, _10987_, _11164_);
  or _69760_ (_18980_, _18979_, _18978_);
  nand _69761_ (_18982_, _10732_, _06544_);
  or _69762_ (_18983_, _18982_, _11164_);
  and _69763_ (_18984_, _18983_, _17401_);
  and _69764_ (_18985_, _18984_, _18980_);
  and _69765_ (_18986_, _10983_, _11208_);
  or _69766_ (_18987_, _18986_, _06542_);
  or _69767_ (_18988_, _18987_, _18985_);
  and _69768_ (_18989_, _18988_, _18752_);
  and _69769_ (_18990_, _11290_, _10496_);
  or _69770_ (_18991_, _18990_, _18989_);
  and _69771_ (_18993_, _18991_, _07242_);
  nand _69772_ (_18994_, _18931_, _06375_);
  nor _69773_ (_18995_, _18994_, _11249_);
  or _69774_ (_18996_, _18995_, _17507_);
  or _69775_ (_18997_, _18996_, _18993_);
  nand _69776_ (_18998_, _17507_, _11165_);
  and _69777_ (_18999_, _18998_, _18997_);
  or _69778_ (_19000_, _18999_, _17506_);
  nand _69779_ (_19001_, _17506_, _11165_);
  and _69780_ (_19002_, _19001_, _17430_);
  and _69781_ (_19004_, _19002_, _19000_);
  nor _69782_ (_19005_, _11165_, _17430_);
  or _69783_ (_19006_, _19005_, _11014_);
  or _69784_ (_19007_, _19006_, _19004_);
  or _69785_ (_19008_, _11013_, \oc8051_golden_model_1.ACC [5]);
  or _69786_ (_19009_, _19008_, _09447_);
  and _69787_ (_19010_, _19009_, _06531_);
  and _69788_ (_19011_, _19010_, _19007_);
  nand _69789_ (_19012_, _11024_, _11249_);
  and _69790_ (_19013_, _19012_, _11023_);
  or _69791_ (_19015_, _19013_, _19011_);
  nand _69792_ (_19016_, _11021_, _11291_);
  and _69793_ (_19017_, _19016_, _09056_);
  and _69794_ (_19018_, _19017_, _19015_);
  and _69795_ (_19019_, _15350_, _07939_);
  or _69796_ (_19020_, _19019_, _18758_);
  and _69797_ (_19021_, _19020_, _06366_);
  or _69798_ (_19022_, _19021_, _14283_);
  or _69799_ (_19023_, _19022_, _19018_);
  and _69800_ (_19024_, _19023_, _18749_);
  or _69801_ (_19026_, _19024_, _11041_);
  and _69802_ (_19027_, _11086_, _10610_);
  nor _69803_ (_19028_, _19027_, _11087_);
  or _69804_ (_19029_, _19028_, _11069_);
  and _69805_ (_19030_, _19029_, _06541_);
  and _69806_ (_19031_, _19030_, _19026_);
  nand _69807_ (_19032_, _11114_, _10860_);
  nor _69808_ (_19033_, _11115_, _06541_);
  and _69809_ (_19034_, _19033_, _19032_);
  or _69810_ (_19035_, _19034_, _11097_);
  or _69811_ (_19037_, _19035_, _19031_);
  and _69812_ (_19038_, _11142_, _10542_);
  nor _69813_ (_19039_, _19038_, _11143_);
  or _69814_ (_19040_, _19039_, _11127_);
  and _69815_ (_19041_, _19040_, _11126_);
  and _69816_ (_19042_, _19041_, _19037_);
  nand _69817_ (_19043_, _11125_, \oc8051_golden_model_1.ACC [4]);
  nand _69818_ (_19044_, _19043_, _12151_);
  or _69819_ (_19045_, _19044_, _19042_);
  and _69820_ (_19046_, _11232_, _11210_);
  nor _69821_ (_19048_, _19046_, _11233_);
  or _69822_ (_19049_, _19048_, _11203_);
  nor _69823_ (_19050_, _11189_, _11166_);
  nor _69824_ (_19051_, _19050_, _11190_);
  or _69825_ (_19052_, _19051_, _11157_);
  and _69826_ (_19053_, _19052_, _06285_);
  and _69827_ (_19054_, _19053_, _19049_);
  and _69828_ (_19055_, _19054_, _19045_);
  not _69829_ (_19056_, _13012_);
  nor _69830_ (_19057_, _11273_, _11250_);
  nor _69831_ (_19059_, _19057_, _11274_);
  or _69832_ (_19060_, _19059_, _11243_);
  and _69833_ (_19061_, _19060_, _19056_);
  or _69834_ (_19062_, _19061_, _19055_);
  and _69835_ (_19063_, _11315_, _12600_);
  nor _69836_ (_19064_, _11315_, _12600_);
  or _69837_ (_19065_, _19064_, _11321_);
  or _69838_ (_19066_, _19065_, _19063_);
  and _69839_ (_19067_, _19066_, _11285_);
  and _69840_ (_19068_, _19067_, _19062_);
  and _69841_ (_19070_, _11284_, \oc8051_golden_model_1.ACC [4]);
  or _69842_ (_19071_, _19070_, _06568_);
  or _69843_ (_19072_, _19071_, _19068_);
  or _69844_ (_19073_, _18814_, _06926_);
  and _69845_ (_19074_, _19073_, _11331_);
  and _69846_ (_19075_, _19074_, _19072_);
  nor _69847_ (_19076_, _11338_, _10170_);
  or _69848_ (_19077_, _19076_, _11339_);
  and _69849_ (_19078_, _19077_, _11330_);
  or _69850_ (_19079_, _19078_, _11335_);
  or _69851_ (_19081_, _19079_, _19075_);
  nand _69852_ (_19082_, _11335_, _10116_);
  and _69853_ (_19083_, _19082_, _05928_);
  and _69854_ (_19084_, _19083_, _19081_);
  and _69855_ (_19085_, _18844_, _05927_);
  or _69856_ (_19086_, _19085_, _06278_);
  or _69857_ (_19087_, _19086_, _19084_);
  and _69858_ (_19088_, _15532_, _07939_);
  or _69859_ (_19089_, _19088_, _18758_);
  or _69860_ (_19090_, _19089_, _06279_);
  and _69861_ (_19092_, _19090_, _11354_);
  and _69862_ (_19093_, _19092_, _19087_);
  nor _69863_ (_19094_, _11364_, \oc8051_golden_model_1.ACC [5]);
  nor _69864_ (_19095_, _19094_, _11365_);
  and _69865_ (_19096_, _19095_, _11353_);
  or _69866_ (_19097_, _19096_, _11360_);
  or _69867_ (_19098_, _19097_, _19093_);
  nand _69868_ (_19099_, _11360_, _10116_);
  and _69869_ (_19100_, _19099_, _01347_);
  and _69870_ (_19101_, _19100_, _19098_);
  or _69871_ (_19103_, _19101_, _18746_);
  and _69872_ (_43167_, _19103_, _42618_);
  nor _69873_ (_19104_, _01347_, _10116_);
  or _69874_ (_19105_, _11116_, _10893_);
  and _69875_ (_19106_, _11117_, _06540_);
  and _69876_ (_19107_, _19106_, _19105_);
  nand _69877_ (_19108_, _11021_, _11288_);
  or _69878_ (_19109_, _17401_, _11204_);
  or _69879_ (_19110_, _11207_, _10502_);
  nor _69880_ (_19111_, _07939_, _10116_);
  and _69881_ (_19113_, _15657_, _07939_);
  or _69882_ (_19114_, _19113_, _19111_);
  and _69883_ (_19115_, _19114_, _10094_);
  nor _69884_ (_19116_, _08142_, _10490_);
  or _69885_ (_19117_, _19116_, _19111_);
  or _69886_ (_19118_, _19117_, _07215_);
  or _69887_ (_19119_, _09447_, _10170_);
  and _69888_ (_19120_, _09447_, _10170_);
  or _69889_ (_19121_, _18867_, _19120_);
  and _69890_ (_19122_, _19121_, _19119_);
  nor _69891_ (_19124_, _19122_, _11207_);
  and _69892_ (_19125_, _19122_, _11207_);
  nor _69893_ (_19126_, _19125_, _19124_);
  nor _69894_ (_19127_, _18877_, _18871_);
  and _69895_ (_19128_, _19127_, \oc8051_golden_model_1.PSW [7]);
  or _69896_ (_19129_, _19128_, _19126_);
  nand _69897_ (_19130_, _19128_, _19126_);
  and _69898_ (_19131_, _19130_, _19129_);
  or _69899_ (_19132_, _19131_, _10588_);
  nand _69900_ (_19133_, _10744_, _08142_);
  nand _69901_ (_19135_, _10756_, _08142_);
  nor _69902_ (_19136_, _06781_, _10116_);
  and _69903_ (_19137_, _06781_, _10116_);
  nor _69904_ (_19138_, _19137_, _19136_);
  nand _69905_ (_19139_, _19138_, _10755_);
  and _69906_ (_19140_, _19139_, _10759_);
  and _69907_ (_19141_, _19140_, _19135_);
  and _69908_ (_19142_, _10758_, _09446_);
  or _69909_ (_19143_, _19142_, _19141_);
  and _69910_ (_19144_, _19143_, _10769_);
  and _69911_ (_19146_, _15554_, _07939_);
  or _69912_ (_19147_, _19146_, _19111_);
  and _69913_ (_19148_, _19147_, _06341_);
  or _69914_ (_19149_, _19148_, _10775_);
  or _69915_ (_19150_, _19149_, _19144_);
  not _69916_ (_19151_, _18819_);
  nor _69917_ (_19152_, _19151_, _10789_);
  and _69918_ (_19153_, _19151_, _10789_);
  or _69919_ (_19154_, _19153_, _19152_);
  or _69920_ (_19155_, _19154_, _10776_);
  and _69921_ (_19157_, _19155_, _06466_);
  and _69922_ (_19158_, _19157_, _19150_);
  nor _69923_ (_19159_, _08636_, _10116_);
  and _69924_ (_19160_, _15570_, _08636_);
  or _69925_ (_19161_, _19160_, _19159_);
  and _69926_ (_19162_, _19161_, _06272_);
  and _69927_ (_19163_, _19117_, _06461_);
  or _69928_ (_19164_, _19163_, _10744_);
  or _69929_ (_19165_, _19164_, _19162_);
  or _69930_ (_19166_, _19165_, _19158_);
  and _69931_ (_19168_, _19166_, _19133_);
  or _69932_ (_19169_, _19168_, _07174_);
  or _69933_ (_19170_, _09446_, _07175_);
  and _69934_ (_19171_, _19170_, _06465_);
  and _69935_ (_19172_, _19171_, _19169_);
  nor _69936_ (_19173_, _08144_, _06465_);
  or _69937_ (_19174_, _19173_, _10811_);
  or _69938_ (_19175_, _19174_, _19172_);
  nand _69939_ (_19176_, _10811_, _10213_);
  and _69940_ (_19177_, _19176_, _19175_);
  or _69941_ (_19179_, _19177_, _06268_);
  and _69942_ (_19180_, _15551_, _08636_);
  or _69943_ (_19181_, _19180_, _19159_);
  or _69944_ (_19182_, _19181_, _06269_);
  and _69945_ (_19183_, _19182_, _06262_);
  and _69946_ (_19184_, _19183_, _19179_);
  or _69947_ (_19185_, _19159_, _15585_);
  and _69948_ (_19186_, _19185_, _06261_);
  and _69949_ (_19187_, _19186_, _19161_);
  or _69950_ (_19188_, _19187_, _09531_);
  or _69951_ (_19190_, _19188_, _19184_);
  nor _69952_ (_19191_, _10046_, _10044_);
  nor _69953_ (_19192_, _19191_, _10047_);
  or _69954_ (_19193_, _19192_, _09537_);
  and _69955_ (_19194_, _19193_, _10735_);
  and _69956_ (_19195_, _19194_, _19190_);
  nand _69957_ (_19196_, _08244_, \oc8051_golden_model_1.ACC [5]);
  nor _69958_ (_19197_, _08244_, \oc8051_golden_model_1.ACC [5]);
  or _69959_ (_19198_, _18780_, _19197_);
  and _69960_ (_19199_, _19198_, _19196_);
  nor _69961_ (_19201_, _19199_, _11163_);
  and _69962_ (_19202_, _19199_, _11163_);
  nor _69963_ (_19203_, _19202_, _19201_);
  nor _69964_ (_19204_, _18790_, _18785_);
  and _69965_ (_19205_, _19204_, \oc8051_golden_model_1.PSW [7]);
  or _69966_ (_19206_, _19205_, _19203_);
  nand _69967_ (_19207_, _19205_, _19203_);
  and _69968_ (_19208_, _19207_, _10737_);
  and _69969_ (_19209_, _19208_, _19206_);
  or _69970_ (_19210_, _19209_, _10656_);
  or _69971_ (_19212_, _19210_, _19195_);
  and _69972_ (_19213_, _19212_, _06517_);
  and _69973_ (_19214_, _19213_, _19132_);
  or _69974_ (_19215_, _18885_, _14129_);
  and _69975_ (_19216_, _19215_, _14128_);
  nor _69976_ (_19217_, _19216_, _11247_);
  and _69977_ (_19218_, _19216_, _11247_);
  nor _69978_ (_19219_, _19218_, _19217_);
  nor _69979_ (_19220_, _18895_, _18889_);
  and _69980_ (_19221_, _19220_, \oc8051_golden_model_1.PSW [7]);
  nand _69981_ (_19223_, _19221_, _19219_);
  or _69982_ (_19224_, _19221_, _19219_);
  and _69983_ (_19225_, _19224_, _06512_);
  and _69984_ (_19226_, _19225_, _19223_);
  or _69985_ (_19227_, _19226_, _19214_);
  and _69986_ (_19228_, _19227_, _10517_);
  or _69987_ (_19229_, _18763_, _14168_);
  and _69988_ (_19230_, _19229_, _14167_);
  nor _69989_ (_19231_, _19230_, _11289_);
  and _69990_ (_19232_, _19230_, _11289_);
  nor _69991_ (_19234_, _19232_, _19231_);
  nor _69992_ (_19235_, _18774_, _18767_);
  and _69993_ (_19236_, _19235_, \oc8051_golden_model_1.PSW [7]);
  or _69994_ (_19237_, _19236_, _19234_);
  nand _69995_ (_19238_, _19236_, _19234_);
  and _69996_ (_19239_, _19238_, _10516_);
  and _69997_ (_19240_, _19239_, _19237_);
  or _69998_ (_19241_, _19240_, _10515_);
  or _69999_ (_19242_, _19241_, _19228_);
  nand _70000_ (_19243_, _06317_, _10515_);
  and _70001_ (_19245_, _19243_, _06258_);
  and _70002_ (_19246_, _19245_, _19242_);
  and _70003_ (_19247_, _15602_, _08636_);
  or _70004_ (_19248_, _19247_, _19159_);
  and _70005_ (_19249_, _19248_, _06257_);
  or _70006_ (_19250_, _19249_, _10080_);
  or _70007_ (_19251_, _19250_, _19246_);
  and _70008_ (_19252_, _19251_, _19118_);
  or _70009_ (_19253_, _19252_, _07460_);
  and _70010_ (_19254_, _09446_, _07939_);
  or _70011_ (_19256_, _19111_, _07208_);
  or _70012_ (_19257_, _19256_, _19254_);
  and _70013_ (_19258_, _19257_, _05982_);
  and _70014_ (_19259_, _19258_, _19253_);
  or _70015_ (_19260_, _19259_, _19115_);
  and _70016_ (_19261_, _19260_, _12172_);
  nor _70017_ (_19262_, _06317_, _05975_);
  not _70018_ (_19263_, _10122_);
  nor _70019_ (_19264_, _19263_, _10117_);
  and _70020_ (_19265_, _19264_, _05973_);
  and _70021_ (_19267_, _19265_, _10093_);
  or _70022_ (_19268_, _19267_, _19262_);
  or _70023_ (_19269_, _19268_, _19261_);
  and _70024_ (_19270_, _19269_, _06219_);
  and _70025_ (_19271_, _15664_, _07939_);
  or _70026_ (_19272_, _19271_, _19111_);
  and _70027_ (_19273_, _19272_, _06218_);
  or _70028_ (_19274_, _19273_, _10929_);
  or _70029_ (_19275_, _19274_, _19270_);
  nand _70030_ (_19276_, _10929_, _06317_);
  and _70031_ (_19278_, _19276_, _17962_);
  and _70032_ (_19279_, _19278_, _19275_);
  and _70033_ (_19280_, _17965_, _11163_);
  or _70034_ (_19281_, _19280_, _10506_);
  or _70035_ (_19282_, _19281_, _19279_);
  or _70036_ (_19283_, _11163_, _17969_);
  and _70037_ (_19284_, _19283_, _18952_);
  and _70038_ (_19285_, _19284_, _19282_);
  or _70039_ (_19286_, _17511_, _11163_);
  and _70040_ (_19287_, _19286_, _18286_);
  or _70041_ (_19289_, _19287_, _19285_);
  or _70042_ (_19290_, _17512_, _11163_);
  and _70043_ (_19291_, _19290_, _17510_);
  and _70044_ (_19292_, _19291_, _19289_);
  and _70045_ (_19293_, _11163_, _06888_);
  or _70046_ (_19294_, _19293_, _10948_);
  or _70047_ (_19295_, _19294_, _19292_);
  and _70048_ (_19296_, _19295_, _19110_);
  or _70049_ (_19297_, _19296_, _06533_);
  or _70050_ (_19298_, _11247_, _06534_);
  and _70051_ (_19300_, _19298_, _10955_);
  and _70052_ (_19301_, _19300_, _19297_);
  and _70053_ (_19302_, _10954_, _11289_);
  or _70054_ (_19303_, _19302_, _06369_);
  or _70055_ (_19304_, _19303_, _19301_);
  and _70056_ (_19305_, _15549_, _07939_);
  or _70057_ (_19306_, _19305_, _19111_);
  or _70058_ (_19307_, _19306_, _07237_);
  and _70059_ (_19308_, _19307_, _19304_);
  or _70060_ (_19309_, _19308_, _06536_);
  or _70061_ (_19311_, _19111_, _07240_);
  and _70062_ (_19312_, _19311_, _10986_);
  and _70063_ (_19313_, _19312_, _19309_);
  and _70064_ (_19314_, _10987_, _11160_);
  or _70065_ (_19315_, _19314_, _10983_);
  or _70066_ (_19316_, _19315_, _19313_);
  and _70067_ (_19317_, _19316_, _19109_);
  or _70068_ (_19318_, _19317_, _06542_);
  or _70069_ (_19319_, _11244_, _06543_);
  and _70070_ (_19320_, _19319_, _10497_);
  and _70071_ (_19322_, _19320_, _19318_);
  and _70072_ (_19323_, _11286_, _10496_);
  or _70073_ (_19324_, _19323_, _19322_);
  and _70074_ (_19325_, _19324_, _07242_);
  and _70075_ (_19326_, _10998_, _07043_);
  nand _70076_ (_19327_, _19272_, _06375_);
  or _70077_ (_19328_, _19327_, _11246_);
  nand _70078_ (_19329_, _19328_, _19326_);
  or _70079_ (_19330_, _19329_, _19325_);
  or _70080_ (_19331_, _19326_, _11162_);
  and _70081_ (_19333_, _19331_, _11009_);
  and _70082_ (_19334_, _19333_, _19330_);
  and _70083_ (_19335_, _11008_, _11162_);
  or _70084_ (_19336_, _19335_, _11014_);
  or _70085_ (_19337_, _19336_, _19334_);
  or _70086_ (_19338_, _11013_, _11205_);
  and _70087_ (_19339_, _19338_, _06531_);
  and _70088_ (_19340_, _19339_, _19337_);
  nand _70089_ (_19341_, _11024_, _11246_);
  and _70090_ (_19342_, _19341_, _11023_);
  or _70091_ (_19344_, _19342_, _19340_);
  and _70092_ (_19345_, _19344_, _19108_);
  or _70093_ (_19346_, _19345_, _06366_);
  and _70094_ (_19347_, _15546_, _07939_);
  or _70095_ (_19348_, _19111_, _09056_);
  or _70096_ (_19349_, _19348_, _19347_);
  and _70097_ (_19350_, _19349_, _11037_);
  and _70098_ (_19351_, _19350_, _19346_);
  nor _70099_ (_19352_, _11060_, _10722_);
  nor _70100_ (_19353_, _19352_, _11061_);
  and _70101_ (_19355_, _19353_, _14283_);
  or _70102_ (_19356_, _19355_, _11041_);
  or _70103_ (_19357_, _19356_, _19351_);
  or _70104_ (_19358_, _11088_, _10649_);
  and _70105_ (_19359_, _19358_, _11089_);
  or _70106_ (_19360_, _19359_, _11069_);
  and _70107_ (_19361_, _19360_, _06541_);
  and _70108_ (_19362_, _19361_, _19357_);
  or _70109_ (_19363_, _19362_, _19107_);
  and _70110_ (_19364_, _19363_, _11127_);
  or _70111_ (_19366_, _11144_, _10579_);
  nor _70112_ (_19367_, _11145_, _11127_);
  and _70113_ (_19368_, _19367_, _19366_);
  or _70114_ (_19369_, _19368_, _11125_);
  or _70115_ (_19370_, _19369_, _19364_);
  nand _70116_ (_19371_, _11125_, _10170_);
  and _70117_ (_19372_, _19371_, _11157_);
  and _70118_ (_19373_, _19372_, _19370_);
  nor _70119_ (_19374_, _11191_, _11163_);
  nor _70120_ (_19375_, _19374_, _11192_);
  and _70121_ (_19377_, _19375_, _18059_);
  or _70122_ (_19378_, _19377_, _11201_);
  or _70123_ (_19379_, _19378_, _19373_);
  nor _70124_ (_19380_, _11234_, _11207_);
  nor _70125_ (_19381_, _19380_, _11235_);
  or _70126_ (_19382_, _19381_, _11203_);
  and _70127_ (_19383_, _19382_, _06285_);
  and _70128_ (_19384_, _19383_, _19379_);
  or _70129_ (_19385_, _11275_, _11247_);
  and _70130_ (_19386_, _19385_, _11276_);
  or _70131_ (_19388_, _19386_, _11243_);
  and _70132_ (_19389_, _19388_, _19056_);
  or _70133_ (_19390_, _19389_, _19384_);
  or _70134_ (_19391_, _11317_, _11289_);
  and _70135_ (_19392_, _19391_, _11318_);
  or _70136_ (_19393_, _19392_, _11321_);
  and _70137_ (_19394_, _19393_, _11285_);
  and _70138_ (_19395_, _19394_, _19390_);
  and _70139_ (_19396_, _11284_, \oc8051_golden_model_1.ACC [5]);
  or _70140_ (_19397_, _19396_, _06568_);
  or _70141_ (_19399_, _19397_, _19395_);
  or _70142_ (_19400_, _19147_, _06926_);
  and _70143_ (_19401_, _19400_, _11331_);
  and _70144_ (_19402_, _19401_, _19399_);
  nor _70145_ (_19403_, _11339_, _10116_);
  or _70146_ (_19404_, _19403_, _11340_);
  and _70147_ (_19405_, _19404_, _11330_);
  or _70148_ (_19406_, _19405_, _11335_);
  or _70149_ (_19407_, _19406_, _19402_);
  nand _70150_ (_19408_, _11335_, _08572_);
  and _70151_ (_19410_, _19408_, _05928_);
  and _70152_ (_19411_, _19410_, _19407_);
  and _70153_ (_19412_, _19181_, _05927_);
  or _70154_ (_19413_, _19412_, _06278_);
  or _70155_ (_19414_, _19413_, _19411_);
  and _70156_ (_19415_, _15734_, _07939_);
  or _70157_ (_19416_, _19415_, _19111_);
  or _70158_ (_19417_, _19416_, _06279_);
  and _70159_ (_19418_, _19417_, _11354_);
  and _70160_ (_19419_, _19418_, _19414_);
  nor _70161_ (_19421_, _11365_, \oc8051_golden_model_1.ACC [6]);
  nor _70162_ (_19422_, _19421_, _11366_);
  and _70163_ (_19423_, _19422_, _11353_);
  or _70164_ (_19424_, _19423_, _11360_);
  or _70165_ (_19425_, _19424_, _19419_);
  nand _70166_ (_19426_, _11360_, _08572_);
  and _70167_ (_19427_, _19426_, _01347_);
  and _70168_ (_19428_, _19427_, _19425_);
  or _70169_ (_19429_, _19428_, _19104_);
  and _70170_ (_43168_, _19429_, _42618_);
  not _70171_ (_19431_, \oc8051_golden_model_1.PCON [0]);
  nor _70172_ (_19432_, _01347_, _19431_);
  nand _70173_ (_19433_, _11263_, _07951_);
  nor _70174_ (_19434_, _07951_, _19431_);
  nor _70175_ (_19435_, _19434_, _07234_);
  nand _70176_ (_19436_, _19435_, _19433_);
  and _70177_ (_19437_, _07951_, _07133_);
  or _70178_ (_19438_, _19437_, _19434_);
  or _70179_ (_19439_, _19438_, _07215_);
  nor _70180_ (_19440_, _08390_, _11380_);
  or _70181_ (_19442_, _19440_, _19434_);
  or _70182_ (_19443_, _19442_, _07151_);
  and _70183_ (_19444_, _07951_, \oc8051_golden_model_1.ACC [0]);
  or _70184_ (_19445_, _19444_, _19434_);
  and _70185_ (_19446_, _19445_, _07141_);
  nor _70186_ (_19447_, _07141_, _19431_);
  or _70187_ (_19448_, _19447_, _06341_);
  or _70188_ (_19449_, _19448_, _19446_);
  and _70189_ (_19450_, _19449_, _07166_);
  and _70190_ (_19451_, _19450_, _19443_);
  and _70191_ (_19453_, _19438_, _06461_);
  or _70192_ (_19454_, _19453_, _19451_);
  and _70193_ (_19455_, _19454_, _06465_);
  and _70194_ (_19456_, _19445_, _06464_);
  or _70195_ (_19457_, _19456_, _10080_);
  or _70196_ (_19458_, _19457_, _19455_);
  and _70197_ (_19459_, _19458_, _19439_);
  or _70198_ (_19460_, _19459_, _07460_);
  and _70199_ (_19461_, _09392_, _07951_);
  or _70200_ (_19462_, _19434_, _07208_);
  or _70201_ (_19464_, _19462_, _19461_);
  and _70202_ (_19465_, _19464_, _19460_);
  or _70203_ (_19466_, _19465_, _10094_);
  and _70204_ (_19467_, _14467_, _07951_);
  or _70205_ (_19468_, _19434_, _05982_);
  or _70206_ (_19469_, _19468_, _19467_);
  and _70207_ (_19470_, _19469_, _06219_);
  and _70208_ (_19471_, _19470_, _19466_);
  and _70209_ (_19472_, _07951_, _08954_);
  or _70210_ (_19473_, _19472_, _19434_);
  and _70211_ (_19475_, _19473_, _06218_);
  or _70212_ (_19476_, _19475_, _06369_);
  or _70213_ (_19477_, _19476_, _19471_);
  and _70214_ (_19478_, _14366_, _07951_);
  or _70215_ (_19479_, _19478_, _19434_);
  or _70216_ (_19480_, _19479_, _07237_);
  and _70217_ (_19481_, _19480_, _07240_);
  and _70218_ (_19482_, _19481_, _19477_);
  nor _70219_ (_19483_, _12580_, _11380_);
  or _70220_ (_19484_, _19483_, _19434_);
  and _70221_ (_19486_, _19433_, _06536_);
  and _70222_ (_19487_, _19486_, _19484_);
  or _70223_ (_19488_, _19487_, _19482_);
  and _70224_ (_19489_, _19488_, _07242_);
  nand _70225_ (_19490_, _19473_, _06375_);
  nor _70226_ (_19491_, _19490_, _19440_);
  or _70227_ (_19492_, _19491_, _06545_);
  or _70228_ (_19493_, _19492_, _19489_);
  and _70229_ (_19494_, _19493_, _19436_);
  or _70230_ (_19495_, _19494_, _06366_);
  and _70231_ (_19497_, _14363_, _07951_);
  or _70232_ (_19498_, _19497_, _19434_);
  or _70233_ (_19499_, _19498_, _09056_);
  and _70234_ (_19500_, _19499_, _09061_);
  and _70235_ (_19501_, _19500_, _19495_);
  not _70236_ (_19502_, _06661_);
  and _70237_ (_19503_, _19484_, _06528_);
  or _70238_ (_19504_, _19503_, _19502_);
  or _70239_ (_19505_, _19504_, _19501_);
  or _70240_ (_19506_, _19442_, _06661_);
  and _70241_ (_19508_, _19506_, _01347_);
  and _70242_ (_19509_, _19508_, _19505_);
  or _70243_ (_19510_, _19509_, _19432_);
  and _70244_ (_43170_, _19510_, _42618_);
  not _70245_ (_19511_, \oc8051_golden_model_1.PCON [1]);
  nor _70246_ (_19512_, _01347_, _19511_);
  nand _70247_ (_19513_, _07951_, _07038_);
  or _70248_ (_19514_, _07951_, \oc8051_golden_model_1.PCON [1]);
  and _70249_ (_19515_, _19514_, _06218_);
  and _70250_ (_19516_, _19515_, _19513_);
  nor _70251_ (_19518_, _07951_, _19511_);
  nor _70252_ (_19519_, _11380_, _07357_);
  or _70253_ (_19520_, _19519_, _19518_);
  or _70254_ (_19521_, _19520_, _07215_);
  and _70255_ (_19522_, _14562_, _07951_);
  not _70256_ (_19523_, _19522_);
  and _70257_ (_19524_, _19523_, _19514_);
  or _70258_ (_19525_, _19524_, _07151_);
  and _70259_ (_19526_, _07951_, \oc8051_golden_model_1.ACC [1]);
  or _70260_ (_19527_, _19526_, _19518_);
  and _70261_ (_19529_, _19527_, _07141_);
  nor _70262_ (_19530_, _07141_, _19511_);
  or _70263_ (_19531_, _19530_, _06341_);
  or _70264_ (_19532_, _19531_, _19529_);
  and _70265_ (_19533_, _19532_, _07166_);
  and _70266_ (_19534_, _19533_, _19525_);
  and _70267_ (_19535_, _19520_, _06461_);
  or _70268_ (_19536_, _19535_, _19534_);
  and _70269_ (_19537_, _19536_, _06465_);
  and _70270_ (_19538_, _19527_, _06464_);
  or _70271_ (_19540_, _19538_, _10080_);
  or _70272_ (_19541_, _19540_, _19537_);
  and _70273_ (_19542_, _19541_, _19521_);
  or _70274_ (_19543_, _19542_, _07460_);
  and _70275_ (_19544_, _09451_, _07951_);
  or _70276_ (_19545_, _19518_, _07208_);
  or _70277_ (_19546_, _19545_, _19544_);
  and _70278_ (_19547_, _19546_, _05982_);
  and _70279_ (_19548_, _19547_, _19543_);
  or _70280_ (_19549_, _14653_, _11380_);
  and _70281_ (_19551_, _19514_, _10094_);
  and _70282_ (_19552_, _19551_, _19549_);
  or _70283_ (_19553_, _19552_, _19548_);
  and _70284_ (_19554_, _19553_, _06219_);
  or _70285_ (_19555_, _19554_, _19516_);
  and _70286_ (_19556_, _19555_, _07237_);
  or _70287_ (_19557_, _14668_, _11380_);
  and _70288_ (_19558_, _19514_, _06369_);
  and _70289_ (_19559_, _19558_, _19557_);
  or _70290_ (_19560_, _19559_, _06536_);
  or _70291_ (_19562_, _19560_, _19556_);
  nor _70292_ (_19563_, _11261_, _11380_);
  or _70293_ (_19564_, _19563_, _19518_);
  nand _70294_ (_19565_, _11260_, _07951_);
  and _70295_ (_19566_, _19565_, _19564_);
  or _70296_ (_19567_, _19566_, _07240_);
  and _70297_ (_19568_, _19567_, _07242_);
  and _70298_ (_19569_, _19568_, _19562_);
  or _70299_ (_19570_, _14666_, _11380_);
  and _70300_ (_19571_, _19514_, _06375_);
  and _70301_ (_19573_, _19571_, _19570_);
  or _70302_ (_19574_, _19573_, _06545_);
  or _70303_ (_19575_, _19574_, _19569_);
  nor _70304_ (_19576_, _19518_, _07234_);
  nand _70305_ (_19577_, _19576_, _19565_);
  and _70306_ (_19578_, _19577_, _09056_);
  and _70307_ (_19579_, _19578_, _19575_);
  or _70308_ (_19580_, _19513_, _08341_);
  and _70309_ (_19581_, _19514_, _06366_);
  and _70310_ (_19582_, _19581_, _19580_);
  or _70311_ (_19584_, _19582_, _06528_);
  or _70312_ (_19585_, _19584_, _19579_);
  or _70313_ (_19586_, _19564_, _09061_);
  and _70314_ (_19587_, _19586_, _06926_);
  and _70315_ (_19588_, _19587_, _19585_);
  and _70316_ (_19589_, _19524_, _06568_);
  or _70317_ (_19590_, _19589_, _06278_);
  or _70318_ (_19591_, _19590_, _19588_);
  or _70319_ (_19592_, _19518_, _06279_);
  or _70320_ (_19593_, _19592_, _19522_);
  and _70321_ (_19595_, _19593_, _01347_);
  and _70322_ (_19596_, _19595_, _19591_);
  or _70323_ (_19597_, _19596_, _19512_);
  and _70324_ (_43171_, _19597_, _42618_);
  not _70325_ (_19598_, \oc8051_golden_model_1.PCON [2]);
  nor _70326_ (_19599_, _01347_, _19598_);
  nor _70327_ (_19600_, _07951_, _19598_);
  nor _70328_ (_19601_, _11380_, _07776_);
  or _70329_ (_19602_, _19601_, _19600_);
  or _70330_ (_19603_, _19602_, _07215_);
  and _70331_ (_19605_, _14770_, _07951_);
  or _70332_ (_19606_, _19605_, _19600_);
  and _70333_ (_19607_, _19606_, _06341_);
  nor _70334_ (_19608_, _07141_, _19598_);
  and _70335_ (_19609_, _07951_, \oc8051_golden_model_1.ACC [2]);
  or _70336_ (_19610_, _19609_, _19600_);
  and _70337_ (_19611_, _19610_, _07141_);
  or _70338_ (_19612_, _19611_, _19608_);
  and _70339_ (_19613_, _19612_, _07151_);
  or _70340_ (_19614_, _19613_, _06461_);
  or _70341_ (_19616_, _19614_, _19607_);
  or _70342_ (_19617_, _19602_, _07166_);
  and _70343_ (_19618_, _19617_, _06465_);
  and _70344_ (_19619_, _19618_, _19616_);
  and _70345_ (_19620_, _19610_, _06464_);
  or _70346_ (_19621_, _19620_, _10080_);
  or _70347_ (_19622_, _19621_, _19619_);
  and _70348_ (_19623_, _19622_, _19603_);
  or _70349_ (_19624_, _19623_, _07460_);
  and _70350_ (_19625_, _09450_, _07951_);
  or _70351_ (_19627_, _19600_, _07208_);
  or _70352_ (_19628_, _19627_, _19625_);
  and _70353_ (_19629_, _19628_, _19624_);
  or _70354_ (_19630_, _19629_, _10094_);
  and _70355_ (_19631_, _14859_, _07951_);
  or _70356_ (_19632_, _19600_, _05982_);
  or _70357_ (_19633_, _19632_, _19631_);
  and _70358_ (_19634_, _19633_, _06219_);
  and _70359_ (_19635_, _19634_, _19630_);
  and _70360_ (_19636_, _07951_, _08973_);
  or _70361_ (_19638_, _19636_, _19600_);
  and _70362_ (_19639_, _19638_, _06218_);
  or _70363_ (_19640_, _19639_, _06369_);
  or _70364_ (_19641_, _19640_, _19635_);
  and _70365_ (_19642_, _14751_, _07951_);
  or _70366_ (_19643_, _19642_, _19600_);
  or _70367_ (_19644_, _19643_, _07237_);
  and _70368_ (_19645_, _19644_, _07240_);
  and _70369_ (_19646_, _19645_, _19641_);
  and _70370_ (_19647_, _11259_, _07951_);
  or _70371_ (_19649_, _19647_, _19600_);
  and _70372_ (_19650_, _19649_, _06536_);
  or _70373_ (_19651_, _19650_, _19646_);
  and _70374_ (_19652_, _19651_, _07242_);
  or _70375_ (_19653_, _19600_, _08440_);
  and _70376_ (_19654_, _19638_, _06375_);
  and _70377_ (_19655_, _19654_, _19653_);
  or _70378_ (_19656_, _19655_, _19652_);
  and _70379_ (_19657_, _19656_, _07234_);
  and _70380_ (_19658_, _19610_, _06545_);
  and _70381_ (_19660_, _19658_, _19653_);
  or _70382_ (_19661_, _19660_, _06366_);
  or _70383_ (_19662_, _19661_, _19657_);
  and _70384_ (_19663_, _14748_, _07951_);
  or _70385_ (_19664_, _19600_, _09056_);
  or _70386_ (_19665_, _19664_, _19663_);
  and _70387_ (_19666_, _19665_, _09061_);
  and _70388_ (_19667_, _19666_, _19662_);
  nor _70389_ (_19668_, _11258_, _11380_);
  or _70390_ (_19669_, _19668_, _19600_);
  and _70391_ (_19671_, _19669_, _06528_);
  or _70392_ (_19672_, _19671_, _19667_);
  and _70393_ (_19673_, _19672_, _06926_);
  and _70394_ (_19674_, _19606_, _06568_);
  or _70395_ (_19675_, _19674_, _06278_);
  or _70396_ (_19676_, _19675_, _19673_);
  and _70397_ (_19677_, _14926_, _07951_);
  or _70398_ (_19678_, _19600_, _06279_);
  or _70399_ (_19679_, _19678_, _19677_);
  and _70400_ (_19680_, _19679_, _01347_);
  and _70401_ (_19682_, _19680_, _19676_);
  or _70402_ (_19683_, _19682_, _19599_);
  and _70403_ (_43172_, _19683_, _42618_);
  not _70404_ (_19684_, \oc8051_golden_model_1.PCON [3]);
  nor _70405_ (_19685_, _01347_, _19684_);
  nor _70406_ (_19686_, _07951_, _19684_);
  and _70407_ (_19687_, _14953_, _07951_);
  or _70408_ (_19688_, _19687_, _19686_);
  or _70409_ (_19689_, _19688_, _07151_);
  and _70410_ (_19690_, _07951_, \oc8051_golden_model_1.ACC [3]);
  or _70411_ (_19692_, _19690_, _19686_);
  and _70412_ (_19693_, _19692_, _07141_);
  nor _70413_ (_19694_, _07141_, _19684_);
  or _70414_ (_19695_, _19694_, _06341_);
  or _70415_ (_19696_, _19695_, _19693_);
  and _70416_ (_19697_, _19696_, _07166_);
  and _70417_ (_19698_, _19697_, _19689_);
  nor _70418_ (_19699_, _11380_, _07594_);
  or _70419_ (_19700_, _19699_, _19686_);
  and _70420_ (_19701_, _19700_, _06461_);
  or _70421_ (_19703_, _19701_, _19698_);
  and _70422_ (_19704_, _19703_, _06465_);
  and _70423_ (_19705_, _19692_, _06464_);
  or _70424_ (_19706_, _19705_, _10080_);
  or _70425_ (_19707_, _19706_, _19704_);
  or _70426_ (_19708_, _19700_, _07215_);
  and _70427_ (_19709_, _19708_, _07208_);
  and _70428_ (_19710_, _19709_, _19707_);
  and _70429_ (_19711_, _09449_, _07951_);
  or _70430_ (_19712_, _19711_, _19686_);
  and _70431_ (_19714_, _19712_, _07460_);
  or _70432_ (_19715_, _19714_, _10094_);
  or _70433_ (_19716_, _19715_, _19710_);
  and _70434_ (_19717_, _15048_, _07951_);
  or _70435_ (_19718_, _19686_, _05982_);
  or _70436_ (_19719_, _19718_, _19717_);
  and _70437_ (_19720_, _19719_, _06219_);
  and _70438_ (_19721_, _19720_, _19716_);
  and _70439_ (_19722_, _07951_, _08930_);
  or _70440_ (_19723_, _19722_, _19686_);
  and _70441_ (_19725_, _19723_, _06218_);
  or _70442_ (_19726_, _19725_, _06369_);
  or _70443_ (_19727_, _19726_, _19721_);
  and _70444_ (_19728_, _14943_, _07951_);
  or _70445_ (_19729_, _19728_, _19686_);
  or _70446_ (_19730_, _19729_, _07237_);
  and _70447_ (_19731_, _19730_, _07240_);
  and _70448_ (_19732_, _19731_, _19727_);
  and _70449_ (_19733_, _12577_, _07951_);
  or _70450_ (_19734_, _19733_, _19686_);
  and _70451_ (_19736_, _19734_, _06536_);
  or _70452_ (_19737_, _19736_, _19732_);
  and _70453_ (_19738_, _19737_, _07242_);
  or _70454_ (_19739_, _19686_, _08292_);
  and _70455_ (_19740_, _19723_, _06375_);
  and _70456_ (_19741_, _19740_, _19739_);
  or _70457_ (_19742_, _19741_, _19738_);
  and _70458_ (_19743_, _19742_, _07234_);
  and _70459_ (_19744_, _19692_, _06545_);
  and _70460_ (_19745_, _19744_, _19739_);
  or _70461_ (_19747_, _19745_, _06366_);
  or _70462_ (_19748_, _19747_, _19743_);
  and _70463_ (_19749_, _14940_, _07951_);
  or _70464_ (_19750_, _19686_, _09056_);
  or _70465_ (_19751_, _19750_, _19749_);
  and _70466_ (_19752_, _19751_, _09061_);
  and _70467_ (_19753_, _19752_, _19748_);
  nor _70468_ (_19754_, _11256_, _11380_);
  or _70469_ (_19755_, _19754_, _19686_);
  and _70470_ (_19756_, _19755_, _06528_);
  or _70471_ (_19758_, _19756_, _19753_);
  and _70472_ (_19759_, _19758_, _06926_);
  and _70473_ (_19760_, _19688_, _06568_);
  or _70474_ (_19761_, _19760_, _06278_);
  or _70475_ (_19762_, _19761_, _19759_);
  and _70476_ (_19763_, _15128_, _07951_);
  or _70477_ (_19764_, _19686_, _06279_);
  or _70478_ (_19765_, _19764_, _19763_);
  and _70479_ (_19766_, _19765_, _01347_);
  and _70480_ (_19767_, _19766_, _19762_);
  or _70481_ (_19770_, _19767_, _19685_);
  and _70482_ (_43173_, _19770_, _42618_);
  not _70483_ (_19771_, \oc8051_golden_model_1.PCON [4]);
  nor _70484_ (_19772_, _01347_, _19771_);
  nor _70485_ (_19773_, _07951_, _19771_);
  nor _70486_ (_19774_, _08541_, _11380_);
  or _70487_ (_19775_, _19774_, _19773_);
  or _70488_ (_19776_, _19775_, _07215_);
  and _70489_ (_19777_, _15162_, _07951_);
  or _70490_ (_19778_, _19777_, _19773_);
  or _70491_ (_19781_, _19778_, _07151_);
  and _70492_ (_19782_, _07951_, \oc8051_golden_model_1.ACC [4]);
  or _70493_ (_19783_, _19782_, _19773_);
  and _70494_ (_19784_, _19783_, _07141_);
  nor _70495_ (_19785_, _07141_, _19771_);
  or _70496_ (_19786_, _19785_, _06341_);
  or _70497_ (_19787_, _19786_, _19784_);
  and _70498_ (_19788_, _19787_, _07166_);
  and _70499_ (_19789_, _19788_, _19781_);
  and _70500_ (_19790_, _19775_, _06461_);
  or _70501_ (_19793_, _19790_, _19789_);
  and _70502_ (_19794_, _19793_, _06465_);
  and _70503_ (_19795_, _19783_, _06464_);
  or _70504_ (_19796_, _19795_, _10080_);
  or _70505_ (_19797_, _19796_, _19794_);
  and _70506_ (_19798_, _19797_, _19776_);
  or _70507_ (_19799_, _19798_, _07460_);
  and _70508_ (_19800_, _09448_, _07951_);
  or _70509_ (_19801_, _19773_, _07208_);
  or _70510_ (_19802_, _19801_, _19800_);
  and _70511_ (_19805_, _19802_, _19799_);
  or _70512_ (_19806_, _19805_, _10094_);
  and _70513_ (_19807_, _15254_, _07951_);
  or _70514_ (_19808_, _19773_, _05982_);
  or _70515_ (_19809_, _19808_, _19807_);
  and _70516_ (_19810_, _19809_, _06219_);
  and _70517_ (_19811_, _19810_, _19806_);
  and _70518_ (_19812_, _08959_, _07951_);
  or _70519_ (_19813_, _19812_, _19773_);
  and _70520_ (_19814_, _19813_, _06218_);
  or _70521_ (_19817_, _19814_, _06369_);
  or _70522_ (_19818_, _19817_, _19811_);
  and _70523_ (_19819_, _15269_, _07951_);
  or _70524_ (_19820_, _19819_, _19773_);
  or _70525_ (_19821_, _19820_, _07237_);
  and _70526_ (_19822_, _19821_, _07240_);
  and _70527_ (_19823_, _19822_, _19818_);
  and _70528_ (_19824_, _11254_, _07951_);
  or _70529_ (_19825_, _19824_, _19773_);
  and _70530_ (_19826_, _19825_, _06536_);
  or _70531_ (_19829_, _19826_, _19823_);
  and _70532_ (_19830_, _19829_, _07242_);
  or _70533_ (_19831_, _19773_, _08544_);
  and _70534_ (_19832_, _19813_, _06375_);
  and _70535_ (_19833_, _19832_, _19831_);
  or _70536_ (_19834_, _19833_, _19830_);
  and _70537_ (_19835_, _19834_, _07234_);
  and _70538_ (_19836_, _19783_, _06545_);
  and _70539_ (_19837_, _19836_, _19831_);
  or _70540_ (_19838_, _19837_, _06366_);
  or _70541_ (_19841_, _19838_, _19835_);
  and _70542_ (_19842_, _15266_, _07951_);
  or _70543_ (_19843_, _19773_, _09056_);
  or _70544_ (_19844_, _19843_, _19842_);
  and _70545_ (_19845_, _19844_, _09061_);
  and _70546_ (_19846_, _19845_, _19841_);
  nor _70547_ (_19847_, _11253_, _11380_);
  or _70548_ (_19848_, _19847_, _19773_);
  and _70549_ (_19849_, _19848_, _06528_);
  or _70550_ (_19850_, _19849_, _19846_);
  and _70551_ (_19852_, _19850_, _06926_);
  and _70552_ (_19853_, _19778_, _06568_);
  or _70553_ (_19854_, _19853_, _06278_);
  or _70554_ (_19855_, _19854_, _19852_);
  and _70555_ (_19856_, _15329_, _07951_);
  or _70556_ (_19857_, _19773_, _06279_);
  or _70557_ (_19858_, _19857_, _19856_);
  and _70558_ (_19859_, _19858_, _01347_);
  and _70559_ (_19860_, _19859_, _19855_);
  or _70560_ (_19861_, _19860_, _19772_);
  and _70561_ (_43174_, _19861_, _42618_);
  not _70562_ (_19863_, \oc8051_golden_model_1.PCON [5]);
  nor _70563_ (_19864_, _01347_, _19863_);
  nor _70564_ (_19865_, _07951_, _19863_);
  nor _70565_ (_19866_, _08244_, _11380_);
  or _70566_ (_19867_, _19866_, _19865_);
  or _70567_ (_19868_, _19867_, _07215_);
  and _70568_ (_19869_, _15358_, _07951_);
  or _70569_ (_19870_, _19869_, _19865_);
  or _70570_ (_19871_, _19870_, _07151_);
  and _70571_ (_19873_, _07951_, \oc8051_golden_model_1.ACC [5]);
  or _70572_ (_19874_, _19873_, _19865_);
  and _70573_ (_19875_, _19874_, _07141_);
  nor _70574_ (_19876_, _07141_, _19863_);
  or _70575_ (_19877_, _19876_, _06341_);
  or _70576_ (_19878_, _19877_, _19875_);
  and _70577_ (_19879_, _19878_, _07166_);
  and _70578_ (_19880_, _19879_, _19871_);
  and _70579_ (_19881_, _19867_, _06461_);
  or _70580_ (_19882_, _19881_, _19880_);
  and _70581_ (_19884_, _19882_, _06465_);
  and _70582_ (_19885_, _19874_, _06464_);
  or _70583_ (_19886_, _19885_, _10080_);
  or _70584_ (_19887_, _19886_, _19884_);
  and _70585_ (_19888_, _19887_, _19868_);
  or _70586_ (_19889_, _19888_, _07460_);
  and _70587_ (_19890_, _09447_, _07951_);
  or _70588_ (_19891_, _19865_, _07208_);
  or _70589_ (_19892_, _19891_, _19890_);
  and _70590_ (_19893_, _19892_, _05982_);
  and _70591_ (_19895_, _19893_, _19889_);
  and _70592_ (_19896_, _15459_, _07951_);
  or _70593_ (_19897_, _19896_, _19865_);
  and _70594_ (_19898_, _19897_, _10094_);
  or _70595_ (_19899_, _19898_, _06218_);
  or _70596_ (_19900_, _19899_, _19895_);
  and _70597_ (_19901_, _08946_, _07951_);
  or _70598_ (_19902_, _19901_, _19865_);
  or _70599_ (_19903_, _19902_, _06219_);
  and _70600_ (_19904_, _19903_, _19900_);
  or _70601_ (_19906_, _19904_, _06369_);
  and _70602_ (_19907_, _15353_, _07951_);
  or _70603_ (_19908_, _19907_, _19865_);
  or _70604_ (_19909_, _19908_, _07237_);
  and _70605_ (_19910_, _19909_, _07240_);
  and _70606_ (_19911_, _19910_, _19906_);
  and _70607_ (_19912_, _11250_, _07951_);
  or _70608_ (_19913_, _19912_, _19865_);
  and _70609_ (_19914_, _19913_, _06536_);
  or _70610_ (_19915_, _19914_, _19911_);
  and _70611_ (_19917_, _19915_, _07242_);
  or _70612_ (_19918_, _19865_, _08247_);
  and _70613_ (_19919_, _19902_, _06375_);
  and _70614_ (_19920_, _19919_, _19918_);
  or _70615_ (_19921_, _19920_, _19917_);
  and _70616_ (_19922_, _19921_, _07234_);
  and _70617_ (_19923_, _19874_, _06545_);
  and _70618_ (_19924_, _19923_, _19918_);
  or _70619_ (_19925_, _19924_, _06366_);
  or _70620_ (_19926_, _19925_, _19922_);
  and _70621_ (_19928_, _15350_, _07951_);
  or _70622_ (_19929_, _19865_, _09056_);
  or _70623_ (_19930_, _19929_, _19928_);
  and _70624_ (_19931_, _19930_, _09061_);
  and _70625_ (_19932_, _19931_, _19926_);
  nor _70626_ (_19933_, _11249_, _11380_);
  or _70627_ (_19934_, _19933_, _19865_);
  and _70628_ (_19935_, _19934_, _06528_);
  or _70629_ (_19936_, _19935_, _19932_);
  and _70630_ (_19937_, _19936_, _06926_);
  and _70631_ (_19939_, _19870_, _06568_);
  or _70632_ (_19940_, _19939_, _06278_);
  or _70633_ (_19941_, _19940_, _19937_);
  and _70634_ (_19942_, _15532_, _07951_);
  or _70635_ (_19943_, _19865_, _06279_);
  or _70636_ (_19944_, _19943_, _19942_);
  and _70637_ (_19945_, _19944_, _01347_);
  and _70638_ (_19946_, _19945_, _19941_);
  or _70639_ (_19947_, _19946_, _19864_);
  and _70640_ (_43175_, _19947_, _42618_);
  not _70641_ (_19949_, \oc8051_golden_model_1.PCON [6]);
  nor _70642_ (_19950_, _01347_, _19949_);
  nor _70643_ (_19951_, _07951_, _19949_);
  nor _70644_ (_19952_, _08142_, _11380_);
  or _70645_ (_19953_, _19952_, _19951_);
  or _70646_ (_19954_, _19953_, _07215_);
  and _70647_ (_19955_, _15554_, _07951_);
  or _70648_ (_19956_, _19955_, _19951_);
  or _70649_ (_19957_, _19956_, _07151_);
  and _70650_ (_19958_, _07951_, \oc8051_golden_model_1.ACC [6]);
  or _70651_ (_19960_, _19958_, _19951_);
  and _70652_ (_19961_, _19960_, _07141_);
  nor _70653_ (_19962_, _07141_, _19949_);
  or _70654_ (_19963_, _19962_, _06341_);
  or _70655_ (_19964_, _19963_, _19961_);
  and _70656_ (_19965_, _19964_, _07166_);
  and _70657_ (_19966_, _19965_, _19957_);
  and _70658_ (_19967_, _19953_, _06461_);
  or _70659_ (_19968_, _19967_, _19966_);
  and _70660_ (_19969_, _19968_, _06465_);
  and _70661_ (_19971_, _19960_, _06464_);
  or _70662_ (_19972_, _19971_, _10080_);
  or _70663_ (_19973_, _19972_, _19969_);
  and _70664_ (_19974_, _19973_, _19954_);
  or _70665_ (_19975_, _19974_, _07460_);
  and _70666_ (_19976_, _09446_, _07951_);
  or _70667_ (_19977_, _19951_, _07208_);
  or _70668_ (_19978_, _19977_, _19976_);
  and _70669_ (_19979_, _19978_, _05982_);
  and _70670_ (_19980_, _19979_, _19975_);
  and _70671_ (_19982_, _15657_, _07951_);
  or _70672_ (_19983_, _19982_, _19951_);
  and _70673_ (_19984_, _19983_, _10094_);
  or _70674_ (_19985_, _19984_, _06218_);
  or _70675_ (_19986_, _19985_, _19980_);
  and _70676_ (_19987_, _15664_, _07951_);
  or _70677_ (_19988_, _19987_, _19951_);
  or _70678_ (_19989_, _19988_, _06219_);
  and _70679_ (_19990_, _19989_, _19986_);
  or _70680_ (_19991_, _19990_, _06369_);
  and _70681_ (_19993_, _15549_, _07951_);
  or _70682_ (_19994_, _19993_, _19951_);
  or _70683_ (_19995_, _19994_, _07237_);
  and _70684_ (_19996_, _19995_, _07240_);
  and _70685_ (_19997_, _19996_, _19991_);
  and _70686_ (_19998_, _11247_, _07951_);
  or _70687_ (_19999_, _19998_, _19951_);
  and _70688_ (_20000_, _19999_, _06536_);
  or _70689_ (_20001_, _20000_, _19997_);
  and _70690_ (_20002_, _20001_, _07242_);
  or _70691_ (_20004_, _19951_, _08145_);
  and _70692_ (_20005_, _19988_, _06375_);
  and _70693_ (_20006_, _20005_, _20004_);
  or _70694_ (_20007_, _20006_, _20002_);
  and _70695_ (_20008_, _20007_, _07234_);
  and _70696_ (_20009_, _19960_, _06545_);
  and _70697_ (_20010_, _20009_, _20004_);
  or _70698_ (_20011_, _20010_, _06366_);
  or _70699_ (_20012_, _20011_, _20008_);
  and _70700_ (_20013_, _15546_, _07951_);
  or _70701_ (_20015_, _19951_, _09056_);
  or _70702_ (_20016_, _20015_, _20013_);
  and _70703_ (_20017_, _20016_, _09061_);
  and _70704_ (_20018_, _20017_, _20012_);
  nor _70705_ (_20019_, _11246_, _11380_);
  or _70706_ (_20020_, _20019_, _19951_);
  and _70707_ (_20021_, _20020_, _06528_);
  or _70708_ (_20022_, _20021_, _20018_);
  and _70709_ (_20023_, _20022_, _06926_);
  and _70710_ (_20024_, _19956_, _06568_);
  or _70711_ (_20026_, _20024_, _06278_);
  or _70712_ (_20027_, _20026_, _20023_);
  and _70713_ (_20028_, _15734_, _07951_);
  or _70714_ (_20029_, _19951_, _06279_);
  or _70715_ (_20030_, _20029_, _20028_);
  and _70716_ (_20031_, _20030_, _01347_);
  and _70717_ (_20032_, _20031_, _20027_);
  or _70718_ (_20033_, _20032_, _19950_);
  and _70719_ (_43176_, _20033_, _42618_);
  not _70720_ (_20034_, \oc8051_golden_model_1.TMOD [0]);
  nor _70721_ (_20036_, _01347_, _20034_);
  nand _70722_ (_20037_, _11263_, _07914_);
  nor _70723_ (_20038_, _07914_, _20034_);
  nor _70724_ (_20039_, _20038_, _07234_);
  nand _70725_ (_20040_, _20039_, _20037_);
  and _70726_ (_20041_, _07914_, _07133_);
  or _70727_ (_20042_, _20041_, _20038_);
  or _70728_ (_20043_, _20042_, _07215_);
  nor _70729_ (_20044_, _08390_, _11457_);
  or _70730_ (_20045_, _20044_, _20038_);
  or _70731_ (_20047_, _20045_, _07151_);
  and _70732_ (_20048_, _07914_, \oc8051_golden_model_1.ACC [0]);
  or _70733_ (_20049_, _20048_, _20038_);
  and _70734_ (_20050_, _20049_, _07141_);
  nor _70735_ (_20051_, _07141_, _20034_);
  or _70736_ (_20052_, _20051_, _06341_);
  or _70737_ (_20053_, _20052_, _20050_);
  and _70738_ (_20054_, _20053_, _07166_);
  and _70739_ (_20055_, _20054_, _20047_);
  and _70740_ (_20056_, _20042_, _06461_);
  or _70741_ (_20058_, _20056_, _20055_);
  and _70742_ (_20059_, _20058_, _06465_);
  and _70743_ (_20060_, _20049_, _06464_);
  or _70744_ (_20061_, _20060_, _10080_);
  or _70745_ (_20062_, _20061_, _20059_);
  and _70746_ (_20063_, _20062_, _20043_);
  or _70747_ (_20064_, _20063_, _07460_);
  and _70748_ (_20065_, _09392_, _07914_);
  or _70749_ (_20066_, _20038_, _07208_);
  or _70750_ (_20067_, _20066_, _20065_);
  and _70751_ (_20069_, _20067_, _20064_);
  or _70752_ (_20070_, _20069_, _10094_);
  and _70753_ (_20071_, _14467_, _07914_);
  or _70754_ (_20072_, _20038_, _05982_);
  or _70755_ (_20073_, _20072_, _20071_);
  and _70756_ (_20074_, _20073_, _06219_);
  and _70757_ (_20075_, _20074_, _20070_);
  and _70758_ (_20076_, _07914_, _08954_);
  or _70759_ (_20077_, _20076_, _20038_);
  and _70760_ (_20078_, _20077_, _06218_);
  or _70761_ (_20080_, _20078_, _06369_);
  or _70762_ (_20081_, _20080_, _20075_);
  and _70763_ (_20082_, _14366_, _07914_);
  or _70764_ (_20083_, _20082_, _20038_);
  or _70765_ (_20084_, _20083_, _07237_);
  and _70766_ (_20085_, _20084_, _07240_);
  and _70767_ (_20086_, _20085_, _20081_);
  nor _70768_ (_20087_, _12580_, _11457_);
  or _70769_ (_20088_, _20087_, _20038_);
  and _70770_ (_20089_, _20037_, _06536_);
  and _70771_ (_20091_, _20089_, _20088_);
  or _70772_ (_20092_, _20091_, _20086_);
  and _70773_ (_20093_, _20092_, _07242_);
  nand _70774_ (_20094_, _20077_, _06375_);
  nor _70775_ (_20095_, _20094_, _20044_);
  or _70776_ (_20096_, _20095_, _06545_);
  or _70777_ (_20097_, _20096_, _20093_);
  and _70778_ (_20098_, _20097_, _20040_);
  or _70779_ (_20099_, _20098_, _06366_);
  and _70780_ (_20100_, _14363_, _07914_);
  or _70781_ (_20102_, _20038_, _09056_);
  or _70782_ (_20103_, _20102_, _20100_);
  and _70783_ (_20104_, _20103_, _09061_);
  and _70784_ (_20105_, _20104_, _20099_);
  and _70785_ (_20106_, _20088_, _06528_);
  or _70786_ (_20107_, _20106_, _19502_);
  or _70787_ (_20108_, _20107_, _20105_);
  or _70788_ (_20109_, _20045_, _06661_);
  and _70789_ (_20110_, _20109_, _01347_);
  and _70790_ (_20111_, _20110_, _20108_);
  or _70791_ (_20113_, _20111_, _20036_);
  and _70792_ (_43178_, _20113_, _42618_);
  and _70793_ (_20114_, _01351_, \oc8051_golden_model_1.TMOD [1]);
  nand _70794_ (_20115_, _07914_, _07038_);
  or _70795_ (_20116_, _07914_, \oc8051_golden_model_1.TMOD [1]);
  and _70796_ (_20117_, _20116_, _06218_);
  and _70797_ (_20118_, _20117_, _20115_);
  and _70798_ (_20119_, _11457_, \oc8051_golden_model_1.TMOD [1]);
  nor _70799_ (_20120_, _11457_, _07357_);
  or _70800_ (_20121_, _20120_, _20119_);
  or _70801_ (_20123_, _20121_, _07215_);
  and _70802_ (_20124_, _14562_, _07914_);
  not _70803_ (_20125_, _20124_);
  and _70804_ (_20126_, _20125_, _20116_);
  or _70805_ (_20127_, _20126_, _07151_);
  and _70806_ (_20128_, _07914_, \oc8051_golden_model_1.ACC [1]);
  or _70807_ (_20129_, _20128_, _20119_);
  and _70808_ (_20130_, _20129_, _07141_);
  and _70809_ (_20131_, _07142_, \oc8051_golden_model_1.TMOD [1]);
  or _70810_ (_20132_, _20131_, _06341_);
  or _70811_ (_20134_, _20132_, _20130_);
  and _70812_ (_20135_, _20134_, _07166_);
  and _70813_ (_20136_, _20135_, _20127_);
  and _70814_ (_20137_, _20121_, _06461_);
  or _70815_ (_20138_, _20137_, _20136_);
  and _70816_ (_20139_, _20138_, _06465_);
  and _70817_ (_20140_, _20129_, _06464_);
  or _70818_ (_20141_, _20140_, _10080_);
  or _70819_ (_20142_, _20141_, _20139_);
  and _70820_ (_20143_, _20142_, _20123_);
  or _70821_ (_20145_, _20143_, _07460_);
  and _70822_ (_20146_, _09451_, _07914_);
  or _70823_ (_20147_, _20119_, _07208_);
  or _70824_ (_20148_, _20147_, _20146_);
  and _70825_ (_20149_, _20148_, _05982_);
  and _70826_ (_20150_, _20149_, _20145_);
  or _70827_ (_20151_, _14653_, _11457_);
  and _70828_ (_20152_, _20116_, _10094_);
  and _70829_ (_20153_, _20152_, _20151_);
  or _70830_ (_20154_, _20153_, _20150_);
  and _70831_ (_20156_, _20154_, _06219_);
  or _70832_ (_20157_, _20156_, _20118_);
  and _70833_ (_20158_, _20157_, _07237_);
  or _70834_ (_20159_, _14668_, _11457_);
  and _70835_ (_20160_, _20116_, _06369_);
  and _70836_ (_20161_, _20160_, _20159_);
  or _70837_ (_20162_, _20161_, _06536_);
  or _70838_ (_20163_, _20162_, _20158_);
  and _70839_ (_20164_, _11262_, _07914_);
  or _70840_ (_20165_, _20164_, _20119_);
  or _70841_ (_20167_, _20165_, _07240_);
  and _70842_ (_20168_, _20167_, _07242_);
  and _70843_ (_20169_, _20168_, _20163_);
  or _70844_ (_20170_, _14666_, _11457_);
  and _70845_ (_20171_, _20116_, _06375_);
  and _70846_ (_20172_, _20171_, _20170_);
  or _70847_ (_20173_, _20172_, _06545_);
  or _70848_ (_20174_, _20173_, _20169_);
  and _70849_ (_20175_, _20128_, _08341_);
  or _70850_ (_20176_, _20119_, _07234_);
  or _70851_ (_20178_, _20176_, _20175_);
  and _70852_ (_20179_, _20178_, _09056_);
  and _70853_ (_20180_, _20179_, _20174_);
  or _70854_ (_20181_, _20115_, _08341_);
  and _70855_ (_20182_, _20116_, _06366_);
  and _70856_ (_20183_, _20182_, _20181_);
  or _70857_ (_20184_, _20183_, _06528_);
  or _70858_ (_20185_, _20184_, _20180_);
  nor _70859_ (_20186_, _11261_, _11457_);
  or _70860_ (_20187_, _20186_, _20119_);
  or _70861_ (_20189_, _20187_, _09061_);
  and _70862_ (_20190_, _20189_, _06926_);
  and _70863_ (_20191_, _20190_, _20185_);
  and _70864_ (_20192_, _20126_, _06568_);
  or _70865_ (_20193_, _20192_, _06278_);
  or _70866_ (_20194_, _20193_, _20191_);
  or _70867_ (_20195_, _20119_, _06279_);
  or _70868_ (_20196_, _20195_, _20124_);
  and _70869_ (_20197_, _20196_, _01347_);
  and _70870_ (_20198_, _20197_, _20194_);
  or _70871_ (_20200_, _20198_, _20114_);
  and _70872_ (_43179_, _20200_, _42618_);
  and _70873_ (_20201_, _01351_, \oc8051_golden_model_1.TMOD [2]);
  and _70874_ (_20202_, _11457_, \oc8051_golden_model_1.TMOD [2]);
  and _70875_ (_20203_, _09450_, _07914_);
  or _70876_ (_20204_, _20203_, _20202_);
  and _70877_ (_20205_, _20204_, _07460_);
  and _70878_ (_20206_, _14770_, _07914_);
  or _70879_ (_20207_, _20206_, _20202_);
  or _70880_ (_20208_, _20207_, _07151_);
  and _70881_ (_20210_, _07914_, \oc8051_golden_model_1.ACC [2]);
  or _70882_ (_20211_, _20210_, _20202_);
  and _70883_ (_20212_, _20211_, _07141_);
  and _70884_ (_20213_, _07142_, \oc8051_golden_model_1.TMOD [2]);
  or _70885_ (_20214_, _20213_, _06341_);
  or _70886_ (_20215_, _20214_, _20212_);
  and _70887_ (_20216_, _20215_, _07166_);
  and _70888_ (_20217_, _20216_, _20208_);
  nor _70889_ (_20218_, _11457_, _07776_);
  or _70890_ (_20219_, _20218_, _20202_);
  and _70891_ (_20221_, _20219_, _06461_);
  or _70892_ (_20222_, _20221_, _20217_);
  and _70893_ (_20223_, _20222_, _06465_);
  and _70894_ (_20224_, _20211_, _06464_);
  or _70895_ (_20225_, _20224_, _10080_);
  or _70896_ (_20226_, _20225_, _20223_);
  or _70897_ (_20227_, _20219_, _07215_);
  and _70898_ (_20228_, _20227_, _07208_);
  and _70899_ (_20229_, _20228_, _20226_);
  or _70900_ (_20230_, _20229_, _10094_);
  or _70901_ (_20232_, _20230_, _20205_);
  and _70902_ (_20233_, _14859_, _07914_);
  or _70903_ (_20234_, _20202_, _05982_);
  or _70904_ (_20235_, _20234_, _20233_);
  and _70905_ (_20236_, _20235_, _06219_);
  and _70906_ (_20237_, _20236_, _20232_);
  and _70907_ (_20238_, _07914_, _08973_);
  or _70908_ (_20239_, _20238_, _20202_);
  and _70909_ (_20240_, _20239_, _06218_);
  or _70910_ (_20241_, _20240_, _06369_);
  or _70911_ (_20243_, _20241_, _20237_);
  and _70912_ (_20244_, _14751_, _07914_);
  or _70913_ (_20245_, _20244_, _20202_);
  or _70914_ (_20246_, _20245_, _07237_);
  and _70915_ (_20247_, _20246_, _07240_);
  and _70916_ (_20248_, _20247_, _20243_);
  and _70917_ (_20249_, _11259_, _07914_);
  or _70918_ (_20250_, _20249_, _20202_);
  and _70919_ (_20251_, _20250_, _06536_);
  or _70920_ (_20252_, _20251_, _20248_);
  and _70921_ (_20254_, _20252_, _07242_);
  or _70922_ (_20255_, _20202_, _08440_);
  and _70923_ (_20256_, _20239_, _06375_);
  and _70924_ (_20257_, _20256_, _20255_);
  or _70925_ (_20258_, _20257_, _20254_);
  and _70926_ (_20259_, _20258_, _07234_);
  and _70927_ (_20260_, _20211_, _06545_);
  and _70928_ (_20261_, _20260_, _20255_);
  or _70929_ (_20262_, _20261_, _06366_);
  or _70930_ (_20263_, _20262_, _20259_);
  and _70931_ (_20265_, _14748_, _07914_);
  or _70932_ (_20266_, _20202_, _09056_);
  or _70933_ (_20267_, _20266_, _20265_);
  and _70934_ (_20268_, _20267_, _09061_);
  and _70935_ (_20269_, _20268_, _20263_);
  nor _70936_ (_20270_, _11258_, _11457_);
  or _70937_ (_20271_, _20270_, _20202_);
  and _70938_ (_20272_, _20271_, _06528_);
  or _70939_ (_20273_, _20272_, _20269_);
  and _70940_ (_20274_, _20273_, _06926_);
  and _70941_ (_20276_, _20207_, _06568_);
  or _70942_ (_20277_, _20276_, _06278_);
  or _70943_ (_20278_, _20277_, _20274_);
  and _70944_ (_20279_, _14926_, _07914_);
  or _70945_ (_20280_, _20202_, _06279_);
  or _70946_ (_20281_, _20280_, _20279_);
  and _70947_ (_20282_, _20281_, _01347_);
  and _70948_ (_20283_, _20282_, _20278_);
  or _70949_ (_20284_, _20283_, _20201_);
  and _70950_ (_43180_, _20284_, _42618_);
  and _70951_ (_20286_, _01351_, \oc8051_golden_model_1.TMOD [3]);
  and _70952_ (_20287_, _11457_, \oc8051_golden_model_1.TMOD [3]);
  and _70953_ (_20288_, _14953_, _07914_);
  or _70954_ (_20289_, _20288_, _20287_);
  or _70955_ (_20290_, _20289_, _07151_);
  and _70956_ (_20291_, _07914_, \oc8051_golden_model_1.ACC [3]);
  or _70957_ (_20292_, _20291_, _20287_);
  and _70958_ (_20293_, _20292_, _07141_);
  and _70959_ (_20294_, _07142_, \oc8051_golden_model_1.TMOD [3]);
  or _70960_ (_20295_, _20294_, _06341_);
  or _70961_ (_20297_, _20295_, _20293_);
  and _70962_ (_20298_, _20297_, _07166_);
  and _70963_ (_20299_, _20298_, _20290_);
  nor _70964_ (_20300_, _11457_, _07594_);
  or _70965_ (_20301_, _20300_, _20287_);
  and _70966_ (_20302_, _20301_, _06461_);
  or _70967_ (_20303_, _20302_, _20299_);
  and _70968_ (_20304_, _20303_, _06465_);
  and _70969_ (_20305_, _20292_, _06464_);
  or _70970_ (_20306_, _20305_, _10080_);
  or _70971_ (_20308_, _20306_, _20304_);
  or _70972_ (_20309_, _20301_, _07215_);
  and _70973_ (_20310_, _20309_, _07208_);
  and _70974_ (_20311_, _20310_, _20308_);
  and _70975_ (_20312_, _09449_, _07914_);
  or _70976_ (_20313_, _20312_, _20287_);
  and _70977_ (_20314_, _20313_, _07460_);
  or _70978_ (_20315_, _20314_, _10094_);
  or _70979_ (_20316_, _20315_, _20311_);
  and _70980_ (_20317_, _15048_, _07914_);
  or _70981_ (_20319_, _20287_, _05982_);
  or _70982_ (_20320_, _20319_, _20317_);
  and _70983_ (_20321_, _20320_, _06219_);
  and _70984_ (_20322_, _20321_, _20316_);
  and _70985_ (_20323_, _07914_, _08930_);
  or _70986_ (_20324_, _20323_, _20287_);
  and _70987_ (_20325_, _20324_, _06218_);
  or _70988_ (_20326_, _20325_, _06369_);
  or _70989_ (_20327_, _20326_, _20322_);
  and _70990_ (_20328_, _14943_, _07914_);
  or _70991_ (_20330_, _20328_, _20287_);
  or _70992_ (_20331_, _20330_, _07237_);
  and _70993_ (_20332_, _20331_, _07240_);
  and _70994_ (_20333_, _20332_, _20327_);
  and _70995_ (_20334_, _12577_, _07914_);
  or _70996_ (_20335_, _20334_, _20287_);
  and _70997_ (_20336_, _20335_, _06536_);
  or _70998_ (_20337_, _20336_, _20333_);
  and _70999_ (_20338_, _20337_, _07242_);
  or _71000_ (_20339_, _20287_, _08292_);
  and _71001_ (_20341_, _20324_, _06375_);
  and _71002_ (_20342_, _20341_, _20339_);
  or _71003_ (_20343_, _20342_, _20338_);
  and _71004_ (_20344_, _20343_, _07234_);
  and _71005_ (_20345_, _20292_, _06545_);
  and _71006_ (_20346_, _20345_, _20339_);
  or _71007_ (_20347_, _20346_, _06366_);
  or _71008_ (_20348_, _20347_, _20344_);
  and _71009_ (_20349_, _14940_, _07914_);
  or _71010_ (_20350_, _20287_, _09056_);
  or _71011_ (_20352_, _20350_, _20349_);
  and _71012_ (_20353_, _20352_, _09061_);
  and _71013_ (_20354_, _20353_, _20348_);
  nor _71014_ (_20355_, _11256_, _11457_);
  or _71015_ (_20356_, _20355_, _20287_);
  and _71016_ (_20357_, _20356_, _06528_);
  or _71017_ (_20358_, _20357_, _20354_);
  and _71018_ (_20359_, _20358_, _06926_);
  and _71019_ (_20360_, _20289_, _06568_);
  or _71020_ (_20361_, _20360_, _06278_);
  or _71021_ (_20363_, _20361_, _20359_);
  and _71022_ (_20364_, _15128_, _07914_);
  or _71023_ (_20365_, _20287_, _06279_);
  or _71024_ (_20366_, _20365_, _20364_);
  and _71025_ (_20367_, _20366_, _01347_);
  and _71026_ (_20368_, _20367_, _20363_);
  or _71027_ (_20369_, _20368_, _20286_);
  and _71028_ (_43182_, _20369_, _42618_);
  and _71029_ (_20370_, _01351_, \oc8051_golden_model_1.TMOD [4]);
  and _71030_ (_20371_, _11457_, \oc8051_golden_model_1.TMOD [4]);
  nor _71031_ (_20373_, _08541_, _11457_);
  or _71032_ (_20374_, _20373_, _20371_);
  or _71033_ (_20375_, _20374_, _07215_);
  and _71034_ (_20376_, _15162_, _07914_);
  or _71035_ (_20377_, _20376_, _20371_);
  or _71036_ (_20378_, _20377_, _07151_);
  and _71037_ (_20379_, _07914_, \oc8051_golden_model_1.ACC [4]);
  or _71038_ (_20380_, _20379_, _20371_);
  and _71039_ (_20381_, _20380_, _07141_);
  and _71040_ (_20382_, _07142_, \oc8051_golden_model_1.TMOD [4]);
  or _71041_ (_20384_, _20382_, _06341_);
  or _71042_ (_20385_, _20384_, _20381_);
  and _71043_ (_20386_, _20385_, _07166_);
  and _71044_ (_20387_, _20386_, _20378_);
  and _71045_ (_20388_, _20374_, _06461_);
  or _71046_ (_20389_, _20388_, _20387_);
  and _71047_ (_20390_, _20389_, _06465_);
  and _71048_ (_20391_, _20380_, _06464_);
  or _71049_ (_20392_, _20391_, _10080_);
  or _71050_ (_20393_, _20392_, _20390_);
  and _71051_ (_20395_, _20393_, _20375_);
  or _71052_ (_20396_, _20395_, _07460_);
  and _71053_ (_20397_, _09448_, _07914_);
  or _71054_ (_20398_, _20371_, _07208_);
  or _71055_ (_20399_, _20398_, _20397_);
  and _71056_ (_20400_, _20399_, _20396_);
  or _71057_ (_20401_, _20400_, _10094_);
  and _71058_ (_20402_, _15254_, _07914_);
  or _71059_ (_20403_, _20371_, _05982_);
  or _71060_ (_20404_, _20403_, _20402_);
  and _71061_ (_20406_, _20404_, _06219_);
  and _71062_ (_20407_, _20406_, _20401_);
  and _71063_ (_20408_, _08959_, _07914_);
  or _71064_ (_20409_, _20408_, _20371_);
  and _71065_ (_20410_, _20409_, _06218_);
  or _71066_ (_20411_, _20410_, _06369_);
  or _71067_ (_20412_, _20411_, _20407_);
  and _71068_ (_20413_, _15269_, _07914_);
  or _71069_ (_20414_, _20413_, _20371_);
  or _71070_ (_20415_, _20414_, _07237_);
  and _71071_ (_20417_, _20415_, _07240_);
  and _71072_ (_20418_, _20417_, _20412_);
  and _71073_ (_20419_, _11254_, _07914_);
  or _71074_ (_20420_, _20419_, _20371_);
  and _71075_ (_20421_, _20420_, _06536_);
  or _71076_ (_20422_, _20421_, _20418_);
  and _71077_ (_20423_, _20422_, _07242_);
  or _71078_ (_20424_, _20371_, _08544_);
  and _71079_ (_20425_, _20409_, _06375_);
  and _71080_ (_20426_, _20425_, _20424_);
  or _71081_ (_20428_, _20426_, _20423_);
  and _71082_ (_20429_, _20428_, _07234_);
  and _71083_ (_20430_, _20380_, _06545_);
  and _71084_ (_20431_, _20430_, _20424_);
  or _71085_ (_20432_, _20431_, _06366_);
  or _71086_ (_20433_, _20432_, _20429_);
  and _71087_ (_20434_, _15266_, _07914_);
  or _71088_ (_20435_, _20371_, _09056_);
  or _71089_ (_20436_, _20435_, _20434_);
  and _71090_ (_20437_, _20436_, _09061_);
  and _71091_ (_20439_, _20437_, _20433_);
  nor _71092_ (_20440_, _11253_, _11457_);
  or _71093_ (_20441_, _20440_, _20371_);
  and _71094_ (_20442_, _20441_, _06528_);
  or _71095_ (_20443_, _20442_, _20439_);
  and _71096_ (_20444_, _20443_, _06926_);
  and _71097_ (_20445_, _20377_, _06568_);
  or _71098_ (_20446_, _20445_, _06278_);
  or _71099_ (_20447_, _20446_, _20444_);
  and _71100_ (_20448_, _15329_, _07914_);
  or _71101_ (_20450_, _20371_, _06279_);
  or _71102_ (_20451_, _20450_, _20448_);
  and _71103_ (_20452_, _20451_, _01347_);
  and _71104_ (_20453_, _20452_, _20447_);
  or _71105_ (_20454_, _20453_, _20370_);
  and _71106_ (_43183_, _20454_, _42618_);
  and _71107_ (_20455_, _01351_, \oc8051_golden_model_1.TMOD [5]);
  and _71108_ (_20456_, _11457_, \oc8051_golden_model_1.TMOD [5]);
  nor _71109_ (_20457_, _08244_, _11457_);
  or _71110_ (_20458_, _20457_, _20456_);
  or _71111_ (_20460_, _20458_, _07215_);
  and _71112_ (_20461_, _15358_, _07914_);
  or _71113_ (_20462_, _20461_, _20456_);
  or _71114_ (_20463_, _20462_, _07151_);
  and _71115_ (_20464_, _07914_, \oc8051_golden_model_1.ACC [5]);
  or _71116_ (_20465_, _20464_, _20456_);
  and _71117_ (_20466_, _20465_, _07141_);
  and _71118_ (_20467_, _07142_, \oc8051_golden_model_1.TMOD [5]);
  or _71119_ (_20468_, _20467_, _06341_);
  or _71120_ (_20469_, _20468_, _20466_);
  and _71121_ (_20471_, _20469_, _07166_);
  and _71122_ (_20472_, _20471_, _20463_);
  and _71123_ (_20473_, _20458_, _06461_);
  or _71124_ (_20474_, _20473_, _20472_);
  and _71125_ (_20475_, _20474_, _06465_);
  and _71126_ (_20476_, _20465_, _06464_);
  or _71127_ (_20477_, _20476_, _10080_);
  or _71128_ (_20478_, _20477_, _20475_);
  and _71129_ (_20479_, _20478_, _20460_);
  or _71130_ (_20480_, _20479_, _07460_);
  and _71131_ (_20482_, _09447_, _07914_);
  or _71132_ (_20483_, _20456_, _07208_);
  or _71133_ (_20484_, _20483_, _20482_);
  and _71134_ (_20485_, _20484_, _05982_);
  and _71135_ (_20486_, _20485_, _20480_);
  and _71136_ (_20487_, _15459_, _07914_);
  or _71137_ (_20488_, _20487_, _20456_);
  and _71138_ (_20489_, _20488_, _10094_);
  or _71139_ (_20490_, _20489_, _06218_);
  or _71140_ (_20491_, _20490_, _20486_);
  and _71141_ (_20493_, _08946_, _07914_);
  or _71142_ (_20494_, _20493_, _20456_);
  or _71143_ (_20495_, _20494_, _06219_);
  and _71144_ (_20496_, _20495_, _20491_);
  or _71145_ (_20497_, _20496_, _06369_);
  and _71146_ (_20498_, _15353_, _07914_);
  or _71147_ (_20499_, _20498_, _20456_);
  or _71148_ (_20500_, _20499_, _07237_);
  and _71149_ (_20501_, _20500_, _07240_);
  and _71150_ (_20502_, _20501_, _20497_);
  and _71151_ (_20504_, _11250_, _07914_);
  or _71152_ (_20505_, _20504_, _20456_);
  and _71153_ (_20506_, _20505_, _06536_);
  or _71154_ (_20507_, _20506_, _20502_);
  and _71155_ (_20508_, _20507_, _07242_);
  or _71156_ (_20509_, _20456_, _08247_);
  and _71157_ (_20510_, _20494_, _06375_);
  and _71158_ (_20511_, _20510_, _20509_);
  or _71159_ (_20512_, _20511_, _20508_);
  and _71160_ (_20513_, _20512_, _07234_);
  and _71161_ (_20515_, _20465_, _06545_);
  and _71162_ (_20516_, _20515_, _20509_);
  or _71163_ (_20517_, _20516_, _06366_);
  or _71164_ (_20518_, _20517_, _20513_);
  and _71165_ (_20519_, _15350_, _07914_);
  or _71166_ (_20520_, _20456_, _09056_);
  or _71167_ (_20521_, _20520_, _20519_);
  and _71168_ (_20522_, _20521_, _09061_);
  and _71169_ (_20523_, _20522_, _20518_);
  nor _71170_ (_20524_, _11249_, _11457_);
  or _71171_ (_20526_, _20524_, _20456_);
  and _71172_ (_20527_, _20526_, _06528_);
  or _71173_ (_20528_, _20527_, _20523_);
  and _71174_ (_20529_, _20528_, _06926_);
  and _71175_ (_20530_, _20462_, _06568_);
  or _71176_ (_20531_, _20530_, _06278_);
  or _71177_ (_20532_, _20531_, _20529_);
  and _71178_ (_20533_, _15532_, _07914_);
  or _71179_ (_20534_, _20456_, _06279_);
  or _71180_ (_20535_, _20534_, _20533_);
  and _71181_ (_20537_, _20535_, _01347_);
  and _71182_ (_20538_, _20537_, _20532_);
  or _71183_ (_20539_, _20538_, _20455_);
  and _71184_ (_43184_, _20539_, _42618_);
  and _71185_ (_20540_, _01351_, \oc8051_golden_model_1.TMOD [6]);
  and _71186_ (_20541_, _11457_, \oc8051_golden_model_1.TMOD [6]);
  and _71187_ (_20542_, _15554_, _07914_);
  or _71188_ (_20543_, _20542_, _20541_);
  or _71189_ (_20544_, _20543_, _07151_);
  and _71190_ (_20545_, _07914_, \oc8051_golden_model_1.ACC [6]);
  or _71191_ (_20547_, _20545_, _20541_);
  and _71192_ (_20548_, _20547_, _07141_);
  and _71193_ (_20549_, _07142_, \oc8051_golden_model_1.TMOD [6]);
  or _71194_ (_20550_, _20549_, _06341_);
  or _71195_ (_20551_, _20550_, _20548_);
  and _71196_ (_20552_, _20551_, _07166_);
  and _71197_ (_20553_, _20552_, _20544_);
  nor _71198_ (_20554_, _08142_, _11457_);
  or _71199_ (_20555_, _20554_, _20541_);
  and _71200_ (_20556_, _20555_, _06461_);
  or _71201_ (_20558_, _20556_, _20553_);
  and _71202_ (_20559_, _20558_, _06465_);
  and _71203_ (_20560_, _20547_, _06464_);
  or _71204_ (_20561_, _20560_, _10080_);
  or _71205_ (_20562_, _20561_, _20559_);
  or _71206_ (_20563_, _20555_, _07215_);
  and _71207_ (_20564_, _20563_, _20562_);
  or _71208_ (_20565_, _20564_, _07460_);
  and _71209_ (_20566_, _09446_, _07914_);
  or _71210_ (_20567_, _20541_, _07208_);
  or _71211_ (_20569_, _20567_, _20566_);
  and _71212_ (_20570_, _20569_, _05982_);
  and _71213_ (_20571_, _20570_, _20565_);
  and _71214_ (_20572_, _15657_, _07914_);
  or _71215_ (_20573_, _20572_, _20541_);
  and _71216_ (_20574_, _20573_, _10094_);
  or _71217_ (_20575_, _20574_, _06218_);
  or _71218_ (_20576_, _20575_, _20571_);
  and _71219_ (_20577_, _15664_, _07914_);
  or _71220_ (_20578_, _20577_, _20541_);
  or _71221_ (_20580_, _20578_, _06219_);
  and _71222_ (_20581_, _20580_, _20576_);
  or _71223_ (_20582_, _20581_, _06369_);
  and _71224_ (_20583_, _15549_, _07914_);
  or _71225_ (_20584_, _20583_, _20541_);
  or _71226_ (_20585_, _20584_, _07237_);
  and _71227_ (_20586_, _20585_, _07240_);
  and _71228_ (_20587_, _20586_, _20582_);
  and _71229_ (_20588_, _11247_, _07914_);
  or _71230_ (_20589_, _20588_, _20541_);
  and _71231_ (_20591_, _20589_, _06536_);
  or _71232_ (_20592_, _20591_, _20587_);
  and _71233_ (_20593_, _20592_, _07242_);
  or _71234_ (_20594_, _20541_, _08145_);
  and _71235_ (_20595_, _20578_, _06375_);
  and _71236_ (_20596_, _20595_, _20594_);
  or _71237_ (_20597_, _20596_, _20593_);
  and _71238_ (_20598_, _20597_, _07234_);
  and _71239_ (_20599_, _20547_, _06545_);
  and _71240_ (_20600_, _20599_, _20594_);
  or _71241_ (_20602_, _20600_, _06366_);
  or _71242_ (_20603_, _20602_, _20598_);
  and _71243_ (_20604_, _15546_, _07914_);
  or _71244_ (_20605_, _20541_, _09056_);
  or _71245_ (_20606_, _20605_, _20604_);
  and _71246_ (_20607_, _20606_, _09061_);
  and _71247_ (_20608_, _20607_, _20603_);
  nor _71248_ (_20609_, _11246_, _11457_);
  or _71249_ (_20610_, _20609_, _20541_);
  and _71250_ (_20611_, _20610_, _06528_);
  or _71251_ (_20613_, _20611_, _20608_);
  and _71252_ (_20614_, _20613_, _06926_);
  and _71253_ (_20615_, _20543_, _06568_);
  or _71254_ (_20616_, _20615_, _06278_);
  or _71255_ (_20617_, _20616_, _20614_);
  and _71256_ (_20618_, _15734_, _07914_);
  or _71257_ (_20619_, _20541_, _06279_);
  or _71258_ (_20620_, _20619_, _20618_);
  and _71259_ (_20621_, _20620_, _01347_);
  and _71260_ (_20622_, _20621_, _20617_);
  or _71261_ (_20624_, _20622_, _20540_);
  and _71262_ (_43185_, _20624_, _42618_);
  not _71263_ (_20625_, \oc8051_golden_model_1.DPL [0]);
  nor _71264_ (_20626_, _01347_, _20625_);
  and _71265_ (_20627_, _07960_, \oc8051_golden_model_1.ACC [0]);
  and _71266_ (_20628_, _20627_, _08390_);
  nor _71267_ (_20629_, _07960_, _20625_);
  or _71268_ (_20630_, _20629_, _07234_);
  or _71269_ (_20631_, _20630_, _20628_);
  and _71270_ (_20632_, _09392_, _07960_);
  or _71271_ (_20634_, _20632_, _20629_);
  and _71272_ (_20635_, _20634_, _07460_);
  and _71273_ (_20636_, _07960_, _07133_);
  or _71274_ (_20637_, _20636_, _20629_);
  or _71275_ (_20638_, _20637_, _07166_);
  nor _71276_ (_20639_, _08390_, _11537_);
  or _71277_ (_20640_, _20639_, _20629_);
  and _71278_ (_20641_, _20640_, _06341_);
  nor _71279_ (_20642_, _07141_, _20625_);
  or _71280_ (_20643_, _20629_, _20627_);
  and _71281_ (_20645_, _20643_, _07141_);
  or _71282_ (_20646_, _20645_, _20642_);
  and _71283_ (_20647_, _20646_, _07151_);
  or _71284_ (_20648_, _20647_, _06461_);
  or _71285_ (_20649_, _20648_, _20641_);
  and _71286_ (_20650_, _20649_, _20638_);
  or _71287_ (_20651_, _20650_, _06464_);
  or _71288_ (_20652_, _20643_, _06465_);
  and _71289_ (_20653_, _20652_, _11562_);
  and _71290_ (_20654_, _20653_, _20651_);
  and _71291_ (_20656_, _11561_, _20625_);
  or _71292_ (_20657_, _20656_, _20654_);
  and _71293_ (_20658_, _20657_, _06374_);
  nor _71294_ (_20659_, _06872_, _06374_);
  or _71295_ (_20660_, _20659_, _10080_);
  or _71296_ (_20661_, _20660_, _20658_);
  or _71297_ (_20662_, _20637_, _07215_);
  and _71298_ (_20663_, _20662_, _07208_);
  and _71299_ (_20664_, _20663_, _20661_);
  or _71300_ (_20665_, _20664_, _10094_);
  or _71301_ (_20666_, _20665_, _20635_);
  and _71302_ (_20667_, _14467_, _07960_);
  or _71303_ (_20668_, _20629_, _05982_);
  or _71304_ (_20669_, _20668_, _20667_);
  and _71305_ (_20670_, _20669_, _06219_);
  and _71306_ (_20671_, _20670_, _20666_);
  and _71307_ (_20672_, _07960_, _08954_);
  or _71308_ (_20673_, _20672_, _20629_);
  and _71309_ (_20674_, _20673_, _06218_);
  or _71310_ (_20675_, _20674_, _06369_);
  or _71311_ (_20677_, _20675_, _20671_);
  and _71312_ (_20678_, _14366_, _07960_);
  or _71313_ (_20679_, _20678_, _20629_);
  or _71314_ (_20680_, _20679_, _07237_);
  and _71315_ (_20681_, _20680_, _07240_);
  and _71316_ (_20682_, _20681_, _20677_);
  nor _71317_ (_20683_, _12580_, _11537_);
  or _71318_ (_20684_, _20683_, _20629_);
  nor _71319_ (_20685_, _20628_, _07240_);
  and _71320_ (_20686_, _20685_, _20684_);
  or _71321_ (_20689_, _20686_, _20682_);
  and _71322_ (_20690_, _20689_, _07242_);
  nand _71323_ (_20691_, _20673_, _06375_);
  nor _71324_ (_20692_, _20691_, _20639_);
  or _71325_ (_20693_, _20692_, _06545_);
  or _71326_ (_20694_, _20693_, _20690_);
  and _71327_ (_20695_, _20694_, _20631_);
  or _71328_ (_20696_, _20695_, _06366_);
  and _71329_ (_20697_, _14363_, _07960_);
  or _71330_ (_20698_, _20697_, _20629_);
  or _71331_ (_20700_, _20698_, _09056_);
  and _71332_ (_20701_, _20700_, _09061_);
  and _71333_ (_20702_, _20701_, _20696_);
  and _71334_ (_20703_, _20684_, _06528_);
  or _71335_ (_20704_, _20703_, _19502_);
  or _71336_ (_20705_, _20704_, _20702_);
  or _71337_ (_20706_, _20640_, _06661_);
  and _71338_ (_20707_, _20706_, _01347_);
  and _71339_ (_20708_, _20707_, _20705_);
  or _71340_ (_20709_, _20708_, _20626_);
  and _71341_ (_43187_, _20709_, _42618_);
  not _71342_ (_20710_, \oc8051_golden_model_1.DPL [1]);
  nor _71343_ (_20711_, _01347_, _20710_);
  or _71344_ (_20712_, _09451_, _11537_);
  or _71345_ (_20713_, _07960_, \oc8051_golden_model_1.DPL [1]);
  and _71346_ (_20714_, _20713_, _07460_);
  and _71347_ (_20715_, _20714_, _20712_);
  nor _71348_ (_20716_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor _71349_ (_20717_, _20716_, _11566_);
  and _71350_ (_20718_, _20717_, _11561_);
  and _71351_ (_20720_, _14562_, _07960_);
  not _71352_ (_20721_, _20720_);
  and _71353_ (_20722_, _20721_, _20713_);
  or _71354_ (_20723_, _20722_, _07151_);
  nor _71355_ (_20724_, _07960_, _20710_);
  and _71356_ (_20725_, _07960_, \oc8051_golden_model_1.ACC [1]);
  or _71357_ (_20726_, _20725_, _20724_);
  and _71358_ (_20727_, _20726_, _07141_);
  nor _71359_ (_20728_, _07141_, _20710_);
  or _71360_ (_20729_, _20728_, _06341_);
  or _71361_ (_20732_, _20729_, _20727_);
  and _71362_ (_20733_, _20732_, _07166_);
  and _71363_ (_20734_, _20733_, _20723_);
  nor _71364_ (_20735_, _11537_, _07357_);
  or _71365_ (_20736_, _20735_, _20724_);
  and _71366_ (_20737_, _20736_, _06461_);
  or _71367_ (_20738_, _20737_, _06464_);
  or _71368_ (_20739_, _20738_, _20734_);
  or _71369_ (_20740_, _20726_, _06465_);
  and _71370_ (_20741_, _20740_, _11562_);
  and _71371_ (_20742_, _20741_, _20739_);
  or _71372_ (_20743_, _20742_, _20718_);
  and _71373_ (_20744_, _20743_, _06374_);
  nor _71374_ (_20745_, _07038_, _06374_);
  or _71375_ (_20746_, _20745_, _10080_);
  or _71376_ (_20747_, _20746_, _20744_);
  or _71377_ (_20748_, _20736_, _07215_);
  and _71378_ (_20749_, _20748_, _07208_);
  and _71379_ (_20750_, _20749_, _20747_);
  or _71380_ (_20751_, _20750_, _20715_);
  and _71381_ (_20753_, _20751_, _05982_);
  or _71382_ (_20754_, _14653_, _11537_);
  and _71383_ (_20755_, _20713_, _10094_);
  and _71384_ (_20756_, _20755_, _20754_);
  or _71385_ (_20757_, _20756_, _20753_);
  and _71386_ (_20758_, _20757_, _06219_);
  nand _71387_ (_20759_, _07960_, _07038_);
  and _71388_ (_20760_, _20713_, _06218_);
  and _71389_ (_20761_, _20760_, _20759_);
  or _71390_ (_20762_, _20761_, _20758_);
  and _71391_ (_20765_, _20762_, _07237_);
  or _71392_ (_20766_, _14668_, _11537_);
  and _71393_ (_20767_, _20713_, _06369_);
  and _71394_ (_20768_, _20767_, _20766_);
  or _71395_ (_20769_, _20768_, _06536_);
  or _71396_ (_20770_, _20769_, _20765_);
  nor _71397_ (_20771_, _11261_, _11537_);
  or _71398_ (_20772_, _20771_, _20724_);
  nand _71399_ (_20773_, _11260_, _07960_);
  and _71400_ (_20774_, _20773_, _20772_);
  or _71401_ (_20776_, _20774_, _07240_);
  and _71402_ (_20777_, _20776_, _07242_);
  and _71403_ (_20778_, _20777_, _20770_);
  or _71404_ (_20779_, _14666_, _11537_);
  and _71405_ (_20780_, _20713_, _06375_);
  and _71406_ (_20781_, _20780_, _20779_);
  or _71407_ (_20782_, _20781_, _06545_);
  or _71408_ (_20783_, _20782_, _20778_);
  nor _71409_ (_20784_, _20724_, _07234_);
  nand _71410_ (_20785_, _20784_, _20773_);
  and _71411_ (_20787_, _20785_, _09056_);
  and _71412_ (_20788_, _20787_, _20783_);
  or _71413_ (_20789_, _20759_, _08341_);
  and _71414_ (_20790_, _20713_, _06366_);
  and _71415_ (_20791_, _20790_, _20789_);
  or _71416_ (_20792_, _20791_, _06528_);
  or _71417_ (_20793_, _20792_, _20788_);
  or _71418_ (_20794_, _20772_, _09061_);
  and _71419_ (_20795_, _20794_, _06926_);
  and _71420_ (_20796_, _20795_, _20793_);
  and _71421_ (_20798_, _20722_, _06568_);
  or _71422_ (_20799_, _20798_, _06278_);
  or _71423_ (_20800_, _20799_, _20796_);
  or _71424_ (_20801_, _20724_, _06279_);
  or _71425_ (_20802_, _20801_, _20720_);
  and _71426_ (_20803_, _20802_, _01347_);
  and _71427_ (_20804_, _20803_, _20800_);
  or _71428_ (_20805_, _20804_, _20711_);
  and _71429_ (_43188_, _20805_, _42618_);
  not _71430_ (_20806_, \oc8051_golden_model_1.DPL [2]);
  nor _71431_ (_20807_, _01347_, _20806_);
  nor _71432_ (_20808_, _07960_, _20806_);
  nor _71433_ (_20809_, _11537_, _07776_);
  or _71434_ (_20810_, _20809_, _20808_);
  or _71435_ (_20811_, _20810_, _07215_);
  or _71436_ (_20812_, _20810_, _07166_);
  and _71437_ (_20813_, _14770_, _07960_);
  or _71438_ (_20814_, _20813_, _20808_);
  and _71439_ (_20815_, _20814_, _06341_);
  nor _71440_ (_20816_, _07141_, _20806_);
  and _71441_ (_20819_, _07960_, \oc8051_golden_model_1.ACC [2]);
  or _71442_ (_20820_, _20819_, _20808_);
  and _71443_ (_20821_, _20820_, _07141_);
  or _71444_ (_20822_, _20821_, _20816_);
  and _71445_ (_20823_, _20822_, _07151_);
  or _71446_ (_20824_, _20823_, _06461_);
  or _71447_ (_20825_, _20824_, _20815_);
  and _71448_ (_20826_, _20825_, _20812_);
  or _71449_ (_20827_, _20826_, _06464_);
  or _71450_ (_20828_, _20820_, _06465_);
  and _71451_ (_20830_, _20828_, _11562_);
  and _71452_ (_20831_, _20830_, _20827_);
  nor _71453_ (_20832_, _11566_, \oc8051_golden_model_1.DPL [2]);
  nor _71454_ (_20833_, _20832_, _11567_);
  and _71455_ (_20834_, _20833_, _11561_);
  or _71456_ (_20835_, _20834_, _20831_);
  and _71457_ (_20836_, _20835_, _06374_);
  nor _71458_ (_20837_, _06697_, _06374_);
  or _71459_ (_20838_, _20837_, _10080_);
  or _71460_ (_20839_, _20838_, _20836_);
  and _71461_ (_20841_, _20839_, _20811_);
  or _71462_ (_20842_, _20841_, _07460_);
  and _71463_ (_20843_, _09450_, _07960_);
  or _71464_ (_20844_, _20808_, _07208_);
  or _71465_ (_20845_, _20844_, _20843_);
  and _71466_ (_20846_, _20845_, _05982_);
  and _71467_ (_20847_, _20846_, _20842_);
  and _71468_ (_20848_, _14859_, _07960_);
  or _71469_ (_20849_, _20848_, _20808_);
  and _71470_ (_20850_, _20849_, _10094_);
  or _71471_ (_20852_, _20850_, _06218_);
  or _71472_ (_20853_, _20852_, _20847_);
  and _71473_ (_20854_, _07960_, _08973_);
  or _71474_ (_20855_, _20854_, _20808_);
  or _71475_ (_20856_, _20855_, _06219_);
  and _71476_ (_20857_, _20856_, _20853_);
  or _71477_ (_20858_, _20857_, _06369_);
  and _71478_ (_20859_, _14751_, _07960_);
  or _71479_ (_20860_, _20859_, _20808_);
  or _71480_ (_20861_, _20860_, _07237_);
  and _71481_ (_20863_, _20861_, _07240_);
  and _71482_ (_20864_, _20863_, _20858_);
  and _71483_ (_20865_, _11259_, _07960_);
  or _71484_ (_20866_, _20865_, _20808_);
  and _71485_ (_20867_, _20866_, _06536_);
  or _71486_ (_20868_, _20867_, _20864_);
  and _71487_ (_20869_, _20868_, _07242_);
  or _71488_ (_20870_, _20808_, _08440_);
  and _71489_ (_20871_, _20855_, _06375_);
  and _71490_ (_20872_, _20871_, _20870_);
  or _71491_ (_20874_, _20872_, _20869_);
  and _71492_ (_20875_, _20874_, _07234_);
  and _71493_ (_20876_, _20820_, _06545_);
  and _71494_ (_20877_, _20876_, _20870_);
  or _71495_ (_20878_, _20877_, _06366_);
  or _71496_ (_20879_, _20878_, _20875_);
  and _71497_ (_20880_, _14748_, _07960_);
  or _71498_ (_20881_, _20808_, _09056_);
  or _71499_ (_20882_, _20881_, _20880_);
  and _71500_ (_20883_, _20882_, _09061_);
  and _71501_ (_20885_, _20883_, _20879_);
  nor _71502_ (_20886_, _11258_, _11537_);
  or _71503_ (_20887_, _20886_, _20808_);
  and _71504_ (_20888_, _20887_, _06528_);
  or _71505_ (_20889_, _20888_, _20885_);
  and _71506_ (_20890_, _20889_, _06926_);
  and _71507_ (_20891_, _20814_, _06568_);
  or _71508_ (_20892_, _20891_, _06278_);
  or _71509_ (_20893_, _20892_, _20890_);
  and _71510_ (_20894_, _14926_, _07960_);
  or _71511_ (_20896_, _20808_, _06279_);
  or _71512_ (_20897_, _20896_, _20894_);
  and _71513_ (_20898_, _20897_, _01347_);
  and _71514_ (_20899_, _20898_, _20893_);
  or _71515_ (_20900_, _20899_, _20807_);
  and _71516_ (_43189_, _20900_, _42618_);
  not _71517_ (_20901_, \oc8051_golden_model_1.DPL [3]);
  nor _71518_ (_20902_, _01347_, _20901_);
  nor _71519_ (_20903_, _07960_, _20901_);
  nor _71520_ (_20904_, _11537_, _07594_);
  or _71521_ (_20906_, _20904_, _20903_);
  or _71522_ (_20907_, _20906_, _07215_);
  and _71523_ (_20908_, _14953_, _07960_);
  or _71524_ (_20909_, _20908_, _20903_);
  or _71525_ (_20910_, _20909_, _07151_);
  and _71526_ (_20911_, _07960_, \oc8051_golden_model_1.ACC [3]);
  or _71527_ (_20912_, _20911_, _20903_);
  and _71528_ (_20913_, _20912_, _07141_);
  nor _71529_ (_20914_, _07141_, _20901_);
  or _71530_ (_20915_, _20914_, _06341_);
  or _71531_ (_20917_, _20915_, _20913_);
  and _71532_ (_20918_, _20917_, _07166_);
  and _71533_ (_20919_, _20918_, _20910_);
  and _71534_ (_20920_, _20906_, _06461_);
  or _71535_ (_20921_, _20920_, _06464_);
  or _71536_ (_20922_, _20921_, _20919_);
  or _71537_ (_20923_, _20912_, _06465_);
  and _71538_ (_20924_, _20923_, _11562_);
  and _71539_ (_20925_, _20924_, _20922_);
  nor _71540_ (_20926_, _11567_, \oc8051_golden_model_1.DPL [3]);
  nor _71541_ (_20928_, _20926_, _11568_);
  and _71542_ (_20929_, _20928_, _11561_);
  or _71543_ (_20930_, _20929_, _20925_);
  and _71544_ (_20931_, _20930_, _06374_);
  nor _71545_ (_20932_, _06452_, _06374_);
  or _71546_ (_20933_, _20932_, _10080_);
  or _71547_ (_20934_, _20933_, _20931_);
  and _71548_ (_20935_, _20934_, _20907_);
  or _71549_ (_20936_, _20935_, _07460_);
  and _71550_ (_20937_, _09449_, _07960_);
  or _71551_ (_20938_, _20903_, _07208_);
  or _71552_ (_20939_, _20938_, _20937_);
  and _71553_ (_20940_, _20939_, _05982_);
  and _71554_ (_20941_, _20940_, _20936_);
  and _71555_ (_20942_, _15048_, _07960_);
  or _71556_ (_20943_, _20942_, _20903_);
  and _71557_ (_20944_, _20943_, _10094_);
  or _71558_ (_20945_, _20944_, _06218_);
  or _71559_ (_20946_, _20945_, _20941_);
  and _71560_ (_20947_, _07960_, _08930_);
  or _71561_ (_20950_, _20947_, _20903_);
  or _71562_ (_20951_, _20950_, _06219_);
  and _71563_ (_20952_, _20951_, _20946_);
  or _71564_ (_20953_, _20952_, _06369_);
  and _71565_ (_20954_, _14943_, _07960_);
  or _71566_ (_20955_, _20954_, _20903_);
  or _71567_ (_20956_, _20955_, _07237_);
  and _71568_ (_20957_, _20956_, _07240_);
  and _71569_ (_20958_, _20957_, _20953_);
  and _71570_ (_20959_, _12577_, _07960_);
  or _71571_ (_20961_, _20959_, _20903_);
  and _71572_ (_20962_, _20961_, _06536_);
  or _71573_ (_20963_, _20962_, _20958_);
  and _71574_ (_20964_, _20963_, _07242_);
  or _71575_ (_20965_, _20903_, _08292_);
  and _71576_ (_20966_, _20950_, _06375_);
  and _71577_ (_20967_, _20966_, _20965_);
  or _71578_ (_20968_, _20967_, _20964_);
  and _71579_ (_20969_, _20968_, _07234_);
  and _71580_ (_20970_, _20912_, _06545_);
  and _71581_ (_20972_, _20970_, _20965_);
  or _71582_ (_20973_, _20972_, _06366_);
  or _71583_ (_20974_, _20973_, _20969_);
  and _71584_ (_20975_, _14940_, _07960_);
  or _71585_ (_20976_, _20903_, _09056_);
  or _71586_ (_20977_, _20976_, _20975_);
  and _71587_ (_20978_, _20977_, _09061_);
  and _71588_ (_20979_, _20978_, _20974_);
  nor _71589_ (_20980_, _11256_, _11537_);
  or _71590_ (_20981_, _20980_, _20903_);
  and _71591_ (_20983_, _20981_, _06528_);
  or _71592_ (_20984_, _20983_, _20979_);
  and _71593_ (_20985_, _20984_, _06926_);
  and _71594_ (_20986_, _20909_, _06568_);
  or _71595_ (_20987_, _20986_, _06278_);
  or _71596_ (_20988_, _20987_, _20985_);
  and _71597_ (_20989_, _15128_, _07960_);
  or _71598_ (_20990_, _20903_, _06279_);
  or _71599_ (_20991_, _20990_, _20989_);
  and _71600_ (_20992_, _20991_, _01347_);
  and _71601_ (_20994_, _20992_, _20988_);
  or _71602_ (_20995_, _20994_, _20902_);
  and _71603_ (_43190_, _20995_, _42618_);
  not _71604_ (_20996_, \oc8051_golden_model_1.DPL [4]);
  nor _71605_ (_20997_, _01347_, _20996_);
  nor _71606_ (_20998_, _07960_, _20996_);
  nor _71607_ (_20999_, _08541_, _11537_);
  or _71608_ (_21000_, _20999_, _20998_);
  or _71609_ (_21001_, _21000_, _07215_);
  and _71610_ (_21002_, _15162_, _07960_);
  or _71611_ (_21004_, _21002_, _20998_);
  or _71612_ (_21005_, _21004_, _07151_);
  and _71613_ (_21006_, _07960_, \oc8051_golden_model_1.ACC [4]);
  or _71614_ (_21007_, _21006_, _20998_);
  and _71615_ (_21008_, _21007_, _07141_);
  nor _71616_ (_21009_, _07141_, _20996_);
  or _71617_ (_21010_, _21009_, _06341_);
  or _71618_ (_21011_, _21010_, _21008_);
  and _71619_ (_21012_, _21011_, _07166_);
  and _71620_ (_21013_, _21012_, _21005_);
  and _71621_ (_21015_, _21000_, _06461_);
  or _71622_ (_21016_, _21015_, _06464_);
  or _71623_ (_21017_, _21016_, _21013_);
  or _71624_ (_21018_, _21007_, _06465_);
  and _71625_ (_21019_, _21018_, _11562_);
  and _71626_ (_21020_, _21019_, _21017_);
  nor _71627_ (_21021_, _11568_, \oc8051_golden_model_1.DPL [4]);
  nor _71628_ (_21022_, _21021_, _11569_);
  and _71629_ (_21023_, _21022_, _11561_);
  or _71630_ (_21024_, _21023_, _21020_);
  and _71631_ (_21026_, _21024_, _06374_);
  nor _71632_ (_21027_, _08892_, _06374_);
  or _71633_ (_21028_, _21027_, _10080_);
  or _71634_ (_21029_, _21028_, _21026_);
  and _71635_ (_21030_, _21029_, _21001_);
  or _71636_ (_21031_, _21030_, _07460_);
  and _71637_ (_21032_, _09448_, _07960_);
  or _71638_ (_21033_, _20998_, _07208_);
  or _71639_ (_21034_, _21033_, _21032_);
  and _71640_ (_21035_, _21034_, _05982_);
  and _71641_ (_21037_, _21035_, _21031_);
  and _71642_ (_21038_, _15254_, _07960_);
  or _71643_ (_21039_, _21038_, _20998_);
  and _71644_ (_21040_, _21039_, _10094_);
  or _71645_ (_21041_, _21040_, _06218_);
  or _71646_ (_21042_, _21041_, _21037_);
  and _71647_ (_21043_, _08959_, _07960_);
  or _71648_ (_21044_, _21043_, _20998_);
  or _71649_ (_21045_, _21044_, _06219_);
  and _71650_ (_21046_, _21045_, _21042_);
  or _71651_ (_21048_, _21046_, _06369_);
  and _71652_ (_21049_, _15269_, _07960_);
  or _71653_ (_21050_, _21049_, _20998_);
  or _71654_ (_21051_, _21050_, _07237_);
  and _71655_ (_21052_, _21051_, _07240_);
  and _71656_ (_21053_, _21052_, _21048_);
  and _71657_ (_21054_, _11254_, _07960_);
  or _71658_ (_21055_, _21054_, _20998_);
  and _71659_ (_21056_, _21055_, _06536_);
  or _71660_ (_21057_, _21056_, _21053_);
  and _71661_ (_21059_, _21057_, _07242_);
  or _71662_ (_21060_, _20998_, _08544_);
  and _71663_ (_21061_, _21044_, _06375_);
  and _71664_ (_21062_, _21061_, _21060_);
  or _71665_ (_21063_, _21062_, _21059_);
  and _71666_ (_21064_, _21063_, _07234_);
  and _71667_ (_21065_, _21007_, _06545_);
  and _71668_ (_21066_, _21065_, _21060_);
  or _71669_ (_21067_, _21066_, _06366_);
  or _71670_ (_21068_, _21067_, _21064_);
  and _71671_ (_21070_, _15266_, _07960_);
  or _71672_ (_21071_, _20998_, _09056_);
  or _71673_ (_21072_, _21071_, _21070_);
  and _71674_ (_21073_, _21072_, _09061_);
  and _71675_ (_21074_, _21073_, _21068_);
  nor _71676_ (_21075_, _11253_, _11537_);
  or _71677_ (_21076_, _21075_, _20998_);
  and _71678_ (_21077_, _21076_, _06528_);
  or _71679_ (_21078_, _21077_, _21074_);
  and _71680_ (_21079_, _21078_, _06926_);
  and _71681_ (_21081_, _21004_, _06568_);
  or _71682_ (_21082_, _21081_, _06278_);
  or _71683_ (_21083_, _21082_, _21079_);
  and _71684_ (_21084_, _15329_, _07960_);
  or _71685_ (_21085_, _20998_, _06279_);
  or _71686_ (_21086_, _21085_, _21084_);
  and _71687_ (_21087_, _21086_, _01347_);
  and _71688_ (_21088_, _21087_, _21083_);
  or _71689_ (_21089_, _21088_, _20997_);
  and _71690_ (_43191_, _21089_, _42618_);
  not _71691_ (_21091_, \oc8051_golden_model_1.DPL [5]);
  nor _71692_ (_21092_, _01347_, _21091_);
  nor _71693_ (_21093_, _07960_, _21091_);
  nor _71694_ (_21094_, _08244_, _11537_);
  or _71695_ (_21095_, _21094_, _21093_);
  or _71696_ (_21096_, _21095_, _07215_);
  and _71697_ (_21097_, _15358_, _07960_);
  or _71698_ (_21098_, _21097_, _21093_);
  or _71699_ (_21099_, _21098_, _07151_);
  and _71700_ (_21100_, _07960_, \oc8051_golden_model_1.ACC [5]);
  or _71701_ (_21102_, _21100_, _21093_);
  and _71702_ (_21103_, _21102_, _07141_);
  nor _71703_ (_21104_, _07141_, _21091_);
  or _71704_ (_21105_, _21104_, _06341_);
  or _71705_ (_21106_, _21105_, _21103_);
  and _71706_ (_21107_, _21106_, _07166_);
  and _71707_ (_21108_, _21107_, _21099_);
  and _71708_ (_21109_, _21095_, _06461_);
  or _71709_ (_21110_, _21109_, _06464_);
  or _71710_ (_21111_, _21110_, _21108_);
  or _71711_ (_21112_, _21102_, _06465_);
  and _71712_ (_21113_, _21112_, _11562_);
  and _71713_ (_21114_, _21113_, _21111_);
  nor _71714_ (_21115_, _11569_, \oc8051_golden_model_1.DPL [5]);
  nor _71715_ (_21116_, _21115_, _11570_);
  and _71716_ (_21117_, _21116_, _11561_);
  or _71717_ (_21118_, _21117_, _21114_);
  and _71718_ (_21119_, _21118_, _06374_);
  nor _71719_ (_21120_, _08926_, _06374_);
  or _71720_ (_21121_, _21120_, _10080_);
  or _71721_ (_21124_, _21121_, _21119_);
  and _71722_ (_21125_, _21124_, _21096_);
  or _71723_ (_21126_, _21125_, _07460_);
  and _71724_ (_21127_, _09447_, _07960_);
  or _71725_ (_21128_, _21093_, _07208_);
  or _71726_ (_21129_, _21128_, _21127_);
  and _71727_ (_21130_, _21129_, _05982_);
  and _71728_ (_21131_, _21130_, _21126_);
  and _71729_ (_21132_, _15459_, _07960_);
  or _71730_ (_21133_, _21132_, _21093_);
  and _71731_ (_21135_, _21133_, _10094_);
  or _71732_ (_21136_, _21135_, _06218_);
  or _71733_ (_21137_, _21136_, _21131_);
  and _71734_ (_21138_, _08946_, _07960_);
  or _71735_ (_21139_, _21138_, _21093_);
  or _71736_ (_21140_, _21139_, _06219_);
  and _71737_ (_21141_, _21140_, _21137_);
  or _71738_ (_21142_, _21141_, _06369_);
  and _71739_ (_21143_, _15353_, _07960_);
  or _71740_ (_21144_, _21143_, _21093_);
  or _71741_ (_21146_, _21144_, _07237_);
  and _71742_ (_21147_, _21146_, _07240_);
  and _71743_ (_21148_, _21147_, _21142_);
  and _71744_ (_21149_, _11250_, _07960_);
  or _71745_ (_21150_, _21149_, _21093_);
  and _71746_ (_21151_, _21150_, _06536_);
  or _71747_ (_21152_, _21151_, _21148_);
  and _71748_ (_21153_, _21152_, _07242_);
  or _71749_ (_21154_, _21093_, _08247_);
  and _71750_ (_21155_, _21139_, _06375_);
  and _71751_ (_21157_, _21155_, _21154_);
  or _71752_ (_21158_, _21157_, _21153_);
  and _71753_ (_21159_, _21158_, _07234_);
  and _71754_ (_21160_, _21102_, _06545_);
  and _71755_ (_21161_, _21160_, _21154_);
  or _71756_ (_21162_, _21161_, _06366_);
  or _71757_ (_21163_, _21162_, _21159_);
  and _71758_ (_21164_, _15350_, _07960_);
  or _71759_ (_21165_, _21093_, _09056_);
  or _71760_ (_21166_, _21165_, _21164_);
  and _71761_ (_21168_, _21166_, _09061_);
  and _71762_ (_21169_, _21168_, _21163_);
  nor _71763_ (_21170_, _11249_, _11537_);
  or _71764_ (_21171_, _21170_, _21093_);
  and _71765_ (_21172_, _21171_, _06528_);
  or _71766_ (_21173_, _21172_, _21169_);
  and _71767_ (_21174_, _21173_, _06926_);
  and _71768_ (_21175_, _21098_, _06568_);
  or _71769_ (_21176_, _21175_, _06278_);
  or _71770_ (_21177_, _21176_, _21174_);
  and _71771_ (_21179_, _15532_, _07960_);
  or _71772_ (_21180_, _21093_, _06279_);
  or _71773_ (_21181_, _21180_, _21179_);
  and _71774_ (_21182_, _21181_, _01347_);
  and _71775_ (_21183_, _21182_, _21177_);
  or _71776_ (_21184_, _21183_, _21092_);
  and _71777_ (_43192_, _21184_, _42618_);
  not _71778_ (_21185_, \oc8051_golden_model_1.DPL [6]);
  nor _71779_ (_21186_, _01347_, _21185_);
  nor _71780_ (_21187_, _07960_, _21185_);
  nor _71781_ (_21189_, _08142_, _11537_);
  or _71782_ (_21190_, _21189_, _21187_);
  or _71783_ (_21191_, _21190_, _07215_);
  and _71784_ (_21192_, _15554_, _07960_);
  or _71785_ (_21193_, _21192_, _21187_);
  or _71786_ (_21194_, _21193_, _07151_);
  and _71787_ (_21195_, _07960_, \oc8051_golden_model_1.ACC [6]);
  or _71788_ (_21196_, _21195_, _21187_);
  and _71789_ (_21197_, _21196_, _07141_);
  nor _71790_ (_21198_, _07141_, _21185_);
  or _71791_ (_21200_, _21198_, _06341_);
  or _71792_ (_21201_, _21200_, _21197_);
  and _71793_ (_21202_, _21201_, _07166_);
  and _71794_ (_21203_, _21202_, _21194_);
  and _71795_ (_21204_, _21190_, _06461_);
  or _71796_ (_21205_, _21204_, _06464_);
  or _71797_ (_21206_, _21205_, _21203_);
  or _71798_ (_21207_, _21196_, _06465_);
  and _71799_ (_21208_, _21207_, _11562_);
  and _71800_ (_21209_, _21208_, _21206_);
  nor _71801_ (_21211_, _11570_, \oc8051_golden_model_1.DPL [6]);
  nor _71802_ (_21212_, _21211_, _11571_);
  and _71803_ (_21213_, _21212_, _11561_);
  or _71804_ (_21214_, _21213_, _21209_);
  and _71805_ (_21215_, _21214_, _06374_);
  nor _71806_ (_21216_, _08857_, _06374_);
  or _71807_ (_21217_, _21216_, _10080_);
  or _71808_ (_21218_, _21217_, _21215_);
  and _71809_ (_21219_, _21218_, _21191_);
  or _71810_ (_21220_, _21219_, _07460_);
  and _71811_ (_21222_, _09446_, _07960_);
  or _71812_ (_21223_, _21187_, _07208_);
  or _71813_ (_21224_, _21223_, _21222_);
  and _71814_ (_21225_, _21224_, _05982_);
  and _71815_ (_21226_, _21225_, _21220_);
  and _71816_ (_21227_, _15657_, _07960_);
  or _71817_ (_21228_, _21227_, _21187_);
  and _71818_ (_21229_, _21228_, _10094_);
  or _71819_ (_21230_, _21229_, _06218_);
  or _71820_ (_21231_, _21230_, _21226_);
  and _71821_ (_21233_, _15664_, _07960_);
  or _71822_ (_21234_, _21233_, _21187_);
  or _71823_ (_21235_, _21234_, _06219_);
  and _71824_ (_21236_, _21235_, _21231_);
  or _71825_ (_21237_, _21236_, _06369_);
  and _71826_ (_21238_, _15549_, _07960_);
  or _71827_ (_21239_, _21238_, _21187_);
  or _71828_ (_21240_, _21239_, _07237_);
  and _71829_ (_21241_, _21240_, _07240_);
  and _71830_ (_21242_, _21241_, _21237_);
  and _71831_ (_21244_, _11247_, _07960_);
  or _71832_ (_21245_, _21244_, _21187_);
  and _71833_ (_21246_, _21245_, _06536_);
  or _71834_ (_21247_, _21246_, _21242_);
  and _71835_ (_21248_, _21247_, _07242_);
  or _71836_ (_21249_, _21187_, _08145_);
  and _71837_ (_21250_, _21234_, _06375_);
  and _71838_ (_21251_, _21250_, _21249_);
  or _71839_ (_21252_, _21251_, _21248_);
  and _71840_ (_21253_, _21252_, _07234_);
  and _71841_ (_21255_, _21196_, _06545_);
  and _71842_ (_21256_, _21255_, _21249_);
  or _71843_ (_21257_, _21256_, _06366_);
  or _71844_ (_21258_, _21257_, _21253_);
  and _71845_ (_21259_, _15546_, _07960_);
  or _71846_ (_21260_, _21187_, _09056_);
  or _71847_ (_21261_, _21260_, _21259_);
  and _71848_ (_21262_, _21261_, _09061_);
  and _71849_ (_21263_, _21262_, _21258_);
  nor _71850_ (_21264_, _11246_, _11537_);
  or _71851_ (_21266_, _21264_, _21187_);
  and _71852_ (_21267_, _21266_, _06528_);
  or _71853_ (_21268_, _21267_, _21263_);
  and _71854_ (_21269_, _21268_, _06926_);
  and _71855_ (_21270_, _21193_, _06568_);
  or _71856_ (_21271_, _21270_, _06278_);
  or _71857_ (_21272_, _21271_, _21269_);
  and _71858_ (_21273_, _15734_, _07960_);
  or _71859_ (_21274_, _21187_, _06279_);
  or _71860_ (_21275_, _21274_, _21273_);
  and _71861_ (_21277_, _21275_, _01347_);
  and _71862_ (_21278_, _21277_, _21272_);
  or _71863_ (_21279_, _21278_, _21186_);
  and _71864_ (_43193_, _21279_, _42618_);
  nor _71865_ (_21280_, _01347_, _12693_);
  nor _71866_ (_21281_, _07963_, _12693_);
  and _71867_ (_21282_, _07963_, \oc8051_golden_model_1.ACC [0]);
  and _71868_ (_21283_, _21282_, _08390_);
  or _71869_ (_21284_, _21283_, _21281_);
  or _71870_ (_21285_, _21284_, _07234_);
  and _71871_ (_21287_, _09392_, _07963_);
  or _71872_ (_21288_, _21287_, _21281_);
  and _71873_ (_21289_, _21288_, _07460_);
  and _71874_ (_21290_, _08186_, _07133_);
  or _71875_ (_21291_, _21290_, _21281_);
  or _71876_ (_21292_, _21291_, _07166_);
  nor _71877_ (_21293_, _08390_, _11633_);
  or _71878_ (_21294_, _21293_, _21281_);
  and _71879_ (_21295_, _21294_, _06341_);
  nor _71880_ (_21296_, _07141_, _12693_);
  or _71881_ (_21298_, _21282_, _21281_);
  and _71882_ (_21299_, _21298_, _07141_);
  or _71883_ (_21300_, _21299_, _21296_);
  and _71884_ (_21301_, _21300_, _07151_);
  or _71885_ (_21302_, _21301_, _06461_);
  or _71886_ (_21303_, _21302_, _21295_);
  and _71887_ (_21304_, _21303_, _21292_);
  or _71888_ (_21305_, _21304_, _06464_);
  or _71889_ (_21306_, _21298_, _06465_);
  and _71890_ (_21307_, _21306_, _11562_);
  and _71891_ (_21308_, _21307_, _21305_);
  or _71892_ (_21309_, _11573_, \oc8051_golden_model_1.DPH [0]);
  nor _71893_ (_21310_, _11660_, _11562_);
  and _71894_ (_21311_, _21310_, _21309_);
  or _71895_ (_21312_, _21311_, _21308_);
  and _71896_ (_21313_, _21312_, _06374_);
  nor _71897_ (_21314_, _06374_, _06251_);
  or _71898_ (_21315_, _21314_, _10080_);
  or _71899_ (_21316_, _21315_, _21313_);
  or _71900_ (_21317_, _21291_, _07215_);
  and _71901_ (_21320_, _21317_, _07208_);
  and _71902_ (_21321_, _21320_, _21316_);
  or _71903_ (_21322_, _21321_, _10094_);
  or _71904_ (_21323_, _21322_, _21289_);
  and _71905_ (_21324_, _14467_, _08186_);
  or _71906_ (_21325_, _21281_, _05982_);
  or _71907_ (_21326_, _21325_, _21324_);
  and _71908_ (_21327_, _21326_, _06219_);
  and _71909_ (_21328_, _21327_, _21323_);
  and _71910_ (_21329_, _07963_, _08954_);
  or _71911_ (_21331_, _21329_, _21281_);
  and _71912_ (_21332_, _21331_, _06218_);
  or _71913_ (_21333_, _21332_, _06369_);
  or _71914_ (_21334_, _21333_, _21328_);
  and _71915_ (_21335_, _14366_, _07963_);
  or _71916_ (_21336_, _21335_, _21281_);
  or _71917_ (_21337_, _21336_, _07237_);
  and _71918_ (_21338_, _21337_, _07240_);
  and _71919_ (_21339_, _21338_, _21334_);
  nor _71920_ (_21340_, _12580_, _11633_);
  or _71921_ (_21342_, _21340_, _21281_);
  nor _71922_ (_21343_, _21283_, _07240_);
  and _71923_ (_21344_, _21343_, _21342_);
  or _71924_ (_21345_, _21344_, _21339_);
  and _71925_ (_21346_, _21345_, _07242_);
  nand _71926_ (_21347_, _21331_, _06375_);
  nor _71927_ (_21348_, _21347_, _21293_);
  or _71928_ (_21349_, _21348_, _06545_);
  or _71929_ (_21350_, _21349_, _21346_);
  and _71930_ (_21351_, _21350_, _21285_);
  or _71931_ (_21353_, _21351_, _06366_);
  and _71932_ (_21354_, _14363_, _07963_);
  or _71933_ (_21355_, _21354_, _21281_);
  or _71934_ (_21356_, _21355_, _09056_);
  and _71935_ (_21357_, _21356_, _09061_);
  and _71936_ (_21358_, _21357_, _21353_);
  and _71937_ (_21359_, _21342_, _06528_);
  or _71938_ (_21360_, _21359_, _19502_);
  or _71939_ (_21361_, _21360_, _21358_);
  or _71940_ (_21362_, _21294_, _06661_);
  and _71941_ (_21364_, _21362_, _01347_);
  and _71942_ (_21365_, _21364_, _21361_);
  or _71943_ (_21366_, _21365_, _21280_);
  and _71944_ (_43195_, _21366_, _42618_);
  not _71945_ (_21367_, \oc8051_golden_model_1.DPH [1]);
  nor _71946_ (_21368_, _01347_, _21367_);
  or _71947_ (_21369_, _07963_, \oc8051_golden_model_1.DPH [1]);
  and _71948_ (_21370_, _21369_, _06218_);
  nand _71949_ (_21371_, _08186_, _07038_);
  and _71950_ (_21372_, _21371_, _21370_);
  or _71951_ (_21374_, _09451_, _11633_);
  and _71952_ (_21375_, _21369_, _07460_);
  and _71953_ (_21376_, _21375_, _21374_);
  nor _71954_ (_21377_, _11660_, \oc8051_golden_model_1.DPH [1]);
  nor _71955_ (_21378_, _21377_, _11661_);
  and _71956_ (_21379_, _21378_, _11561_);
  and _71957_ (_21380_, _14562_, _08186_);
  not _71958_ (_21381_, _21380_);
  and _71959_ (_21382_, _21381_, _21369_);
  or _71960_ (_21383_, _21382_, _07151_);
  nor _71961_ (_21385_, _07963_, _21367_);
  and _71962_ (_21386_, _07963_, \oc8051_golden_model_1.ACC [1]);
  or _71963_ (_21387_, _21386_, _21385_);
  and _71964_ (_21388_, _21387_, _07141_);
  nor _71965_ (_21389_, _07141_, _21367_);
  or _71966_ (_21390_, _21389_, _06341_);
  or _71967_ (_21391_, _21390_, _21388_);
  and _71968_ (_21392_, _21391_, _07166_);
  and _71969_ (_21393_, _21392_, _21383_);
  nor _71970_ (_21394_, _11633_, _07357_);
  or _71971_ (_21396_, _21394_, _21385_);
  and _71972_ (_21397_, _21396_, _06461_);
  or _71973_ (_21398_, _21397_, _06464_);
  or _71974_ (_21399_, _21398_, _21393_);
  or _71975_ (_21400_, _21387_, _06465_);
  and _71976_ (_21401_, _21400_, _11562_);
  and _71977_ (_21402_, _21401_, _21399_);
  or _71978_ (_21403_, _21402_, _21379_);
  and _71979_ (_21404_, _21403_, _06374_);
  nor _71980_ (_21405_, _07004_, _06374_);
  or _71981_ (_21407_, _21405_, _10080_);
  or _71982_ (_21408_, _21407_, _21404_);
  or _71983_ (_21409_, _21396_, _07215_);
  and _71984_ (_21410_, _21409_, _07208_);
  and _71985_ (_21411_, _21410_, _21408_);
  or _71986_ (_21412_, _21411_, _21376_);
  and _71987_ (_21413_, _21412_, _05982_);
  and _71988_ (_21414_, _14653_, _07963_);
  or _71989_ (_21415_, _21414_, _21385_);
  and _71990_ (_21416_, _21415_, _10094_);
  or _71991_ (_21418_, _21416_, _21413_);
  and _71992_ (_21419_, _21418_, _06219_);
  or _71993_ (_21420_, _21419_, _21372_);
  and _71994_ (_21421_, _21420_, _07237_);
  or _71995_ (_21422_, _14668_, _11633_);
  and _71996_ (_21423_, _21369_, _06369_);
  and _71997_ (_21424_, _21423_, _21422_);
  or _71998_ (_21425_, _21424_, _06536_);
  or _71999_ (_21426_, _21425_, _21421_);
  nor _72000_ (_21427_, _11261_, _11633_);
  or _72001_ (_21429_, _21427_, _21385_);
  nand _72002_ (_21430_, _11260_, _08186_);
  and _72003_ (_21431_, _21430_, _21429_);
  or _72004_ (_21432_, _21431_, _07240_);
  and _72005_ (_21433_, _21432_, _07242_);
  and _72006_ (_21434_, _21433_, _21426_);
  or _72007_ (_21435_, _14666_, _11633_);
  and _72008_ (_21436_, _21369_, _06375_);
  and _72009_ (_21437_, _21436_, _21435_);
  or _72010_ (_21438_, _21437_, _06545_);
  or _72011_ (_21440_, _21438_, _21434_);
  nor _72012_ (_21441_, _21385_, _07234_);
  nand _72013_ (_21442_, _21441_, _21430_);
  and _72014_ (_21443_, _21442_, _09056_);
  and _72015_ (_21444_, _21443_, _21440_);
  or _72016_ (_21445_, _21371_, _08341_);
  and _72017_ (_21446_, _21369_, _06366_);
  and _72018_ (_21447_, _21446_, _21445_);
  or _72019_ (_21448_, _21447_, _06528_);
  or _72020_ (_21449_, _21448_, _21444_);
  or _72021_ (_21451_, _21429_, _09061_);
  and _72022_ (_21452_, _21451_, _06926_);
  and _72023_ (_21453_, _21452_, _21449_);
  and _72024_ (_21454_, _21382_, _06568_);
  or _72025_ (_21455_, _21454_, _06278_);
  or _72026_ (_21456_, _21455_, _21453_);
  or _72027_ (_21457_, _21385_, _06279_);
  or _72028_ (_21458_, _21457_, _21380_);
  and _72029_ (_21459_, _21458_, _01347_);
  and _72030_ (_21460_, _21459_, _21456_);
  or _72031_ (_21462_, _21460_, _21368_);
  and _72032_ (_43196_, _21462_, _42618_);
  and _72033_ (_21463_, _01351_, \oc8051_golden_model_1.DPH [2]);
  and _72034_ (_21464_, _11633_, \oc8051_golden_model_1.DPH [2]);
  nor _72035_ (_21465_, _11633_, _07776_);
  or _72036_ (_21466_, _21465_, _21464_);
  or _72037_ (_21467_, _21466_, _07215_);
  or _72038_ (_21468_, _11661_, \oc8051_golden_model_1.DPH [2]);
  nor _72039_ (_21469_, _11662_, _11562_);
  and _72040_ (_21470_, _21469_, _21468_);
  and _72041_ (_21472_, _14770_, _08186_);
  or _72042_ (_21473_, _21472_, _21464_);
  or _72043_ (_21474_, _21473_, _07151_);
  and _72044_ (_21475_, _07963_, \oc8051_golden_model_1.ACC [2]);
  or _72045_ (_21476_, _21475_, _21464_);
  and _72046_ (_21477_, _21476_, _07141_);
  and _72047_ (_21478_, _07142_, \oc8051_golden_model_1.DPH [2]);
  or _72048_ (_21479_, _21478_, _06341_);
  or _72049_ (_21480_, _21479_, _21477_);
  and _72050_ (_21481_, _21480_, _07166_);
  and _72051_ (_21483_, _21481_, _21474_);
  and _72052_ (_21484_, _21466_, _06461_);
  or _72053_ (_21485_, _21484_, _06464_);
  or _72054_ (_21486_, _21485_, _21483_);
  or _72055_ (_21487_, _21476_, _06465_);
  and _72056_ (_21488_, _21487_, _11562_);
  and _72057_ (_21489_, _21488_, _21486_);
  or _72058_ (_21490_, _21489_, _21470_);
  and _72059_ (_21491_, _21490_, _06374_);
  nor _72060_ (_21492_, _06656_, _06374_);
  or _72061_ (_21494_, _21492_, _10080_);
  or _72062_ (_21495_, _21494_, _21491_);
  and _72063_ (_21496_, _21495_, _21467_);
  or _72064_ (_21497_, _21496_, _07460_);
  or _72065_ (_21498_, _21464_, _07208_);
  and _72066_ (_21499_, _09450_, _07963_);
  or _72067_ (_21500_, _21499_, _21498_);
  and _72068_ (_21501_, _21500_, _05982_);
  and _72069_ (_21502_, _21501_, _21497_);
  and _72070_ (_21503_, _14859_, _07963_);
  or _72071_ (_21505_, _21503_, _21464_);
  and _72072_ (_21506_, _21505_, _10094_);
  or _72073_ (_21507_, _21506_, _06218_);
  or _72074_ (_21508_, _21507_, _21502_);
  and _72075_ (_21509_, _07963_, _08973_);
  or _72076_ (_21510_, _21509_, _21464_);
  or _72077_ (_21511_, _21510_, _06219_);
  and _72078_ (_21512_, _21511_, _21508_);
  or _72079_ (_21513_, _21512_, _06369_);
  and _72080_ (_21514_, _14751_, _07963_);
  or _72081_ (_21516_, _21514_, _21464_);
  or _72082_ (_21517_, _21516_, _07237_);
  and _72083_ (_21518_, _21517_, _07240_);
  and _72084_ (_21519_, _21518_, _21513_);
  and _72085_ (_21520_, _11259_, _07963_);
  or _72086_ (_21521_, _21520_, _21464_);
  and _72087_ (_21522_, _21521_, _06536_);
  or _72088_ (_21523_, _21522_, _21519_);
  and _72089_ (_21524_, _21523_, _07242_);
  or _72090_ (_21525_, _21464_, _08440_);
  and _72091_ (_21527_, _21510_, _06375_);
  and _72092_ (_21528_, _21527_, _21525_);
  or _72093_ (_21529_, _21528_, _21524_);
  and _72094_ (_21530_, _21529_, _07234_);
  and _72095_ (_21531_, _21476_, _06545_);
  and _72096_ (_21532_, _21531_, _21525_);
  or _72097_ (_21533_, _21532_, _06366_);
  or _72098_ (_21534_, _21533_, _21530_);
  and _72099_ (_21535_, _14748_, _08186_);
  or _72100_ (_21536_, _21464_, _09056_);
  or _72101_ (_21538_, _21536_, _21535_);
  and _72102_ (_21539_, _21538_, _09061_);
  and _72103_ (_21540_, _21539_, _21534_);
  nor _72104_ (_21541_, _11258_, _11633_);
  or _72105_ (_21542_, _21541_, _21464_);
  and _72106_ (_21543_, _21542_, _06528_);
  or _72107_ (_21544_, _21543_, _21540_);
  and _72108_ (_21545_, _21544_, _06926_);
  and _72109_ (_21546_, _21473_, _06568_);
  or _72110_ (_21547_, _21546_, _06278_);
  or _72111_ (_21549_, _21547_, _21545_);
  and _72112_ (_21550_, _14926_, _08186_);
  or _72113_ (_21551_, _21464_, _06279_);
  or _72114_ (_21552_, _21551_, _21550_);
  and _72115_ (_21553_, _21552_, _01347_);
  and _72116_ (_21554_, _21553_, _21549_);
  or _72117_ (_21555_, _21554_, _21463_);
  and _72118_ (_43197_, _21555_, _42618_);
  and _72119_ (_21556_, _01351_, \oc8051_golden_model_1.DPH [3]);
  and _72120_ (_21557_, _11633_, \oc8051_golden_model_1.DPH [3]);
  nor _72121_ (_21559_, _11633_, _07594_);
  or _72122_ (_21560_, _21559_, _21557_);
  or _72123_ (_21561_, _21560_, _07215_);
  or _72124_ (_21562_, _11662_, \oc8051_golden_model_1.DPH [3]);
  nor _72125_ (_21563_, _11663_, _11562_);
  and _72126_ (_21564_, _21563_, _21562_);
  and _72127_ (_21565_, _14953_, _08186_);
  or _72128_ (_21566_, _21565_, _21557_);
  or _72129_ (_21567_, _21566_, _07151_);
  and _72130_ (_21568_, _07963_, \oc8051_golden_model_1.ACC [3]);
  or _72131_ (_21570_, _21568_, _21557_);
  and _72132_ (_21571_, _21570_, _07141_);
  and _72133_ (_21572_, _07142_, \oc8051_golden_model_1.DPH [3]);
  or _72134_ (_21573_, _21572_, _06341_);
  or _72135_ (_21574_, _21573_, _21571_);
  and _72136_ (_21575_, _21574_, _07166_);
  and _72137_ (_21576_, _21575_, _21567_);
  and _72138_ (_21577_, _21560_, _06461_);
  or _72139_ (_21578_, _21577_, _06464_);
  or _72140_ (_21579_, _21578_, _21576_);
  or _72141_ (_21581_, _21570_, _06465_);
  and _72142_ (_21582_, _21581_, _11562_);
  and _72143_ (_21583_, _21582_, _21579_);
  or _72144_ (_21584_, _21583_, _21564_);
  and _72145_ (_21585_, _21584_, _06374_);
  nor _72146_ (_21586_, _06374_, _06213_);
  or _72147_ (_21587_, _21586_, _10080_);
  or _72148_ (_21588_, _21587_, _21585_);
  and _72149_ (_21589_, _21588_, _21561_);
  or _72150_ (_21590_, _21589_, _07460_);
  or _72151_ (_21592_, _21557_, _07208_);
  and _72152_ (_21593_, _09449_, _07963_);
  or _72153_ (_21594_, _21593_, _21592_);
  and _72154_ (_21595_, _21594_, _05982_);
  and _72155_ (_21596_, _21595_, _21590_);
  and _72156_ (_21597_, _15048_, _07963_);
  or _72157_ (_21598_, _21597_, _21557_);
  and _72158_ (_21599_, _21598_, _10094_);
  or _72159_ (_21600_, _21599_, _06218_);
  or _72160_ (_21601_, _21600_, _21596_);
  and _72161_ (_21603_, _07963_, _08930_);
  or _72162_ (_21604_, _21603_, _21557_);
  or _72163_ (_21605_, _21604_, _06219_);
  and _72164_ (_21606_, _21605_, _21601_);
  or _72165_ (_21607_, _21606_, _06369_);
  and _72166_ (_21608_, _14943_, _07963_);
  or _72167_ (_21609_, _21608_, _21557_);
  or _72168_ (_21610_, _21609_, _07237_);
  and _72169_ (_21611_, _21610_, _07240_);
  and _72170_ (_21612_, _21611_, _21607_);
  and _72171_ (_21614_, _12577_, _07963_);
  or _72172_ (_21615_, _21614_, _21557_);
  and _72173_ (_21616_, _21615_, _06536_);
  or _72174_ (_21617_, _21616_, _21612_);
  and _72175_ (_21618_, _21617_, _07242_);
  or _72176_ (_21619_, _21557_, _08292_);
  and _72177_ (_21620_, _21604_, _06375_);
  and _72178_ (_21621_, _21620_, _21619_);
  or _72179_ (_21622_, _21621_, _21618_);
  and _72180_ (_21623_, _21622_, _07234_);
  and _72181_ (_21625_, _21570_, _06545_);
  and _72182_ (_21626_, _21625_, _21619_);
  or _72183_ (_21627_, _21626_, _06366_);
  or _72184_ (_21628_, _21627_, _21623_);
  and _72185_ (_21629_, _14940_, _08186_);
  or _72186_ (_21630_, _21557_, _09056_);
  or _72187_ (_21631_, _21630_, _21629_);
  and _72188_ (_21632_, _21631_, _09061_);
  and _72189_ (_21633_, _21632_, _21628_);
  nor _72190_ (_21634_, _11256_, _11633_);
  or _72191_ (_21636_, _21634_, _21557_);
  and _72192_ (_21637_, _21636_, _06528_);
  or _72193_ (_21638_, _21637_, _21633_);
  and _72194_ (_21639_, _21638_, _06926_);
  and _72195_ (_21640_, _21566_, _06568_);
  or _72196_ (_21641_, _21640_, _06278_);
  or _72197_ (_21642_, _21641_, _21639_);
  and _72198_ (_21643_, _15128_, _08186_);
  or _72199_ (_21644_, _21557_, _06279_);
  or _72200_ (_21645_, _21644_, _21643_);
  and _72201_ (_21647_, _21645_, _01347_);
  and _72202_ (_21648_, _21647_, _21642_);
  or _72203_ (_21649_, _21648_, _21556_);
  and _72204_ (_43198_, _21649_, _42618_);
  not _72205_ (_21650_, \oc8051_golden_model_1.DPH [4]);
  nor _72206_ (_21651_, _01347_, _21650_);
  nor _72207_ (_21652_, _07963_, _21650_);
  nor _72208_ (_21653_, _08541_, _11633_);
  or _72209_ (_21654_, _21653_, _21652_);
  or _72210_ (_21655_, _21654_, _07215_);
  and _72211_ (_21656_, _15162_, _08186_);
  or _72212_ (_21657_, _21656_, _21652_);
  or _72213_ (_21658_, _21657_, _07151_);
  and _72214_ (_21659_, _07963_, \oc8051_golden_model_1.ACC [4]);
  or _72215_ (_21660_, _21659_, _21652_);
  and _72216_ (_21661_, _21660_, _07141_);
  nor _72217_ (_21662_, _07141_, _21650_);
  or _72218_ (_21663_, _21662_, _06341_);
  or _72219_ (_21664_, _21663_, _21661_);
  and _72220_ (_21665_, _21664_, _07166_);
  and _72221_ (_21668_, _21665_, _21658_);
  and _72222_ (_21669_, _21654_, _06461_);
  or _72223_ (_21670_, _21669_, _06464_);
  or _72224_ (_21671_, _21670_, _21668_);
  or _72225_ (_21672_, _21660_, _06465_);
  and _72226_ (_21673_, _21672_, _11562_);
  and _72227_ (_21674_, _21673_, _21671_);
  or _72228_ (_21675_, _11663_, \oc8051_golden_model_1.DPH [4]);
  nor _72229_ (_21676_, _11664_, _11562_);
  and _72230_ (_21677_, _21676_, _21675_);
  or _72231_ (_21679_, _21677_, _21674_);
  and _72232_ (_21680_, _21679_, _06374_);
  nor _72233_ (_21681_, _06968_, _06374_);
  or _72234_ (_21682_, _21681_, _10080_);
  or _72235_ (_21683_, _21682_, _21680_);
  and _72236_ (_21684_, _21683_, _21655_);
  or _72237_ (_21685_, _21684_, _07460_);
  or _72238_ (_21686_, _21652_, _07208_);
  and _72239_ (_21687_, _09448_, _07963_);
  or _72240_ (_21688_, _21687_, _21686_);
  and _72241_ (_21690_, _21688_, _05982_);
  and _72242_ (_21691_, _21690_, _21685_);
  and _72243_ (_21692_, _15254_, _07963_);
  or _72244_ (_21693_, _21692_, _21652_);
  and _72245_ (_21694_, _21693_, _10094_);
  or _72246_ (_21695_, _21694_, _06218_);
  or _72247_ (_21696_, _21695_, _21691_);
  and _72248_ (_21697_, _08959_, _07963_);
  or _72249_ (_21698_, _21697_, _21652_);
  or _72250_ (_21699_, _21698_, _06219_);
  and _72251_ (_21701_, _21699_, _21696_);
  or _72252_ (_21702_, _21701_, _06369_);
  and _72253_ (_21703_, _15269_, _07963_);
  or _72254_ (_21704_, _21703_, _21652_);
  or _72255_ (_21705_, _21704_, _07237_);
  and _72256_ (_21706_, _21705_, _07240_);
  and _72257_ (_21707_, _21706_, _21702_);
  and _72258_ (_21708_, _11254_, _07963_);
  or _72259_ (_21709_, _21708_, _21652_);
  and _72260_ (_21710_, _21709_, _06536_);
  or _72261_ (_21712_, _21710_, _21707_);
  and _72262_ (_21713_, _21712_, _07242_);
  or _72263_ (_21714_, _21652_, _08544_);
  and _72264_ (_21715_, _21698_, _06375_);
  and _72265_ (_21716_, _21715_, _21714_);
  or _72266_ (_21717_, _21716_, _21713_);
  and _72267_ (_21718_, _21717_, _07234_);
  and _72268_ (_21719_, _21660_, _06545_);
  and _72269_ (_21720_, _21719_, _21714_);
  or _72270_ (_21721_, _21720_, _06366_);
  or _72271_ (_21723_, _21721_, _21718_);
  and _72272_ (_21724_, _15266_, _08186_);
  or _72273_ (_21725_, _21652_, _09056_);
  or _72274_ (_21726_, _21725_, _21724_);
  and _72275_ (_21727_, _21726_, _09061_);
  and _72276_ (_21728_, _21727_, _21723_);
  nor _72277_ (_21729_, _11253_, _11633_);
  or _72278_ (_21730_, _21729_, _21652_);
  and _72279_ (_21731_, _21730_, _06528_);
  or _72280_ (_21732_, _21731_, _21728_);
  and _72281_ (_21734_, _21732_, _06926_);
  and _72282_ (_21735_, _21657_, _06568_);
  or _72283_ (_21736_, _21735_, _06278_);
  or _72284_ (_21737_, _21736_, _21734_);
  and _72285_ (_21738_, _15329_, _08186_);
  or _72286_ (_21739_, _21652_, _06279_);
  or _72287_ (_21740_, _21739_, _21738_);
  and _72288_ (_21741_, _21740_, _01347_);
  and _72289_ (_21742_, _21741_, _21737_);
  or _72290_ (_21743_, _21742_, _21651_);
  and _72291_ (_43199_, _21743_, _42618_);
  and _72292_ (_21745_, _01351_, \oc8051_golden_model_1.DPH [5]);
  and _72293_ (_21746_, _11633_, \oc8051_golden_model_1.DPH [5]);
  nor _72294_ (_21747_, _08244_, _11633_);
  or _72295_ (_21748_, _21747_, _21746_);
  or _72296_ (_21749_, _21748_, _07215_);
  and _72297_ (_21750_, _15358_, _08186_);
  or _72298_ (_21751_, _21750_, _21746_);
  or _72299_ (_21752_, _21751_, _07151_);
  and _72300_ (_21753_, _07963_, \oc8051_golden_model_1.ACC [5]);
  or _72301_ (_21755_, _21753_, _21746_);
  and _72302_ (_21756_, _21755_, _07141_);
  and _72303_ (_21757_, _07142_, \oc8051_golden_model_1.DPH [5]);
  or _72304_ (_21758_, _21757_, _06341_);
  or _72305_ (_21759_, _21758_, _21756_);
  and _72306_ (_21760_, _21759_, _07166_);
  and _72307_ (_21761_, _21760_, _21752_);
  and _72308_ (_21762_, _21748_, _06461_);
  or _72309_ (_21763_, _21762_, _06464_);
  or _72310_ (_21764_, _21763_, _21761_);
  or _72311_ (_21765_, _21755_, _06465_);
  and _72312_ (_21766_, _21765_, _11562_);
  and _72313_ (_21767_, _21766_, _21764_);
  or _72314_ (_21768_, _11664_, \oc8051_golden_model_1.DPH [5]);
  nor _72315_ (_21769_, _11665_, _11562_);
  and _72316_ (_21770_, _21769_, _21768_);
  or _72317_ (_21771_, _21770_, _21767_);
  and _72318_ (_21772_, _21771_, _06374_);
  nor _72319_ (_21773_, _06611_, _06374_);
  or _72320_ (_21774_, _21773_, _10080_);
  or _72321_ (_21777_, _21774_, _21772_);
  and _72322_ (_21778_, _21777_, _21749_);
  or _72323_ (_21779_, _21778_, _07460_);
  or _72324_ (_21780_, _21746_, _07208_);
  and _72325_ (_21781_, _09447_, _07963_);
  or _72326_ (_21782_, _21781_, _21780_);
  and _72327_ (_21783_, _21782_, _05982_);
  and _72328_ (_21784_, _21783_, _21779_);
  and _72329_ (_21785_, _15459_, _07963_);
  or _72330_ (_21786_, _21785_, _21746_);
  and _72331_ (_21788_, _21786_, _10094_);
  or _72332_ (_21789_, _21788_, _06218_);
  or _72333_ (_21790_, _21789_, _21784_);
  and _72334_ (_21791_, _08946_, _07963_);
  or _72335_ (_21792_, _21791_, _21746_);
  or _72336_ (_21793_, _21792_, _06219_);
  and _72337_ (_21794_, _21793_, _21790_);
  or _72338_ (_21795_, _21794_, _06369_);
  and _72339_ (_21796_, _15353_, _07963_);
  or _72340_ (_21797_, _21796_, _21746_);
  or _72341_ (_21799_, _21797_, _07237_);
  and _72342_ (_21800_, _21799_, _07240_);
  and _72343_ (_21801_, _21800_, _21795_);
  and _72344_ (_21802_, _11250_, _07963_);
  or _72345_ (_21803_, _21802_, _21746_);
  and _72346_ (_21804_, _21803_, _06536_);
  or _72347_ (_21805_, _21804_, _21801_);
  and _72348_ (_21806_, _21805_, _07242_);
  or _72349_ (_21807_, _21746_, _08247_);
  and _72350_ (_21808_, _21792_, _06375_);
  and _72351_ (_21810_, _21808_, _21807_);
  or _72352_ (_21811_, _21810_, _21806_);
  and _72353_ (_21812_, _21811_, _07234_);
  and _72354_ (_21813_, _21755_, _06545_);
  and _72355_ (_21814_, _21813_, _21807_);
  or _72356_ (_21815_, _21814_, _06366_);
  or _72357_ (_21816_, _21815_, _21812_);
  and _72358_ (_21817_, _15350_, _08186_);
  or _72359_ (_21818_, _21746_, _09056_);
  or _72360_ (_21819_, _21818_, _21817_);
  and _72361_ (_21821_, _21819_, _09061_);
  and _72362_ (_21822_, _21821_, _21816_);
  nor _72363_ (_21823_, _11249_, _11633_);
  or _72364_ (_21824_, _21823_, _21746_);
  and _72365_ (_21825_, _21824_, _06528_);
  or _72366_ (_21826_, _21825_, _21822_);
  and _72367_ (_21827_, _21826_, _06926_);
  and _72368_ (_21828_, _21751_, _06568_);
  or _72369_ (_21829_, _21828_, _06278_);
  or _72370_ (_21830_, _21829_, _21827_);
  and _72371_ (_21832_, _15532_, _08186_);
  or _72372_ (_21833_, _21746_, _06279_);
  or _72373_ (_21834_, _21833_, _21832_);
  and _72374_ (_21835_, _21834_, _01347_);
  and _72375_ (_21836_, _21835_, _21830_);
  or _72376_ (_21837_, _21836_, _21745_);
  and _72377_ (_43200_, _21837_, _42618_);
  not _72378_ (_21838_, \oc8051_golden_model_1.DPH [6]);
  nor _72379_ (_21839_, _01347_, _21838_);
  nor _72380_ (_21840_, _07963_, _21838_);
  nor _72381_ (_21842_, _08142_, _11633_);
  or _72382_ (_21843_, _21842_, _21840_);
  or _72383_ (_21844_, _21843_, _07215_);
  and _72384_ (_21845_, _15554_, _08186_);
  or _72385_ (_21846_, _21845_, _21840_);
  or _72386_ (_21847_, _21846_, _07151_);
  and _72387_ (_21848_, _07963_, \oc8051_golden_model_1.ACC [6]);
  or _72388_ (_21849_, _21848_, _21840_);
  and _72389_ (_21850_, _21849_, _07141_);
  nor _72390_ (_21851_, _07141_, _21838_);
  or _72391_ (_21853_, _21851_, _06341_);
  or _72392_ (_21854_, _21853_, _21850_);
  and _72393_ (_21855_, _21854_, _07166_);
  and _72394_ (_21856_, _21855_, _21847_);
  and _72395_ (_21857_, _21843_, _06461_);
  or _72396_ (_21858_, _21857_, _06464_);
  or _72397_ (_21859_, _21858_, _21856_);
  or _72398_ (_21860_, _21849_, _06465_);
  and _72399_ (_21861_, _21860_, _11562_);
  and _72400_ (_21862_, _21861_, _21859_);
  or _72401_ (_21864_, _11665_, \oc8051_golden_model_1.DPH [6]);
  nor _72402_ (_21865_, _11666_, _11562_);
  and _72403_ (_21866_, _21865_, _21864_);
  or _72404_ (_21867_, _21866_, _21862_);
  and _72405_ (_21868_, _21867_, _06374_);
  nor _72406_ (_21869_, _06374_, _06317_);
  or _72407_ (_21870_, _21869_, _10080_);
  or _72408_ (_21871_, _21870_, _21868_);
  and _72409_ (_21872_, _21871_, _21844_);
  or _72410_ (_21873_, _21872_, _07460_);
  or _72411_ (_21875_, _21840_, _07208_);
  and _72412_ (_21876_, _09446_, _07963_);
  or _72413_ (_21877_, _21876_, _21875_);
  and _72414_ (_21878_, _21877_, _05982_);
  and _72415_ (_21879_, _21878_, _21873_);
  and _72416_ (_21880_, _15657_, _07963_);
  or _72417_ (_21881_, _21880_, _21840_);
  and _72418_ (_21882_, _21881_, _10094_);
  or _72419_ (_21883_, _21882_, _06218_);
  or _72420_ (_21884_, _21883_, _21879_);
  and _72421_ (_21886_, _15664_, _07963_);
  or _72422_ (_21887_, _21886_, _21840_);
  or _72423_ (_21888_, _21887_, _06219_);
  and _72424_ (_21889_, _21888_, _21884_);
  or _72425_ (_21890_, _21889_, _06369_);
  and _72426_ (_21891_, _15549_, _07963_);
  or _72427_ (_21892_, _21891_, _21840_);
  or _72428_ (_21893_, _21892_, _07237_);
  and _72429_ (_21894_, _21893_, _07240_);
  and _72430_ (_21895_, _21894_, _21890_);
  and _72431_ (_21897_, _11247_, _07963_);
  or _72432_ (_21898_, _21897_, _21840_);
  and _72433_ (_21899_, _21898_, _06536_);
  or _72434_ (_21900_, _21899_, _21895_);
  and _72435_ (_21901_, _21900_, _07242_);
  or _72436_ (_21902_, _21840_, _08145_);
  and _72437_ (_21903_, _21887_, _06375_);
  and _72438_ (_21904_, _21903_, _21902_);
  or _72439_ (_21905_, _21904_, _21901_);
  and _72440_ (_21906_, _21905_, _07234_);
  and _72441_ (_21908_, _21849_, _06545_);
  and _72442_ (_21909_, _21908_, _21902_);
  or _72443_ (_21910_, _21909_, _06366_);
  or _72444_ (_21911_, _21910_, _21906_);
  and _72445_ (_21912_, _15546_, _08186_);
  or _72446_ (_21913_, _21840_, _09056_);
  or _72447_ (_21914_, _21913_, _21912_);
  and _72448_ (_21915_, _21914_, _09061_);
  and _72449_ (_21916_, _21915_, _21911_);
  nor _72450_ (_21917_, _11246_, _11633_);
  or _72451_ (_21919_, _21917_, _21840_);
  and _72452_ (_21920_, _21919_, _06528_);
  or _72453_ (_21921_, _21920_, _21916_);
  and _72454_ (_21922_, _21921_, _06926_);
  and _72455_ (_21923_, _21846_, _06568_);
  or _72456_ (_21924_, _21923_, _06278_);
  or _72457_ (_21925_, _21924_, _21922_);
  and _72458_ (_21926_, _15734_, _08186_);
  or _72459_ (_21927_, _21840_, _06279_);
  or _72460_ (_21928_, _21927_, _21926_);
  and _72461_ (_21930_, _21928_, _01347_);
  and _72462_ (_21931_, _21930_, _21925_);
  or _72463_ (_21932_, _21931_, _21839_);
  and _72464_ (_43201_, _21932_, _42618_);
  not _72465_ (_21933_, \oc8051_golden_model_1.TL1 [0]);
  nor _72466_ (_21934_, _01347_, _21933_);
  nand _72467_ (_21935_, _11263_, _07968_);
  nor _72468_ (_21936_, _07968_, _21933_);
  nor _72469_ (_21937_, _21936_, _07234_);
  nand _72470_ (_21938_, _21937_, _21935_);
  and _72471_ (_21940_, _07968_, _07133_);
  or _72472_ (_21941_, _21940_, _21936_);
  or _72473_ (_21942_, _21941_, _07215_);
  nor _72474_ (_21943_, _08390_, _11726_);
  or _72475_ (_21944_, _21943_, _21936_);
  or _72476_ (_21945_, _21944_, _07151_);
  and _72477_ (_21946_, _07968_, \oc8051_golden_model_1.ACC [0]);
  or _72478_ (_21947_, _21946_, _21936_);
  and _72479_ (_21948_, _21947_, _07141_);
  nor _72480_ (_21949_, _07141_, _21933_);
  or _72481_ (_21951_, _21949_, _06341_);
  or _72482_ (_21952_, _21951_, _21948_);
  and _72483_ (_21953_, _21952_, _07166_);
  and _72484_ (_21954_, _21953_, _21945_);
  and _72485_ (_21955_, _21941_, _06461_);
  or _72486_ (_21956_, _21955_, _21954_);
  and _72487_ (_21957_, _21956_, _06465_);
  and _72488_ (_21958_, _21947_, _06464_);
  or _72489_ (_21959_, _21958_, _10080_);
  or _72490_ (_21960_, _21959_, _21957_);
  and _72491_ (_21962_, _21960_, _21942_);
  or _72492_ (_21963_, _21962_, _07460_);
  and _72493_ (_21964_, _09392_, _07968_);
  or _72494_ (_21965_, _21936_, _07208_);
  or _72495_ (_21966_, _21965_, _21964_);
  and _72496_ (_21967_, _21966_, _21963_);
  or _72497_ (_21968_, _21967_, _10094_);
  and _72498_ (_21969_, _14467_, _07968_);
  or _72499_ (_21970_, _21936_, _05982_);
  or _72500_ (_21971_, _21970_, _21969_);
  and _72501_ (_21973_, _21971_, _06219_);
  and _72502_ (_21974_, _21973_, _21968_);
  and _72503_ (_21975_, _07968_, _08954_);
  or _72504_ (_21976_, _21975_, _21936_);
  and _72505_ (_21977_, _21976_, _06218_);
  or _72506_ (_21978_, _21977_, _06369_);
  or _72507_ (_21979_, _21978_, _21974_);
  and _72508_ (_21980_, _14366_, _07968_);
  or _72509_ (_21981_, _21980_, _21936_);
  or _72510_ (_21982_, _21981_, _07237_);
  and _72511_ (_21984_, _21982_, _07240_);
  and _72512_ (_21985_, _21984_, _21979_);
  nor _72513_ (_21986_, _12580_, _11726_);
  or _72514_ (_21987_, _21986_, _21936_);
  and _72515_ (_21988_, _21935_, _06536_);
  and _72516_ (_21989_, _21988_, _21987_);
  or _72517_ (_21990_, _21989_, _21985_);
  and _72518_ (_21991_, _21990_, _07242_);
  nand _72519_ (_21992_, _21976_, _06375_);
  nor _72520_ (_21993_, _21992_, _21943_);
  or _72521_ (_21995_, _21993_, _06545_);
  or _72522_ (_21996_, _21995_, _21991_);
  and _72523_ (_21997_, _21996_, _21938_);
  or _72524_ (_21998_, _21997_, _06366_);
  and _72525_ (_21999_, _14363_, _07968_);
  or _72526_ (_22000_, _21936_, _09056_);
  or _72527_ (_22001_, _22000_, _21999_);
  and _72528_ (_22002_, _22001_, _09061_);
  and _72529_ (_22003_, _22002_, _21998_);
  and _72530_ (_22004_, _21987_, _06528_);
  or _72531_ (_22006_, _22004_, _19502_);
  or _72532_ (_22007_, _22006_, _22003_);
  or _72533_ (_22008_, _21944_, _06661_);
  and _72534_ (_22009_, _22008_, _01347_);
  and _72535_ (_22010_, _22009_, _22007_);
  or _72536_ (_22011_, _22010_, _21934_);
  and _72537_ (_43202_, _22011_, _42618_);
  not _72538_ (_22012_, \oc8051_golden_model_1.TL1 [1]);
  nor _72539_ (_22013_, _01347_, _22012_);
  or _72540_ (_22014_, _07968_, \oc8051_golden_model_1.TL1 [1]);
  and _72541_ (_22016_, _14562_, _07968_);
  not _72542_ (_22017_, _22016_);
  and _72543_ (_22018_, _22017_, _22014_);
  or _72544_ (_22019_, _22018_, _07151_);
  nor _72545_ (_22020_, _07968_, _22012_);
  and _72546_ (_22021_, _07968_, \oc8051_golden_model_1.ACC [1]);
  or _72547_ (_22022_, _22021_, _22020_);
  and _72548_ (_22023_, _22022_, _07141_);
  nor _72549_ (_22024_, _07141_, _22012_);
  or _72550_ (_22025_, _22024_, _06341_);
  or _72551_ (_22027_, _22025_, _22023_);
  and _72552_ (_22028_, _22027_, _07166_);
  and _72553_ (_22029_, _22028_, _22019_);
  nor _72554_ (_22030_, _11726_, _07357_);
  or _72555_ (_22031_, _22030_, _22020_);
  and _72556_ (_22032_, _22031_, _06461_);
  or _72557_ (_22033_, _22032_, _22029_);
  and _72558_ (_22034_, _22033_, _06465_);
  and _72559_ (_22035_, _22022_, _06464_);
  or _72560_ (_22036_, _22035_, _10080_);
  or _72561_ (_22038_, _22036_, _22034_);
  or _72562_ (_22039_, _22031_, _07215_);
  and _72563_ (_22040_, _22039_, _22038_);
  or _72564_ (_22041_, _22040_, _07460_);
  and _72565_ (_22042_, _09451_, _07968_);
  or _72566_ (_22043_, _22020_, _07208_);
  or _72567_ (_22044_, _22043_, _22042_);
  and _72568_ (_22045_, _22044_, _05982_);
  and _72569_ (_22046_, _22045_, _22041_);
  or _72570_ (_22047_, _14653_, _11726_);
  and _72571_ (_22049_, _22014_, _10094_);
  and _72572_ (_22050_, _22049_, _22047_);
  or _72573_ (_22051_, _22050_, _22046_);
  and _72574_ (_22052_, _22051_, _06219_);
  nand _72575_ (_22053_, _07968_, _07038_);
  and _72576_ (_22054_, _22014_, _06218_);
  and _72577_ (_22055_, _22054_, _22053_);
  or _72578_ (_22056_, _22055_, _22052_);
  and _72579_ (_22057_, _22056_, _07237_);
  or _72580_ (_22058_, _14668_, _11726_);
  and _72581_ (_22060_, _22014_, _06369_);
  and _72582_ (_22061_, _22060_, _22058_);
  or _72583_ (_22062_, _22061_, _06536_);
  or _72584_ (_22063_, _22062_, _22057_);
  nor _72585_ (_22064_, _11261_, _11726_);
  or _72586_ (_22065_, _22064_, _22020_);
  nand _72587_ (_22066_, _11260_, _07968_);
  and _72588_ (_22067_, _22066_, _22065_);
  or _72589_ (_22068_, _22067_, _07240_);
  and _72590_ (_22069_, _22068_, _07242_);
  and _72591_ (_22071_, _22069_, _22063_);
  or _72592_ (_22072_, _14666_, _11726_);
  and _72593_ (_22073_, _22014_, _06375_);
  and _72594_ (_22074_, _22073_, _22072_);
  or _72595_ (_22075_, _22074_, _06545_);
  or _72596_ (_22076_, _22075_, _22071_);
  nor _72597_ (_22077_, _22020_, _07234_);
  nand _72598_ (_22078_, _22077_, _22066_);
  and _72599_ (_22079_, _22078_, _09056_);
  and _72600_ (_22080_, _22079_, _22076_);
  or _72601_ (_22082_, _22053_, _08341_);
  and _72602_ (_22083_, _22014_, _06366_);
  and _72603_ (_22084_, _22083_, _22082_);
  or _72604_ (_22085_, _22084_, _06528_);
  or _72605_ (_22086_, _22085_, _22080_);
  or _72606_ (_22087_, _22065_, _09061_);
  and _72607_ (_22088_, _22087_, _06926_);
  and _72608_ (_22089_, _22088_, _22086_);
  and _72609_ (_22090_, _22018_, _06568_);
  or _72610_ (_22091_, _22090_, _06278_);
  or _72611_ (_22093_, _22091_, _22089_);
  or _72612_ (_22094_, _22020_, _06279_);
  or _72613_ (_22095_, _22094_, _22016_);
  and _72614_ (_22096_, _22095_, _01347_);
  and _72615_ (_22097_, _22096_, _22093_);
  or _72616_ (_22098_, _22097_, _22013_);
  and _72617_ (_43204_, _22098_, _42618_);
  and _72618_ (_22099_, _01351_, \oc8051_golden_model_1.TL1 [2]);
  and _72619_ (_22100_, _11726_, \oc8051_golden_model_1.TL1 [2]);
  nor _72620_ (_22101_, _11726_, _07776_);
  or _72621_ (_22103_, _22101_, _22100_);
  or _72622_ (_22104_, _22103_, _07215_);
  and _72623_ (_22105_, _14770_, _07968_);
  or _72624_ (_22106_, _22105_, _22100_);
  and _72625_ (_22107_, _22106_, _06341_);
  and _72626_ (_22108_, _07142_, \oc8051_golden_model_1.TL1 [2]);
  and _72627_ (_22109_, _07968_, \oc8051_golden_model_1.ACC [2]);
  or _72628_ (_22110_, _22109_, _22100_);
  and _72629_ (_22111_, _22110_, _07141_);
  or _72630_ (_22112_, _22111_, _22108_);
  and _72631_ (_22114_, _22112_, _07151_);
  or _72632_ (_22115_, _22114_, _06461_);
  or _72633_ (_22116_, _22115_, _22107_);
  or _72634_ (_22117_, _22103_, _07166_);
  and _72635_ (_22118_, _22117_, _06465_);
  and _72636_ (_22119_, _22118_, _22116_);
  and _72637_ (_22120_, _22110_, _06464_);
  or _72638_ (_22121_, _22120_, _10080_);
  or _72639_ (_22122_, _22121_, _22119_);
  and _72640_ (_22123_, _22122_, _22104_);
  or _72641_ (_22126_, _22123_, _07460_);
  and _72642_ (_22127_, _09450_, _07968_);
  or _72643_ (_22128_, _22100_, _07208_);
  or _72644_ (_22129_, _22128_, _22127_);
  and _72645_ (_22130_, _22129_, _22126_);
  or _72646_ (_22131_, _22130_, _10094_);
  and _72647_ (_22132_, _14859_, _07968_);
  or _72648_ (_22133_, _22100_, _05982_);
  or _72649_ (_22134_, _22133_, _22132_);
  and _72650_ (_22135_, _22134_, _06219_);
  and _72651_ (_22137_, _22135_, _22131_);
  and _72652_ (_22138_, _07968_, _08973_);
  or _72653_ (_22139_, _22138_, _22100_);
  and _72654_ (_22140_, _22139_, _06218_);
  or _72655_ (_22141_, _22140_, _06369_);
  or _72656_ (_22142_, _22141_, _22137_);
  and _72657_ (_22143_, _14751_, _07968_);
  or _72658_ (_22144_, _22143_, _22100_);
  or _72659_ (_22145_, _22144_, _07237_);
  and _72660_ (_22146_, _22145_, _07240_);
  and _72661_ (_22148_, _22146_, _22142_);
  and _72662_ (_22149_, _11259_, _07968_);
  or _72663_ (_22150_, _22149_, _22100_);
  and _72664_ (_22151_, _22150_, _06536_);
  or _72665_ (_22152_, _22151_, _22148_);
  and _72666_ (_22153_, _22152_, _07242_);
  or _72667_ (_22154_, _22100_, _08440_);
  and _72668_ (_22155_, _22139_, _06375_);
  and _72669_ (_22156_, _22155_, _22154_);
  or _72670_ (_22157_, _22156_, _22153_);
  and _72671_ (_22159_, _22157_, _07234_);
  and _72672_ (_22160_, _22110_, _06545_);
  and _72673_ (_22161_, _22160_, _22154_);
  or _72674_ (_22162_, _22161_, _06366_);
  or _72675_ (_22163_, _22162_, _22159_);
  and _72676_ (_22164_, _14748_, _07968_);
  or _72677_ (_22165_, _22100_, _09056_);
  or _72678_ (_22166_, _22165_, _22164_);
  and _72679_ (_22167_, _22166_, _09061_);
  and _72680_ (_22168_, _22167_, _22163_);
  nor _72681_ (_22170_, _11258_, _11726_);
  or _72682_ (_22171_, _22170_, _22100_);
  and _72683_ (_22172_, _22171_, _06528_);
  or _72684_ (_22173_, _22172_, _22168_);
  and _72685_ (_22174_, _22173_, _06926_);
  and _72686_ (_22175_, _22106_, _06568_);
  or _72687_ (_22176_, _22175_, _06278_);
  or _72688_ (_22177_, _22176_, _22174_);
  and _72689_ (_22178_, _14926_, _07968_);
  or _72690_ (_22179_, _22100_, _06279_);
  or _72691_ (_22181_, _22179_, _22178_);
  and _72692_ (_22182_, _22181_, _01347_);
  and _72693_ (_22183_, _22182_, _22177_);
  or _72694_ (_22184_, _22183_, _22099_);
  and _72695_ (_43205_, _22184_, _42618_);
  and _72696_ (_22185_, _01351_, \oc8051_golden_model_1.TL1 [3]);
  and _72697_ (_22186_, _11726_, \oc8051_golden_model_1.TL1 [3]);
  and _72698_ (_22187_, _14953_, _07968_);
  or _72699_ (_22188_, _22187_, _22186_);
  or _72700_ (_22189_, _22188_, _07151_);
  and _72701_ (_22191_, _07968_, \oc8051_golden_model_1.ACC [3]);
  or _72702_ (_22192_, _22191_, _22186_);
  and _72703_ (_22193_, _22192_, _07141_);
  and _72704_ (_22194_, _07142_, \oc8051_golden_model_1.TL1 [3]);
  or _72705_ (_22195_, _22194_, _06341_);
  or _72706_ (_22196_, _22195_, _22193_);
  and _72707_ (_22197_, _22196_, _07166_);
  and _72708_ (_22198_, _22197_, _22189_);
  nor _72709_ (_22199_, _11726_, _07594_);
  or _72710_ (_22200_, _22199_, _22186_);
  and _72711_ (_22202_, _22200_, _06461_);
  or _72712_ (_22203_, _22202_, _22198_);
  and _72713_ (_22204_, _22203_, _06465_);
  and _72714_ (_22205_, _22192_, _06464_);
  or _72715_ (_22206_, _22205_, _10080_);
  or _72716_ (_22207_, _22206_, _22204_);
  or _72717_ (_22208_, _22200_, _07215_);
  and _72718_ (_22209_, _22208_, _22207_);
  or _72719_ (_22210_, _22209_, _07460_);
  and _72720_ (_22211_, _09449_, _07968_);
  or _72721_ (_22212_, _22186_, _07208_);
  or _72722_ (_22213_, _22212_, _22211_);
  and _72723_ (_22214_, _22213_, _05982_);
  and _72724_ (_22215_, _22214_, _22210_);
  and _72725_ (_22216_, _15048_, _07968_);
  or _72726_ (_22217_, _22216_, _22186_);
  and _72727_ (_22218_, _22217_, _10094_);
  or _72728_ (_22219_, _22218_, _06218_);
  or _72729_ (_22220_, _22219_, _22215_);
  and _72730_ (_22221_, _07968_, _08930_);
  or _72731_ (_22224_, _22221_, _22186_);
  or _72732_ (_22225_, _22224_, _06219_);
  and _72733_ (_22226_, _22225_, _22220_);
  or _72734_ (_22227_, _22226_, _06369_);
  and _72735_ (_22228_, _14943_, _07968_);
  or _72736_ (_22229_, _22228_, _22186_);
  or _72737_ (_22230_, _22229_, _07237_);
  and _72738_ (_22231_, _22230_, _07240_);
  and _72739_ (_22232_, _22231_, _22227_);
  and _72740_ (_22233_, _12577_, _07968_);
  or _72741_ (_22235_, _22233_, _22186_);
  and _72742_ (_22236_, _22235_, _06536_);
  or _72743_ (_22237_, _22236_, _22232_);
  and _72744_ (_22238_, _22237_, _07242_);
  or _72745_ (_22239_, _22186_, _08292_);
  and _72746_ (_22240_, _22224_, _06375_);
  and _72747_ (_22241_, _22240_, _22239_);
  or _72748_ (_22242_, _22241_, _22238_);
  and _72749_ (_22243_, _22242_, _07234_);
  and _72750_ (_22244_, _22192_, _06545_);
  and _72751_ (_22246_, _22244_, _22239_);
  or _72752_ (_22247_, _22246_, _06366_);
  or _72753_ (_22248_, _22247_, _22243_);
  and _72754_ (_22249_, _14940_, _07968_);
  or _72755_ (_22250_, _22186_, _09056_);
  or _72756_ (_22251_, _22250_, _22249_);
  and _72757_ (_22252_, _22251_, _09061_);
  and _72758_ (_22253_, _22252_, _22248_);
  nor _72759_ (_22254_, _11256_, _11726_);
  or _72760_ (_22255_, _22254_, _22186_);
  and _72761_ (_22257_, _22255_, _06528_);
  or _72762_ (_22258_, _22257_, _22253_);
  and _72763_ (_22259_, _22258_, _06926_);
  and _72764_ (_22260_, _22188_, _06568_);
  or _72765_ (_22261_, _22260_, _06278_);
  or _72766_ (_22262_, _22261_, _22259_);
  and _72767_ (_22263_, _15128_, _07968_);
  or _72768_ (_22264_, _22186_, _06279_);
  or _72769_ (_22265_, _22264_, _22263_);
  and _72770_ (_22266_, _22265_, _01347_);
  and _72771_ (_22268_, _22266_, _22262_);
  or _72772_ (_22269_, _22268_, _22185_);
  and _72773_ (_43206_, _22269_, _42618_);
  and _72774_ (_22270_, _01351_, \oc8051_golden_model_1.TL1 [4]);
  and _72775_ (_22271_, _11726_, \oc8051_golden_model_1.TL1 [4]);
  and _72776_ (_22272_, _15162_, _07968_);
  or _72777_ (_22273_, _22272_, _22271_);
  or _72778_ (_22274_, _22273_, _07151_);
  and _72779_ (_22275_, _07968_, \oc8051_golden_model_1.ACC [4]);
  or _72780_ (_22276_, _22275_, _22271_);
  and _72781_ (_22278_, _22276_, _07141_);
  and _72782_ (_22279_, _07142_, \oc8051_golden_model_1.TL1 [4]);
  or _72783_ (_22280_, _22279_, _06341_);
  or _72784_ (_22281_, _22280_, _22278_);
  and _72785_ (_22282_, _22281_, _07166_);
  and _72786_ (_22283_, _22282_, _22274_);
  nor _72787_ (_22284_, _08541_, _11726_);
  or _72788_ (_22285_, _22284_, _22271_);
  and _72789_ (_22286_, _22285_, _06461_);
  or _72790_ (_22287_, _22286_, _22283_);
  and _72791_ (_22289_, _22287_, _06465_);
  and _72792_ (_22290_, _22276_, _06464_);
  or _72793_ (_22291_, _22290_, _10080_);
  or _72794_ (_22292_, _22291_, _22289_);
  or _72795_ (_22293_, _22285_, _07215_);
  and _72796_ (_22294_, _22293_, _22292_);
  or _72797_ (_22295_, _22294_, _07460_);
  and _72798_ (_22296_, _09448_, _07968_);
  or _72799_ (_22297_, _22271_, _07208_);
  or _72800_ (_22298_, _22297_, _22296_);
  and _72801_ (_22300_, _22298_, _22295_);
  or _72802_ (_22301_, _22300_, _10094_);
  and _72803_ (_22302_, _15254_, _07968_);
  or _72804_ (_22303_, _22271_, _05982_);
  or _72805_ (_22304_, _22303_, _22302_);
  and _72806_ (_22305_, _22304_, _06219_);
  and _72807_ (_22306_, _22305_, _22301_);
  and _72808_ (_22307_, _08959_, _07968_);
  or _72809_ (_22308_, _22307_, _22271_);
  and _72810_ (_22309_, _22308_, _06218_);
  or _72811_ (_22311_, _22309_, _06369_);
  or _72812_ (_22312_, _22311_, _22306_);
  and _72813_ (_22313_, _15269_, _07968_);
  or _72814_ (_22314_, _22313_, _22271_);
  or _72815_ (_22315_, _22314_, _07237_);
  and _72816_ (_22316_, _22315_, _07240_);
  and _72817_ (_22317_, _22316_, _22312_);
  and _72818_ (_22318_, _11254_, _07968_);
  or _72819_ (_22319_, _22318_, _22271_);
  and _72820_ (_22320_, _22319_, _06536_);
  or _72821_ (_22322_, _22320_, _22317_);
  and _72822_ (_22323_, _22322_, _07242_);
  or _72823_ (_22324_, _22271_, _08544_);
  and _72824_ (_22325_, _22308_, _06375_);
  and _72825_ (_22326_, _22325_, _22324_);
  or _72826_ (_22327_, _22326_, _22323_);
  and _72827_ (_22328_, _22327_, _07234_);
  and _72828_ (_22329_, _22276_, _06545_);
  and _72829_ (_22330_, _22329_, _22324_);
  or _72830_ (_22331_, _22330_, _06366_);
  or _72831_ (_22333_, _22331_, _22328_);
  and _72832_ (_22334_, _15266_, _07968_);
  or _72833_ (_22335_, _22271_, _09056_);
  or _72834_ (_22336_, _22335_, _22334_);
  and _72835_ (_22337_, _22336_, _09061_);
  and _72836_ (_22338_, _22337_, _22333_);
  nor _72837_ (_22339_, _11253_, _11726_);
  or _72838_ (_22340_, _22339_, _22271_);
  and _72839_ (_22341_, _22340_, _06528_);
  or _72840_ (_22342_, _22341_, _22338_);
  and _72841_ (_22344_, _22342_, _06926_);
  and _72842_ (_22345_, _22273_, _06568_);
  or _72843_ (_22346_, _22345_, _06278_);
  or _72844_ (_22347_, _22346_, _22344_);
  and _72845_ (_22348_, _15329_, _07968_);
  or _72846_ (_22349_, _22271_, _06279_);
  or _72847_ (_22350_, _22349_, _22348_);
  and _72848_ (_22351_, _22350_, _01347_);
  and _72849_ (_22352_, _22351_, _22347_);
  or _72850_ (_22353_, _22352_, _22270_);
  and _72851_ (_43207_, _22353_, _42618_);
  and _72852_ (_22355_, _01351_, \oc8051_golden_model_1.TL1 [5]);
  and _72853_ (_22356_, _11726_, \oc8051_golden_model_1.TL1 [5]);
  nor _72854_ (_22357_, _08244_, _11726_);
  or _72855_ (_22358_, _22357_, _22356_);
  or _72856_ (_22359_, _22358_, _07215_);
  and _72857_ (_22360_, _15358_, _07968_);
  or _72858_ (_22361_, _22360_, _22356_);
  or _72859_ (_22362_, _22361_, _07151_);
  and _72860_ (_22363_, _07968_, \oc8051_golden_model_1.ACC [5]);
  or _72861_ (_22365_, _22363_, _22356_);
  and _72862_ (_22366_, _22365_, _07141_);
  and _72863_ (_22367_, _07142_, \oc8051_golden_model_1.TL1 [5]);
  or _72864_ (_22368_, _22367_, _06341_);
  or _72865_ (_22369_, _22368_, _22366_);
  and _72866_ (_22370_, _22369_, _07166_);
  and _72867_ (_22371_, _22370_, _22362_);
  and _72868_ (_22372_, _22358_, _06461_);
  or _72869_ (_22373_, _22372_, _22371_);
  and _72870_ (_22374_, _22373_, _06465_);
  and _72871_ (_22376_, _22365_, _06464_);
  or _72872_ (_22377_, _22376_, _10080_);
  or _72873_ (_22378_, _22377_, _22374_);
  and _72874_ (_22379_, _22378_, _22359_);
  or _72875_ (_22380_, _22379_, _07460_);
  and _72876_ (_22381_, _09447_, _07968_);
  or _72877_ (_22382_, _22356_, _07208_);
  or _72878_ (_22383_, _22382_, _22381_);
  and _72879_ (_22384_, _22383_, _05982_);
  and _72880_ (_22385_, _22384_, _22380_);
  and _72881_ (_22387_, _15459_, _07968_);
  or _72882_ (_22388_, _22387_, _22356_);
  and _72883_ (_22389_, _22388_, _10094_);
  or _72884_ (_22390_, _22389_, _06218_);
  or _72885_ (_22391_, _22390_, _22385_);
  and _72886_ (_22392_, _08946_, _07968_);
  or _72887_ (_22393_, _22392_, _22356_);
  or _72888_ (_22394_, _22393_, _06219_);
  and _72889_ (_22395_, _22394_, _22391_);
  or _72890_ (_22396_, _22395_, _06369_);
  and _72891_ (_22398_, _15353_, _07968_);
  or _72892_ (_22399_, _22398_, _22356_);
  or _72893_ (_22400_, _22399_, _07237_);
  and _72894_ (_22401_, _22400_, _07240_);
  and _72895_ (_22402_, _22401_, _22396_);
  and _72896_ (_22403_, _11250_, _07968_);
  or _72897_ (_22404_, _22403_, _22356_);
  and _72898_ (_22405_, _22404_, _06536_);
  or _72899_ (_22406_, _22405_, _22402_);
  and _72900_ (_22407_, _22406_, _07242_);
  or _72901_ (_22409_, _22356_, _08247_);
  and _72902_ (_22410_, _22393_, _06375_);
  and _72903_ (_22411_, _22410_, _22409_);
  or _72904_ (_22412_, _22411_, _22407_);
  and _72905_ (_22413_, _22412_, _07234_);
  and _72906_ (_22414_, _22365_, _06545_);
  and _72907_ (_22415_, _22414_, _22409_);
  or _72908_ (_22416_, _22415_, _06366_);
  or _72909_ (_22417_, _22416_, _22413_);
  and _72910_ (_22418_, _15350_, _07968_);
  or _72911_ (_22420_, _22356_, _09056_);
  or _72912_ (_22421_, _22420_, _22418_);
  and _72913_ (_22422_, _22421_, _09061_);
  and _72914_ (_22423_, _22422_, _22417_);
  nor _72915_ (_22424_, _11249_, _11726_);
  or _72916_ (_22425_, _22424_, _22356_);
  and _72917_ (_22426_, _22425_, _06528_);
  or _72918_ (_22427_, _22426_, _22423_);
  and _72919_ (_22428_, _22427_, _06926_);
  and _72920_ (_22429_, _22361_, _06568_);
  or _72921_ (_22431_, _22429_, _06278_);
  or _72922_ (_22432_, _22431_, _22428_);
  and _72923_ (_22433_, _15532_, _07968_);
  or _72924_ (_22434_, _22356_, _06279_);
  or _72925_ (_22435_, _22434_, _22433_);
  and _72926_ (_22436_, _22435_, _01347_);
  and _72927_ (_22437_, _22436_, _22432_);
  or _72928_ (_22438_, _22437_, _22355_);
  and _72929_ (_43208_, _22438_, _42618_);
  and _72930_ (_22439_, _01351_, \oc8051_golden_model_1.TL1 [6]);
  and _72931_ (_22441_, _11726_, \oc8051_golden_model_1.TL1 [6]);
  and _72932_ (_22442_, _15554_, _07968_);
  or _72933_ (_22443_, _22442_, _22441_);
  or _72934_ (_22444_, _22443_, _07151_);
  and _72935_ (_22445_, _07968_, \oc8051_golden_model_1.ACC [6]);
  or _72936_ (_22446_, _22445_, _22441_);
  and _72937_ (_22447_, _22446_, _07141_);
  and _72938_ (_22448_, _07142_, \oc8051_golden_model_1.TL1 [6]);
  or _72939_ (_22449_, _22448_, _06341_);
  or _72940_ (_22450_, _22449_, _22447_);
  and _72941_ (_22452_, _22450_, _07166_);
  and _72942_ (_22453_, _22452_, _22444_);
  nor _72943_ (_22454_, _08142_, _11726_);
  or _72944_ (_22455_, _22454_, _22441_);
  and _72945_ (_22456_, _22455_, _06461_);
  or _72946_ (_22457_, _22456_, _22453_);
  and _72947_ (_22458_, _22457_, _06465_);
  and _72948_ (_22459_, _22446_, _06464_);
  or _72949_ (_22460_, _22459_, _10080_);
  or _72950_ (_22461_, _22460_, _22458_);
  or _72951_ (_22463_, _22455_, _07215_);
  and _72952_ (_22464_, _22463_, _22461_);
  or _72953_ (_22465_, _22464_, _07460_);
  and _72954_ (_22466_, _09446_, _07968_);
  or _72955_ (_22467_, _22441_, _07208_);
  or _72956_ (_22468_, _22467_, _22466_);
  and _72957_ (_22469_, _22468_, _05982_);
  and _72958_ (_22470_, _22469_, _22465_);
  and _72959_ (_22471_, _15657_, _07968_);
  or _72960_ (_22472_, _22471_, _22441_);
  and _72961_ (_22474_, _22472_, _10094_);
  or _72962_ (_22475_, _22474_, _06218_);
  or _72963_ (_22476_, _22475_, _22470_);
  and _72964_ (_22477_, _15664_, _07968_);
  or _72965_ (_22478_, _22477_, _22441_);
  or _72966_ (_22479_, _22478_, _06219_);
  and _72967_ (_22480_, _22479_, _22476_);
  or _72968_ (_22481_, _22480_, _06369_);
  and _72969_ (_22482_, _15549_, _07968_);
  or _72970_ (_22483_, _22482_, _22441_);
  or _72971_ (_22485_, _22483_, _07237_);
  and _72972_ (_22486_, _22485_, _07240_);
  and _72973_ (_22487_, _22486_, _22481_);
  and _72974_ (_22488_, _11247_, _07968_);
  or _72975_ (_22489_, _22488_, _22441_);
  and _72976_ (_22490_, _22489_, _06536_);
  or _72977_ (_22491_, _22490_, _22487_);
  and _72978_ (_22492_, _22491_, _07242_);
  or _72979_ (_22493_, _22441_, _08145_);
  and _72980_ (_22494_, _22478_, _06375_);
  and _72981_ (_22496_, _22494_, _22493_);
  or _72982_ (_22497_, _22496_, _22492_);
  and _72983_ (_22498_, _22497_, _07234_);
  and _72984_ (_22499_, _22446_, _06545_);
  and _72985_ (_22500_, _22499_, _22493_);
  or _72986_ (_22501_, _22500_, _06366_);
  or _72987_ (_22502_, _22501_, _22498_);
  and _72988_ (_22503_, _15546_, _07968_);
  or _72989_ (_22504_, _22441_, _09056_);
  or _72990_ (_22505_, _22504_, _22503_);
  and _72991_ (_22506_, _22505_, _09061_);
  and _72992_ (_22507_, _22506_, _22502_);
  nor _72993_ (_22508_, _11246_, _11726_);
  or _72994_ (_22509_, _22508_, _22441_);
  and _72995_ (_22510_, _22509_, _06528_);
  or _72996_ (_22511_, _22510_, _22507_);
  and _72997_ (_22512_, _22511_, _06926_);
  and _72998_ (_22513_, _22443_, _06568_);
  or _72999_ (_22514_, _22513_, _06278_);
  or _73000_ (_22515_, _22514_, _22512_);
  and _73001_ (_22518_, _15734_, _07968_);
  or _73002_ (_22519_, _22441_, _06279_);
  or _73003_ (_22520_, _22519_, _22518_);
  and _73004_ (_22521_, _22520_, _01347_);
  and _73005_ (_22522_, _22521_, _22515_);
  or _73006_ (_22523_, _22522_, _22439_);
  and _73007_ (_43209_, _22523_, _42618_);
  not _73008_ (_22524_, \oc8051_golden_model_1.TL0 [0]);
  nor _73009_ (_22525_, _01347_, _22524_);
  nand _73010_ (_22526_, _11263_, _07919_);
  nor _73011_ (_22528_, _07919_, _22524_);
  nor _73012_ (_22529_, _22528_, _07234_);
  nand _73013_ (_22530_, _22529_, _22526_);
  nor _73014_ (_22531_, _08390_, _11804_);
  or _73015_ (_22532_, _22531_, _22528_);
  or _73016_ (_22533_, _22532_, _07151_);
  and _73017_ (_22534_, _07919_, \oc8051_golden_model_1.ACC [0]);
  or _73018_ (_22535_, _22534_, _22528_);
  and _73019_ (_22536_, _22535_, _07141_);
  nor _73020_ (_22537_, _07141_, _22524_);
  or _73021_ (_22539_, _22537_, _06341_);
  or _73022_ (_22540_, _22539_, _22536_);
  and _73023_ (_22541_, _22540_, _07166_);
  and _73024_ (_22542_, _22541_, _22533_);
  and _73025_ (_22543_, _07919_, _07133_);
  or _73026_ (_22544_, _22543_, _22528_);
  and _73027_ (_22545_, _22544_, _06461_);
  or _73028_ (_22546_, _22545_, _22542_);
  and _73029_ (_22547_, _22546_, _06465_);
  and _73030_ (_22548_, _22535_, _06464_);
  or _73031_ (_22550_, _22548_, _10080_);
  or _73032_ (_22551_, _22550_, _22547_);
  or _73033_ (_22552_, _22544_, _07215_);
  and _73034_ (_22553_, _22552_, _22551_);
  or _73035_ (_22554_, _22553_, _07460_);
  and _73036_ (_22555_, _09392_, _07919_);
  or _73037_ (_22556_, _22528_, _07208_);
  or _73038_ (_22557_, _22556_, _22555_);
  and _73039_ (_22558_, _22557_, _22554_);
  or _73040_ (_22559_, _22558_, _10094_);
  and _73041_ (_22561_, _14467_, _07919_);
  or _73042_ (_22562_, _22528_, _05982_);
  or _73043_ (_22563_, _22562_, _22561_);
  and _73044_ (_22564_, _22563_, _06219_);
  and _73045_ (_22565_, _22564_, _22559_);
  and _73046_ (_22566_, _07919_, _08954_);
  or _73047_ (_22567_, _22566_, _22528_);
  and _73048_ (_22568_, _22567_, _06218_);
  or _73049_ (_22569_, _22568_, _06369_);
  or _73050_ (_22570_, _22569_, _22565_);
  and _73051_ (_22572_, _14366_, _07919_);
  or _73052_ (_22573_, _22572_, _22528_);
  or _73053_ (_22574_, _22573_, _07237_);
  and _73054_ (_22575_, _22574_, _07240_);
  and _73055_ (_22576_, _22575_, _22570_);
  nor _73056_ (_22577_, _12580_, _11804_);
  or _73057_ (_22578_, _22577_, _22528_);
  and _73058_ (_22579_, _22526_, _06536_);
  and _73059_ (_22580_, _22579_, _22578_);
  or _73060_ (_22581_, _22580_, _22576_);
  and _73061_ (_22583_, _22581_, _07242_);
  nand _73062_ (_22584_, _22567_, _06375_);
  nor _73063_ (_22585_, _22584_, _22531_);
  or _73064_ (_22586_, _22585_, _06545_);
  or _73065_ (_22587_, _22586_, _22583_);
  and _73066_ (_22588_, _22587_, _22530_);
  or _73067_ (_22589_, _22588_, _06366_);
  and _73068_ (_22590_, _14363_, _07919_);
  or _73069_ (_22591_, _22528_, _09056_);
  or _73070_ (_22592_, _22591_, _22590_);
  and _73071_ (_22594_, _22592_, _09061_);
  and _73072_ (_22595_, _22594_, _22589_);
  and _73073_ (_22596_, _22578_, _06528_);
  or _73074_ (_22597_, _22596_, _19502_);
  or _73075_ (_22598_, _22597_, _22595_);
  or _73076_ (_22599_, _22532_, _06661_);
  and _73077_ (_22600_, _22599_, _01347_);
  and _73078_ (_22601_, _22600_, _22598_);
  or _73079_ (_22602_, _22601_, _22525_);
  and _73080_ (_43211_, _22602_, _42618_);
  not _73081_ (_22604_, \oc8051_golden_model_1.TL0 [1]);
  nor _73082_ (_22605_, _01347_, _22604_);
  and _73083_ (_22606_, _09451_, _07919_);
  nor _73084_ (_22607_, _07919_, _22604_);
  or _73085_ (_22608_, _22607_, _07208_);
  or _73086_ (_22609_, _22608_, _22606_);
  nor _73087_ (_22610_, _11804_, _07357_);
  and _73088_ (_22611_, _07215_, _07166_);
  or _73089_ (_22612_, _22611_, _22607_);
  or _73090_ (_22613_, _22612_, _22610_);
  and _73091_ (_22614_, _07919_, \oc8051_golden_model_1.ACC [1]);
  or _73092_ (_22615_, _22614_, _22607_);
  and _73093_ (_22616_, _22615_, _06464_);
  or _73094_ (_22617_, _22616_, _10080_);
  or _73095_ (_22618_, _07919_, \oc8051_golden_model_1.TL0 [1]);
  and _73096_ (_22619_, _14562_, _07919_);
  not _73097_ (_22620_, _22619_);
  and _73098_ (_22621_, _22620_, _22618_);
  and _73099_ (_22622_, _22621_, _06341_);
  nor _73100_ (_22623_, _07141_, _22604_);
  and _73101_ (_22626_, _22615_, _07141_);
  or _73102_ (_22627_, _22626_, _22623_);
  and _73103_ (_22628_, _22627_, _07151_);
  or _73104_ (_22629_, _22628_, _06461_);
  or _73105_ (_22630_, _22629_, _22622_);
  and _73106_ (_22631_, _22630_, _06465_);
  or _73107_ (_22632_, _22631_, _22617_);
  and _73108_ (_22633_, _22632_, _22613_);
  or _73109_ (_22634_, _22633_, _07460_);
  and _73110_ (_22635_, _22634_, _05982_);
  and _73111_ (_22637_, _22635_, _22609_);
  or _73112_ (_22638_, _14653_, _11804_);
  and _73113_ (_22639_, _22618_, _10094_);
  and _73114_ (_22640_, _22639_, _22638_);
  or _73115_ (_22641_, _22640_, _22637_);
  and _73116_ (_22642_, _22641_, _06219_);
  nand _73117_ (_22643_, _07919_, _07038_);
  and _73118_ (_22644_, _22618_, _06218_);
  and _73119_ (_22645_, _22644_, _22643_);
  or _73120_ (_22646_, _22645_, _22642_);
  and _73121_ (_22648_, _22646_, _07237_);
  or _73122_ (_22649_, _14668_, _11804_);
  and _73123_ (_22650_, _22618_, _06369_);
  and _73124_ (_22651_, _22650_, _22649_);
  or _73125_ (_22652_, _22651_, _06536_);
  or _73126_ (_22653_, _22652_, _22648_);
  nor _73127_ (_22654_, _11261_, _11804_);
  or _73128_ (_22655_, _22654_, _22607_);
  nand _73129_ (_22656_, _11260_, _07919_);
  and _73130_ (_22657_, _22656_, _22655_);
  or _73131_ (_22659_, _22657_, _07240_);
  and _73132_ (_22660_, _22659_, _07242_);
  and _73133_ (_22661_, _22660_, _22653_);
  or _73134_ (_22662_, _14666_, _11804_);
  and _73135_ (_22663_, _22618_, _06375_);
  and _73136_ (_22664_, _22663_, _22662_);
  or _73137_ (_22665_, _22664_, _06545_);
  or _73138_ (_22666_, _22665_, _22661_);
  nor _73139_ (_22667_, _22607_, _07234_);
  nand _73140_ (_22668_, _22667_, _22656_);
  and _73141_ (_22670_, _22668_, _09056_);
  and _73142_ (_22671_, _22670_, _22666_);
  or _73143_ (_22672_, _22643_, _08341_);
  and _73144_ (_22673_, _22618_, _06366_);
  and _73145_ (_22674_, _22673_, _22672_);
  or _73146_ (_22675_, _22674_, _06528_);
  or _73147_ (_22676_, _22675_, _22671_);
  or _73148_ (_22677_, _22655_, _09061_);
  and _73149_ (_22678_, _22677_, _06926_);
  and _73150_ (_22679_, _22678_, _22676_);
  and _73151_ (_22681_, _22621_, _06568_);
  or _73152_ (_22682_, _22681_, _06278_);
  or _73153_ (_22683_, _22682_, _22679_);
  or _73154_ (_22684_, _22607_, _06279_);
  or _73155_ (_22685_, _22684_, _22619_);
  and _73156_ (_22686_, _22685_, _01347_);
  and _73157_ (_22687_, _22686_, _22683_);
  or _73158_ (_22688_, _22687_, _22605_);
  and _73159_ (_43212_, _22688_, _42618_);
  and _73160_ (_22689_, _01351_, \oc8051_golden_model_1.TL0 [2]);
  and _73161_ (_22691_, _11804_, \oc8051_golden_model_1.TL0 [2]);
  nor _73162_ (_22692_, _11804_, _07776_);
  or _73163_ (_22693_, _22692_, _22691_);
  or _73164_ (_22694_, _22693_, _07215_);
  and _73165_ (_22695_, _14770_, _07919_);
  or _73166_ (_22696_, _22695_, _22691_);
  and _73167_ (_22697_, _22696_, _06341_);
  and _73168_ (_22698_, _07142_, \oc8051_golden_model_1.TL0 [2]);
  and _73169_ (_22699_, _07919_, \oc8051_golden_model_1.ACC [2]);
  or _73170_ (_22700_, _22699_, _22691_);
  and _73171_ (_22702_, _22700_, _07141_);
  or _73172_ (_22703_, _22702_, _22698_);
  and _73173_ (_22704_, _22703_, _07151_);
  or _73174_ (_22705_, _22704_, _06461_);
  or _73175_ (_22706_, _22705_, _22697_);
  or _73176_ (_22707_, _22693_, _07166_);
  and _73177_ (_22708_, _22707_, _06465_);
  and _73178_ (_22709_, _22708_, _22706_);
  and _73179_ (_22710_, _22700_, _06464_);
  or _73180_ (_22711_, _22710_, _10080_);
  or _73181_ (_22713_, _22711_, _22709_);
  and _73182_ (_22714_, _22713_, _22694_);
  or _73183_ (_22715_, _22714_, _07460_);
  and _73184_ (_22716_, _09450_, _07919_);
  or _73185_ (_22717_, _22691_, _07208_);
  or _73186_ (_22718_, _22717_, _22716_);
  and _73187_ (_22719_, _22718_, _22715_);
  or _73188_ (_22720_, _22719_, _10094_);
  and _73189_ (_22721_, _14859_, _07919_);
  or _73190_ (_22722_, _22691_, _05982_);
  or _73191_ (_22724_, _22722_, _22721_);
  and _73192_ (_22725_, _22724_, _06219_);
  and _73193_ (_22726_, _22725_, _22720_);
  and _73194_ (_22727_, _07919_, _08973_);
  or _73195_ (_22728_, _22727_, _22691_);
  and _73196_ (_22729_, _22728_, _06218_);
  or _73197_ (_22730_, _22729_, _06369_);
  or _73198_ (_22731_, _22730_, _22726_);
  and _73199_ (_22732_, _14751_, _07919_);
  or _73200_ (_22733_, _22732_, _22691_);
  or _73201_ (_22735_, _22733_, _07237_);
  and _73202_ (_22736_, _22735_, _07240_);
  and _73203_ (_22737_, _22736_, _22731_);
  and _73204_ (_22738_, _11259_, _07919_);
  or _73205_ (_22739_, _22738_, _22691_);
  and _73206_ (_22740_, _22739_, _06536_);
  or _73207_ (_22741_, _22740_, _22737_);
  and _73208_ (_22742_, _22741_, _07242_);
  or _73209_ (_22743_, _22691_, _08440_);
  and _73210_ (_22744_, _22728_, _06375_);
  and _73211_ (_22746_, _22744_, _22743_);
  or _73212_ (_22747_, _22746_, _22742_);
  and _73213_ (_22748_, _22747_, _07234_);
  and _73214_ (_22749_, _22700_, _06545_);
  and _73215_ (_22750_, _22749_, _22743_);
  or _73216_ (_22751_, _22750_, _06366_);
  or _73217_ (_22752_, _22751_, _22748_);
  and _73218_ (_22753_, _14748_, _07919_);
  or _73219_ (_22754_, _22691_, _09056_);
  or _73220_ (_22755_, _22754_, _22753_);
  and _73221_ (_22757_, _22755_, _09061_);
  and _73222_ (_22758_, _22757_, _22752_);
  nor _73223_ (_22759_, _11258_, _11804_);
  or _73224_ (_22760_, _22759_, _22691_);
  and _73225_ (_22761_, _22760_, _06528_);
  or _73226_ (_22762_, _22761_, _22758_);
  and _73227_ (_22763_, _22762_, _06926_);
  and _73228_ (_22764_, _22696_, _06568_);
  or _73229_ (_22765_, _22764_, _06278_);
  or _73230_ (_22766_, _22765_, _22763_);
  and _73231_ (_22768_, _14926_, _07919_);
  or _73232_ (_22769_, _22691_, _06279_);
  or _73233_ (_22770_, _22769_, _22768_);
  and _73234_ (_22771_, _22770_, _01347_);
  and _73235_ (_22772_, _22771_, _22766_);
  or _73236_ (_22773_, _22772_, _22689_);
  and _73237_ (_43213_, _22773_, _42618_);
  and _73238_ (_22774_, _01351_, \oc8051_golden_model_1.TL0 [3]);
  and _73239_ (_22775_, _11804_, \oc8051_golden_model_1.TL0 [3]);
  and _73240_ (_22776_, _14953_, _07919_);
  or _73241_ (_22778_, _22776_, _22775_);
  or _73242_ (_22779_, _22778_, _07151_);
  and _73243_ (_22780_, _07919_, \oc8051_golden_model_1.ACC [3]);
  or _73244_ (_22781_, _22780_, _22775_);
  and _73245_ (_22782_, _22781_, _07141_);
  and _73246_ (_22783_, _07142_, \oc8051_golden_model_1.TL0 [3]);
  or _73247_ (_22784_, _22783_, _06341_);
  or _73248_ (_22785_, _22784_, _22782_);
  and _73249_ (_22786_, _22785_, _07166_);
  and _73250_ (_22787_, _22786_, _22779_);
  nor _73251_ (_22789_, _11804_, _07594_);
  or _73252_ (_22790_, _22789_, _22775_);
  and _73253_ (_22791_, _22790_, _06461_);
  or _73254_ (_22792_, _22791_, _22787_);
  and _73255_ (_22793_, _22792_, _06465_);
  and _73256_ (_22794_, _22781_, _06464_);
  or _73257_ (_22795_, _22794_, _10080_);
  or _73258_ (_22796_, _22795_, _22793_);
  or _73259_ (_22797_, _22790_, _07215_);
  and _73260_ (_22798_, _22797_, _22796_);
  or _73261_ (_22800_, _22798_, _07460_);
  and _73262_ (_22801_, _09449_, _07919_);
  or _73263_ (_22802_, _22775_, _07208_);
  or _73264_ (_22803_, _22802_, _22801_);
  and _73265_ (_22804_, _22803_, _05982_);
  and _73266_ (_22805_, _22804_, _22800_);
  and _73267_ (_22806_, _15048_, _07919_);
  or _73268_ (_22807_, _22806_, _22775_);
  and _73269_ (_22808_, _22807_, _10094_);
  or _73270_ (_22809_, _22808_, _06218_);
  or _73271_ (_22811_, _22809_, _22805_);
  and _73272_ (_22812_, _07919_, _08930_);
  or _73273_ (_22813_, _22812_, _22775_);
  or _73274_ (_22814_, _22813_, _06219_);
  and _73275_ (_22815_, _22814_, _22811_);
  or _73276_ (_22816_, _22815_, _06369_);
  and _73277_ (_22817_, _14943_, _07919_);
  or _73278_ (_22818_, _22817_, _22775_);
  or _73279_ (_22819_, _22818_, _07237_);
  and _73280_ (_22820_, _22819_, _07240_);
  and _73281_ (_22822_, _22820_, _22816_);
  and _73282_ (_22823_, _12577_, _07919_);
  or _73283_ (_22824_, _22823_, _22775_);
  and _73284_ (_22825_, _22824_, _06536_);
  or _73285_ (_22826_, _22825_, _22822_);
  and _73286_ (_22827_, _22826_, _07242_);
  or _73287_ (_22828_, _22775_, _08292_);
  and _73288_ (_22829_, _22813_, _06375_);
  and _73289_ (_22830_, _22829_, _22828_);
  or _73290_ (_22831_, _22830_, _22827_);
  and _73291_ (_22832_, _22831_, _07234_);
  and _73292_ (_22833_, _22781_, _06545_);
  and _73293_ (_22834_, _22833_, _22828_);
  or _73294_ (_22835_, _22834_, _06366_);
  or _73295_ (_22836_, _22835_, _22832_);
  and _73296_ (_22837_, _14940_, _07919_);
  or _73297_ (_22838_, _22775_, _09056_);
  or _73298_ (_22839_, _22838_, _22837_);
  and _73299_ (_22840_, _22839_, _09061_);
  and _73300_ (_22841_, _22840_, _22836_);
  nor _73301_ (_22844_, _11256_, _11804_);
  or _73302_ (_22845_, _22844_, _22775_);
  and _73303_ (_22846_, _22845_, _06528_);
  or _73304_ (_22847_, _22846_, _22841_);
  and _73305_ (_22848_, _22847_, _06926_);
  and _73306_ (_22849_, _22778_, _06568_);
  or _73307_ (_22850_, _22849_, _06278_);
  or _73308_ (_22851_, _22850_, _22848_);
  and _73309_ (_22852_, _15128_, _07919_);
  or _73310_ (_22853_, _22775_, _06279_);
  or _73311_ (_22855_, _22853_, _22852_);
  and _73312_ (_22856_, _22855_, _01347_);
  and _73313_ (_22857_, _22856_, _22851_);
  or _73314_ (_22858_, _22857_, _22774_);
  and _73315_ (_43214_, _22858_, _42618_);
  and _73316_ (_22859_, _01351_, \oc8051_golden_model_1.TL0 [4]);
  and _73317_ (_22860_, _11804_, \oc8051_golden_model_1.TL0 [4]);
  nor _73318_ (_22861_, _08541_, _11804_);
  or _73319_ (_22862_, _22861_, _22860_);
  or _73320_ (_22863_, _22862_, _07215_);
  and _73321_ (_22865_, _15162_, _07919_);
  or _73322_ (_22866_, _22865_, _22860_);
  or _73323_ (_22867_, _22866_, _07151_);
  and _73324_ (_22868_, _07919_, \oc8051_golden_model_1.ACC [4]);
  or _73325_ (_22869_, _22868_, _22860_);
  and _73326_ (_22870_, _22869_, _07141_);
  and _73327_ (_22871_, _07142_, \oc8051_golden_model_1.TL0 [4]);
  or _73328_ (_22872_, _22871_, _06341_);
  or _73329_ (_22873_, _22872_, _22870_);
  and _73330_ (_22874_, _22873_, _07166_);
  and _73331_ (_22876_, _22874_, _22867_);
  and _73332_ (_22877_, _22862_, _06461_);
  or _73333_ (_22878_, _22877_, _22876_);
  and _73334_ (_22879_, _22878_, _06465_);
  and _73335_ (_22880_, _22869_, _06464_);
  or _73336_ (_22881_, _22880_, _10080_);
  or _73337_ (_22882_, _22881_, _22879_);
  and _73338_ (_22883_, _22882_, _22863_);
  or _73339_ (_22884_, _22883_, _07460_);
  and _73340_ (_22885_, _09448_, _07919_);
  or _73341_ (_22887_, _22860_, _07208_);
  or _73342_ (_22888_, _22887_, _22885_);
  and _73343_ (_22889_, _22888_, _22884_);
  or _73344_ (_22890_, _22889_, _10094_);
  and _73345_ (_22891_, _15254_, _07919_);
  or _73346_ (_22892_, _22860_, _05982_);
  or _73347_ (_22893_, _22892_, _22891_);
  and _73348_ (_22894_, _22893_, _06219_);
  and _73349_ (_22895_, _22894_, _22890_);
  and _73350_ (_22896_, _08959_, _07919_);
  or _73351_ (_22898_, _22896_, _22860_);
  and _73352_ (_22899_, _22898_, _06218_);
  or _73353_ (_22900_, _22899_, _06369_);
  or _73354_ (_22901_, _22900_, _22895_);
  and _73355_ (_22902_, _15269_, _07919_);
  or _73356_ (_22903_, _22902_, _22860_);
  or _73357_ (_22904_, _22903_, _07237_);
  and _73358_ (_22905_, _22904_, _07240_);
  and _73359_ (_22906_, _22905_, _22901_);
  and _73360_ (_22907_, _11254_, _07919_);
  or _73361_ (_22909_, _22907_, _22860_);
  and _73362_ (_22910_, _22909_, _06536_);
  or _73363_ (_22911_, _22910_, _22906_);
  and _73364_ (_22912_, _22911_, _07242_);
  or _73365_ (_22913_, _22860_, _08544_);
  and _73366_ (_22914_, _22898_, _06375_);
  and _73367_ (_22915_, _22914_, _22913_);
  or _73368_ (_22916_, _22915_, _22912_);
  and _73369_ (_22917_, _22916_, _07234_);
  and _73370_ (_22918_, _22869_, _06545_);
  and _73371_ (_22920_, _22918_, _22913_);
  or _73372_ (_22921_, _22920_, _06366_);
  or _73373_ (_22922_, _22921_, _22917_);
  and _73374_ (_22923_, _15266_, _07919_);
  or _73375_ (_22924_, _22860_, _09056_);
  or _73376_ (_22925_, _22924_, _22923_);
  and _73377_ (_22926_, _22925_, _09061_);
  and _73378_ (_22927_, _22926_, _22922_);
  nor _73379_ (_22928_, _11253_, _11804_);
  or _73380_ (_22929_, _22928_, _22860_);
  and _73381_ (_22931_, _22929_, _06528_);
  or _73382_ (_22932_, _22931_, _22927_);
  and _73383_ (_22933_, _22932_, _06926_);
  and _73384_ (_22934_, _22866_, _06568_);
  or _73385_ (_22935_, _22934_, _06278_);
  or _73386_ (_22936_, _22935_, _22933_);
  and _73387_ (_22937_, _15329_, _07919_);
  or _73388_ (_22938_, _22860_, _06279_);
  or _73389_ (_22939_, _22938_, _22937_);
  and _73390_ (_22940_, _22939_, _01347_);
  and _73391_ (_22942_, _22940_, _22936_);
  or _73392_ (_22943_, _22942_, _22859_);
  and _73393_ (_43215_, _22943_, _42618_);
  and _73394_ (_22944_, _01351_, \oc8051_golden_model_1.TL0 [5]);
  and _73395_ (_22945_, _11804_, \oc8051_golden_model_1.TL0 [5]);
  nor _73396_ (_22946_, _08244_, _11804_);
  or _73397_ (_22947_, _22946_, _22945_);
  or _73398_ (_22948_, _22947_, _07215_);
  and _73399_ (_22949_, _15358_, _07919_);
  or _73400_ (_22950_, _22949_, _22945_);
  or _73401_ (_22952_, _22950_, _07151_);
  and _73402_ (_22953_, _07919_, \oc8051_golden_model_1.ACC [5]);
  or _73403_ (_22954_, _22953_, _22945_);
  and _73404_ (_22955_, _22954_, _07141_);
  and _73405_ (_22956_, _07142_, \oc8051_golden_model_1.TL0 [5]);
  or _73406_ (_22957_, _22956_, _06341_);
  or _73407_ (_22958_, _22957_, _22955_);
  and _73408_ (_22959_, _22958_, _07166_);
  and _73409_ (_22960_, _22959_, _22952_);
  and _73410_ (_22961_, _22947_, _06461_);
  or _73411_ (_22963_, _22961_, _22960_);
  and _73412_ (_22964_, _22963_, _06465_);
  and _73413_ (_22965_, _22954_, _06464_);
  or _73414_ (_22966_, _22965_, _10080_);
  or _73415_ (_22967_, _22966_, _22964_);
  and _73416_ (_22968_, _22967_, _22948_);
  or _73417_ (_22969_, _22968_, _07460_);
  and _73418_ (_22970_, _09447_, _07919_);
  or _73419_ (_22971_, _22945_, _07208_);
  or _73420_ (_22972_, _22971_, _22970_);
  and _73421_ (_22974_, _22972_, _05982_);
  and _73422_ (_22975_, _22974_, _22969_);
  and _73423_ (_22976_, _15459_, _07919_);
  or _73424_ (_22977_, _22976_, _22945_);
  and _73425_ (_22978_, _22977_, _10094_);
  or _73426_ (_22979_, _22978_, _06218_);
  or _73427_ (_22980_, _22979_, _22975_);
  and _73428_ (_22981_, _08946_, _07919_);
  or _73429_ (_22982_, _22981_, _22945_);
  or _73430_ (_22983_, _22982_, _06219_);
  and _73431_ (_22985_, _22983_, _22980_);
  or _73432_ (_22986_, _22985_, _06369_);
  and _73433_ (_22987_, _15353_, _07919_);
  or _73434_ (_22988_, _22987_, _22945_);
  or _73435_ (_22989_, _22988_, _07237_);
  and _73436_ (_22990_, _22989_, _07240_);
  and _73437_ (_22991_, _22990_, _22986_);
  and _73438_ (_22992_, _11250_, _07919_);
  or _73439_ (_22993_, _22992_, _22945_);
  and _73440_ (_22994_, _22993_, _06536_);
  or _73441_ (_22996_, _22994_, _22991_);
  and _73442_ (_22997_, _22996_, _07242_);
  or _73443_ (_22998_, _22945_, _08247_);
  and _73444_ (_22999_, _22982_, _06375_);
  and _73445_ (_23000_, _22999_, _22998_);
  or _73446_ (_23001_, _23000_, _22997_);
  and _73447_ (_23002_, _23001_, _07234_);
  and _73448_ (_23003_, _22954_, _06545_);
  and _73449_ (_23004_, _23003_, _22998_);
  or _73450_ (_23005_, _23004_, _06366_);
  or _73451_ (_23007_, _23005_, _23002_);
  and _73452_ (_23008_, _15350_, _07919_);
  or _73453_ (_23009_, _22945_, _09056_);
  or _73454_ (_23010_, _23009_, _23008_);
  and _73455_ (_23011_, _23010_, _09061_);
  and _73456_ (_23012_, _23011_, _23007_);
  nor _73457_ (_23013_, _11249_, _11804_);
  or _73458_ (_23014_, _23013_, _22945_);
  and _73459_ (_23015_, _23014_, _06528_);
  or _73460_ (_23016_, _23015_, _23012_);
  and _73461_ (_23018_, _23016_, _06926_);
  and _73462_ (_23019_, _22950_, _06568_);
  or _73463_ (_23020_, _23019_, _06278_);
  or _73464_ (_23021_, _23020_, _23018_);
  and _73465_ (_23022_, _15532_, _07919_);
  or _73466_ (_23023_, _22945_, _06279_);
  or _73467_ (_23024_, _23023_, _23022_);
  and _73468_ (_23025_, _23024_, _01347_);
  and _73469_ (_23026_, _23025_, _23021_);
  or _73470_ (_23027_, _23026_, _22944_);
  and _73471_ (_43216_, _23027_, _42618_);
  and _73472_ (_23029_, _01351_, \oc8051_golden_model_1.TL0 [6]);
  and _73473_ (_23030_, _11804_, \oc8051_golden_model_1.TL0 [6]);
  nor _73474_ (_23031_, _08142_, _11804_);
  or _73475_ (_23032_, _23031_, _23030_);
  or _73476_ (_23033_, _23032_, _07215_);
  and _73477_ (_23034_, _15554_, _07919_);
  or _73478_ (_23035_, _23034_, _23030_);
  or _73479_ (_23036_, _23035_, _07151_);
  and _73480_ (_23037_, _07919_, \oc8051_golden_model_1.ACC [6]);
  or _73481_ (_23039_, _23037_, _23030_);
  and _73482_ (_23040_, _23039_, _07141_);
  and _73483_ (_23041_, _07142_, \oc8051_golden_model_1.TL0 [6]);
  or _73484_ (_23042_, _23041_, _06341_);
  or _73485_ (_23043_, _23042_, _23040_);
  and _73486_ (_23044_, _23043_, _07166_);
  and _73487_ (_23045_, _23044_, _23036_);
  and _73488_ (_23046_, _23032_, _06461_);
  or _73489_ (_23047_, _23046_, _23045_);
  and _73490_ (_23048_, _23047_, _06465_);
  and _73491_ (_23050_, _23039_, _06464_);
  or _73492_ (_23051_, _23050_, _10080_);
  or _73493_ (_23052_, _23051_, _23048_);
  and _73494_ (_23053_, _23052_, _23033_);
  or _73495_ (_23054_, _23053_, _07460_);
  and _73496_ (_23055_, _09446_, _07919_);
  or _73497_ (_23056_, _23030_, _07208_);
  or _73498_ (_23057_, _23056_, _23055_);
  and _73499_ (_23058_, _23057_, _05982_);
  and _73500_ (_23059_, _23058_, _23054_);
  and _73501_ (_23061_, _15657_, _07919_);
  or _73502_ (_23062_, _23061_, _23030_);
  and _73503_ (_23063_, _23062_, _10094_);
  or _73504_ (_23064_, _23063_, _06218_);
  or _73505_ (_23065_, _23064_, _23059_);
  and _73506_ (_23066_, _15664_, _07919_);
  or _73507_ (_23067_, _23066_, _23030_);
  or _73508_ (_23068_, _23067_, _06219_);
  and _73509_ (_23069_, _23068_, _23065_);
  or _73510_ (_23070_, _23069_, _06369_);
  and _73511_ (_23072_, _15549_, _07919_);
  or _73512_ (_23073_, _23072_, _23030_);
  or _73513_ (_23074_, _23073_, _07237_);
  and _73514_ (_23075_, _23074_, _07240_);
  and _73515_ (_23076_, _23075_, _23070_);
  and _73516_ (_23077_, _11247_, _07919_);
  or _73517_ (_23078_, _23077_, _23030_);
  and _73518_ (_23079_, _23078_, _06536_);
  or _73519_ (_23080_, _23079_, _23076_);
  and _73520_ (_23081_, _23080_, _07242_);
  or _73521_ (_23083_, _23030_, _08145_);
  and _73522_ (_23084_, _23067_, _06375_);
  and _73523_ (_23085_, _23084_, _23083_);
  or _73524_ (_23086_, _23085_, _23081_);
  and _73525_ (_23087_, _23086_, _07234_);
  and _73526_ (_23088_, _23039_, _06545_);
  and _73527_ (_23089_, _23088_, _23083_);
  or _73528_ (_23090_, _23089_, _06366_);
  or _73529_ (_23091_, _23090_, _23087_);
  and _73530_ (_23092_, _15546_, _07919_);
  or _73531_ (_23093_, _23030_, _09056_);
  or _73532_ (_23094_, _23093_, _23092_);
  and _73533_ (_23095_, _23094_, _09061_);
  and _73534_ (_23096_, _23095_, _23091_);
  nor _73535_ (_23097_, _11246_, _11804_);
  or _73536_ (_23098_, _23097_, _23030_);
  and _73537_ (_23099_, _23098_, _06528_);
  or _73538_ (_23100_, _23099_, _23096_);
  and _73539_ (_23101_, _23100_, _06926_);
  and _73540_ (_23102_, _23035_, _06568_);
  or _73541_ (_23105_, _23102_, _06278_);
  or _73542_ (_23106_, _23105_, _23101_);
  and _73543_ (_23107_, _15734_, _07919_);
  or _73544_ (_23108_, _23030_, _06279_);
  or _73545_ (_23109_, _23108_, _23107_);
  and _73546_ (_23110_, _23109_, _01347_);
  and _73547_ (_23111_, _23110_, _23106_);
  or _73548_ (_23112_, _23111_, _23029_);
  and _73549_ (_43217_, _23112_, _42618_);
  not _73550_ (_23113_, \oc8051_golden_model_1.TCON [0]);
  nor _73551_ (_23115_, _01347_, _23113_);
  nand _73552_ (_23116_, _11263_, _07928_);
  nor _73553_ (_23117_, _07928_, _23113_);
  nor _73554_ (_23118_, _23117_, _07234_);
  nand _73555_ (_23119_, _23118_, _23116_);
  and _73556_ (_23120_, _07928_, _07133_);
  or _73557_ (_23121_, _23120_, _23117_);
  or _73558_ (_23122_, _23121_, _07215_);
  nor _73559_ (_23123_, _08390_, _11882_);
  or _73560_ (_23124_, _23123_, _23117_);
  or _73561_ (_23126_, _23124_, _07151_);
  and _73562_ (_23127_, _07928_, \oc8051_golden_model_1.ACC [0]);
  or _73563_ (_23128_, _23127_, _23117_);
  and _73564_ (_23129_, _23128_, _07141_);
  nor _73565_ (_23130_, _07141_, _23113_);
  or _73566_ (_23131_, _23130_, _06341_);
  or _73567_ (_23132_, _23131_, _23129_);
  and _73568_ (_23133_, _23132_, _06273_);
  and _73569_ (_23134_, _23133_, _23126_);
  nor _73570_ (_23135_, _08616_, _23113_);
  and _73571_ (_23137_, _14382_, _08616_);
  or _73572_ (_23138_, _23137_, _23135_);
  and _73573_ (_23139_, _23138_, _06272_);
  or _73574_ (_23140_, _23139_, _23134_);
  and _73575_ (_23141_, _23140_, _07166_);
  and _73576_ (_23142_, _23121_, _06461_);
  or _73577_ (_23143_, _23142_, _06464_);
  or _73578_ (_23144_, _23143_, _23141_);
  or _73579_ (_23145_, _23128_, _06465_);
  and _73580_ (_23146_, _23145_, _06269_);
  and _73581_ (_23148_, _23146_, _23144_);
  and _73582_ (_23149_, _23117_, _06268_);
  or _73583_ (_23150_, _23149_, _06261_);
  or _73584_ (_23151_, _23150_, _23148_);
  or _73585_ (_23152_, _23124_, _06262_);
  and _73586_ (_23153_, _23152_, _06258_);
  and _73587_ (_23154_, _23153_, _23151_);
  and _73588_ (_23155_, _14413_, _08616_);
  or _73589_ (_23156_, _23155_, _23135_);
  and _73590_ (_23157_, _23156_, _06257_);
  or _73591_ (_23159_, _23157_, _10080_);
  or _73592_ (_23160_, _23159_, _23154_);
  and _73593_ (_23161_, _23160_, _23122_);
  or _73594_ (_23162_, _23161_, _07460_);
  and _73595_ (_23163_, _09392_, _07928_);
  or _73596_ (_23164_, _23117_, _07208_);
  or _73597_ (_23165_, _23164_, _23163_);
  and _73598_ (_23166_, _23165_, _23162_);
  or _73599_ (_23167_, _23166_, _10094_);
  and _73600_ (_23168_, _14467_, _07928_);
  or _73601_ (_23170_, _23117_, _05982_);
  or _73602_ (_23171_, _23170_, _23168_);
  and _73603_ (_23172_, _23171_, _06219_);
  and _73604_ (_23173_, _23172_, _23167_);
  and _73605_ (_23174_, _07928_, _08954_);
  or _73606_ (_23175_, _23174_, _23117_);
  and _73607_ (_23176_, _23175_, _06218_);
  or _73608_ (_23177_, _23176_, _06369_);
  or _73609_ (_23178_, _23177_, _23173_);
  and _73610_ (_23179_, _14366_, _07928_);
  or _73611_ (_23181_, _23179_, _23117_);
  or _73612_ (_23182_, _23181_, _07237_);
  and _73613_ (_23183_, _23182_, _07240_);
  and _73614_ (_23184_, _23183_, _23178_);
  nor _73615_ (_23185_, _12580_, _11882_);
  or _73616_ (_23186_, _23185_, _23117_);
  and _73617_ (_23187_, _23116_, _06536_);
  and _73618_ (_23188_, _23187_, _23186_);
  or _73619_ (_23189_, _23188_, _23184_);
  and _73620_ (_23190_, _23189_, _07242_);
  nand _73621_ (_23192_, _23175_, _06375_);
  nor _73622_ (_23193_, _23192_, _23123_);
  or _73623_ (_23194_, _23193_, _06545_);
  or _73624_ (_23195_, _23194_, _23190_);
  and _73625_ (_23196_, _23195_, _23119_);
  or _73626_ (_23197_, _23196_, _06366_);
  and _73627_ (_23198_, _14363_, _07928_);
  or _73628_ (_23199_, _23117_, _09056_);
  or _73629_ (_23200_, _23199_, _23198_);
  and _73630_ (_23201_, _23200_, _09061_);
  and _73631_ (_23203_, _23201_, _23197_);
  and _73632_ (_23204_, _23186_, _06528_);
  or _73633_ (_23205_, _23204_, _06568_);
  or _73634_ (_23206_, _23205_, _23203_);
  or _73635_ (_23207_, _23124_, _06926_);
  and _73636_ (_23208_, _23207_, _23206_);
  or _73637_ (_23209_, _23208_, _05927_);
  or _73638_ (_23210_, _23117_, _05928_);
  and _73639_ (_23211_, _23210_, _23209_);
  or _73640_ (_23212_, _23211_, _06278_);
  or _73641_ (_23214_, _23124_, _06279_);
  and _73642_ (_23215_, _23214_, _01347_);
  and _73643_ (_23216_, _23215_, _23212_);
  or _73644_ (_23217_, _23216_, _23115_);
  and _73645_ (_43219_, _23217_, _42618_);
  not _73646_ (_23218_, \oc8051_golden_model_1.TCON [1]);
  nor _73647_ (_23219_, _01347_, _23218_);
  nor _73648_ (_23220_, _07928_, _23218_);
  nor _73649_ (_23221_, _11261_, _11882_);
  or _73650_ (_23222_, _23221_, _23220_);
  or _73651_ (_23224_, _23222_, _09061_);
  nor _73652_ (_23225_, _11882_, _07357_);
  or _73653_ (_23226_, _23225_, _23220_);
  or _73654_ (_23227_, _23226_, _07166_);
  or _73655_ (_23228_, _07928_, \oc8051_golden_model_1.TCON [1]);
  and _73656_ (_23229_, _14562_, _07928_);
  not _73657_ (_23230_, _23229_);
  and _73658_ (_23231_, _23230_, _23228_);
  or _73659_ (_23232_, _23231_, _07151_);
  and _73660_ (_23233_, _07928_, \oc8051_golden_model_1.ACC [1]);
  or _73661_ (_23235_, _23233_, _23220_);
  and _73662_ (_23236_, _23235_, _07141_);
  nor _73663_ (_23237_, _07141_, _23218_);
  or _73664_ (_23238_, _23237_, _06341_);
  or _73665_ (_23239_, _23238_, _23236_);
  and _73666_ (_23240_, _23239_, _06273_);
  and _73667_ (_23241_, _23240_, _23232_);
  nor _73668_ (_23242_, _08616_, _23218_);
  and _73669_ (_23243_, _14557_, _08616_);
  or _73670_ (_23244_, _23243_, _23242_);
  and _73671_ (_23246_, _23244_, _06272_);
  or _73672_ (_23247_, _23246_, _06461_);
  or _73673_ (_23248_, _23247_, _23241_);
  and _73674_ (_23249_, _23248_, _23227_);
  or _73675_ (_23250_, _23249_, _06464_);
  or _73676_ (_23251_, _23235_, _06465_);
  and _73677_ (_23252_, _23251_, _06269_);
  and _73678_ (_23253_, _23252_, _23250_);
  and _73679_ (_23254_, _14560_, _08616_);
  or _73680_ (_23255_, _23254_, _23242_);
  and _73681_ (_23257_, _23255_, _06268_);
  or _73682_ (_23258_, _23257_, _06261_);
  or _73683_ (_23259_, _23258_, _23253_);
  and _73684_ (_23260_, _23243_, _14556_);
  or _73685_ (_23261_, _23242_, _06262_);
  or _73686_ (_23262_, _23261_, _23260_);
  and _73687_ (_23263_, _23262_, _06258_);
  and _73688_ (_23264_, _23263_, _23259_);
  or _73689_ (_23265_, _23242_, _14597_);
  and _73690_ (_23266_, _23265_, _06257_);
  and _73691_ (_23268_, _23266_, _23244_);
  or _73692_ (_23269_, _23268_, _10080_);
  or _73693_ (_23270_, _23269_, _23264_);
  or _73694_ (_23271_, _23226_, _07215_);
  and _73695_ (_23272_, _23271_, _23270_);
  or _73696_ (_23273_, _23272_, _07460_);
  and _73697_ (_23274_, _09451_, _07928_);
  or _73698_ (_23275_, _23220_, _07208_);
  or _73699_ (_23276_, _23275_, _23274_);
  and _73700_ (_23277_, _23276_, _05982_);
  and _73701_ (_23279_, _23277_, _23273_);
  and _73702_ (_23280_, _14653_, _07928_);
  or _73703_ (_23281_, _23280_, _23220_);
  and _73704_ (_23282_, _23281_, _10094_);
  or _73705_ (_23283_, _23282_, _23279_);
  and _73706_ (_23284_, _23283_, _06219_);
  nand _73707_ (_23285_, _07928_, _07038_);
  and _73708_ (_23286_, _23228_, _06218_);
  and _73709_ (_23287_, _23286_, _23285_);
  or _73710_ (_23288_, _23287_, _23284_);
  and _73711_ (_23290_, _23288_, _07237_);
  or _73712_ (_23291_, _14668_, _11882_);
  and _73713_ (_23292_, _23228_, _06369_);
  and _73714_ (_23293_, _23292_, _23291_);
  or _73715_ (_23294_, _23293_, _06536_);
  or _73716_ (_23295_, _23294_, _23290_);
  nand _73717_ (_23296_, _11260_, _07928_);
  and _73718_ (_23297_, _23296_, _23222_);
  or _73719_ (_23298_, _23297_, _07240_);
  and _73720_ (_23299_, _23298_, _07242_);
  and _73721_ (_23301_, _23299_, _23295_);
  or _73722_ (_23302_, _14666_, _11882_);
  and _73723_ (_23303_, _23228_, _06375_);
  and _73724_ (_23304_, _23303_, _23302_);
  or _73725_ (_23305_, _23304_, _06545_);
  or _73726_ (_23306_, _23305_, _23301_);
  nor _73727_ (_23307_, _23220_, _07234_);
  nand _73728_ (_23308_, _23307_, _23296_);
  and _73729_ (_23309_, _23308_, _09056_);
  and _73730_ (_23310_, _23309_, _23306_);
  or _73731_ (_23312_, _23285_, _08341_);
  and _73732_ (_23313_, _23228_, _06366_);
  and _73733_ (_23314_, _23313_, _23312_);
  or _73734_ (_23315_, _23314_, _06528_);
  or _73735_ (_23316_, _23315_, _23310_);
  and _73736_ (_23317_, _23316_, _23224_);
  or _73737_ (_23318_, _23317_, _06568_);
  or _73738_ (_23319_, _23231_, _06926_);
  and _73739_ (_23320_, _23319_, _05928_);
  and _73740_ (_23321_, _23320_, _23318_);
  and _73741_ (_23323_, _23255_, _05927_);
  or _73742_ (_23324_, _23323_, _06278_);
  or _73743_ (_23325_, _23324_, _23321_);
  or _73744_ (_23326_, _23220_, _06279_);
  or _73745_ (_23327_, _23326_, _23229_);
  and _73746_ (_23328_, _23327_, _01347_);
  and _73747_ (_23329_, _23328_, _23325_);
  or _73748_ (_23330_, _23329_, _23219_);
  and _73749_ (_43220_, _23330_, _42618_);
  and _73750_ (_23331_, _01351_, \oc8051_golden_model_1.TCON [2]);
  and _73751_ (_23333_, _11882_, \oc8051_golden_model_1.TCON [2]);
  nor _73752_ (_23334_, _11882_, _07776_);
  or _73753_ (_23335_, _23334_, _23333_);
  or _73754_ (_23336_, _23335_, _07215_);
  or _73755_ (_23337_, _23335_, _07166_);
  and _73756_ (_23338_, _14770_, _07928_);
  or _73757_ (_23339_, _23338_, _23333_);
  or _73758_ (_23340_, _23339_, _07151_);
  and _73759_ (_23341_, _07928_, \oc8051_golden_model_1.ACC [2]);
  or _73760_ (_23342_, _23341_, _23333_);
  and _73761_ (_23344_, _23342_, _07141_);
  and _73762_ (_23345_, _07142_, \oc8051_golden_model_1.TCON [2]);
  or _73763_ (_23346_, _23345_, _06341_);
  or _73764_ (_23347_, _23346_, _23344_);
  and _73765_ (_23348_, _23347_, _06273_);
  and _73766_ (_23349_, _23348_, _23340_);
  and _73767_ (_23350_, _11890_, \oc8051_golden_model_1.TCON [2]);
  and _73768_ (_23351_, _14774_, _08616_);
  or _73769_ (_23352_, _23351_, _23350_);
  and _73770_ (_23353_, _23352_, _06272_);
  or _73771_ (_23355_, _23353_, _06461_);
  or _73772_ (_23356_, _23355_, _23349_);
  and _73773_ (_23357_, _23356_, _23337_);
  or _73774_ (_23358_, _23357_, _06464_);
  or _73775_ (_23359_, _23342_, _06465_);
  and _73776_ (_23360_, _23359_, _06269_);
  and _73777_ (_23361_, _23360_, _23358_);
  and _73778_ (_23362_, _14756_, _08616_);
  or _73779_ (_23363_, _23362_, _23350_);
  and _73780_ (_23364_, _23363_, _06268_);
  or _73781_ (_23366_, _23364_, _06261_);
  or _73782_ (_23367_, _23366_, _23361_);
  and _73783_ (_23368_, _23351_, _14789_);
  or _73784_ (_23369_, _23350_, _06262_);
  or _73785_ (_23370_, _23369_, _23368_);
  and _73786_ (_23371_, _23370_, _06258_);
  and _73787_ (_23372_, _23371_, _23367_);
  and _73788_ (_23373_, _14804_, _08616_);
  or _73789_ (_23374_, _23373_, _23350_);
  and _73790_ (_23375_, _23374_, _06257_);
  or _73791_ (_23376_, _23375_, _10080_);
  or _73792_ (_23377_, _23376_, _23372_);
  and _73793_ (_23378_, _23377_, _23336_);
  or _73794_ (_23379_, _23378_, _07460_);
  and _73795_ (_23380_, _09450_, _07928_);
  or _73796_ (_23381_, _23333_, _07208_);
  or _73797_ (_23382_, _23381_, _23380_);
  and _73798_ (_23383_, _23382_, _05982_);
  and _73799_ (_23384_, _23383_, _23379_);
  and _73800_ (_23385_, _14859_, _07928_);
  or _73801_ (_23388_, _23385_, _23333_);
  and _73802_ (_23389_, _23388_, _10094_);
  or _73803_ (_23390_, _23389_, _06218_);
  or _73804_ (_23391_, _23390_, _23384_);
  and _73805_ (_23392_, _07928_, _08973_);
  or _73806_ (_23393_, _23392_, _23333_);
  or _73807_ (_23394_, _23393_, _06219_);
  and _73808_ (_23395_, _23394_, _23391_);
  or _73809_ (_23396_, _23395_, _06369_);
  and _73810_ (_23397_, _14751_, _07928_);
  or _73811_ (_23399_, _23397_, _23333_);
  or _73812_ (_23400_, _23399_, _07237_);
  and _73813_ (_23401_, _23400_, _07240_);
  and _73814_ (_23402_, _23401_, _23396_);
  and _73815_ (_23403_, _11259_, _07928_);
  or _73816_ (_23404_, _23403_, _23333_);
  and _73817_ (_23405_, _23404_, _06536_);
  or _73818_ (_23406_, _23405_, _23402_);
  and _73819_ (_23407_, _23406_, _07242_);
  or _73820_ (_23408_, _23333_, _08440_);
  and _73821_ (_23410_, _23393_, _06375_);
  and _73822_ (_23411_, _23410_, _23408_);
  or _73823_ (_23412_, _23411_, _23407_);
  and _73824_ (_23413_, _23412_, _07234_);
  and _73825_ (_23414_, _23342_, _06545_);
  and _73826_ (_23415_, _23414_, _23408_);
  or _73827_ (_23416_, _23415_, _06366_);
  or _73828_ (_23417_, _23416_, _23413_);
  and _73829_ (_23418_, _14748_, _07928_);
  or _73830_ (_23419_, _23333_, _09056_);
  or _73831_ (_23421_, _23419_, _23418_);
  and _73832_ (_23422_, _23421_, _09061_);
  and _73833_ (_23423_, _23422_, _23417_);
  nor _73834_ (_23424_, _11258_, _11882_);
  or _73835_ (_23425_, _23424_, _23333_);
  and _73836_ (_23426_, _23425_, _06528_);
  or _73837_ (_23427_, _23426_, _06568_);
  or _73838_ (_23428_, _23427_, _23423_);
  or _73839_ (_23429_, _23339_, _06926_);
  and _73840_ (_23430_, _23429_, _05928_);
  and _73841_ (_23432_, _23430_, _23428_);
  and _73842_ (_23433_, _23363_, _05927_);
  or _73843_ (_23434_, _23433_, _06278_);
  or _73844_ (_23435_, _23434_, _23432_);
  and _73845_ (_23436_, _14926_, _07928_);
  or _73846_ (_23437_, _23333_, _06279_);
  or _73847_ (_23438_, _23437_, _23436_);
  and _73848_ (_23439_, _23438_, _01347_);
  and _73849_ (_23440_, _23439_, _23435_);
  or _73850_ (_23441_, _23440_, _23331_);
  and _73851_ (_43221_, _23441_, _42618_);
  and _73852_ (_23443_, _01351_, \oc8051_golden_model_1.TCON [3]);
  and _73853_ (_23444_, _11882_, \oc8051_golden_model_1.TCON [3]);
  nor _73854_ (_23445_, _11882_, _07594_);
  or _73855_ (_23446_, _23445_, _23444_);
  or _73856_ (_23447_, _23446_, _07215_);
  and _73857_ (_23448_, _14953_, _07928_);
  or _73858_ (_23449_, _23448_, _23444_);
  or _73859_ (_23450_, _23449_, _07151_);
  and _73860_ (_23451_, _07928_, \oc8051_golden_model_1.ACC [3]);
  or _73861_ (_23453_, _23451_, _23444_);
  and _73862_ (_23454_, _23453_, _07141_);
  and _73863_ (_23455_, _07142_, \oc8051_golden_model_1.TCON [3]);
  or _73864_ (_23456_, _23455_, _06341_);
  or _73865_ (_23457_, _23456_, _23454_);
  and _73866_ (_23458_, _23457_, _06273_);
  and _73867_ (_23459_, _23458_, _23450_);
  and _73868_ (_23460_, _11890_, \oc8051_golden_model_1.TCON [3]);
  and _73869_ (_23461_, _14950_, _08616_);
  or _73870_ (_23462_, _23461_, _23460_);
  and _73871_ (_23464_, _23462_, _06272_);
  or _73872_ (_23465_, _23464_, _06461_);
  or _73873_ (_23466_, _23465_, _23459_);
  or _73874_ (_23467_, _23446_, _07166_);
  and _73875_ (_23468_, _23467_, _23466_);
  or _73876_ (_23469_, _23468_, _06464_);
  or _73877_ (_23470_, _23453_, _06465_);
  and _73878_ (_23471_, _23470_, _06269_);
  and _73879_ (_23472_, _23471_, _23469_);
  and _73880_ (_23473_, _14948_, _08616_);
  or _73881_ (_23475_, _23473_, _23460_);
  and _73882_ (_23476_, _23475_, _06268_);
  or _73883_ (_23477_, _23476_, _06261_);
  or _73884_ (_23478_, _23477_, _23472_);
  or _73885_ (_23479_, _23460_, _14979_);
  and _73886_ (_23480_, _23479_, _23462_);
  or _73887_ (_23481_, _23480_, _06262_);
  and _73888_ (_23482_, _23481_, _06258_);
  and _73889_ (_23483_, _23482_, _23478_);
  or _73890_ (_23484_, _23460_, _14992_);
  and _73891_ (_23486_, _23484_, _06257_);
  and _73892_ (_23487_, _23486_, _23462_);
  or _73893_ (_23488_, _23487_, _10080_);
  or _73894_ (_23489_, _23488_, _23483_);
  and _73895_ (_23490_, _23489_, _23447_);
  or _73896_ (_23491_, _23490_, _07460_);
  and _73897_ (_23492_, _09449_, _07928_);
  or _73898_ (_23493_, _23444_, _07208_);
  or _73899_ (_23494_, _23493_, _23492_);
  and _73900_ (_23495_, _23494_, _05982_);
  and _73901_ (_23497_, _23495_, _23491_);
  and _73902_ (_23498_, _15048_, _07928_);
  or _73903_ (_23499_, _23498_, _23444_);
  and _73904_ (_23500_, _23499_, _10094_);
  or _73905_ (_23501_, _23500_, _06218_);
  or _73906_ (_23502_, _23501_, _23497_);
  and _73907_ (_23503_, _07928_, _08930_);
  or _73908_ (_23504_, _23503_, _23444_);
  or _73909_ (_23505_, _23504_, _06219_);
  and _73910_ (_23506_, _23505_, _23502_);
  or _73911_ (_23508_, _23506_, _06369_);
  and _73912_ (_23509_, _14943_, _07928_);
  or _73913_ (_23510_, _23509_, _23444_);
  or _73914_ (_23511_, _23510_, _07237_);
  and _73915_ (_23512_, _23511_, _07240_);
  and _73916_ (_23513_, _23512_, _23508_);
  and _73917_ (_23514_, _12577_, _07928_);
  or _73918_ (_23515_, _23514_, _23444_);
  and _73919_ (_23516_, _23515_, _06536_);
  or _73920_ (_23517_, _23516_, _23513_);
  and _73921_ (_23519_, _23517_, _07242_);
  or _73922_ (_23520_, _23444_, _08292_);
  and _73923_ (_23521_, _23504_, _06375_);
  and _73924_ (_23522_, _23521_, _23520_);
  or _73925_ (_23523_, _23522_, _23519_);
  and _73926_ (_23524_, _23523_, _07234_);
  and _73927_ (_23525_, _23453_, _06545_);
  and _73928_ (_23526_, _23525_, _23520_);
  or _73929_ (_23527_, _23526_, _06366_);
  or _73930_ (_23528_, _23527_, _23524_);
  and _73931_ (_23530_, _14940_, _07928_);
  or _73932_ (_23531_, _23444_, _09056_);
  or _73933_ (_23532_, _23531_, _23530_);
  and _73934_ (_23533_, _23532_, _09061_);
  and _73935_ (_23534_, _23533_, _23528_);
  nor _73936_ (_23535_, _11256_, _11882_);
  or _73937_ (_23536_, _23535_, _23444_);
  and _73938_ (_23537_, _23536_, _06528_);
  or _73939_ (_23538_, _23537_, _06568_);
  or _73940_ (_23539_, _23538_, _23534_);
  or _73941_ (_23541_, _23449_, _06926_);
  and _73942_ (_23542_, _23541_, _05928_);
  and _73943_ (_23543_, _23542_, _23539_);
  and _73944_ (_23544_, _23475_, _05927_);
  or _73945_ (_23545_, _23544_, _06278_);
  or _73946_ (_23546_, _23545_, _23543_);
  and _73947_ (_23547_, _15128_, _07928_);
  or _73948_ (_23548_, _23444_, _06279_);
  or _73949_ (_23549_, _23548_, _23547_);
  and _73950_ (_23550_, _23549_, _01347_);
  and _73951_ (_23552_, _23550_, _23546_);
  or _73952_ (_23553_, _23552_, _23443_);
  and _73953_ (_43223_, _23553_, _42618_);
  and _73954_ (_23554_, _01351_, \oc8051_golden_model_1.TCON [4]);
  and _73955_ (_23555_, _11882_, \oc8051_golden_model_1.TCON [4]);
  nor _73956_ (_23556_, _08541_, _11882_);
  or _73957_ (_23557_, _23556_, _23555_);
  or _73958_ (_23558_, _23557_, _07215_);
  and _73959_ (_23559_, _11890_, \oc8051_golden_model_1.TCON [4]);
  and _73960_ (_23560_, _15176_, _08616_);
  or _73961_ (_23562_, _23560_, _23559_);
  and _73962_ (_23563_, _23562_, _06268_);
  and _73963_ (_23564_, _15162_, _07928_);
  or _73964_ (_23565_, _23564_, _23555_);
  or _73965_ (_23566_, _23565_, _07151_);
  and _73966_ (_23567_, _07928_, \oc8051_golden_model_1.ACC [4]);
  or _73967_ (_23568_, _23567_, _23555_);
  and _73968_ (_23569_, _23568_, _07141_);
  and _73969_ (_23570_, _07142_, \oc8051_golden_model_1.TCON [4]);
  or _73970_ (_23571_, _23570_, _06341_);
  or _73971_ (_23573_, _23571_, _23569_);
  and _73972_ (_23574_, _23573_, _06273_);
  and _73973_ (_23575_, _23574_, _23566_);
  and _73974_ (_23576_, _15166_, _08616_);
  or _73975_ (_23577_, _23576_, _23559_);
  and _73976_ (_23578_, _23577_, _06272_);
  or _73977_ (_23579_, _23578_, _06461_);
  or _73978_ (_23580_, _23579_, _23575_);
  or _73979_ (_23581_, _23557_, _07166_);
  and _73980_ (_23582_, _23581_, _23580_);
  or _73981_ (_23584_, _23582_, _06464_);
  or _73982_ (_23585_, _23568_, _06465_);
  and _73983_ (_23586_, _23585_, _06269_);
  and _73984_ (_23587_, _23586_, _23584_);
  or _73985_ (_23588_, _23587_, _23563_);
  and _73986_ (_23589_, _23588_, _06262_);
  or _73987_ (_23590_, _23559_, _15183_);
  and _73988_ (_23591_, _23590_, _06261_);
  and _73989_ (_23592_, _23591_, _23577_);
  or _73990_ (_23593_, _23592_, _23589_);
  and _73991_ (_23595_, _23593_, _06258_);
  and _73992_ (_23596_, _15200_, _08616_);
  or _73993_ (_23597_, _23596_, _23559_);
  and _73994_ (_23598_, _23597_, _06257_);
  or _73995_ (_23599_, _23598_, _10080_);
  or _73996_ (_23600_, _23599_, _23595_);
  and _73997_ (_23601_, _23600_, _23558_);
  or _73998_ (_23602_, _23601_, _07460_);
  and _73999_ (_23603_, _09448_, _07928_);
  or _74000_ (_23604_, _23555_, _07208_);
  or _74001_ (_23605_, _23604_, _23603_);
  and _74002_ (_23606_, _23605_, _05982_);
  and _74003_ (_23607_, _23606_, _23602_);
  and _74004_ (_23608_, _15254_, _07928_);
  or _74005_ (_23609_, _23608_, _23555_);
  and _74006_ (_23610_, _23609_, _10094_);
  or _74007_ (_23611_, _23610_, _06218_);
  or _74008_ (_23612_, _23611_, _23607_);
  and _74009_ (_23613_, _08959_, _07928_);
  or _74010_ (_23614_, _23613_, _23555_);
  or _74011_ (_23616_, _23614_, _06219_);
  and _74012_ (_23617_, _23616_, _23612_);
  or _74013_ (_23618_, _23617_, _06369_);
  and _74014_ (_23619_, _15269_, _07928_);
  or _74015_ (_23620_, _23619_, _23555_);
  or _74016_ (_23621_, _23620_, _07237_);
  and _74017_ (_23622_, _23621_, _07240_);
  and _74018_ (_23623_, _23622_, _23618_);
  and _74019_ (_23624_, _11254_, _07928_);
  or _74020_ (_23625_, _23624_, _23555_);
  and _74021_ (_23627_, _23625_, _06536_);
  or _74022_ (_23628_, _23627_, _23623_);
  and _74023_ (_23629_, _23628_, _07242_);
  or _74024_ (_23630_, _23555_, _08544_);
  and _74025_ (_23631_, _23614_, _06375_);
  and _74026_ (_23632_, _23631_, _23630_);
  or _74027_ (_23633_, _23632_, _23629_);
  and _74028_ (_23634_, _23633_, _07234_);
  and _74029_ (_23635_, _23568_, _06545_);
  and _74030_ (_23636_, _23635_, _23630_);
  or _74031_ (_23638_, _23636_, _06366_);
  or _74032_ (_23639_, _23638_, _23634_);
  and _74033_ (_23640_, _15266_, _07928_);
  or _74034_ (_23641_, _23555_, _09056_);
  or _74035_ (_23642_, _23641_, _23640_);
  and _74036_ (_23643_, _23642_, _09061_);
  and _74037_ (_23644_, _23643_, _23639_);
  nor _74038_ (_23645_, _11253_, _11882_);
  or _74039_ (_23646_, _23645_, _23555_);
  and _74040_ (_23647_, _23646_, _06528_);
  or _74041_ (_23648_, _23647_, _06568_);
  or _74042_ (_23649_, _23648_, _23644_);
  or _74043_ (_23650_, _23565_, _06926_);
  and _74044_ (_23651_, _23650_, _05928_);
  and _74045_ (_23652_, _23651_, _23649_);
  and _74046_ (_23653_, _23562_, _05927_);
  or _74047_ (_23654_, _23653_, _06278_);
  or _74048_ (_23655_, _23654_, _23652_);
  and _74049_ (_23656_, _15329_, _07928_);
  or _74050_ (_23657_, _23555_, _06279_);
  or _74051_ (_23659_, _23657_, _23656_);
  and _74052_ (_23660_, _23659_, _01347_);
  and _74053_ (_23661_, _23660_, _23655_);
  or _74054_ (_23662_, _23661_, _23554_);
  and _74055_ (_43224_, _23662_, _42618_);
  and _74056_ (_23663_, _01351_, \oc8051_golden_model_1.TCON [5]);
  and _74057_ (_23664_, _11882_, \oc8051_golden_model_1.TCON [5]);
  and _74058_ (_23665_, _15358_, _07928_);
  or _74059_ (_23666_, _23665_, _23664_);
  or _74060_ (_23667_, _23666_, _07151_);
  and _74061_ (_23668_, _07928_, \oc8051_golden_model_1.ACC [5]);
  or _74062_ (_23669_, _23668_, _23664_);
  and _74063_ (_23670_, _23669_, _07141_);
  and _74064_ (_23671_, _07142_, \oc8051_golden_model_1.TCON [5]);
  or _74065_ (_23672_, _23671_, _06341_);
  or _74066_ (_23673_, _23672_, _23670_);
  and _74067_ (_23674_, _23673_, _06273_);
  and _74068_ (_23675_, _23674_, _23667_);
  and _74069_ (_23676_, _11890_, \oc8051_golden_model_1.TCON [5]);
  and _74070_ (_23677_, _15372_, _08616_);
  or _74071_ (_23679_, _23677_, _23676_);
  and _74072_ (_23680_, _23679_, _06272_);
  or _74073_ (_23681_, _23680_, _06461_);
  or _74074_ (_23682_, _23681_, _23675_);
  nor _74075_ (_23683_, _08244_, _11882_);
  or _74076_ (_23684_, _23683_, _23664_);
  or _74077_ (_23685_, _23684_, _07166_);
  and _74078_ (_23686_, _23685_, _23682_);
  or _74079_ (_23687_, _23686_, _06464_);
  or _74080_ (_23688_, _23669_, _06465_);
  and _74081_ (_23690_, _23688_, _06269_);
  and _74082_ (_23691_, _23690_, _23687_);
  and _74083_ (_23692_, _15355_, _08616_);
  or _74084_ (_23693_, _23692_, _23676_);
  and _74085_ (_23694_, _23693_, _06268_);
  or _74086_ (_23695_, _23694_, _06261_);
  or _74087_ (_23696_, _23695_, _23691_);
  or _74088_ (_23697_, _23676_, _15387_);
  and _74089_ (_23698_, _23697_, _23679_);
  or _74090_ (_23699_, _23698_, _06262_);
  and _74091_ (_23700_, _23699_, _06258_);
  and _74092_ (_23701_, _23700_, _23696_);
  or _74093_ (_23702_, _23676_, _15403_);
  and _74094_ (_23703_, _23702_, _06257_);
  and _74095_ (_23704_, _23703_, _23679_);
  or _74096_ (_23705_, _23704_, _10080_);
  or _74097_ (_23706_, _23705_, _23701_);
  or _74098_ (_23707_, _23684_, _07215_);
  and _74099_ (_23708_, _23707_, _23706_);
  or _74100_ (_23709_, _23708_, _07460_);
  and _74101_ (_23711_, _09447_, _07928_);
  or _74102_ (_23712_, _23664_, _07208_);
  or _74103_ (_23713_, _23712_, _23711_);
  and _74104_ (_23714_, _23713_, _05982_);
  and _74105_ (_23715_, _23714_, _23709_);
  and _74106_ (_23716_, _15459_, _07928_);
  or _74107_ (_23717_, _23716_, _23664_);
  and _74108_ (_23718_, _23717_, _10094_);
  or _74109_ (_23719_, _23718_, _06218_);
  or _74110_ (_23720_, _23719_, _23715_);
  and _74111_ (_23722_, _08946_, _07928_);
  or _74112_ (_23723_, _23722_, _23664_);
  or _74113_ (_23724_, _23723_, _06219_);
  and _74114_ (_23725_, _23724_, _23720_);
  or _74115_ (_23726_, _23725_, _06369_);
  and _74116_ (_23727_, _15353_, _07928_);
  or _74117_ (_23728_, _23727_, _23664_);
  or _74118_ (_23729_, _23728_, _07237_);
  and _74119_ (_23730_, _23729_, _07240_);
  and _74120_ (_23731_, _23730_, _23726_);
  and _74121_ (_23732_, _11250_, _07928_);
  or _74122_ (_23733_, _23732_, _23664_);
  and _74123_ (_23734_, _23733_, _06536_);
  or _74124_ (_23735_, _23734_, _23731_);
  and _74125_ (_23736_, _23735_, _07242_);
  or _74126_ (_23737_, _23664_, _08247_);
  and _74127_ (_23738_, _23723_, _06375_);
  and _74128_ (_23739_, _23738_, _23737_);
  or _74129_ (_23740_, _23739_, _23736_);
  and _74130_ (_23741_, _23740_, _07234_);
  and _74131_ (_23743_, _23669_, _06545_);
  and _74132_ (_23744_, _23743_, _23737_);
  or _74133_ (_23745_, _23744_, _06366_);
  or _74134_ (_23746_, _23745_, _23741_);
  and _74135_ (_23747_, _15350_, _07928_);
  or _74136_ (_23748_, _23664_, _09056_);
  or _74137_ (_23749_, _23748_, _23747_);
  and _74138_ (_23750_, _23749_, _09061_);
  and _74139_ (_23751_, _23750_, _23746_);
  nor _74140_ (_23752_, _11249_, _11882_);
  or _74141_ (_23754_, _23752_, _23664_);
  and _74142_ (_23755_, _23754_, _06528_);
  or _74143_ (_23756_, _23755_, _06568_);
  or _74144_ (_23757_, _23756_, _23751_);
  or _74145_ (_23758_, _23666_, _06926_);
  and _74146_ (_23759_, _23758_, _05928_);
  and _74147_ (_23760_, _23759_, _23757_);
  and _74148_ (_23761_, _23693_, _05927_);
  or _74149_ (_23762_, _23761_, _06278_);
  or _74150_ (_23763_, _23762_, _23760_);
  and _74151_ (_23764_, _15532_, _07928_);
  or _74152_ (_23765_, _23664_, _06279_);
  or _74153_ (_23766_, _23765_, _23764_);
  and _74154_ (_23767_, _23766_, _01347_);
  and _74155_ (_23768_, _23767_, _23763_);
  or _74156_ (_23769_, _23768_, _23663_);
  and _74157_ (_43225_, _23769_, _42618_);
  and _74158_ (_23770_, _01351_, \oc8051_golden_model_1.TCON [6]);
  and _74159_ (_23771_, _11882_, \oc8051_golden_model_1.TCON [6]);
  and _74160_ (_23772_, _15554_, _07928_);
  or _74161_ (_23774_, _23772_, _23771_);
  or _74162_ (_23775_, _23774_, _07151_);
  and _74163_ (_23776_, _07928_, \oc8051_golden_model_1.ACC [6]);
  or _74164_ (_23777_, _23776_, _23771_);
  and _74165_ (_23778_, _23777_, _07141_);
  and _74166_ (_23779_, _07142_, \oc8051_golden_model_1.TCON [6]);
  or _74167_ (_23780_, _23779_, _06341_);
  or _74168_ (_23781_, _23780_, _23778_);
  and _74169_ (_23782_, _23781_, _06273_);
  and _74170_ (_23783_, _23782_, _23775_);
  and _74171_ (_23785_, _11890_, \oc8051_golden_model_1.TCON [6]);
  and _74172_ (_23786_, _15570_, _08616_);
  or _74173_ (_23787_, _23786_, _23785_);
  and _74174_ (_23788_, _23787_, _06272_);
  or _74175_ (_23789_, _23788_, _06461_);
  or _74176_ (_23790_, _23789_, _23783_);
  nor _74177_ (_23791_, _08142_, _11882_);
  or _74178_ (_23792_, _23791_, _23771_);
  or _74179_ (_23793_, _23792_, _07166_);
  and _74180_ (_23794_, _23793_, _23790_);
  or _74181_ (_23795_, _23794_, _06464_);
  or _74182_ (_23796_, _23777_, _06465_);
  and _74183_ (_23797_, _23796_, _06269_);
  and _74184_ (_23798_, _23797_, _23795_);
  and _74185_ (_23799_, _15551_, _08616_);
  or _74186_ (_23800_, _23799_, _23785_);
  and _74187_ (_23801_, _23800_, _06268_);
  or _74188_ (_23802_, _23801_, _06261_);
  or _74189_ (_23803_, _23802_, _23798_);
  or _74190_ (_23804_, _23785_, _15585_);
  and _74191_ (_23805_, _23804_, _23787_);
  or _74192_ (_23806_, _23805_, _06262_);
  and _74193_ (_23807_, _23806_, _06258_);
  and _74194_ (_23808_, _23807_, _23803_);
  and _74195_ (_23809_, _15602_, _08616_);
  or _74196_ (_23810_, _23809_, _23785_);
  and _74197_ (_23811_, _23810_, _06257_);
  or _74198_ (_23812_, _23811_, _10080_);
  or _74199_ (_23813_, _23812_, _23808_);
  or _74200_ (_23814_, _23792_, _07215_);
  and _74201_ (_23817_, _23814_, _23813_);
  or _74202_ (_23818_, _23817_, _07460_);
  and _74203_ (_23819_, _09446_, _07928_);
  or _74204_ (_23820_, _23771_, _07208_);
  or _74205_ (_23821_, _23820_, _23819_);
  and _74206_ (_23822_, _23821_, _05982_);
  and _74207_ (_23823_, _23822_, _23818_);
  and _74208_ (_23824_, _15657_, _07928_);
  or _74209_ (_23825_, _23824_, _23771_);
  and _74210_ (_23826_, _23825_, _10094_);
  or _74211_ (_23827_, _23826_, _06218_);
  or _74212_ (_23828_, _23827_, _23823_);
  and _74213_ (_23829_, _15664_, _07928_);
  or _74214_ (_23830_, _23829_, _23771_);
  or _74215_ (_23831_, _23830_, _06219_);
  and _74216_ (_23832_, _23831_, _23828_);
  or _74217_ (_23833_, _23832_, _06369_);
  and _74218_ (_23834_, _15549_, _07928_);
  or _74219_ (_23835_, _23834_, _23771_);
  or _74220_ (_23836_, _23835_, _07237_);
  and _74221_ (_23838_, _23836_, _07240_);
  and _74222_ (_23839_, _23838_, _23833_);
  and _74223_ (_23840_, _11247_, _07928_);
  or _74224_ (_23841_, _23840_, _23771_);
  and _74225_ (_23842_, _23841_, _06536_);
  or _74226_ (_23843_, _23842_, _23839_);
  and _74227_ (_23844_, _23843_, _07242_);
  or _74228_ (_23845_, _23771_, _08145_);
  and _74229_ (_23846_, _23830_, _06375_);
  and _74230_ (_23847_, _23846_, _23845_);
  or _74231_ (_23849_, _23847_, _23844_);
  and _74232_ (_23850_, _23849_, _07234_);
  and _74233_ (_23851_, _23777_, _06545_);
  and _74234_ (_23852_, _23851_, _23845_);
  or _74235_ (_23853_, _23852_, _06366_);
  or _74236_ (_23854_, _23853_, _23850_);
  and _74237_ (_23855_, _15546_, _07928_);
  or _74238_ (_23856_, _23771_, _09056_);
  or _74239_ (_23857_, _23856_, _23855_);
  and _74240_ (_23858_, _23857_, _09061_);
  and _74241_ (_23859_, _23858_, _23854_);
  nor _74242_ (_23860_, _11246_, _11882_);
  or _74243_ (_23861_, _23860_, _23771_);
  and _74244_ (_23862_, _23861_, _06528_);
  or _74245_ (_23863_, _23862_, _06568_);
  or _74246_ (_23864_, _23863_, _23859_);
  or _74247_ (_23865_, _23774_, _06926_);
  and _74248_ (_23866_, _23865_, _05928_);
  and _74249_ (_23867_, _23866_, _23864_);
  and _74250_ (_23868_, _23800_, _05927_);
  or _74251_ (_23870_, _23868_, _06278_);
  or _74252_ (_23871_, _23870_, _23867_);
  and _74253_ (_23872_, _15734_, _07928_);
  or _74254_ (_23873_, _23771_, _06279_);
  or _74255_ (_23874_, _23873_, _23872_);
  and _74256_ (_23875_, _23874_, _01347_);
  and _74257_ (_23876_, _23875_, _23871_);
  or _74258_ (_23877_, _23876_, _23770_);
  and _74259_ (_43226_, _23877_, _42618_);
  and _74260_ (_23878_, _01351_, \oc8051_golden_model_1.TH1 [0]);
  and _74261_ (_23880_, _07910_, \oc8051_golden_model_1.ACC [0]);
  and _74262_ (_23881_, _23880_, _08390_);
  and _74263_ (_23882_, _11985_, \oc8051_golden_model_1.TH1 [0]);
  or _74264_ (_23883_, _23882_, _07234_);
  or _74265_ (_23884_, _23883_, _23881_);
  and _74266_ (_23885_, _07910_, _07133_);
  or _74267_ (_23886_, _23885_, _23882_);
  or _74268_ (_23887_, _23886_, _07215_);
  nor _74269_ (_23888_, _08390_, _11985_);
  or _74270_ (_23889_, _23888_, _23882_);
  or _74271_ (_23890_, _23889_, _07151_);
  or _74272_ (_23891_, _23882_, _23880_);
  and _74273_ (_23892_, _23891_, _07141_);
  and _74274_ (_23893_, _07142_, \oc8051_golden_model_1.TH1 [0]);
  or _74275_ (_23894_, _23893_, _06341_);
  or _74276_ (_23895_, _23894_, _23892_);
  and _74277_ (_23896_, _23895_, _07166_);
  and _74278_ (_23897_, _23896_, _23890_);
  and _74279_ (_23898_, _23886_, _06461_);
  or _74280_ (_23899_, _23898_, _23897_);
  and _74281_ (_23901_, _23899_, _06465_);
  and _74282_ (_23902_, _23891_, _06464_);
  or _74283_ (_23903_, _23902_, _10080_);
  or _74284_ (_23904_, _23903_, _23901_);
  and _74285_ (_23905_, _23904_, _23887_);
  or _74286_ (_23906_, _23905_, _07460_);
  and _74287_ (_23907_, _09392_, _07910_);
  or _74288_ (_23908_, _23882_, _07208_);
  or _74289_ (_23909_, _23908_, _23907_);
  and _74290_ (_23910_, _23909_, _23906_);
  or _74291_ (_23912_, _23910_, _10094_);
  and _74292_ (_23913_, _14467_, _07910_);
  or _74293_ (_23914_, _23882_, _05982_);
  or _74294_ (_23915_, _23914_, _23913_);
  and _74295_ (_23916_, _23915_, _06219_);
  and _74296_ (_23917_, _23916_, _23912_);
  and _74297_ (_23918_, _07910_, _08954_);
  or _74298_ (_23919_, _23918_, _23882_);
  and _74299_ (_23920_, _23919_, _06218_);
  or _74300_ (_23921_, _23920_, _06369_);
  or _74301_ (_23922_, _23921_, _23917_);
  and _74302_ (_23923_, _14366_, _07910_);
  or _74303_ (_23924_, _23923_, _23882_);
  or _74304_ (_23925_, _23924_, _07237_);
  and _74305_ (_23926_, _23925_, _07240_);
  and _74306_ (_23927_, _23926_, _23922_);
  nor _74307_ (_23928_, _12580_, _11985_);
  or _74308_ (_23929_, _23928_, _23882_);
  nor _74309_ (_23930_, _23881_, _07240_);
  and _74310_ (_23931_, _23930_, _23929_);
  or _74311_ (_23933_, _23931_, _23927_);
  and _74312_ (_23934_, _23933_, _07242_);
  nand _74313_ (_23935_, _23919_, _06375_);
  nor _74314_ (_23936_, _23935_, _23888_);
  or _74315_ (_23937_, _23936_, _06545_);
  or _74316_ (_23938_, _23937_, _23934_);
  and _74317_ (_23939_, _23938_, _23884_);
  or _74318_ (_23940_, _23939_, _06366_);
  and _74319_ (_23941_, _14363_, _07910_);
  or _74320_ (_23942_, _23882_, _09056_);
  or _74321_ (_23944_, _23942_, _23941_);
  and _74322_ (_23945_, _23944_, _09061_);
  and _74323_ (_23946_, _23945_, _23940_);
  and _74324_ (_23947_, _23929_, _06528_);
  or _74325_ (_23948_, _23947_, _19502_);
  or _74326_ (_23949_, _23948_, _23946_);
  or _74327_ (_23950_, _23889_, _06661_);
  and _74328_ (_23951_, _23950_, _01347_);
  and _74329_ (_23952_, _23951_, _23949_);
  or _74330_ (_23953_, _23952_, _23878_);
  and _74331_ (_43228_, _23953_, _42618_);
  and _74332_ (_23954_, _01351_, \oc8051_golden_model_1.TH1 [1]);
  nand _74333_ (_23955_, _07910_, _07038_);
  or _74334_ (_23956_, _07910_, \oc8051_golden_model_1.TH1 [1]);
  and _74335_ (_23957_, _23956_, _06218_);
  and _74336_ (_23958_, _23957_, _23955_);
  and _74337_ (_23959_, _11985_, \oc8051_golden_model_1.TH1 [1]);
  nor _74338_ (_23960_, _11985_, _07357_);
  or _74339_ (_23961_, _23960_, _23959_);
  or _74340_ (_23962_, _23961_, _07215_);
  and _74341_ (_23964_, _14562_, _07910_);
  not _74342_ (_23965_, _23964_);
  and _74343_ (_23966_, _23965_, _23956_);
  or _74344_ (_23967_, _23966_, _07151_);
  and _74345_ (_23968_, _07910_, \oc8051_golden_model_1.ACC [1]);
  or _74346_ (_23969_, _23968_, _23959_);
  and _74347_ (_23970_, _23969_, _07141_);
  and _74348_ (_23971_, _07142_, \oc8051_golden_model_1.TH1 [1]);
  or _74349_ (_23972_, _23971_, _06341_);
  or _74350_ (_23973_, _23972_, _23970_);
  and _74351_ (_23975_, _23973_, _07166_);
  and _74352_ (_23976_, _23975_, _23967_);
  and _74353_ (_23977_, _23961_, _06461_);
  or _74354_ (_23978_, _23977_, _23976_);
  and _74355_ (_23979_, _23978_, _06465_);
  and _74356_ (_23980_, _23969_, _06464_);
  or _74357_ (_23981_, _23980_, _10080_);
  or _74358_ (_23982_, _23981_, _23979_);
  and _74359_ (_23983_, _23982_, _23962_);
  or _74360_ (_23984_, _23983_, _07460_);
  and _74361_ (_23985_, _09451_, _07910_);
  or _74362_ (_23986_, _23959_, _07208_);
  or _74363_ (_23987_, _23986_, _23985_);
  and _74364_ (_23988_, _23987_, _05982_);
  and _74365_ (_23989_, _23988_, _23984_);
  or _74366_ (_23990_, _14653_, _11985_);
  and _74367_ (_23991_, _23956_, _10094_);
  and _74368_ (_23992_, _23991_, _23990_);
  or _74369_ (_23993_, _23992_, _23989_);
  and _74370_ (_23994_, _23993_, _06219_);
  or _74371_ (_23996_, _23994_, _23958_);
  and _74372_ (_23997_, _23996_, _07237_);
  or _74373_ (_23998_, _14668_, _11985_);
  and _74374_ (_23999_, _23956_, _06369_);
  and _74375_ (_24000_, _23999_, _23998_);
  or _74376_ (_24001_, _24000_, _06536_);
  or _74377_ (_24002_, _24001_, _23997_);
  and _74378_ (_24003_, _11262_, _07910_);
  or _74379_ (_24004_, _24003_, _23959_);
  or _74380_ (_24005_, _24004_, _07240_);
  and _74381_ (_24007_, _24005_, _07242_);
  and _74382_ (_24008_, _24007_, _24002_);
  or _74383_ (_24009_, _14666_, _11985_);
  and _74384_ (_24010_, _23956_, _06375_);
  and _74385_ (_24011_, _24010_, _24009_);
  or _74386_ (_24012_, _24011_, _06545_);
  or _74387_ (_24013_, _24012_, _24008_);
  and _74388_ (_24014_, _23968_, _08341_);
  or _74389_ (_24015_, _23959_, _07234_);
  or _74390_ (_24016_, _24015_, _24014_);
  and _74391_ (_24018_, _24016_, _09056_);
  and _74392_ (_24019_, _24018_, _24013_);
  or _74393_ (_24020_, _23955_, _08341_);
  and _74394_ (_24021_, _23956_, _06366_);
  and _74395_ (_24022_, _24021_, _24020_);
  or _74396_ (_24023_, _24022_, _06528_);
  or _74397_ (_24024_, _24023_, _24019_);
  nor _74398_ (_24025_, _11261_, _11985_);
  or _74399_ (_24026_, _24025_, _23959_);
  or _74400_ (_24027_, _24026_, _09061_);
  and _74401_ (_24028_, _24027_, _06926_);
  and _74402_ (_24029_, _24028_, _24024_);
  and _74403_ (_24030_, _23966_, _06568_);
  or _74404_ (_24031_, _24030_, _06278_);
  or _74405_ (_24032_, _24031_, _24029_);
  or _74406_ (_24033_, _23959_, _06279_);
  or _74407_ (_24034_, _24033_, _23964_);
  and _74408_ (_24035_, _24034_, _01347_);
  and _74409_ (_24036_, _24035_, _24032_);
  or _74410_ (_24037_, _24036_, _23954_);
  and _74411_ (_43229_, _24037_, _42618_);
  and _74412_ (_24039_, _01351_, \oc8051_golden_model_1.TH1 [2]);
  and _74413_ (_24040_, _11985_, \oc8051_golden_model_1.TH1 [2]);
  and _74414_ (_24041_, _09450_, _07910_);
  or _74415_ (_24042_, _24041_, _24040_);
  and _74416_ (_24043_, _24042_, _07460_);
  and _74417_ (_24044_, _14770_, _07910_);
  or _74418_ (_24045_, _24044_, _24040_);
  or _74419_ (_24046_, _24045_, _07151_);
  and _74420_ (_24047_, _07910_, \oc8051_golden_model_1.ACC [2]);
  or _74421_ (_24049_, _24047_, _24040_);
  and _74422_ (_24050_, _24049_, _07141_);
  and _74423_ (_24051_, _07142_, \oc8051_golden_model_1.TH1 [2]);
  or _74424_ (_24052_, _24051_, _06341_);
  or _74425_ (_24053_, _24052_, _24050_);
  and _74426_ (_24054_, _24053_, _07166_);
  and _74427_ (_24055_, _24054_, _24046_);
  nor _74428_ (_24056_, _11985_, _07776_);
  or _74429_ (_24057_, _24056_, _24040_);
  and _74430_ (_24058_, _24057_, _06461_);
  or _74431_ (_24059_, _24058_, _24055_);
  and _74432_ (_24060_, _24059_, _06465_);
  and _74433_ (_24061_, _24049_, _06464_);
  or _74434_ (_24062_, _24061_, _10080_);
  or _74435_ (_24063_, _24062_, _24060_);
  or _74436_ (_24064_, _24057_, _07215_);
  and _74437_ (_24065_, _24064_, _07208_);
  and _74438_ (_24066_, _24065_, _24063_);
  or _74439_ (_24067_, _24066_, _10094_);
  or _74440_ (_24068_, _24067_, _24043_);
  and _74441_ (_24070_, _14859_, _07910_);
  or _74442_ (_24071_, _24040_, _05982_);
  or _74443_ (_24072_, _24071_, _24070_);
  and _74444_ (_24073_, _24072_, _06219_);
  and _74445_ (_24074_, _24073_, _24068_);
  and _74446_ (_24075_, _07910_, _08973_);
  or _74447_ (_24076_, _24075_, _24040_);
  and _74448_ (_24077_, _24076_, _06218_);
  or _74449_ (_24078_, _24077_, _06369_);
  or _74450_ (_24079_, _24078_, _24074_);
  and _74451_ (_24081_, _14751_, _07910_);
  or _74452_ (_24082_, _24081_, _24040_);
  or _74453_ (_24083_, _24082_, _07237_);
  and _74454_ (_24084_, _24083_, _07240_);
  and _74455_ (_24085_, _24084_, _24079_);
  and _74456_ (_24086_, _11259_, _07910_);
  or _74457_ (_24087_, _24086_, _24040_);
  and _74458_ (_24088_, _24087_, _06536_);
  or _74459_ (_24089_, _24088_, _24085_);
  and _74460_ (_24090_, _24089_, _07242_);
  or _74461_ (_24092_, _24040_, _08440_);
  and _74462_ (_24093_, _24076_, _06375_);
  and _74463_ (_24094_, _24093_, _24092_);
  or _74464_ (_24095_, _24094_, _24090_);
  and _74465_ (_24096_, _24095_, _07234_);
  and _74466_ (_24097_, _24049_, _06545_);
  and _74467_ (_24098_, _24097_, _24092_);
  or _74468_ (_24099_, _24098_, _06366_);
  or _74469_ (_24100_, _24099_, _24096_);
  and _74470_ (_24101_, _14748_, _07910_);
  or _74471_ (_24102_, _24040_, _09056_);
  or _74472_ (_24103_, _24102_, _24101_);
  and _74473_ (_24104_, _24103_, _09061_);
  and _74474_ (_24105_, _24104_, _24100_);
  nor _74475_ (_24106_, _11258_, _11985_);
  or _74476_ (_24107_, _24106_, _24040_);
  and _74477_ (_24108_, _24107_, _06528_);
  or _74478_ (_24109_, _24108_, _24105_);
  and _74479_ (_24110_, _24109_, _06926_);
  and _74480_ (_24111_, _24045_, _06568_);
  or _74481_ (_24113_, _24111_, _06278_);
  or _74482_ (_24114_, _24113_, _24110_);
  and _74483_ (_24115_, _14926_, _07910_);
  or _74484_ (_24116_, _24040_, _06279_);
  or _74485_ (_24117_, _24116_, _24115_);
  and _74486_ (_24118_, _24117_, _01347_);
  and _74487_ (_24119_, _24118_, _24114_);
  or _74488_ (_24120_, _24119_, _24039_);
  and _74489_ (_43230_, _24120_, _42618_);
  and _74490_ (_24121_, _01351_, \oc8051_golden_model_1.TH1 [3]);
  and _74491_ (_24123_, _11985_, \oc8051_golden_model_1.TH1 [3]);
  and _74492_ (_24124_, _14953_, _07910_);
  or _74493_ (_24125_, _24124_, _24123_);
  or _74494_ (_24126_, _24125_, _07151_);
  and _74495_ (_24127_, _07910_, \oc8051_golden_model_1.ACC [3]);
  or _74496_ (_24128_, _24127_, _24123_);
  and _74497_ (_24129_, _24128_, _07141_);
  and _74498_ (_24130_, _07142_, \oc8051_golden_model_1.TH1 [3]);
  or _74499_ (_24131_, _24130_, _06341_);
  or _74500_ (_24132_, _24131_, _24129_);
  and _74501_ (_24133_, _24132_, _07166_);
  and _74502_ (_24134_, _24133_, _24126_);
  nor _74503_ (_24135_, _11985_, _07594_);
  or _74504_ (_24136_, _24135_, _24123_);
  and _74505_ (_24137_, _24136_, _06461_);
  or _74506_ (_24138_, _24137_, _24134_);
  and _74507_ (_24139_, _24138_, _06465_);
  and _74508_ (_24140_, _24128_, _06464_);
  or _74509_ (_24141_, _24140_, _10080_);
  or _74510_ (_24142_, _24141_, _24139_);
  or _74511_ (_24144_, _24136_, _07215_);
  and _74512_ (_24145_, _24144_, _24142_);
  or _74513_ (_24146_, _24145_, _07460_);
  and _74514_ (_24147_, _09449_, _07910_);
  or _74515_ (_24148_, _24123_, _07208_);
  or _74516_ (_24149_, _24148_, _24147_);
  and _74517_ (_24150_, _24149_, _05982_);
  and _74518_ (_24151_, _24150_, _24146_);
  and _74519_ (_24152_, _15048_, _07910_);
  or _74520_ (_24153_, _24152_, _24123_);
  and _74521_ (_24155_, _24153_, _10094_);
  or _74522_ (_24156_, _24155_, _06218_);
  or _74523_ (_24157_, _24156_, _24151_);
  and _74524_ (_24158_, _07910_, _08930_);
  or _74525_ (_24159_, _24158_, _24123_);
  or _74526_ (_24160_, _24159_, _06219_);
  and _74527_ (_24161_, _24160_, _24157_);
  or _74528_ (_24162_, _24161_, _06369_);
  and _74529_ (_24163_, _14943_, _07910_);
  or _74530_ (_24164_, _24163_, _24123_);
  or _74531_ (_24166_, _24164_, _07237_);
  and _74532_ (_24167_, _24166_, _07240_);
  and _74533_ (_24168_, _24167_, _24162_);
  and _74534_ (_24169_, _12577_, _07910_);
  or _74535_ (_24170_, _24169_, _24123_);
  and _74536_ (_24171_, _24170_, _06536_);
  or _74537_ (_24172_, _24171_, _24168_);
  and _74538_ (_24173_, _24172_, _07242_);
  or _74539_ (_24174_, _24123_, _08292_);
  and _74540_ (_24175_, _24159_, _06375_);
  and _74541_ (_24177_, _24175_, _24174_);
  or _74542_ (_24178_, _24177_, _24173_);
  and _74543_ (_24179_, _24178_, _07234_);
  and _74544_ (_24180_, _24128_, _06545_);
  and _74545_ (_24181_, _24180_, _24174_);
  or _74546_ (_24182_, _24181_, _06366_);
  or _74547_ (_24183_, _24182_, _24179_);
  and _74548_ (_24184_, _14940_, _07910_);
  or _74549_ (_24185_, _24123_, _09056_);
  or _74550_ (_24186_, _24185_, _24184_);
  and _74551_ (_24188_, _24186_, _09061_);
  and _74552_ (_24189_, _24188_, _24183_);
  nor _74553_ (_24190_, _11256_, _11985_);
  or _74554_ (_24191_, _24190_, _24123_);
  and _74555_ (_24192_, _24191_, _06528_);
  or _74556_ (_24193_, _24192_, _24189_);
  and _74557_ (_24194_, _24193_, _06926_);
  and _74558_ (_24195_, _24125_, _06568_);
  or _74559_ (_24196_, _24195_, _06278_);
  or _74560_ (_24197_, _24196_, _24194_);
  and _74561_ (_24199_, _15128_, _07910_);
  or _74562_ (_24200_, _24123_, _06279_);
  or _74563_ (_24201_, _24200_, _24199_);
  and _74564_ (_24202_, _24201_, _01347_);
  and _74565_ (_24203_, _24202_, _24197_);
  or _74566_ (_24204_, _24203_, _24121_);
  and _74567_ (_43231_, _24204_, _42618_);
  and _74568_ (_24205_, _01351_, \oc8051_golden_model_1.TH1 [4]);
  and _74569_ (_24206_, _11985_, \oc8051_golden_model_1.TH1 [4]);
  nor _74570_ (_24207_, _08541_, _11985_);
  or _74571_ (_24209_, _24207_, _24206_);
  or _74572_ (_24210_, _24209_, _07215_);
  and _74573_ (_24211_, _15162_, _07910_);
  or _74574_ (_24212_, _24211_, _24206_);
  or _74575_ (_24213_, _24212_, _07151_);
  and _74576_ (_24214_, _07910_, \oc8051_golden_model_1.ACC [4]);
  or _74577_ (_24215_, _24214_, _24206_);
  and _74578_ (_24216_, _24215_, _07141_);
  and _74579_ (_24217_, _07142_, \oc8051_golden_model_1.TH1 [4]);
  or _74580_ (_24218_, _24217_, _06341_);
  or _74581_ (_24220_, _24218_, _24216_);
  and _74582_ (_24221_, _24220_, _07166_);
  and _74583_ (_24222_, _24221_, _24213_);
  and _74584_ (_24223_, _24209_, _06461_);
  or _74585_ (_24224_, _24223_, _24222_);
  and _74586_ (_24225_, _24224_, _06465_);
  and _74587_ (_24226_, _24215_, _06464_);
  or _74588_ (_24227_, _24226_, _10080_);
  or _74589_ (_24228_, _24227_, _24225_);
  and _74590_ (_24229_, _24228_, _24210_);
  or _74591_ (_24231_, _24229_, _07460_);
  and _74592_ (_24232_, _09448_, _07910_);
  or _74593_ (_24233_, _24206_, _07208_);
  or _74594_ (_24234_, _24233_, _24232_);
  and _74595_ (_24235_, _24234_, _24231_);
  or _74596_ (_24236_, _24235_, _10094_);
  and _74597_ (_24237_, _15254_, _07910_);
  or _74598_ (_24238_, _24206_, _05982_);
  or _74599_ (_24239_, _24238_, _24237_);
  and _74600_ (_24240_, _24239_, _06219_);
  and _74601_ (_24241_, _24240_, _24236_);
  and _74602_ (_24242_, _08959_, _07910_);
  or _74603_ (_24243_, _24242_, _24206_);
  and _74604_ (_24244_, _24243_, _06218_);
  or _74605_ (_24245_, _24244_, _06369_);
  or _74606_ (_24246_, _24245_, _24241_);
  and _74607_ (_24247_, _15269_, _07910_);
  or _74608_ (_24248_, _24247_, _24206_);
  or _74609_ (_24249_, _24248_, _07237_);
  and _74610_ (_24250_, _24249_, _07240_);
  and _74611_ (_24251_, _24250_, _24246_);
  and _74612_ (_24252_, _11254_, _07910_);
  or _74613_ (_24253_, _24252_, _24206_);
  and _74614_ (_24254_, _24253_, _06536_);
  or _74615_ (_24255_, _24254_, _24251_);
  and _74616_ (_24256_, _24255_, _07242_);
  or _74617_ (_24257_, _24206_, _08544_);
  and _74618_ (_24258_, _24243_, _06375_);
  and _74619_ (_24259_, _24258_, _24257_);
  or _74620_ (_24260_, _24259_, _24256_);
  and _74621_ (_24262_, _24260_, _07234_);
  and _74622_ (_24263_, _24215_, _06545_);
  and _74623_ (_24264_, _24263_, _24257_);
  or _74624_ (_24265_, _24264_, _06366_);
  or _74625_ (_24266_, _24265_, _24262_);
  and _74626_ (_24267_, _15266_, _07910_);
  or _74627_ (_24268_, _24206_, _09056_);
  or _74628_ (_24269_, _24268_, _24267_);
  and _74629_ (_24270_, _24269_, _09061_);
  and _74630_ (_24271_, _24270_, _24266_);
  nor _74631_ (_24273_, _11253_, _11985_);
  or _74632_ (_24274_, _24273_, _24206_);
  and _74633_ (_24275_, _24274_, _06528_);
  or _74634_ (_24276_, _24275_, _24271_);
  and _74635_ (_24277_, _24276_, _06926_);
  and _74636_ (_24278_, _24212_, _06568_);
  or _74637_ (_24279_, _24278_, _06278_);
  or _74638_ (_24280_, _24279_, _24277_);
  and _74639_ (_24281_, _15329_, _07910_);
  or _74640_ (_24282_, _24206_, _06279_);
  or _74641_ (_24285_, _24282_, _24281_);
  and _74642_ (_24286_, _24285_, _01347_);
  and _74643_ (_24287_, _24286_, _24280_);
  or _74644_ (_24288_, _24287_, _24205_);
  and _74645_ (_43232_, _24288_, _42618_);
  and _74646_ (_24289_, _01351_, \oc8051_golden_model_1.TH1 [5]);
  and _74647_ (_24290_, _11985_, \oc8051_golden_model_1.TH1 [5]);
  nor _74648_ (_24291_, _08244_, _11985_);
  or _74649_ (_24292_, _24291_, _24290_);
  or _74650_ (_24293_, _24292_, _07215_);
  and _74651_ (_24295_, _15358_, _07910_);
  or _74652_ (_24296_, _24295_, _24290_);
  or _74653_ (_24297_, _24296_, _07151_);
  and _74654_ (_24298_, _07910_, \oc8051_golden_model_1.ACC [5]);
  or _74655_ (_24299_, _24298_, _24290_);
  and _74656_ (_24300_, _24299_, _07141_);
  and _74657_ (_24301_, _07142_, \oc8051_golden_model_1.TH1 [5]);
  or _74658_ (_24302_, _24301_, _06341_);
  or _74659_ (_24303_, _24302_, _24300_);
  and _74660_ (_24304_, _24303_, _07166_);
  and _74661_ (_24306_, _24304_, _24297_);
  and _74662_ (_24307_, _24292_, _06461_);
  or _74663_ (_24308_, _24307_, _24306_);
  and _74664_ (_24309_, _24308_, _06465_);
  and _74665_ (_24310_, _24299_, _06464_);
  or _74666_ (_24311_, _24310_, _10080_);
  or _74667_ (_24312_, _24311_, _24309_);
  and _74668_ (_24313_, _24312_, _24293_);
  or _74669_ (_24314_, _24313_, _07460_);
  and _74670_ (_24315_, _09447_, _07910_);
  or _74671_ (_24317_, _24290_, _07208_);
  or _74672_ (_24318_, _24317_, _24315_);
  and _74673_ (_24319_, _24318_, _05982_);
  and _74674_ (_24320_, _24319_, _24314_);
  and _74675_ (_24321_, _15459_, _07910_);
  or _74676_ (_24322_, _24321_, _24290_);
  and _74677_ (_24323_, _24322_, _10094_);
  or _74678_ (_24324_, _24323_, _06218_);
  or _74679_ (_24325_, _24324_, _24320_);
  and _74680_ (_24326_, _08946_, _07910_);
  or _74681_ (_24328_, _24326_, _24290_);
  or _74682_ (_24329_, _24328_, _06219_);
  and _74683_ (_24330_, _24329_, _24325_);
  or _74684_ (_24331_, _24330_, _06369_);
  and _74685_ (_24332_, _15353_, _07910_);
  or _74686_ (_24333_, _24332_, _24290_);
  or _74687_ (_24334_, _24333_, _07237_);
  and _74688_ (_24335_, _24334_, _07240_);
  and _74689_ (_24336_, _24335_, _24331_);
  and _74690_ (_24337_, _11250_, _07910_);
  or _74691_ (_24339_, _24337_, _24290_);
  and _74692_ (_24340_, _24339_, _06536_);
  or _74693_ (_24341_, _24340_, _24336_);
  and _74694_ (_24342_, _24341_, _07242_);
  or _74695_ (_24343_, _24290_, _08247_);
  and _74696_ (_24344_, _24328_, _06375_);
  and _74697_ (_24345_, _24344_, _24343_);
  or _74698_ (_24346_, _24345_, _24342_);
  and _74699_ (_24347_, _24346_, _07234_);
  and _74700_ (_24348_, _24299_, _06545_);
  and _74701_ (_24350_, _24348_, _24343_);
  or _74702_ (_24351_, _24350_, _06366_);
  or _74703_ (_24352_, _24351_, _24347_);
  and _74704_ (_24353_, _15350_, _07910_);
  or _74705_ (_24354_, _24290_, _09056_);
  or _74706_ (_24355_, _24354_, _24353_);
  and _74707_ (_24356_, _24355_, _09061_);
  and _74708_ (_24357_, _24356_, _24352_);
  nor _74709_ (_24358_, _11249_, _11985_);
  or _74710_ (_24359_, _24358_, _24290_);
  and _74711_ (_24361_, _24359_, _06528_);
  or _74712_ (_24362_, _24361_, _24357_);
  and _74713_ (_24363_, _24362_, _06926_);
  and _74714_ (_24364_, _24296_, _06568_);
  or _74715_ (_24365_, _24364_, _06278_);
  or _74716_ (_24366_, _24365_, _24363_);
  and _74717_ (_24367_, _15532_, _07910_);
  or _74718_ (_24368_, _24290_, _06279_);
  or _74719_ (_24369_, _24368_, _24367_);
  and _74720_ (_24370_, _24369_, _01347_);
  and _74721_ (_24372_, _24370_, _24366_);
  or _74722_ (_24373_, _24372_, _24289_);
  and _74723_ (_43233_, _24373_, _42618_);
  and _74724_ (_24374_, _01351_, \oc8051_golden_model_1.TH1 [6]);
  and _74725_ (_24375_, _11985_, \oc8051_golden_model_1.TH1 [6]);
  and _74726_ (_24376_, _15554_, _07910_);
  or _74727_ (_24377_, _24376_, _24375_);
  or _74728_ (_24378_, _24377_, _07151_);
  and _74729_ (_24379_, _07910_, \oc8051_golden_model_1.ACC [6]);
  or _74730_ (_24380_, _24379_, _24375_);
  and _74731_ (_24382_, _24380_, _07141_);
  and _74732_ (_24383_, _07142_, \oc8051_golden_model_1.TH1 [6]);
  or _74733_ (_24384_, _24383_, _06341_);
  or _74734_ (_24385_, _24384_, _24382_);
  and _74735_ (_24386_, _24385_, _07166_);
  and _74736_ (_24387_, _24386_, _24378_);
  nor _74737_ (_24388_, _08142_, _11985_);
  or _74738_ (_24389_, _24388_, _24375_);
  and _74739_ (_24390_, _24389_, _06461_);
  or _74740_ (_24391_, _24390_, _24387_);
  and _74741_ (_24393_, _24391_, _06465_);
  and _74742_ (_24394_, _24380_, _06464_);
  or _74743_ (_24395_, _24394_, _10080_);
  or _74744_ (_24396_, _24395_, _24393_);
  or _74745_ (_24397_, _24389_, _07215_);
  and _74746_ (_24398_, _24397_, _24396_);
  or _74747_ (_24399_, _24398_, _07460_);
  and _74748_ (_24400_, _09446_, _07910_);
  or _74749_ (_24401_, _24375_, _07208_);
  or _74750_ (_24402_, _24401_, _24400_);
  and _74751_ (_24404_, _24402_, _05982_);
  and _74752_ (_24405_, _24404_, _24399_);
  and _74753_ (_24406_, _15657_, _07910_);
  or _74754_ (_24407_, _24406_, _24375_);
  and _74755_ (_24408_, _24407_, _10094_);
  or _74756_ (_24409_, _24408_, _06218_);
  or _74757_ (_24410_, _24409_, _24405_);
  and _74758_ (_24411_, _15664_, _07910_);
  or _74759_ (_24412_, _24411_, _24375_);
  or _74760_ (_24413_, _24412_, _06219_);
  and _74761_ (_24415_, _24413_, _24410_);
  or _74762_ (_24416_, _24415_, _06369_);
  and _74763_ (_24417_, _15549_, _07910_);
  or _74764_ (_24418_, _24417_, _24375_);
  or _74765_ (_24419_, _24418_, _07237_);
  and _74766_ (_24420_, _24419_, _07240_);
  and _74767_ (_24421_, _24420_, _24416_);
  and _74768_ (_24422_, _11247_, _07910_);
  or _74769_ (_24423_, _24422_, _24375_);
  and _74770_ (_24424_, _24423_, _06536_);
  or _74771_ (_24426_, _24424_, _24421_);
  and _74772_ (_24427_, _24426_, _07242_);
  or _74773_ (_24428_, _24375_, _08145_);
  and _74774_ (_24429_, _24412_, _06375_);
  and _74775_ (_24430_, _24429_, _24428_);
  or _74776_ (_24431_, _24430_, _24427_);
  and _74777_ (_24432_, _24431_, _07234_);
  and _74778_ (_24433_, _24380_, _06545_);
  and _74779_ (_24434_, _24433_, _24428_);
  or _74780_ (_24435_, _24434_, _06366_);
  or _74781_ (_24437_, _24435_, _24432_);
  and _74782_ (_24438_, _15546_, _07910_);
  or _74783_ (_24439_, _24375_, _09056_);
  or _74784_ (_24440_, _24439_, _24438_);
  and _74785_ (_24441_, _24440_, _09061_);
  and _74786_ (_24442_, _24441_, _24437_);
  nor _74787_ (_24443_, _11246_, _11985_);
  or _74788_ (_24444_, _24443_, _24375_);
  and _74789_ (_24445_, _24444_, _06528_);
  or _74790_ (_24446_, _24445_, _24442_);
  and _74791_ (_24448_, _24446_, _06926_);
  and _74792_ (_24449_, _24377_, _06568_);
  or _74793_ (_24450_, _24449_, _06278_);
  or _74794_ (_24451_, _24450_, _24448_);
  and _74795_ (_24452_, _15734_, _07910_);
  or _74796_ (_24453_, _24375_, _06279_);
  or _74797_ (_24454_, _24453_, _24452_);
  and _74798_ (_24455_, _24454_, _01347_);
  and _74799_ (_24456_, _24455_, _24451_);
  or _74800_ (_24457_, _24456_, _24374_);
  and _74801_ (_43234_, _24457_, _42618_);
  and _74802_ (_24459_, _01351_, \oc8051_golden_model_1.TH0 [0]);
  and _74803_ (_24460_, _07922_, \oc8051_golden_model_1.ACC [0]);
  and _74804_ (_24461_, _24460_, _08390_);
  and _74805_ (_24462_, _12063_, \oc8051_golden_model_1.TH0 [0]);
  or _74806_ (_24463_, _24462_, _07234_);
  or _74807_ (_24464_, _24463_, _24461_);
  or _74808_ (_24465_, _24462_, _24460_);
  and _74809_ (_24466_, _24465_, _06464_);
  or _74810_ (_24467_, _24466_, _10080_);
  nor _74811_ (_24469_, _08390_, _12063_);
  or _74812_ (_24470_, _24469_, _24462_);
  and _74813_ (_24471_, _24470_, _06341_);
  and _74814_ (_24472_, _07142_, \oc8051_golden_model_1.TH0 [0]);
  and _74815_ (_24473_, _24465_, _07141_);
  or _74816_ (_24474_, _24473_, _24472_);
  and _74817_ (_24475_, _24474_, _07151_);
  or _74818_ (_24476_, _24475_, _06461_);
  or _74819_ (_24477_, _24476_, _24471_);
  and _74820_ (_24478_, _24477_, _06465_);
  or _74821_ (_24480_, _24478_, _24467_);
  and _74822_ (_24481_, _07922_, _07133_);
  or _74823_ (_24482_, _24462_, _22611_);
  or _74824_ (_24483_, _24482_, _24481_);
  and _74825_ (_24484_, _24483_, _24480_);
  or _74826_ (_24485_, _24484_, _07460_);
  and _74827_ (_24486_, _09392_, _07922_);
  or _74828_ (_24487_, _24462_, _07208_);
  or _74829_ (_24488_, _24487_, _24486_);
  and _74830_ (_24489_, _24488_, _24485_);
  or _74831_ (_24491_, _24489_, _10094_);
  and _74832_ (_24492_, _14467_, _07922_);
  or _74833_ (_24493_, _24462_, _05982_);
  or _74834_ (_24494_, _24493_, _24492_);
  and _74835_ (_24495_, _24494_, _06219_);
  and _74836_ (_24496_, _24495_, _24491_);
  and _74837_ (_24497_, _07922_, _08954_);
  or _74838_ (_24498_, _24497_, _24462_);
  and _74839_ (_24499_, _24498_, _06218_);
  or _74840_ (_24500_, _24499_, _06369_);
  or _74841_ (_24502_, _24500_, _24496_);
  and _74842_ (_24503_, _14366_, _07922_);
  or _74843_ (_24504_, _24503_, _24462_);
  or _74844_ (_24505_, _24504_, _07237_);
  and _74845_ (_24506_, _24505_, _07240_);
  and _74846_ (_24507_, _24506_, _24502_);
  nor _74847_ (_24508_, _12580_, _12063_);
  or _74848_ (_24509_, _24508_, _24462_);
  nor _74849_ (_24510_, _24461_, _07240_);
  and _74850_ (_24511_, _24510_, _24509_);
  or _74851_ (_24512_, _24511_, _24507_);
  and _74852_ (_24513_, _24512_, _07242_);
  nand _74853_ (_24514_, _24498_, _06375_);
  nor _74854_ (_24515_, _24514_, _24469_);
  or _74855_ (_24516_, _24515_, _06545_);
  or _74856_ (_24517_, _24516_, _24513_);
  and _74857_ (_24518_, _24517_, _24464_);
  or _74858_ (_24519_, _24518_, _06366_);
  and _74859_ (_24520_, _14363_, _07922_);
  or _74860_ (_24521_, _24462_, _09056_);
  or _74861_ (_24524_, _24521_, _24520_);
  and _74862_ (_24525_, _24524_, _09061_);
  and _74863_ (_24526_, _24525_, _24519_);
  and _74864_ (_24527_, _24509_, _06528_);
  or _74865_ (_24528_, _24527_, _19502_);
  or _74866_ (_24529_, _24528_, _24526_);
  or _74867_ (_24530_, _24470_, _06661_);
  and _74868_ (_24531_, _24530_, _01347_);
  and _74869_ (_24532_, _24531_, _24529_);
  or _74870_ (_24533_, _24532_, _24459_);
  and _74871_ (_43236_, _24533_, _42618_);
  not _74872_ (_24535_, \oc8051_golden_model_1.TH0 [1]);
  nor _74873_ (_24536_, _01347_, _24535_);
  nor _74874_ (_24537_, _07922_, _24535_);
  nor _74875_ (_24538_, _12063_, _07357_);
  or _74876_ (_24539_, _24538_, _24537_);
  or _74877_ (_24540_, _24539_, _07215_);
  or _74878_ (_24541_, _07922_, \oc8051_golden_model_1.TH0 [1]);
  and _74879_ (_24542_, _14562_, _07922_);
  not _74880_ (_24543_, _24542_);
  and _74881_ (_24545_, _24543_, _24541_);
  or _74882_ (_24546_, _24545_, _07151_);
  and _74883_ (_24547_, _07922_, \oc8051_golden_model_1.ACC [1]);
  or _74884_ (_24548_, _24547_, _24537_);
  and _74885_ (_24549_, _24548_, _07141_);
  nor _74886_ (_24550_, _07141_, _24535_);
  or _74887_ (_24551_, _24550_, _06341_);
  or _74888_ (_24552_, _24551_, _24549_);
  and _74889_ (_24553_, _24552_, _07166_);
  and _74890_ (_24554_, _24553_, _24546_);
  and _74891_ (_24556_, _24539_, _06461_);
  or _74892_ (_24557_, _24556_, _24554_);
  and _74893_ (_24558_, _24557_, _06465_);
  and _74894_ (_24559_, _24548_, _06464_);
  or _74895_ (_24560_, _24559_, _10080_);
  or _74896_ (_24561_, _24560_, _24558_);
  and _74897_ (_24562_, _24561_, _24540_);
  or _74898_ (_24563_, _24562_, _07460_);
  and _74899_ (_24564_, _09451_, _07922_);
  or _74900_ (_24565_, _24537_, _07208_);
  or _74901_ (_24567_, _24565_, _24564_);
  and _74902_ (_24568_, _24567_, _05982_);
  and _74903_ (_24569_, _24568_, _24563_);
  or _74904_ (_24570_, _14653_, _12063_);
  and _74905_ (_24571_, _24541_, _10094_);
  and _74906_ (_24572_, _24571_, _24570_);
  or _74907_ (_24573_, _24572_, _24569_);
  and _74908_ (_24574_, _24573_, _06219_);
  nand _74909_ (_24575_, _07922_, _07038_);
  and _74910_ (_24576_, _24541_, _06218_);
  and _74911_ (_24578_, _24576_, _24575_);
  or _74912_ (_24579_, _24578_, _24574_);
  and _74913_ (_24580_, _24579_, _07237_);
  or _74914_ (_24581_, _14668_, _12063_);
  and _74915_ (_24582_, _24541_, _06369_);
  and _74916_ (_24583_, _24582_, _24581_);
  or _74917_ (_24584_, _24583_, _06536_);
  or _74918_ (_24585_, _24584_, _24580_);
  nor _74919_ (_24586_, _11261_, _12063_);
  or _74920_ (_24587_, _24586_, _24537_);
  nand _74921_ (_24589_, _11260_, _07922_);
  and _74922_ (_24590_, _24589_, _24587_);
  or _74923_ (_24591_, _24590_, _07240_);
  and _74924_ (_24592_, _24591_, _07242_);
  and _74925_ (_24593_, _24592_, _24585_);
  or _74926_ (_24594_, _14666_, _12063_);
  and _74927_ (_24595_, _24541_, _06375_);
  and _74928_ (_24596_, _24595_, _24594_);
  or _74929_ (_24597_, _24596_, _06545_);
  or _74930_ (_24598_, _24597_, _24593_);
  nor _74931_ (_24600_, _24537_, _07234_);
  nand _74932_ (_24601_, _24600_, _24589_);
  and _74933_ (_24602_, _24601_, _09056_);
  and _74934_ (_24603_, _24602_, _24598_);
  or _74935_ (_24604_, _24575_, _08341_);
  and _74936_ (_24605_, _24541_, _06366_);
  and _74937_ (_24606_, _24605_, _24604_);
  or _74938_ (_24607_, _24606_, _06528_);
  or _74939_ (_24608_, _24607_, _24603_);
  or _74940_ (_24609_, _24587_, _09061_);
  and _74941_ (_24611_, _24609_, _06926_);
  and _74942_ (_24612_, _24611_, _24608_);
  and _74943_ (_24613_, _24545_, _06568_);
  or _74944_ (_24614_, _24613_, _06278_);
  or _74945_ (_24615_, _24614_, _24612_);
  or _74946_ (_24616_, _24537_, _06279_);
  or _74947_ (_24617_, _24616_, _24542_);
  and _74948_ (_24618_, _24617_, _01347_);
  and _74949_ (_24619_, _24618_, _24615_);
  or _74950_ (_24620_, _24619_, _24536_);
  and _74951_ (_43237_, _24620_, _42618_);
  and _74952_ (_24622_, _01351_, \oc8051_golden_model_1.TH0 [2]);
  and _74953_ (_24623_, _12063_, \oc8051_golden_model_1.TH0 [2]);
  and _74954_ (_24624_, _09450_, _07922_);
  or _74955_ (_24625_, _24624_, _24623_);
  and _74956_ (_24626_, _24625_, _07460_);
  and _74957_ (_24627_, _14770_, _07922_);
  or _74958_ (_24628_, _24627_, _24623_);
  or _74959_ (_24629_, _24628_, _07151_);
  and _74960_ (_24630_, _07922_, \oc8051_golden_model_1.ACC [2]);
  or _74961_ (_24632_, _24630_, _24623_);
  and _74962_ (_24633_, _24632_, _07141_);
  and _74963_ (_24634_, _07142_, \oc8051_golden_model_1.TH0 [2]);
  or _74964_ (_24635_, _24634_, _06341_);
  or _74965_ (_24636_, _24635_, _24633_);
  and _74966_ (_24637_, _24636_, _07166_);
  and _74967_ (_24638_, _24637_, _24629_);
  nor _74968_ (_24639_, _12063_, _07776_);
  or _74969_ (_24640_, _24639_, _24623_);
  and _74970_ (_24641_, _24640_, _06461_);
  or _74971_ (_24643_, _24641_, _24638_);
  and _74972_ (_24644_, _24643_, _06465_);
  and _74973_ (_24645_, _24632_, _06464_);
  or _74974_ (_24646_, _24645_, _10080_);
  or _74975_ (_24647_, _24646_, _24644_);
  or _74976_ (_24648_, _24640_, _07215_);
  and _74977_ (_24649_, _24648_, _07208_);
  and _74978_ (_24650_, _24649_, _24647_);
  or _74979_ (_24651_, _24650_, _10094_);
  or _74980_ (_24652_, _24651_, _24626_);
  and _74981_ (_24654_, _14859_, _07922_);
  or _74982_ (_24655_, _24623_, _05982_);
  or _74983_ (_24656_, _24655_, _24654_);
  and _74984_ (_24657_, _24656_, _06219_);
  and _74985_ (_24658_, _24657_, _24652_);
  and _74986_ (_24659_, _07922_, _08973_);
  or _74987_ (_24660_, _24659_, _24623_);
  and _74988_ (_24661_, _24660_, _06218_);
  or _74989_ (_24662_, _24661_, _06369_);
  or _74990_ (_24663_, _24662_, _24658_);
  and _74991_ (_24665_, _14751_, _07922_);
  or _74992_ (_24666_, _24665_, _24623_);
  or _74993_ (_24667_, _24666_, _07237_);
  and _74994_ (_24668_, _24667_, _07240_);
  and _74995_ (_24669_, _24668_, _24663_);
  and _74996_ (_24670_, _11259_, _07922_);
  or _74997_ (_24671_, _24670_, _24623_);
  and _74998_ (_24672_, _24671_, _06536_);
  or _74999_ (_24673_, _24672_, _24669_);
  and _75000_ (_24674_, _24673_, _07242_);
  or _75001_ (_24676_, _24623_, _08440_);
  and _75002_ (_24677_, _24660_, _06375_);
  and _75003_ (_24678_, _24677_, _24676_);
  or _75004_ (_24679_, _24678_, _24674_);
  and _75005_ (_24680_, _24679_, _07234_);
  and _75006_ (_24681_, _24632_, _06545_);
  and _75007_ (_24682_, _24681_, _24676_);
  or _75008_ (_24683_, _24682_, _06366_);
  or _75009_ (_24684_, _24683_, _24680_);
  and _75010_ (_24685_, _14748_, _07922_);
  or _75011_ (_24687_, _24623_, _09056_);
  or _75012_ (_24688_, _24687_, _24685_);
  and _75013_ (_24689_, _24688_, _09061_);
  and _75014_ (_24690_, _24689_, _24684_);
  nor _75015_ (_24691_, _11258_, _12063_);
  or _75016_ (_24692_, _24691_, _24623_);
  and _75017_ (_24693_, _24692_, _06528_);
  or _75018_ (_24694_, _24693_, _24690_);
  and _75019_ (_24695_, _24694_, _06926_);
  and _75020_ (_24696_, _24628_, _06568_);
  or _75021_ (_24698_, _24696_, _06278_);
  or _75022_ (_24699_, _24698_, _24695_);
  and _75023_ (_24700_, _14926_, _07922_);
  or _75024_ (_24701_, _24623_, _06279_);
  or _75025_ (_24702_, _24701_, _24700_);
  and _75026_ (_24703_, _24702_, _01347_);
  and _75027_ (_24704_, _24703_, _24699_);
  or _75028_ (_24705_, _24704_, _24622_);
  and _75029_ (_43238_, _24705_, _42618_);
  and _75030_ (_24706_, _01351_, \oc8051_golden_model_1.TH0 [3]);
  and _75031_ (_24708_, _12063_, \oc8051_golden_model_1.TH0 [3]);
  and _75032_ (_24709_, _14953_, _07922_);
  or _75033_ (_24710_, _24709_, _24708_);
  or _75034_ (_24711_, _24710_, _07151_);
  and _75035_ (_24712_, _07922_, \oc8051_golden_model_1.ACC [3]);
  or _75036_ (_24713_, _24712_, _24708_);
  and _75037_ (_24714_, _24713_, _07141_);
  and _75038_ (_24715_, _07142_, \oc8051_golden_model_1.TH0 [3]);
  or _75039_ (_24716_, _24715_, _06341_);
  or _75040_ (_24717_, _24716_, _24714_);
  and _75041_ (_24719_, _24717_, _07166_);
  and _75042_ (_24720_, _24719_, _24711_);
  nor _75043_ (_24721_, _12063_, _07594_);
  or _75044_ (_24722_, _24721_, _24708_);
  and _75045_ (_24723_, _24722_, _06461_);
  or _75046_ (_24724_, _24723_, _24720_);
  and _75047_ (_24725_, _24724_, _06465_);
  and _75048_ (_24726_, _24713_, _06464_);
  or _75049_ (_24727_, _24726_, _10080_);
  or _75050_ (_24728_, _24727_, _24725_);
  or _75051_ (_24730_, _24722_, _07215_);
  and _75052_ (_24731_, _24730_, _24728_);
  or _75053_ (_24732_, _24731_, _07460_);
  and _75054_ (_24733_, _09449_, _07922_);
  or _75055_ (_24734_, _24708_, _07208_);
  or _75056_ (_24735_, _24734_, _24733_);
  and _75057_ (_24736_, _24735_, _05982_);
  and _75058_ (_24737_, _24736_, _24732_);
  and _75059_ (_24738_, _15048_, _07922_);
  or _75060_ (_24739_, _24738_, _24708_);
  and _75061_ (_24741_, _24739_, _10094_);
  or _75062_ (_24742_, _24741_, _06218_);
  or _75063_ (_24743_, _24742_, _24737_);
  and _75064_ (_24744_, _07922_, _08930_);
  or _75065_ (_24745_, _24744_, _24708_);
  or _75066_ (_24746_, _24745_, _06219_);
  and _75067_ (_24747_, _24746_, _24743_);
  or _75068_ (_24748_, _24747_, _06369_);
  and _75069_ (_24749_, _14943_, _07922_);
  or _75070_ (_24750_, _24749_, _24708_);
  or _75071_ (_24752_, _24750_, _07237_);
  and _75072_ (_24753_, _24752_, _07240_);
  and _75073_ (_24754_, _24753_, _24748_);
  and _75074_ (_24755_, _12577_, _07922_);
  or _75075_ (_24756_, _24755_, _24708_);
  and _75076_ (_24757_, _24756_, _06536_);
  or _75077_ (_24758_, _24757_, _24754_);
  and _75078_ (_24759_, _24758_, _07242_);
  or _75079_ (_24760_, _24708_, _08292_);
  and _75080_ (_24761_, _24745_, _06375_);
  and _75081_ (_24763_, _24761_, _24760_);
  or _75082_ (_24764_, _24763_, _24759_);
  and _75083_ (_24765_, _24764_, _07234_);
  and _75084_ (_24766_, _24713_, _06545_);
  and _75085_ (_24767_, _24766_, _24760_);
  or _75086_ (_24768_, _24767_, _06366_);
  or _75087_ (_24769_, _24768_, _24765_);
  and _75088_ (_24770_, _14940_, _07922_);
  or _75089_ (_24771_, _24708_, _09056_);
  or _75090_ (_24772_, _24771_, _24770_);
  and _75091_ (_24774_, _24772_, _09061_);
  and _75092_ (_24775_, _24774_, _24769_);
  nor _75093_ (_24776_, _11256_, _12063_);
  or _75094_ (_24777_, _24776_, _24708_);
  and _75095_ (_24778_, _24777_, _06528_);
  or _75096_ (_24779_, _24778_, _24775_);
  and _75097_ (_24780_, _24779_, _06926_);
  and _75098_ (_24781_, _24710_, _06568_);
  or _75099_ (_24782_, _24781_, _06278_);
  or _75100_ (_24783_, _24782_, _24780_);
  and _75101_ (_24785_, _15128_, _07922_);
  or _75102_ (_24786_, _24708_, _06279_);
  or _75103_ (_24787_, _24786_, _24785_);
  and _75104_ (_24788_, _24787_, _01347_);
  and _75105_ (_24789_, _24788_, _24783_);
  or _75106_ (_24790_, _24789_, _24706_);
  and _75107_ (_43239_, _24790_, _42618_);
  and _75108_ (_24791_, _01351_, \oc8051_golden_model_1.TH0 [4]);
  and _75109_ (_24792_, _12063_, \oc8051_golden_model_1.TH0 [4]);
  and _75110_ (_24793_, _15162_, _07922_);
  or _75111_ (_24795_, _24793_, _24792_);
  or _75112_ (_24796_, _24795_, _07151_);
  and _75113_ (_24797_, _07922_, \oc8051_golden_model_1.ACC [4]);
  or _75114_ (_24798_, _24797_, _24792_);
  and _75115_ (_24799_, _24798_, _07141_);
  and _75116_ (_24800_, _07142_, \oc8051_golden_model_1.TH0 [4]);
  or _75117_ (_24801_, _24800_, _06341_);
  or _75118_ (_24802_, _24801_, _24799_);
  and _75119_ (_24803_, _24802_, _07166_);
  and _75120_ (_24804_, _24803_, _24796_);
  nor _75121_ (_24806_, _08541_, _12063_);
  or _75122_ (_24807_, _24806_, _24792_);
  and _75123_ (_24808_, _24807_, _06461_);
  or _75124_ (_24809_, _24808_, _24804_);
  and _75125_ (_24810_, _24809_, _06465_);
  and _75126_ (_24811_, _24798_, _06464_);
  or _75127_ (_24812_, _24811_, _10080_);
  or _75128_ (_24813_, _24812_, _24810_);
  or _75129_ (_24814_, _24807_, _07215_);
  and _75130_ (_24815_, _24814_, _24813_);
  or _75131_ (_24817_, _24815_, _07460_);
  and _75132_ (_24818_, _09448_, _07922_);
  or _75133_ (_24819_, _24792_, _07208_);
  or _75134_ (_24820_, _24819_, _24818_);
  and _75135_ (_24821_, _24820_, _24817_);
  or _75136_ (_24822_, _24821_, _10094_);
  and _75137_ (_24823_, _15254_, _07922_);
  or _75138_ (_24824_, _24792_, _05982_);
  or _75139_ (_24825_, _24824_, _24823_);
  and _75140_ (_24826_, _24825_, _06219_);
  and _75141_ (_24828_, _24826_, _24822_);
  and _75142_ (_24829_, _08959_, _07922_);
  or _75143_ (_24830_, _24829_, _24792_);
  and _75144_ (_24831_, _24830_, _06218_);
  or _75145_ (_24832_, _24831_, _06369_);
  or _75146_ (_24833_, _24832_, _24828_);
  and _75147_ (_24834_, _15269_, _07922_);
  or _75148_ (_24835_, _24834_, _24792_);
  or _75149_ (_24836_, _24835_, _07237_);
  and _75150_ (_24837_, _24836_, _07240_);
  and _75151_ (_24839_, _24837_, _24833_);
  and _75152_ (_24840_, _11254_, _07922_);
  or _75153_ (_24841_, _24840_, _24792_);
  and _75154_ (_24842_, _24841_, _06536_);
  or _75155_ (_24843_, _24842_, _24839_);
  and _75156_ (_24844_, _24843_, _07242_);
  or _75157_ (_24845_, _24792_, _08544_);
  and _75158_ (_24846_, _24830_, _06375_);
  and _75159_ (_24847_, _24846_, _24845_);
  or _75160_ (_24848_, _24847_, _24844_);
  and _75161_ (_24850_, _24848_, _07234_);
  and _75162_ (_24851_, _24798_, _06545_);
  and _75163_ (_24852_, _24851_, _24845_);
  or _75164_ (_24853_, _24852_, _06366_);
  or _75165_ (_24854_, _24853_, _24850_);
  and _75166_ (_24855_, _15266_, _07922_);
  or _75167_ (_24856_, _24792_, _09056_);
  or _75168_ (_24857_, _24856_, _24855_);
  and _75169_ (_24858_, _24857_, _09061_);
  and _75170_ (_24859_, _24858_, _24854_);
  nor _75171_ (_24861_, _11253_, _12063_);
  or _75172_ (_24862_, _24861_, _24792_);
  and _75173_ (_24863_, _24862_, _06528_);
  or _75174_ (_24864_, _24863_, _24859_);
  and _75175_ (_24865_, _24864_, _06926_);
  and _75176_ (_24866_, _24795_, _06568_);
  or _75177_ (_24867_, _24866_, _06278_);
  or _75178_ (_24868_, _24867_, _24865_);
  and _75179_ (_24869_, _15329_, _07922_);
  or _75180_ (_24870_, _24792_, _06279_);
  or _75181_ (_24872_, _24870_, _24869_);
  and _75182_ (_24873_, _24872_, _01347_);
  and _75183_ (_24874_, _24873_, _24868_);
  or _75184_ (_24875_, _24874_, _24791_);
  and _75185_ (_43240_, _24875_, _42618_);
  and _75186_ (_24876_, _01351_, \oc8051_golden_model_1.TH0 [5]);
  and _75187_ (_24877_, _12063_, \oc8051_golden_model_1.TH0 [5]);
  nor _75188_ (_24878_, _08244_, _12063_);
  or _75189_ (_24879_, _24878_, _24877_);
  or _75190_ (_24880_, _24879_, _07215_);
  and _75191_ (_24882_, _15358_, _07922_);
  or _75192_ (_24883_, _24882_, _24877_);
  or _75193_ (_24884_, _24883_, _07151_);
  and _75194_ (_24885_, _07922_, \oc8051_golden_model_1.ACC [5]);
  or _75195_ (_24886_, _24885_, _24877_);
  and _75196_ (_24887_, _24886_, _07141_);
  and _75197_ (_24888_, _07142_, \oc8051_golden_model_1.TH0 [5]);
  or _75198_ (_24889_, _24888_, _06341_);
  or _75199_ (_24890_, _24889_, _24887_);
  and _75200_ (_24891_, _24890_, _07166_);
  and _75201_ (_24893_, _24891_, _24884_);
  and _75202_ (_24894_, _24879_, _06461_);
  or _75203_ (_24895_, _24894_, _24893_);
  and _75204_ (_24896_, _24895_, _06465_);
  and _75205_ (_24897_, _24886_, _06464_);
  or _75206_ (_24898_, _24897_, _10080_);
  or _75207_ (_24899_, _24898_, _24896_);
  and _75208_ (_24900_, _24899_, _24880_);
  or _75209_ (_24901_, _24900_, _07460_);
  and _75210_ (_24902_, _09447_, _07922_);
  or _75211_ (_24904_, _24877_, _07208_);
  or _75212_ (_24905_, _24904_, _24902_);
  and _75213_ (_24906_, _24905_, _05982_);
  and _75214_ (_24907_, _24906_, _24901_);
  and _75215_ (_24908_, _15459_, _07922_);
  or _75216_ (_24909_, _24908_, _24877_);
  and _75217_ (_24910_, _24909_, _10094_);
  or _75218_ (_24911_, _24910_, _06218_);
  or _75219_ (_24912_, _24911_, _24907_);
  and _75220_ (_24913_, _08946_, _07922_);
  or _75221_ (_24915_, _24913_, _24877_);
  or _75222_ (_24916_, _24915_, _06219_);
  and _75223_ (_24917_, _24916_, _24912_);
  or _75224_ (_24918_, _24917_, _06369_);
  and _75225_ (_24919_, _15353_, _07922_);
  or _75226_ (_24920_, _24919_, _24877_);
  or _75227_ (_24921_, _24920_, _07237_);
  and _75228_ (_24922_, _24921_, _07240_);
  and _75229_ (_24923_, _24922_, _24918_);
  and _75230_ (_24924_, _11250_, _07922_);
  or _75231_ (_24926_, _24924_, _24877_);
  and _75232_ (_24927_, _24926_, _06536_);
  or _75233_ (_24928_, _24927_, _24923_);
  and _75234_ (_24929_, _24928_, _07242_);
  or _75235_ (_24930_, _24877_, _08247_);
  and _75236_ (_24931_, _24915_, _06375_);
  and _75237_ (_24932_, _24931_, _24930_);
  or _75238_ (_24933_, _24932_, _24929_);
  and _75239_ (_24934_, _24933_, _07234_);
  and _75240_ (_24935_, _24886_, _06545_);
  and _75241_ (_24937_, _24935_, _24930_);
  or _75242_ (_24938_, _24937_, _06366_);
  or _75243_ (_24939_, _24938_, _24934_);
  and _75244_ (_24940_, _15350_, _07922_);
  or _75245_ (_24941_, _24877_, _09056_);
  or _75246_ (_24942_, _24941_, _24940_);
  and _75247_ (_24943_, _24942_, _09061_);
  and _75248_ (_24944_, _24943_, _24939_);
  nor _75249_ (_24945_, _11249_, _12063_);
  or _75250_ (_24946_, _24945_, _24877_);
  and _75251_ (_24948_, _24946_, _06528_);
  or _75252_ (_24949_, _24948_, _24944_);
  and _75253_ (_24950_, _24949_, _06926_);
  and _75254_ (_24951_, _24883_, _06568_);
  or _75255_ (_24952_, _24951_, _06278_);
  or _75256_ (_24953_, _24952_, _24950_);
  and _75257_ (_24954_, _15532_, _07922_);
  or _75258_ (_24955_, _24877_, _06279_);
  or _75259_ (_24956_, _24955_, _24954_);
  and _75260_ (_24957_, _24956_, _01347_);
  and _75261_ (_24959_, _24957_, _24953_);
  or _75262_ (_24960_, _24959_, _24876_);
  and _75263_ (_43242_, _24960_, _42618_);
  and _75264_ (_24961_, _01351_, \oc8051_golden_model_1.TH0 [6]);
  and _75265_ (_24962_, _12063_, \oc8051_golden_model_1.TH0 [6]);
  nor _75266_ (_24963_, _08142_, _12063_);
  or _75267_ (_24964_, _24963_, _24962_);
  or _75268_ (_24965_, _24964_, _07215_);
  and _75269_ (_24966_, _15554_, _07922_);
  or _75270_ (_24967_, _24966_, _24962_);
  or _75271_ (_24969_, _24967_, _07151_);
  and _75272_ (_24970_, _07922_, \oc8051_golden_model_1.ACC [6]);
  or _75273_ (_24971_, _24970_, _24962_);
  and _75274_ (_24972_, _24971_, _07141_);
  and _75275_ (_24973_, _07142_, \oc8051_golden_model_1.TH0 [6]);
  or _75276_ (_24974_, _24973_, _06341_);
  or _75277_ (_24975_, _24974_, _24972_);
  and _75278_ (_24976_, _24975_, _07166_);
  and _75279_ (_24977_, _24976_, _24969_);
  and _75280_ (_24978_, _24964_, _06461_);
  or _75281_ (_24980_, _24978_, _24977_);
  and _75282_ (_24981_, _24980_, _06465_);
  and _75283_ (_24982_, _24971_, _06464_);
  or _75284_ (_24983_, _24982_, _10080_);
  or _75285_ (_24984_, _24983_, _24981_);
  and _75286_ (_24985_, _24984_, _24965_);
  or _75287_ (_24986_, _24985_, _07460_);
  and _75288_ (_24987_, _09446_, _07922_);
  or _75289_ (_24988_, _24962_, _07208_);
  or _75290_ (_24989_, _24988_, _24987_);
  and _75291_ (_24991_, _24989_, _05982_);
  and _75292_ (_24992_, _24991_, _24986_);
  and _75293_ (_24993_, _15657_, _07922_);
  or _75294_ (_24994_, _24993_, _24962_);
  and _75295_ (_24995_, _24994_, _10094_);
  or _75296_ (_24996_, _24995_, _06218_);
  or _75297_ (_24997_, _24996_, _24992_);
  and _75298_ (_24998_, _15664_, _07922_);
  or _75299_ (_24999_, _24998_, _24962_);
  or _75300_ (_25000_, _24999_, _06219_);
  and _75301_ (_25002_, _25000_, _24997_);
  or _75302_ (_25003_, _25002_, _06369_);
  and _75303_ (_25004_, _15549_, _07922_);
  or _75304_ (_25005_, _25004_, _24962_);
  or _75305_ (_25006_, _25005_, _07237_);
  and _75306_ (_25007_, _25006_, _07240_);
  and _75307_ (_25008_, _25007_, _25003_);
  and _75308_ (_25009_, _11247_, _07922_);
  or _75309_ (_25010_, _25009_, _24962_);
  and _75310_ (_25011_, _25010_, _06536_);
  or _75311_ (_25013_, _25011_, _25008_);
  and _75312_ (_25014_, _25013_, _07242_);
  or _75313_ (_25015_, _24962_, _08145_);
  and _75314_ (_25016_, _24999_, _06375_);
  and _75315_ (_25017_, _25016_, _25015_);
  or _75316_ (_25018_, _25017_, _25014_);
  and _75317_ (_25019_, _25018_, _07234_);
  and _75318_ (_25020_, _24971_, _06545_);
  and _75319_ (_25021_, _25020_, _25015_);
  or _75320_ (_25022_, _25021_, _06366_);
  or _75321_ (_25024_, _25022_, _25019_);
  and _75322_ (_25025_, _15546_, _07922_);
  or _75323_ (_25026_, _24962_, _09056_);
  or _75324_ (_25027_, _25026_, _25025_);
  and _75325_ (_25028_, _25027_, _09061_);
  and _75326_ (_25029_, _25028_, _25024_);
  nor _75327_ (_25030_, _11246_, _12063_);
  or _75328_ (_25031_, _25030_, _24962_);
  and _75329_ (_25032_, _25031_, _06528_);
  or _75330_ (_25033_, _25032_, _25029_);
  and _75331_ (_25035_, _25033_, _06926_);
  and _75332_ (_25036_, _24967_, _06568_);
  or _75333_ (_25037_, _25036_, _06278_);
  or _75334_ (_25038_, _25037_, _25035_);
  and _75335_ (_25039_, _15734_, _07922_);
  or _75336_ (_25040_, _24962_, _06279_);
  or _75337_ (_25041_, _25040_, _25039_);
  and _75338_ (_25042_, _25041_, _01347_);
  and _75339_ (_25043_, _25042_, _25038_);
  or _75340_ (_25044_, _25043_, _24961_);
  and _75341_ (_43243_, _25044_, _42618_);
  and _75342_ (_25046_, _13052_, _12141_);
  nor _75343_ (_25047_, _25046_, _05630_);
  and _75344_ (_25048_, _13030_, _13037_);
  nor _75345_ (_25049_, _25048_, _05630_);
  and _75346_ (_25050_, _12151_, _11285_);
  nor _75347_ (_25051_, _25050_, _05630_);
  and _75348_ (_25052_, _10559_, \oc8051_golden_model_1.PC [0]);
  nor _75349_ (_25053_, _10559_, \oc8051_golden_model_1.PC [0]);
  nor _75350_ (_25054_, _25053_, _25052_);
  and _75351_ (_25055_, _25054_, _12800_);
  not _75352_ (_25056_, _12800_);
  and _75353_ (_25057_, _12162_, _09056_);
  nor _75354_ (_25058_, _25057_, _05630_);
  and _75355_ (_25059_, _10979_, _07242_);
  nor _75356_ (_25060_, _25059_, _05630_);
  not _75357_ (_25061_, _12755_);
  and _75358_ (_25062_, _12169_, _07237_);
  nor _75359_ (_25063_, _25062_, _05630_);
  not _75360_ (_25064_, _12733_);
  and _75361_ (_25067_, _06218_, _05630_);
  nor _75362_ (_25068_, _06872_, _06007_);
  and _75363_ (_25069_, _12587_, _05630_);
  and _75364_ (_25070_, _06872_, \oc8051_golden_model_1.PC [0]);
  nor _75365_ (_25071_, _25070_, _12251_);
  not _75366_ (_25072_, _25071_);
  nor _75367_ (_25073_, _25072_, _12587_);
  nor _75368_ (_25074_, _25073_, _25069_);
  nor _75369_ (_25075_, _25074_, _06774_);
  and _75370_ (_25076_, _12333_, _05630_);
  not _75371_ (_25078_, _25076_);
  and _75372_ (_25079_, _25071_, _12335_);
  nor _75373_ (_25080_, _25079_, _12177_);
  and _75374_ (_25081_, _25080_, _25078_);
  nor _75375_ (_25082_, _06872_, _06013_);
  and _75376_ (_25083_, _12513_, _05630_);
  nor _75377_ (_25084_, _12513_, _05630_);
  nor _75378_ (_25085_, _25084_, _25083_);
  and _75379_ (_25086_, _25085_, _07504_);
  nor _75380_ (_25087_, _06872_, _07504_);
  or _75381_ (_25089_, _25087_, _12516_);
  nor _75382_ (_25090_, _25089_, _25086_);
  nor _75383_ (_25091_, _12512_, _05630_);
  nor _75384_ (_25092_, _25091_, _25090_);
  nor _75385_ (_25093_, _25092_, _12387_);
  and _75386_ (_25094_, _12507_, \oc8051_golden_model_1.PC [0]);
  and _75387_ (_25095_, _06251_, _05630_);
  nor _75388_ (_25096_, _25095_, _12458_);
  and _75389_ (_25097_, _25096_, _12393_);
  or _75390_ (_25098_, _25097_, _25094_);
  nor _75391_ (_25100_, _25098_, _08654_);
  nor _75392_ (_25101_, _25100_, _25093_);
  nor _75393_ (_25102_, _25101_, _07154_);
  and _75394_ (_25103_, _07154_, \oc8051_golden_model_1.PC [0]);
  nor _75395_ (_25104_, _25103_, _06341_);
  not _75396_ (_25105_, _25104_);
  nor _75397_ (_25106_, _25105_, _25102_);
  not _75398_ (_25107_, _25106_);
  and _75399_ (_25108_, _25072_, _12534_);
  and _75400_ (_25109_, _12536_, \oc8051_golden_model_1.PC [0]);
  or _75401_ (_25111_, _25109_, _07151_);
  nor _75402_ (_25112_, _25111_, _25108_);
  nor _75403_ (_25113_, _25112_, _12542_);
  and _75404_ (_25114_, _25113_, _25107_);
  nor _75405_ (_25115_, _12541_, _05630_);
  nor _75406_ (_25116_, _25115_, _07611_);
  not _75407_ (_25117_, _25116_);
  nor _75408_ (_25118_, _25117_, _25114_);
  nor _75409_ (_25119_, _06872_, _06010_);
  and _75410_ (_25120_, _12560_, _12550_);
  not _75411_ (_25122_, _25120_);
  nor _75412_ (_25123_, _25122_, _25119_);
  not _75413_ (_25124_, _25123_);
  nor _75414_ (_25125_, _25124_, _25118_);
  nor _75415_ (_25126_, _25120_, _05630_);
  nor _75416_ (_25127_, _25126_, _12563_);
  not _75417_ (_25128_, _25127_);
  nor _75418_ (_25129_, _25128_, _25125_);
  or _75419_ (_25130_, _25129_, _12379_);
  nor _75420_ (_25131_, _25130_, _25082_);
  and _75421_ (_25133_, _12371_, _05630_);
  not _75422_ (_25134_, _25133_);
  nor _75423_ (_25135_, _25072_, _12371_);
  nor _75424_ (_25136_, _25135_, _12378_);
  and _75425_ (_25137_, _25136_, _25134_);
  nor _75426_ (_25138_, _25137_, _25131_);
  nor _75427_ (_25139_, _25138_, _06347_);
  nor _75428_ (_25140_, _25139_, _06480_);
  not _75429_ (_25141_, _25140_);
  nor _75430_ (_25142_, _25141_, _25081_);
  nor _75431_ (_25144_, _25142_, _25075_);
  nor _75432_ (_25145_, _25144_, _06371_);
  and _75433_ (_25146_, _12604_, _05630_);
  nor _75434_ (_25147_, _25072_, _12604_);
  or _75435_ (_25148_, _25147_, _25146_);
  and _75436_ (_25149_, _25148_, _06371_);
  or _75437_ (_25150_, _25149_, _25145_);
  and _75438_ (_25151_, _25150_, _12175_);
  and _75439_ (_25152_, _12174_, _05630_);
  or _75440_ (_25153_, _25152_, _25151_);
  and _75441_ (_25155_, _25153_, _06007_);
  or _75442_ (_25156_, _25155_, _12631_);
  nor _75443_ (_25157_, _25156_, _25068_);
  not _75444_ (_25158_, _06020_);
  nor _75445_ (_25159_, _12630_, _05630_);
  nor _75446_ (_25160_, _25159_, _25158_);
  not _75447_ (_25161_, _25160_);
  nor _75448_ (_25162_, _25161_, _25157_);
  nor _75449_ (_25163_, _06872_, _06020_);
  and _75450_ (_25164_, _12639_, _05984_);
  not _75451_ (_25166_, _25164_);
  nor _75452_ (_25167_, _25166_, _25163_);
  not _75453_ (_25168_, _25167_);
  nor _75454_ (_25169_, _25168_, _25162_);
  nor _75455_ (_25170_, _25164_, _05630_);
  nor _75456_ (_25171_, _25170_, _06254_);
  not _75457_ (_25172_, _25171_);
  nor _75458_ (_25173_, _25172_, _25169_);
  nor _75459_ (_25174_, _06872_, _05978_);
  nor _75460_ (_25175_, _06373_, _10094_);
  and _75461_ (_25177_, _25175_, _12172_);
  not _75462_ (_25178_, _25177_);
  nor _75463_ (_25179_, _25178_, _25174_);
  not _75464_ (_25180_, _25179_);
  nor _75465_ (_25181_, _25180_, _25173_);
  nor _75466_ (_25182_, _25177_, _05630_);
  nor _75467_ (_25183_, _25182_, _12668_);
  not _75468_ (_25184_, _25183_);
  nor _75469_ (_25185_, _25184_, _25181_);
  nor _75470_ (_25186_, _06872_, _05946_);
  or _75471_ (_25188_, _25186_, _12674_);
  or _75472_ (_25189_, _25188_, _25185_);
  or _75473_ (_25190_, _25096_, _12679_);
  and _75474_ (_25191_, _25190_, _25189_);
  and _75475_ (_25192_, _25191_, _06219_);
  or _75476_ (_25193_, _25192_, _25067_);
  and _75477_ (_25194_, _25193_, _12691_);
  and _75478_ (_25195_, _12690_, _06090_);
  or _75479_ (_25196_, _25195_, _25194_);
  and _75480_ (_25197_, _25196_, _05952_);
  nor _75481_ (_25199_, _06872_, _05952_);
  or _75482_ (_25200_, _25199_, _25197_);
  and _75483_ (_25201_, _25200_, _25064_);
  not _75484_ (_25202_, _25062_);
  nor _75485_ (_25203_, _25096_, _11342_);
  and _75486_ (_25204_, _11342_, _05630_);
  nor _75487_ (_25205_, _25204_, _25064_);
  not _75488_ (_25206_, _25205_);
  nor _75489_ (_25207_, _25206_, _25203_);
  nor _75490_ (_25208_, _25207_, _25202_);
  not _75491_ (_25210_, _25208_);
  nor _75492_ (_25211_, _25210_, _25201_);
  nor _75493_ (_25212_, _25211_, _25063_);
  and _75494_ (_25213_, _25212_, _05955_);
  nor _75495_ (_25214_, _06872_, _05955_);
  or _75496_ (_25215_, _25214_, _25213_);
  and _75497_ (_25216_, _25215_, _25061_);
  not _75498_ (_25217_, _25059_);
  nor _75499_ (_25218_, _11342_, _05630_);
  and _75500_ (_25219_, _25096_, _11342_);
  or _75501_ (_25221_, _25219_, _25218_);
  and _75502_ (_25222_, _25221_, _12755_);
  nor _75503_ (_25223_, _25222_, _25217_);
  not _75504_ (_25224_, _25223_);
  nor _75505_ (_25225_, _25224_, _25216_);
  nor _75506_ (_25226_, _25225_, _25060_);
  and _75507_ (_25227_, _25226_, _05961_);
  nor _75508_ (_25228_, _06872_, _05961_);
  or _75509_ (_25229_, _25228_, _25227_);
  and _75510_ (_25230_, _25229_, _12782_);
  not _75511_ (_25232_, _25057_);
  and _75512_ (_25233_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [0]);
  and _75513_ (_25234_, _25096_, _10558_);
  or _75514_ (_25235_, _25234_, _25233_);
  and _75515_ (_25236_, _25235_, _12776_);
  nor _75516_ (_25237_, _25236_, _25232_);
  not _75517_ (_25238_, _25237_);
  nor _75518_ (_25239_, _25238_, _25230_);
  nor _75519_ (_25240_, _25239_, _25058_);
  and _75520_ (_25241_, _25240_, _05966_);
  nor _75521_ (_25243_, _06872_, _05966_);
  or _75522_ (_25244_, _25243_, _25241_);
  and _75523_ (_25245_, _25244_, _25056_);
  and _75524_ (_25246_, _12154_, _11126_);
  not _75525_ (_25247_, _25246_);
  or _75526_ (_25248_, _25247_, _25245_);
  nor _75527_ (_25249_, _25248_, _25055_);
  nor _75528_ (_25250_, _25246_, _05630_);
  nor _75529_ (_25251_, _25250_, _06551_);
  not _75530_ (_25252_, _25251_);
  nor _75531_ (_25254_, _25252_, _25249_);
  and _75532_ (_25255_, _09392_, _06551_);
  or _75533_ (_25256_, _25255_, _25254_);
  and _75534_ (_25257_, _25256_, _05959_);
  nor _75535_ (_25258_, _06872_, _05959_);
  or _75536_ (_25259_, _25258_, _25257_);
  and _75537_ (_25260_, _25259_, _06558_);
  and _75538_ (_25261_, _25072_, _13004_);
  nor _75539_ (_25262_, _13004_, _05630_);
  or _75540_ (_25263_, _25262_, _06558_);
  or _75541_ (_25265_, _25263_, _25261_);
  and _75542_ (_25266_, _25265_, _25050_);
  not _75543_ (_25267_, _25266_);
  nor _75544_ (_25268_, _25267_, _25260_);
  nor _75545_ (_25269_, _25268_, _25051_);
  and _75546_ (_25270_, _25269_, _06282_);
  and _75547_ (_25271_, _09392_, _06281_);
  or _75548_ (_25272_, _25271_, _25270_);
  and _75549_ (_25273_, _25272_, _05964_);
  nor _75550_ (_25274_, _06872_, _05964_);
  nor _75551_ (_25276_, _25274_, _25273_);
  nor _75552_ (_25277_, _25276_, _06362_);
  not _75553_ (_25278_, _25048_);
  and _75554_ (_25279_, _13004_, \oc8051_golden_model_1.PC [0]);
  nor _75555_ (_25280_, _25071_, _13004_);
  nor _75556_ (_25281_, _25280_, _25279_);
  and _75557_ (_25282_, _25281_, _06362_);
  nor _75558_ (_25283_, _25282_, _25278_);
  not _75559_ (_25284_, _25283_);
  nor _75560_ (_25285_, _25284_, _25277_);
  nor _75561_ (_25287_, _25285_, _25049_);
  nor _75562_ (_25288_, _25287_, _07695_);
  and _75563_ (_25289_, _07695_, _06872_);
  nor _75564_ (_25290_, _25289_, _05927_);
  not _75565_ (_25291_, _25290_);
  or _75566_ (_25292_, _25291_, _25288_);
  not _75567_ (_25293_, _25046_);
  and _75568_ (_25294_, _25281_, _05927_);
  nor _75569_ (_25295_, _25294_, _25293_);
  and _75570_ (_25296_, _25295_, _25292_);
  or _75571_ (_25298_, _25296_, _25047_);
  nor _75572_ (_25299_, _06379_, _05939_);
  nand _75573_ (_25300_, _25299_, _25298_);
  not _75574_ (_25301_, _25299_);
  and _75575_ (_25302_, _25301_, _06872_);
  nor _75576_ (_25303_, _25302_, _13068_);
  and _75577_ (_25304_, _25303_, _25300_);
  and _75578_ (_25305_, _13068_, _05630_);
  or _75579_ (_25306_, _25305_, _25304_);
  or _75580_ (_25307_, _25306_, _01351_);
  or _75581_ (_25309_, _01347_, \oc8051_golden_model_1.PC [0]);
  and _75582_ (_25310_, _25309_, _42618_);
  and _75583_ (_43245_, _25310_, _25307_);
  and _75584_ (_25311_, _06278_, _05597_);
  nor _75585_ (_25312_, _13037_, _06111_);
  nor _75586_ (_25313_, _08568_, _06111_);
  nor _75587_ (_25314_, _12151_, _06111_);
  nor _75588_ (_25315_, _12154_, _06111_);
  nor _75589_ (_25316_, _12157_, _06111_);
  nor _75590_ (_25317_, _10979_, _06111_);
  nor _75591_ (_25318_, _12169_, _06111_);
  nor _75592_ (_25319_, _09030_, _05597_);
  nor _75593_ (_25320_, _12639_, _06111_);
  and _75594_ (_25321_, _12621_, _12616_);
  and _75595_ (_25322_, _25321_, _12620_);
  nor _75596_ (_25323_, _25322_, _05597_);
  and _75597_ (_25324_, _12174_, _06043_);
  and _75598_ (_25325_, _12371_, _06043_);
  nor _75599_ (_25326_, _12253_, _12251_);
  nor _75600_ (_25327_, _25326_, _12254_);
  not _75601_ (_25330_, _25327_);
  nor _75602_ (_25331_, _25330_, _12371_);
  or _75603_ (_25332_, _25331_, _25325_);
  nor _75604_ (_25333_, _25332_, _12378_);
  nor _75605_ (_25334_, _12560_, _06111_);
  and _75606_ (_25335_, _10759_, _06784_);
  nor _75607_ (_25336_, _25335_, _06111_);
  and _75608_ (_25337_, _10754_, _06043_);
  nor _75609_ (_25338_, _07038_, _07504_);
  and _75610_ (_25339_, _07486_, \oc8051_golden_model_1.PC [0]);
  nor _75611_ (_25341_, _25339_, _07141_);
  nor _75612_ (_25342_, _25341_, \oc8051_golden_model_1.PC [1]);
  and _75613_ (_25343_, _25341_, \oc8051_golden_model_1.PC [1]);
  nor _75614_ (_25344_, _25343_, _25342_);
  and _75615_ (_25345_, _25344_, _06782_);
  and _75616_ (_25346_, _06781_, _06043_);
  nor _75617_ (_25347_, _25346_, _25345_);
  and _75618_ (_25348_, _25347_, _07504_);
  nor _75619_ (_25349_, _25348_, _10754_);
  not _75620_ (_25350_, _25349_);
  nor _75621_ (_25352_, _25350_, _25338_);
  nor _75622_ (_25353_, _25352_, _25337_);
  not _75623_ (_25354_, _25335_);
  nor _75624_ (_25355_, _25354_, _25353_);
  or _75625_ (_25356_, _25355_, _10768_);
  nor _75626_ (_25357_, _25356_, _25336_);
  nor _75627_ (_25358_, _06043_, _06015_);
  nor _75628_ (_25359_, _25358_, _12387_);
  not _75629_ (_25360_, _25359_);
  nor _75630_ (_25361_, _25360_, _25357_);
  or _75631_ (_25363_, _12393_, \oc8051_golden_model_1.PC [1]);
  and _75632_ (_25364_, _12389_, _12391_);
  and _75633_ (_25365_, _08554_, _08553_);
  nand _75634_ (_25366_, _25365_, _25364_);
  nor _75635_ (_25367_, _12460_, _12458_);
  nor _75636_ (_25368_, _25367_, _12461_);
  nand _75637_ (_25369_, _25368_, _25366_);
  and _75638_ (_25370_, _25369_, _12387_);
  and _75639_ (_25371_, _25370_, _25363_);
  or _75640_ (_25372_, _25371_, _25361_);
  nand _75641_ (_25374_, _25372_, _07155_);
  and _75642_ (_25375_, _07154_, _06043_);
  nor _75643_ (_25376_, _25375_, _06341_);
  nand _75644_ (_25377_, _25376_, _25374_);
  or _75645_ (_25378_, _25327_, _12536_);
  or _75646_ (_25379_, _12534_, _06043_);
  and _75647_ (_25380_, _25379_, _06341_);
  nand _75648_ (_25381_, _25380_, _25378_);
  and _75649_ (_25382_, _25381_, _12541_);
  nand _75650_ (_25383_, _25382_, _25377_);
  nor _75651_ (_25385_, _12541_, _06111_);
  nor _75652_ (_25386_, _25385_, _06272_);
  nand _75653_ (_25387_, _25386_, _25383_);
  and _75654_ (_25388_, _06272_, _05597_);
  nor _75655_ (_25389_, _25388_, _07611_);
  nand _75656_ (_25390_, _25389_, _25387_);
  and _75657_ (_25391_, _07038_, _07611_);
  nor _75658_ (_25392_, _25391_, _06461_);
  nand _75659_ (_25393_, _25392_, _25390_);
  and _75660_ (_25394_, _06461_, _05597_);
  nor _75661_ (_25396_, _25394_, _12551_);
  nand _75662_ (_25397_, _25396_, _25393_);
  nor _75663_ (_25398_, _12550_, _06111_);
  nor _75664_ (_25399_, _25398_, _06464_);
  nand _75665_ (_25400_, _25399_, _25397_);
  not _75666_ (_25401_, _12560_);
  and _75667_ (_25402_, _06464_, _05597_);
  nor _75668_ (_25403_, _25402_, _25401_);
  and _75669_ (_25404_, _25403_, _25400_);
  or _75670_ (_25405_, _25404_, _25334_);
  nand _75671_ (_25407_, _25405_, _06269_);
  and _75672_ (_25408_, _06268_, \oc8051_golden_model_1.PC [1]);
  nor _75673_ (_25409_, _25408_, _12563_);
  and _75674_ (_25410_, _25409_, _25407_);
  nor _75675_ (_25411_, _07038_, _06013_);
  or _75676_ (_25412_, _25411_, _25410_);
  nand _75677_ (_25413_, _25412_, _07303_);
  and _75678_ (_25414_, _06267_, _05597_);
  nor _75679_ (_25415_, _25414_, _12379_);
  and _75680_ (_25416_, _25415_, _25413_);
  or _75681_ (_25418_, _25416_, _25333_);
  nand _75682_ (_25419_, _25418_, _12177_);
  or _75683_ (_25420_, _25330_, _12333_);
  or _75684_ (_25421_, _12335_, _06111_);
  and _75685_ (_25422_, _25421_, _06347_);
  nand _75686_ (_25423_, _25422_, _25420_);
  and _75687_ (_25424_, _25423_, _06774_);
  nand _75688_ (_25425_, _25424_, _25419_);
  and _75689_ (_25426_, _12587_, _06111_);
  nor _75690_ (_25427_, _25327_, _12587_);
  or _75691_ (_25429_, _25427_, _06774_);
  or _75692_ (_25430_, _25429_, _25426_);
  nand _75693_ (_25431_, _25430_, _25425_);
  nand _75694_ (_25432_, _25431_, _12176_);
  and _75695_ (_25433_, _12604_, _06043_);
  nor _75696_ (_25434_, _25330_, _12604_);
  or _75697_ (_25435_, _25434_, _25433_);
  and _75698_ (_25436_, _25435_, _06371_);
  nor _75699_ (_25437_, _25436_, _12174_);
  and _75700_ (_25438_, _25437_, _25432_);
  or _75701_ (_25440_, _25438_, _25324_);
  nand _75702_ (_25441_, _25440_, _06262_);
  and _75703_ (_25442_, _06261_, \oc8051_golden_model_1.PC [1]);
  nor _75704_ (_25443_, _25442_, _12613_);
  nand _75705_ (_25444_, _25443_, _25441_);
  not _75706_ (_25445_, _25322_);
  nor _75707_ (_25446_, _07038_, _06007_);
  nor _75708_ (_25447_, _25446_, _25445_);
  and _75709_ (_25448_, _25447_, _25444_);
  or _75710_ (_25449_, _25448_, _25323_);
  nand _75711_ (_25451_, _25449_, _12630_);
  nor _75712_ (_25452_, _12630_, _06111_);
  nor _75713_ (_25453_, _25452_, _06505_);
  nand _75714_ (_25454_, _25453_, _25451_);
  and _75715_ (_25455_, _06505_, _05597_);
  nor _75716_ (_25456_, _25455_, _25158_);
  nand _75717_ (_25457_, _25456_, _25454_);
  and _75718_ (_25458_, _07038_, _25158_);
  nor _75719_ (_25459_, _25458_, _06504_);
  nand _75720_ (_25460_, _25459_, _25457_);
  not _75721_ (_25462_, _17307_);
  and _75722_ (_25463_, _10588_, _14204_);
  and _75723_ (_25464_, _06504_, _05597_);
  not _75724_ (_25465_, _25464_);
  and _75725_ (_25466_, _25465_, _17311_);
  and _75726_ (_25467_, _25466_, _25463_);
  and _75727_ (_25468_, _25467_, _25462_);
  and _75728_ (_25469_, _25468_, _25460_);
  or _75729_ (_25470_, _25469_, _25320_);
  nand _75730_ (_25471_, _25470_, _12643_);
  nor _75731_ (_25473_, _12643_, _05597_);
  nor _75732_ (_25474_, _25473_, _10515_);
  nand _75733_ (_25475_, _25474_, _25471_);
  nor _75734_ (_25476_, _06043_, _05984_);
  nor _75735_ (_25477_, _25476_, _06257_);
  and _75736_ (_25478_, _25477_, _25475_);
  and _75737_ (_25479_, _06257_, \oc8051_golden_model_1.PC [1]);
  or _75738_ (_25480_, _25479_, _25478_);
  nand _75739_ (_25481_, _25480_, _05978_);
  and _75740_ (_25482_, _07038_, _06254_);
  nor _75741_ (_25484_, _25482_, _06373_);
  nand _75742_ (_25485_, _25484_, _25481_);
  and _75743_ (_25486_, _06373_, _06043_);
  nor _75744_ (_25487_, _25486_, _12659_);
  nand _75745_ (_25488_, _25487_, _25485_);
  nor _75746_ (_25489_, _07216_, _05597_);
  nor _75747_ (_25490_, _25489_, _10094_);
  nand _75748_ (_25491_, _25490_, _25488_);
  not _75749_ (_25492_, _12172_);
  nor _75750_ (_25493_, _06111_, _05982_);
  nor _75751_ (_25495_, _25493_, _25492_);
  nand _75752_ (_25496_, _25495_, _25491_);
  nor _75753_ (_25497_, _12172_, _06111_);
  nor _75754_ (_25498_, _25497_, _06323_);
  nand _75755_ (_25499_, _25498_, _25496_);
  and _75756_ (_25500_, _06323_, _05597_);
  nor _75757_ (_25501_, _25500_, _12668_);
  nand _75758_ (_25502_, _25501_, _25499_);
  and _75759_ (_25503_, _07038_, _12668_);
  nor _75760_ (_25504_, _25503_, _12674_);
  nand _75761_ (_25506_, _25504_, _25502_);
  and _75762_ (_25507_, _25368_, _12674_);
  nor _75763_ (_25508_, _25507_, _09031_);
  and _75764_ (_25509_, _25508_, _25506_);
  or _75765_ (_25510_, _25509_, _25319_);
  nand _75766_ (_25511_, _25510_, _06219_);
  and _75767_ (_25512_, _06218_, _06111_);
  nor _75768_ (_25513_, _25512_, _10929_);
  nand _75769_ (_25514_, _25513_, _25511_);
  and _75770_ (_25515_, _10929_, _05597_);
  nor _75771_ (_25517_, _25515_, _12690_);
  nand _75772_ (_25518_, _25517_, _25514_);
  and _75773_ (_25519_, _12690_, _06109_);
  nor _75774_ (_25520_, _25519_, _06322_);
  nand _75775_ (_25521_, _25520_, _25518_);
  and _75776_ (_25522_, _06322_, _05597_);
  nor _75777_ (_25523_, _25522_, _06217_);
  nand _75778_ (_25524_, _25523_, _25521_);
  and _75779_ (_25525_, _07038_, _06217_);
  nor _75780_ (_25526_, _25525_, _12733_);
  nand _75781_ (_25528_, _25526_, _25524_);
  and _75782_ (_25529_, _11342_, _05597_);
  and _75783_ (_25530_, _25368_, _12759_);
  or _75784_ (_25531_, _25530_, _25529_);
  and _75785_ (_25532_, _25531_, _12733_);
  nor _75786_ (_25533_, _25532_, _12737_);
  and _75787_ (_25534_, _25533_, _25528_);
  or _75788_ (_25535_, _25534_, _25318_);
  nand _75789_ (_25536_, _25535_, _12166_);
  nor _75790_ (_25537_, _12166_, _05597_);
  nor _75791_ (_25539_, _25537_, _06369_);
  nand _75792_ (_25540_, _25539_, _25536_);
  and _75793_ (_25541_, _06369_, _06043_);
  nor _75794_ (_25542_, _25541_, _06536_);
  and _75795_ (_25543_, _25542_, _25540_);
  and _75796_ (_25544_, _06536_, \oc8051_golden_model_1.PC [1]);
  or _75797_ (_25545_, _25544_, _25543_);
  nand _75798_ (_25546_, _25545_, _05955_);
  and _75799_ (_25547_, _07038_, _12750_);
  nor _75800_ (_25548_, _25547_, _12755_);
  nand _75801_ (_25550_, _25548_, _25546_);
  nor _75802_ (_25551_, _25368_, _12759_);
  nor _75803_ (_25552_, _11342_, _05597_);
  nor _75804_ (_25553_, _25552_, _25061_);
  not _75805_ (_25554_, _25553_);
  nor _75806_ (_25555_, _25554_, _25551_);
  nor _75807_ (_25556_, _25555_, _10980_);
  and _75808_ (_25557_, _25556_, _25550_);
  or _75809_ (_25558_, _25557_, _25317_);
  nand _75810_ (_25559_, _25558_, _12164_);
  nor _75811_ (_25561_, _12164_, _05597_);
  nor _75812_ (_25562_, _25561_, _06375_);
  nand _75813_ (_25563_, _25562_, _25559_);
  and _75814_ (_25564_, _06375_, _06043_);
  nor _75815_ (_25565_, _25564_, _06545_);
  and _75816_ (_25566_, _25565_, _25563_);
  and _75817_ (_25567_, _06545_, \oc8051_golden_model_1.PC [1]);
  or _75818_ (_25568_, _25567_, _25566_);
  nand _75819_ (_25569_, _25568_, _05961_);
  and _75820_ (_25570_, _07038_, _07233_);
  nor _75821_ (_25572_, _25570_, _12776_);
  nand _75822_ (_25573_, _25572_, _25569_);
  nor _75823_ (_25574_, _25368_, \oc8051_golden_model_1.PSW [7]);
  and _75824_ (_25575_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor _75825_ (_25576_, _25575_, _12782_);
  not _75826_ (_25577_, _25576_);
  nor _75827_ (_25578_, _25577_, _25574_);
  nor _75828_ (_25579_, _25578_, _17507_);
  and _75829_ (_25580_, _25579_, _25573_);
  nor _75830_ (_25581_, _25580_, _25316_);
  or _75831_ (_25583_, _25581_, _12160_);
  and _75832_ (_25584_, _12160_, _06043_);
  nor _75833_ (_25585_, _25584_, _11011_);
  nand _75834_ (_25586_, _25585_, _25583_);
  and _75835_ (_25587_, _11011_, _06111_);
  nor _75836_ (_25588_, _25587_, _11023_);
  nand _75837_ (_25589_, _25588_, _25586_);
  nor _75838_ (_25590_, _11022_, _05597_);
  nor _75839_ (_25591_, _25590_, _06366_);
  nand _75840_ (_25592_, _25591_, _25589_);
  and _75841_ (_25594_, _06366_, _06043_);
  nor _75842_ (_25595_, _25594_, _06528_);
  and _75843_ (_25596_, _25595_, _25592_);
  and _75844_ (_25597_, _06528_, \oc8051_golden_model_1.PC [1]);
  or _75845_ (_25598_, _25597_, _25596_);
  nand _75846_ (_25599_, _25598_, _05966_);
  and _75847_ (_25600_, _07038_, _12795_);
  nor _75848_ (_25601_, _25600_, _12800_);
  nand _75849_ (_25602_, _25601_, _25599_);
  nor _75850_ (_25603_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and _75851_ (_25605_, _25368_, \oc8051_golden_model_1.PSW [7]);
  or _75852_ (_25606_, _25605_, _25603_);
  and _75853_ (_25607_, _25606_, _12800_);
  nor _75854_ (_25608_, _25607_, _12804_);
  and _75855_ (_25609_, _25608_, _25602_);
  or _75856_ (_25610_, _25609_, _25315_);
  nand _75857_ (_25611_, _25610_, _12153_);
  nor _75858_ (_25612_, _12153_, _05597_);
  nor _75859_ (_25613_, _25612_, _11125_);
  nand _75860_ (_25614_, _25613_, _25611_);
  and _75861_ (_25616_, _11125_, _06111_);
  nor _75862_ (_25617_, _25616_, _06551_);
  and _75863_ (_25618_, _25617_, _25614_);
  and _75864_ (_25619_, _09347_, _06551_);
  or _75865_ (_25620_, _25619_, _25618_);
  nand _75866_ (_25621_, _25620_, _05959_);
  and _75867_ (_25622_, _07038_, _07253_);
  nor _75868_ (_25623_, _25622_, _06365_);
  nand _75869_ (_25624_, _25623_, _25621_);
  not _75870_ (_25625_, _12151_);
  and _75871_ (_25626_, _25330_, _13004_);
  not _75872_ (_25627_, _25626_);
  nor _75873_ (_25628_, _13004_, _06043_);
  nor _75874_ (_25629_, _25628_, _06558_);
  and _75875_ (_25630_, _25629_, _25627_);
  nor _75876_ (_25631_, _25630_, _25625_);
  and _75877_ (_25632_, _25631_, _25624_);
  or _75878_ (_25633_, _25632_, _25314_);
  nand _75879_ (_25634_, _25633_, _13012_);
  nor _75880_ (_25635_, _13012_, _05597_);
  nor _75881_ (_25638_, _25635_, _11284_);
  nand _75882_ (_25639_, _25638_, _25634_);
  and _75883_ (_25640_, _11284_, _06111_);
  nor _75884_ (_25641_, _25640_, _06281_);
  and _75885_ (_25642_, _25641_, _25639_);
  and _75886_ (_25643_, _09347_, _06281_);
  or _75887_ (_25644_, _25643_, _25642_);
  nand _75888_ (_25645_, _25644_, _05964_);
  not _75889_ (_25646_, _05964_);
  and _75890_ (_25647_, _07038_, _25646_);
  nor _75891_ (_25649_, _25647_, _06362_);
  nand _75892_ (_25650_, _25649_, _25645_);
  and _75893_ (_25651_, _13004_, _06111_);
  nor _75894_ (_25652_, _25327_, _13004_);
  nor _75895_ (_25653_, _25652_, _25651_);
  and _75896_ (_25654_, _25653_, _06362_);
  nor _75897_ (_25655_, _25654_, _15693_);
  and _75898_ (_25656_, _25655_, _25650_);
  nor _75899_ (_25657_, _25656_, _25313_);
  nor _75900_ (_25658_, _07482_, _06567_);
  or _75901_ (_25660_, _25658_, _25657_);
  and _75902_ (_25661_, _25658_, _06043_);
  nor _75903_ (_25662_, _25661_, _06568_);
  nand _75904_ (_25663_, _25662_, _25660_);
  and _75905_ (_25664_, _06568_, _05597_);
  nor _75906_ (_25665_, _25664_, _13038_);
  and _75907_ (_25666_, _25665_, _25663_);
  or _75908_ (_25667_, _25666_, _25312_);
  nand _75909_ (_25668_, _25667_, _07271_);
  and _75910_ (_25669_, _07695_, _07038_);
  nor _75911_ (_25671_, _25669_, _05927_);
  nand _75912_ (_25672_, _25671_, _25668_);
  and _75913_ (_25673_, _25653_, _05927_);
  nor _75914_ (_25674_, _25673_, _15111_);
  nand _75915_ (_25675_, _25674_, _25672_);
  nor _75916_ (_25676_, _15107_, _06111_);
  nor _75917_ (_25677_, _25676_, _15115_);
  nand _75918_ (_25678_, _25677_, _25675_);
  and _75919_ (_25679_, _15115_, _06111_);
  nor _75920_ (_25680_, _25679_, _07281_);
  nand _75921_ (_25682_, _25680_, _25678_);
  and _75922_ (_25683_, _07281_, _06043_);
  nor _75923_ (_25684_, _25683_, _06278_);
  and _75924_ (_25685_, _25684_, _25682_);
  or _75925_ (_25686_, _25685_, _25311_);
  nand _75926_ (_25687_, _25686_, _12141_);
  nor _75927_ (_25688_, _12141_, _06043_);
  nor _75928_ (_25689_, _25688_, _25301_);
  nand _75929_ (_25690_, _25689_, _25687_);
  and _75930_ (_25691_, _25301_, _07038_);
  nor _75931_ (_25693_, _25691_, _13068_);
  and _75932_ (_25694_, _25693_, _25690_);
  and _75933_ (_25695_, _13068_, _06111_);
  or _75934_ (_25696_, _25695_, _25694_);
  or _75935_ (_25697_, _25696_, _01351_);
  or _75936_ (_25698_, _01347_, \oc8051_golden_model_1.PC [1]);
  and _75937_ (_25699_, _25698_, _42618_);
  and _75938_ (_43246_, _25699_, _25697_);
  and _75939_ (_25700_, _13068_, _06040_);
  and _75940_ (_25701_, _06278_, _06079_);
  and _75941_ (_25703_, _06568_, _06079_);
  nor _75942_ (_25704_, _12151_, _06040_);
  nor _75943_ (_25705_, _12154_, _06040_);
  nor _75944_ (_25706_, _12162_, _06040_);
  nor _75945_ (_25707_, _10979_, _06040_);
  nor _75946_ (_25708_, _12169_, _06040_);
  and _75947_ (_25709_, _06332_, _06321_);
  nor _75948_ (_25710_, _06699_, _05951_);
  nand _75949_ (_25711_, _25710_, _06079_);
  and _75950_ (_25712_, _07214_, _06085_);
  nor _75951_ (_25714_, _25322_, _06079_);
  and _75952_ (_25715_, _12174_, _06074_);
  and _75953_ (_25716_, _12258_, _12255_);
  nor _75954_ (_25717_, _25716_, _12259_);
  not _75955_ (_25718_, _25717_);
  and _75956_ (_25719_, _25718_, _12335_);
  and _75957_ (_25720_, _12333_, _12248_);
  or _75958_ (_25721_, _25720_, _25719_);
  and _75959_ (_25722_, _25721_, _06347_);
  or _75960_ (_25723_, _12393_, _06085_);
  and _75961_ (_25725_, _12465_, _12462_);
  nor _75962_ (_25726_, _25725_, _12466_);
  nand _75963_ (_25727_, _25726_, _12393_);
  and _75964_ (_25728_, _25727_, _12387_);
  and _75965_ (_25729_, _25728_, _25723_);
  or _75966_ (_25730_, _07504_, _06697_);
  nor _75967_ (_25731_, _07486_, \oc8051_golden_model_1.PC [2]);
  or _75968_ (_25732_, _25731_, _07141_);
  nand _75969_ (_25733_, _07141_, _06079_);
  and _75970_ (_25734_, _25733_, _06782_);
  and _75971_ (_25736_, _25734_, _25732_);
  nor _75972_ (_25737_, _12513_, _06040_);
  or _75973_ (_25738_, _25737_, _06758_);
  or _75974_ (_25739_, _25738_, _25736_);
  and _75975_ (_25740_, _25739_, _12512_);
  and _75976_ (_25741_, _25740_, _25730_);
  nor _75977_ (_25742_, _12512_, _06040_);
  or _75978_ (_25743_, _25742_, _25741_);
  and _75979_ (_25744_, _25743_, _08654_);
  or _75980_ (_25745_, _25744_, _25729_);
  and _75981_ (_25747_, _25745_, _07155_);
  and _75982_ (_25748_, _07154_, _06074_);
  or _75983_ (_25749_, _25748_, _06341_);
  or _75984_ (_25750_, _25749_, _25747_);
  and _75985_ (_25751_, _25718_, _12534_);
  and _75986_ (_25752_, _12536_, _12248_);
  or _75987_ (_25753_, _25752_, _07151_);
  or _75988_ (_25754_, _25753_, _25751_);
  and _75989_ (_25755_, _25754_, _12541_);
  and _75990_ (_25756_, _25755_, _25750_);
  nor _75991_ (_25758_, _12541_, _06040_);
  or _75992_ (_25759_, _25758_, _06272_);
  or _75993_ (_25760_, _25759_, _25756_);
  nand _75994_ (_25761_, _06272_, _06079_);
  and _75995_ (_25762_, _25761_, _06010_);
  and _75996_ (_25763_, _25762_, _25760_);
  and _75997_ (_25764_, _06697_, _07611_);
  or _75998_ (_25765_, _25764_, _06461_);
  or _75999_ (_25766_, _25765_, _25763_);
  nand _76000_ (_25767_, _06461_, _06079_);
  and _76001_ (_25769_, _25767_, _12550_);
  and _76002_ (_25770_, _25769_, _25766_);
  nor _76003_ (_25771_, _12550_, _06040_);
  or _76004_ (_25772_, _25771_, _06464_);
  or _76005_ (_25773_, _25772_, _25770_);
  nand _76006_ (_25774_, _06464_, _06079_);
  and _76007_ (_25775_, _25774_, _12560_);
  and _76008_ (_25776_, _25775_, _25773_);
  nor _76009_ (_25777_, _12560_, _06040_);
  or _76010_ (_25778_, _25777_, _06268_);
  or _76011_ (_25780_, _25778_, _25776_);
  nand _76012_ (_25781_, _06268_, _06079_);
  and _76013_ (_25782_, _25781_, _06013_);
  and _76014_ (_25783_, _25782_, _25780_);
  and _76015_ (_25784_, _06697_, _12563_);
  or _76016_ (_25785_, _25784_, _06267_);
  or _76017_ (_25786_, _25785_, _25783_);
  nand _76018_ (_25787_, _06267_, _06079_);
  and _76019_ (_25788_, _25787_, _12378_);
  and _76020_ (_25789_, _25788_, _25786_);
  nand _76021_ (_25791_, _12371_, _12247_);
  or _76022_ (_25792_, _25718_, _12371_);
  and _76023_ (_25793_, _25792_, _12379_);
  and _76024_ (_25794_, _25793_, _25791_);
  or _76025_ (_25795_, _25794_, _25789_);
  and _76026_ (_25796_, _25795_, _12177_);
  or _76027_ (_25797_, _25796_, _25722_);
  and _76028_ (_25798_, _25797_, _06774_);
  or _76029_ (_25799_, _25718_, _12587_);
  nand _76030_ (_25800_, _12587_, _12247_);
  and _76031_ (_25802_, _25800_, _06480_);
  and _76032_ (_25803_, _25802_, _25799_);
  or _76033_ (_25804_, _25803_, _06371_);
  or _76034_ (_25805_, _25804_, _25798_);
  nor _76035_ (_25806_, _25717_, _12604_);
  and _76036_ (_25807_, _12604_, _12248_);
  or _76037_ (_25808_, _25807_, _12176_);
  or _76038_ (_25809_, _25808_, _25806_);
  and _76039_ (_25810_, _25809_, _12175_);
  and _76040_ (_25811_, _25810_, _25805_);
  or _76041_ (_25813_, _25811_, _25715_);
  and _76042_ (_25814_, _25813_, _06262_);
  and _76043_ (_25815_, _06261_, _06085_);
  or _76044_ (_25816_, _25815_, _12613_);
  or _76045_ (_25817_, _25816_, _25814_);
  or _76046_ (_25818_, _06697_, _06007_);
  and _76047_ (_25819_, _25818_, _25322_);
  and _76048_ (_25820_, _25819_, _25817_);
  or _76049_ (_25821_, _25820_, _25714_);
  and _76050_ (_25822_, _25821_, _12630_);
  nor _76051_ (_25824_, _12630_, _06040_);
  or _76052_ (_25825_, _25824_, _06505_);
  or _76053_ (_25826_, _25825_, _25822_);
  nand _76054_ (_25827_, _06505_, _06079_);
  and _76055_ (_25828_, _25827_, _06020_);
  and _76056_ (_25829_, _25828_, _25826_);
  and _76057_ (_25830_, _06697_, _25158_);
  or _76058_ (_25831_, _25830_, _06504_);
  or _76059_ (_25832_, _25831_, _25829_);
  nand _76060_ (_25833_, _06504_, _06079_);
  and _76061_ (_25835_, _25833_, _12639_);
  and _76062_ (_25836_, _25835_, _25832_);
  nor _76063_ (_25837_, _12639_, _06040_);
  or _76064_ (_25838_, _25837_, _25836_);
  and _76065_ (_25839_, _25838_, _12643_);
  nor _76066_ (_25840_, _12643_, _06079_);
  or _76067_ (_25841_, _25840_, _10515_);
  or _76068_ (_25842_, _25841_, _25839_);
  or _76069_ (_25843_, _06074_, _05984_);
  and _76070_ (_25844_, _25843_, _06258_);
  and _76071_ (_25846_, _25844_, _25842_);
  and _76072_ (_25847_, _06257_, _06085_);
  or _76073_ (_25848_, _25847_, _25846_);
  and _76074_ (_25849_, _25848_, _05978_);
  and _76075_ (_25850_, _06697_, _06254_);
  or _76076_ (_25851_, _25850_, _06373_);
  or _76077_ (_25852_, _25851_, _25849_);
  nor _76078_ (_25853_, _07461_, _06759_);
  nand _76079_ (_25854_, _12247_, _06373_);
  nand _76080_ (_25855_, _25854_, _25853_);
  nor _76081_ (_25857_, _25855_, _07455_);
  and _76082_ (_25858_, _25857_, _25852_);
  nor _76083_ (_25859_, _25858_, _25712_);
  nor _76084_ (_25860_, _07482_, _05945_);
  nor _76085_ (_25861_, _25860_, _25859_);
  and _76086_ (_25862_, _25860_, _06085_);
  or _76087_ (_25863_, _25862_, _10094_);
  or _76088_ (_25864_, _25863_, _25861_);
  or _76089_ (_25865_, _12248_, _05982_);
  and _76090_ (_25866_, _25865_, _12172_);
  and _76091_ (_25868_, _25866_, _25864_);
  nor _76092_ (_25869_, _12172_, _06040_);
  or _76093_ (_25870_, _25869_, _06323_);
  or _76094_ (_25871_, _25870_, _25868_);
  nand _76095_ (_25872_, _06323_, _06079_);
  and _76096_ (_25873_, _25872_, _05946_);
  and _76097_ (_25874_, _25873_, _25871_);
  and _76098_ (_25875_, _06697_, _12668_);
  or _76099_ (_25876_, _25875_, _25874_);
  and _76100_ (_25877_, _25876_, _12679_);
  nor _76101_ (_25879_, _25726_, _12679_);
  or _76102_ (_25880_, _25879_, _25710_);
  or _76103_ (_25881_, _25880_, _25877_);
  and _76104_ (_25882_, _25881_, _25711_);
  or _76105_ (_25883_, _25882_, _25709_);
  nand _76106_ (_25884_, _25709_, _06079_);
  and _76107_ (_25885_, _25884_, _09029_);
  and _76108_ (_25886_, _25885_, _25883_);
  nor _76109_ (_25887_, _09029_, _06079_);
  or _76110_ (_25888_, _25887_, _06218_);
  or _76111_ (_25890_, _25888_, _25886_);
  and _76112_ (_25891_, _12247_, _06218_);
  nor _76113_ (_25892_, _25891_, _10929_);
  and _76114_ (_25893_, _25892_, _25890_);
  and _76115_ (_25894_, _10929_, _06085_);
  or _76116_ (_25895_, _25894_, _25893_);
  nand _76117_ (_25896_, _25895_, _12691_);
  and _76118_ (_25897_, _12690_, _06071_);
  nor _76119_ (_25898_, _25897_, _06322_);
  nand _76120_ (_25899_, _25898_, _25896_);
  and _76121_ (_25901_, _06322_, _06079_);
  nor _76122_ (_25902_, _25901_, _06217_);
  nand _76123_ (_25903_, _25902_, _25899_);
  and _76124_ (_25904_, _06697_, _06217_);
  nor _76125_ (_25905_, _25904_, _12733_);
  nand _76126_ (_25906_, _25905_, _25903_);
  nor _76127_ (_25907_, _25726_, _11342_);
  and _76128_ (_25908_, _11342_, _06085_);
  nor _76129_ (_25909_, _25908_, _25064_);
  not _76130_ (_25910_, _25909_);
  nor _76131_ (_25912_, _25910_, _25907_);
  nor _76132_ (_25913_, _25912_, _12737_);
  and _76133_ (_25914_, _25913_, _25906_);
  or _76134_ (_25915_, _25914_, _25708_);
  nand _76135_ (_25916_, _25915_, _12166_);
  nor _76136_ (_25917_, _12166_, _06079_);
  nor _76137_ (_25918_, _25917_, _06369_);
  nand _76138_ (_25919_, _25918_, _25916_);
  and _76139_ (_25920_, _12247_, _06369_);
  nor _76140_ (_25921_, _25920_, _06536_);
  and _76141_ (_25923_, _25921_, _25919_);
  and _76142_ (_25924_, _06536_, _06085_);
  or _76143_ (_25925_, _25924_, _25923_);
  nand _76144_ (_25926_, _25925_, _05955_);
  and _76145_ (_25927_, _06697_, _12750_);
  nor _76146_ (_25928_, _25927_, _12755_);
  nand _76147_ (_25929_, _25928_, _25926_);
  nor _76148_ (_25930_, _11342_, _06085_);
  and _76149_ (_25931_, _25726_, _11342_);
  or _76150_ (_25932_, _25931_, _25930_);
  and _76151_ (_25934_, _25932_, _12755_);
  nor _76152_ (_25935_, _25934_, _10980_);
  and _76153_ (_25936_, _25935_, _25929_);
  or _76154_ (_25937_, _25936_, _25707_);
  nand _76155_ (_25938_, _25937_, _12164_);
  nor _76156_ (_25939_, _12164_, _06079_);
  nor _76157_ (_25940_, _25939_, _06375_);
  nand _76158_ (_25941_, _25940_, _25938_);
  and _76159_ (_25942_, _12247_, _06375_);
  nor _76160_ (_25943_, _25942_, _06545_);
  and _76161_ (_25945_, _25943_, _25941_);
  and _76162_ (_25946_, _06545_, _06085_);
  or _76163_ (_25947_, _25946_, _25945_);
  nand _76164_ (_25948_, _25947_, _05961_);
  and _76165_ (_25949_, _06697_, _07233_);
  nor _76166_ (_25950_, _25949_, _12776_);
  nand _76167_ (_25951_, _25950_, _25948_);
  nor _76168_ (_25952_, _25726_, \oc8051_golden_model_1.PSW [7]);
  nor _76169_ (_25953_, _06079_, _10558_);
  nor _76170_ (_25954_, _25953_, _12782_);
  not _76171_ (_25955_, _25954_);
  nor _76172_ (_25956_, _25955_, _25952_);
  nor _76173_ (_25957_, _25956_, _12780_);
  and _76174_ (_25958_, _25957_, _25951_);
  or _76175_ (_25959_, _25958_, _25706_);
  nand _76176_ (_25960_, _25959_, _11022_);
  nor _76177_ (_25961_, _11022_, _06079_);
  nor _76178_ (_25962_, _25961_, _06366_);
  nand _76179_ (_25963_, _25962_, _25960_);
  and _76180_ (_25964_, _12247_, _06366_);
  nor _76181_ (_25967_, _25964_, _06528_);
  and _76182_ (_25968_, _25967_, _25963_);
  and _76183_ (_25969_, _06528_, _06085_);
  or _76184_ (_25970_, _25969_, _25968_);
  nand _76185_ (_25971_, _25970_, _05966_);
  and _76186_ (_25972_, _06697_, _12795_);
  nor _76187_ (_25973_, _25972_, _12800_);
  nand _76188_ (_25974_, _25973_, _25971_);
  nor _76189_ (_25975_, _25726_, _10558_);
  nor _76190_ (_25976_, _06079_, \oc8051_golden_model_1.PSW [7]);
  nor _76191_ (_25978_, _25976_, _25056_);
  not _76192_ (_25979_, _25978_);
  nor _76193_ (_25980_, _25979_, _25975_);
  nor _76194_ (_25981_, _25980_, _12804_);
  and _76195_ (_25982_, _25981_, _25974_);
  or _76196_ (_25983_, _25982_, _25705_);
  nand _76197_ (_25984_, _25983_, _12153_);
  nor _76198_ (_25985_, _12153_, _06079_);
  nor _76199_ (_25986_, _25985_, _11125_);
  nand _76200_ (_25987_, _25986_, _25984_);
  and _76201_ (_25989_, _11125_, _06040_);
  nor _76202_ (_25990_, _25989_, _06551_);
  and _76203_ (_25991_, _25990_, _25987_);
  and _76204_ (_25992_, _09302_, _06551_);
  or _76205_ (_25993_, _25992_, _25991_);
  nand _76206_ (_25994_, _25993_, _05959_);
  and _76207_ (_25995_, _06697_, _07253_);
  nor _76208_ (_25996_, _25995_, _06365_);
  nand _76209_ (_25997_, _25996_, _25994_);
  nor _76210_ (_25998_, _12247_, _13004_);
  and _76211_ (_26000_, _25718_, _13004_);
  or _76212_ (_26001_, _26000_, _06558_);
  or _76213_ (_26002_, _26001_, _25998_);
  and _76214_ (_26003_, _26002_, _12151_);
  and _76215_ (_26004_, _26003_, _25997_);
  or _76216_ (_26005_, _26004_, _25704_);
  nand _76217_ (_26006_, _26005_, _13012_);
  nor _76218_ (_26007_, _13012_, _06079_);
  nor _76219_ (_26008_, _26007_, _11284_);
  nand _76220_ (_26009_, _26008_, _26006_);
  and _76221_ (_26011_, _11284_, _06040_);
  nor _76222_ (_26012_, _26011_, _06281_);
  and _76223_ (_26013_, _26012_, _26009_);
  and _76224_ (_26014_, _09302_, _06281_);
  or _76225_ (_26015_, _26014_, _26013_);
  nand _76226_ (_26016_, _26015_, _05964_);
  and _76227_ (_26017_, _06697_, _25646_);
  nor _76228_ (_26018_, _26017_, _06362_);
  nand _76229_ (_26019_, _26018_, _26016_);
  nor _76230_ (_26020_, _25717_, _13004_);
  and _76231_ (_26022_, _12248_, _13004_);
  nor _76232_ (_26023_, _26022_, _26020_);
  and _76233_ (_26024_, _26023_, _06362_);
  nor _76234_ (_26025_, _26024_, _13031_);
  nand _76235_ (_26026_, _26025_, _26019_);
  nor _76236_ (_26027_, _13030_, _06040_);
  nor _76237_ (_26028_, _26027_, _06568_);
  and _76238_ (_26029_, _26028_, _26026_);
  or _76239_ (_26030_, _26029_, _25703_);
  nand _76240_ (_26031_, _26030_, _13037_);
  nor _76241_ (_26033_, _13037_, _06074_);
  nor _76242_ (_26034_, _26033_, _07695_);
  nand _76243_ (_26035_, _26034_, _26031_);
  and _76244_ (_26036_, _07695_, _06697_);
  nor _76245_ (_26037_, _26036_, _05927_);
  nand _76246_ (_26038_, _26037_, _26035_);
  and _76247_ (_26039_, _26023_, _05927_);
  nor _76248_ (_26040_, _26039_, _13053_);
  nand _76249_ (_26041_, _26040_, _26038_);
  nor _76250_ (_26042_, _13052_, _06040_);
  nor _76251_ (_26044_, _26042_, _06278_);
  and _76252_ (_26045_, _26044_, _26041_);
  or _76253_ (_26046_, _26045_, _25701_);
  nand _76254_ (_26047_, _26046_, _12141_);
  nor _76255_ (_26048_, _12141_, _06074_);
  nor _76256_ (_26049_, _26048_, _25301_);
  nand _76257_ (_26050_, _26049_, _26047_);
  and _76258_ (_26051_, _25301_, _06697_);
  nor _76259_ (_26052_, _26051_, _13068_);
  and _76260_ (_26053_, _26052_, _26050_);
  or _76261_ (_26055_, _26053_, _25700_);
  or _76262_ (_26056_, _26055_, _01351_);
  or _76263_ (_26057_, _01347_, \oc8051_golden_model_1.PC [2]);
  and _76264_ (_26058_, _26057_, _42618_);
  and _76265_ (_43247_, _26058_, _26056_);
  and _76266_ (_26059_, _13068_, _06028_);
  and _76267_ (_26060_, _06278_, _05932_);
  and _76268_ (_26061_, _06568_, _05932_);
  nor _76269_ (_26062_, _12151_, _06028_);
  nor _76270_ (_26063_, _12154_, _06028_);
  nor _76271_ (_26065_, _12162_, _06028_);
  nor _76272_ (_26066_, _10979_, _06028_);
  nor _76273_ (_26067_, _12169_, _06028_);
  nor _76274_ (_26068_, _09030_, _05932_);
  nor _76275_ (_26069_, _25322_, _05932_);
  and _76276_ (_26070_, _12174_, _06027_);
  or _76277_ (_26071_, _12534_, _12242_);
  or _76278_ (_26072_, _12245_, _12244_);
  and _76279_ (_26073_, _26072_, _12260_);
  nor _76280_ (_26074_, _26072_, _12260_);
  nor _76281_ (_26076_, _26074_, _26073_);
  or _76282_ (_26077_, _26076_, _12536_);
  and _76283_ (_26078_, _26077_, _26071_);
  or _76284_ (_26079_, _26078_, _07151_);
  and _76285_ (_26080_, _12507_, _05932_);
  or _76286_ (_26081_, _12455_, _12454_);
  and _76287_ (_26082_, _26081_, _12467_);
  nor _76288_ (_26083_, _26081_, _12467_);
  nor _76289_ (_26084_, _26083_, _26082_);
  and _76290_ (_26085_, _26084_, _12393_);
  nor _76291_ (_26087_, _26085_, _26080_);
  nand _76292_ (_26088_, _26087_, _12387_);
  nor _76293_ (_26089_, _12512_, _06028_);
  nor _76294_ (_26090_, _07486_, \oc8051_golden_model_1.PC [3]);
  nor _76295_ (_26091_, _26090_, _07141_);
  and _76296_ (_26092_, _07141_, _05932_);
  nor _76297_ (_26093_, _26092_, _06781_);
  not _76298_ (_26094_, _26093_);
  nor _76299_ (_26095_, _26094_, _26091_);
  not _76300_ (_26096_, _26095_);
  nor _76301_ (_26098_, _12513_, _06028_);
  nor _76302_ (_26099_, _26098_, _06758_);
  and _76303_ (_26100_, _26099_, _26096_);
  nor _76304_ (_26101_, _07504_, _06452_);
  or _76305_ (_26102_, _26101_, _12516_);
  nor _76306_ (_26103_, _26102_, _26100_);
  nor _76307_ (_26104_, _26103_, _26089_);
  nor _76308_ (_26105_, _26104_, _12387_);
  nor _76309_ (_26106_, _26105_, _07154_);
  and _76310_ (_26107_, _26106_, _26088_);
  and _76311_ (_26109_, _07154_, _06028_);
  or _76312_ (_26110_, _26109_, _06341_);
  or _76313_ (_26111_, _26110_, _26107_);
  nand _76314_ (_26112_, _26111_, _26079_);
  nand _76315_ (_26113_, _26112_, _12541_);
  nor _76316_ (_26114_, _12541_, _06028_);
  nor _76317_ (_26115_, _26114_, _06272_);
  nand _76318_ (_26116_, _26115_, _26113_);
  and _76319_ (_26117_, _06272_, _05932_);
  nor _76320_ (_26118_, _26117_, _07611_);
  nand _76321_ (_26120_, _26118_, _26116_);
  and _76322_ (_26121_, _06452_, _07611_);
  nor _76323_ (_26122_, _26121_, _06461_);
  nand _76324_ (_26123_, _26122_, _26120_);
  and _76325_ (_26124_, _06461_, _05932_);
  nor _76326_ (_26125_, _26124_, _12551_);
  nand _76327_ (_26126_, _26125_, _26123_);
  nor _76328_ (_26127_, _12550_, _06028_);
  nor _76329_ (_26128_, _26127_, _06464_);
  nand _76330_ (_26129_, _26128_, _26126_);
  and _76331_ (_26131_, _06464_, _05932_);
  nor _76332_ (_26132_, _26131_, _25401_);
  nand _76333_ (_26133_, _26132_, _26129_);
  nor _76334_ (_26134_, _12560_, _06028_);
  nor _76335_ (_26135_, _26134_, _06268_);
  nand _76336_ (_26136_, _26135_, _26133_);
  and _76337_ (_26137_, _06268_, _05932_);
  nor _76338_ (_26138_, _26137_, _12563_);
  nand _76339_ (_26139_, _26138_, _26136_);
  and _76340_ (_26140_, _06452_, _12563_);
  nor _76341_ (_26142_, _26140_, _06267_);
  nand _76342_ (_26143_, _26142_, _26139_);
  and _76343_ (_26144_, _06267_, _05932_);
  nor _76344_ (_26145_, _26144_, _12379_);
  nand _76345_ (_26146_, _26145_, _26143_);
  and _76346_ (_26147_, _12371_, _12242_);
  not _76347_ (_26148_, _26076_);
  nor _76348_ (_26149_, _26148_, _12371_);
  or _76349_ (_26150_, _26149_, _12378_);
  nor _76350_ (_26151_, _26150_, _26147_);
  nor _76351_ (_26153_, _26151_, _06347_);
  nand _76352_ (_26154_, _26153_, _26146_);
  or _76353_ (_26155_, _26148_, _12333_);
  or _76354_ (_26156_, _12335_, _12243_);
  nand _76355_ (_26157_, _26156_, _26155_);
  nand _76356_ (_26158_, _26157_, _06347_);
  and _76357_ (_26159_, _26158_, _06774_);
  nand _76358_ (_26160_, _26159_, _26154_);
  and _76359_ (_26161_, _12587_, _12242_);
  not _76360_ (_26162_, _26161_);
  nor _76361_ (_26164_, _26148_, _12587_);
  nor _76362_ (_26165_, _26164_, _06774_);
  and _76363_ (_26166_, _26165_, _26162_);
  nor _76364_ (_26167_, _26166_, _06371_);
  nand _76365_ (_26168_, _26167_, _26160_);
  and _76366_ (_26169_, _12604_, _12243_);
  nor _76367_ (_26170_, _26076_, _12604_);
  or _76368_ (_26171_, _26170_, _12176_);
  nor _76369_ (_26172_, _26171_, _26169_);
  nor _76370_ (_26173_, _26172_, _12174_);
  and _76371_ (_26175_, _26173_, _26168_);
  or _76372_ (_26176_, _26175_, _26070_);
  nand _76373_ (_26177_, _26176_, _06262_);
  and _76374_ (_26178_, _06261_, _06033_);
  nor _76375_ (_26179_, _26178_, _12613_);
  nand _76376_ (_26180_, _26179_, _26177_);
  nor _76377_ (_26181_, _06452_, _06007_);
  nor _76378_ (_26182_, _26181_, _25445_);
  and _76379_ (_26183_, _26182_, _26180_);
  or _76380_ (_26184_, _26183_, _26069_);
  nand _76381_ (_26186_, _26184_, _12630_);
  nor _76382_ (_26187_, _12630_, _06028_);
  nor _76383_ (_26188_, _26187_, _06505_);
  nand _76384_ (_26189_, _26188_, _26186_);
  and _76385_ (_26190_, _06505_, _05932_);
  nor _76386_ (_26191_, _26190_, _25158_);
  nand _76387_ (_26192_, _26191_, _26189_);
  and _76388_ (_26193_, _06452_, _25158_);
  nor _76389_ (_26194_, _26193_, _06504_);
  nand _76390_ (_26195_, _26194_, _26192_);
  not _76391_ (_26197_, _12639_);
  and _76392_ (_26198_, _06504_, _05932_);
  nor _76393_ (_26199_, _26198_, _26197_);
  and _76394_ (_26200_, _26199_, _26195_);
  nor _76395_ (_26201_, _12639_, _06028_);
  or _76396_ (_26202_, _26201_, _26200_);
  nand _76397_ (_26203_, _26202_, _12643_);
  nor _76398_ (_26204_, _12643_, _05932_);
  nor _76399_ (_26205_, _26204_, _10515_);
  nand _76400_ (_26206_, _26205_, _26203_);
  nor _76401_ (_26208_, _05984_, _06027_);
  nor _76402_ (_26209_, _26208_, _06257_);
  and _76403_ (_26210_, _26209_, _26206_);
  and _76404_ (_26211_, _06257_, _06033_);
  or _76405_ (_26212_, _26211_, _26210_);
  nand _76406_ (_26213_, _26212_, _05978_);
  and _76407_ (_26214_, _06452_, _06254_);
  nor _76408_ (_26215_, _26214_, _06373_);
  nand _76409_ (_26216_, _26215_, _26213_);
  and _76410_ (_26217_, _12242_, _06373_);
  nor _76411_ (_26219_, _26217_, _12659_);
  nand _76412_ (_26220_, _26219_, _26216_);
  nor _76413_ (_26221_, _07216_, _05932_);
  nor _76414_ (_26222_, _26221_, _10094_);
  nand _76415_ (_26223_, _26222_, _26220_);
  nor _76416_ (_26224_, _12243_, _05982_);
  nor _76417_ (_26225_, _26224_, _25492_);
  nand _76418_ (_26226_, _26225_, _26223_);
  nor _76419_ (_26227_, _12172_, _06028_);
  nor _76420_ (_26228_, _26227_, _06323_);
  nand _76421_ (_26230_, _26228_, _26226_);
  and _76422_ (_26231_, _06323_, _05932_);
  nor _76423_ (_26232_, _26231_, _12668_);
  nand _76424_ (_26233_, _26232_, _26230_);
  and _76425_ (_26234_, _06452_, _12668_);
  nor _76426_ (_26235_, _26234_, _12674_);
  nand _76427_ (_26236_, _26235_, _26233_);
  and _76428_ (_26237_, _26084_, _12674_);
  nor _76429_ (_26238_, _26237_, _09031_);
  and _76430_ (_26239_, _26238_, _26236_);
  or _76431_ (_26241_, _26239_, _26068_);
  nand _76432_ (_26242_, _26241_, _06219_);
  and _76433_ (_26243_, _12243_, _06218_);
  nor _76434_ (_26244_, _26243_, _10929_);
  nand _76435_ (_26245_, _26244_, _26242_);
  and _76436_ (_26246_, _10929_, _05932_);
  nor _76437_ (_26247_, _26246_, _12690_);
  nand _76438_ (_26248_, _26247_, _26245_);
  and _76439_ (_26249_, _12690_, _06004_);
  nor _76440_ (_26250_, _26249_, _06322_);
  and _76441_ (_26252_, _26250_, _26248_);
  and _76442_ (_26253_, _06322_, _05932_);
  or _76443_ (_26254_, _26253_, _06217_);
  or _76444_ (_26255_, _26254_, _26252_);
  and _76445_ (_26256_, _06452_, _06217_);
  nor _76446_ (_26257_, _26256_, _12733_);
  nand _76447_ (_26258_, _26257_, _26255_);
  and _76448_ (_26259_, _11342_, _05932_);
  and _76449_ (_26260_, _26084_, _12759_);
  or _76450_ (_26261_, _26260_, _26259_);
  and _76451_ (_26263_, _26261_, _12733_);
  nor _76452_ (_26264_, _26263_, _12737_);
  and _76453_ (_26265_, _26264_, _26258_);
  or _76454_ (_26266_, _26265_, _26067_);
  nand _76455_ (_26267_, _26266_, _12166_);
  nor _76456_ (_26268_, _12166_, _05932_);
  nor _76457_ (_26269_, _26268_, _06369_);
  and _76458_ (_26270_, _26269_, _26267_);
  and _76459_ (_26271_, _12242_, _06369_);
  or _76460_ (_26272_, _26271_, _06536_);
  nor _76461_ (_26274_, _26272_, _26270_);
  and _76462_ (_26275_, _06536_, _06033_);
  or _76463_ (_26276_, _26275_, _26274_);
  nand _76464_ (_26277_, _26276_, _05955_);
  and _76465_ (_26278_, _06452_, _12750_);
  nor _76466_ (_26279_, _26278_, _12755_);
  nand _76467_ (_26280_, _26279_, _26277_);
  nor _76468_ (_26281_, _11342_, _06033_);
  and _76469_ (_26282_, _26084_, _11342_);
  or _76470_ (_26283_, _26282_, _26281_);
  and _76471_ (_26285_, _26283_, _12755_);
  nor _76472_ (_26286_, _26285_, _10980_);
  and _76473_ (_26287_, _26286_, _26280_);
  or _76474_ (_26288_, _26287_, _26066_);
  nand _76475_ (_26289_, _26288_, _12164_);
  nor _76476_ (_26290_, _12164_, _05932_);
  nor _76477_ (_26291_, _26290_, _06375_);
  nand _76478_ (_26292_, _26291_, _26289_);
  and _76479_ (_26293_, _12242_, _06375_);
  nor _76480_ (_26294_, _26293_, _06545_);
  and _76481_ (_26296_, _26294_, _26292_);
  and _76482_ (_26297_, _06545_, _06033_);
  or _76483_ (_26298_, _26297_, _26296_);
  nand _76484_ (_26299_, _26298_, _05961_);
  and _76485_ (_26300_, _06452_, _07233_);
  nor _76486_ (_26301_, _26300_, _12776_);
  nand _76487_ (_26302_, _26301_, _26299_);
  nor _76488_ (_26303_, _26084_, \oc8051_golden_model_1.PSW [7]);
  nor _76489_ (_26304_, _05932_, _10558_);
  nor _76490_ (_26305_, _26304_, _12782_);
  not _76491_ (_26307_, _26305_);
  nor _76492_ (_26308_, _26307_, _26303_);
  nor _76493_ (_26309_, _26308_, _12780_);
  and _76494_ (_26310_, _26309_, _26302_);
  or _76495_ (_26311_, _26310_, _26065_);
  nand _76496_ (_26312_, _26311_, _11022_);
  nor _76497_ (_26313_, _11022_, _05932_);
  nor _76498_ (_26314_, _26313_, _06366_);
  and _76499_ (_26315_, _26314_, _26312_);
  and _76500_ (_26316_, _12242_, _06366_);
  or _76501_ (_26318_, _26316_, _06528_);
  nor _76502_ (_26319_, _26318_, _26315_);
  and _76503_ (_26320_, _06528_, _06033_);
  or _76504_ (_26321_, _26320_, _26319_);
  nand _76505_ (_26322_, _26321_, _05966_);
  and _76506_ (_26323_, _06452_, _12795_);
  nor _76507_ (_26324_, _26323_, _12800_);
  nand _76508_ (_26325_, _26324_, _26322_);
  and _76509_ (_26326_, _05932_, _10558_);
  and _76510_ (_26327_, _26084_, \oc8051_golden_model_1.PSW [7]);
  or _76511_ (_26329_, _26327_, _26326_);
  and _76512_ (_26330_, _26329_, _12800_);
  nor _76513_ (_26331_, _26330_, _12804_);
  and _76514_ (_26332_, _26331_, _26325_);
  or _76515_ (_26333_, _26332_, _26063_);
  nand _76516_ (_26334_, _26333_, _12153_);
  nor _76517_ (_26335_, _12153_, _05932_);
  nor _76518_ (_26336_, _26335_, _11125_);
  nand _76519_ (_26337_, _26336_, _26334_);
  and _76520_ (_26338_, _11125_, _06028_);
  nor _76521_ (_26340_, _26338_, _06551_);
  and _76522_ (_26341_, _26340_, _26337_);
  and _76523_ (_26342_, _09257_, _06551_);
  or _76524_ (_26343_, _26342_, _26341_);
  nand _76525_ (_26344_, _26343_, _05959_);
  and _76526_ (_26345_, _06452_, _07253_);
  nor _76527_ (_26346_, _26345_, _06365_);
  nand _76528_ (_26347_, _26346_, _26344_);
  and _76529_ (_26348_, _26148_, _13004_);
  nor _76530_ (_26349_, _12242_, _13004_);
  or _76531_ (_26351_, _26349_, _06558_);
  or _76532_ (_26352_, _26351_, _26348_);
  and _76533_ (_26353_, _26352_, _12151_);
  and _76534_ (_26354_, _26353_, _26347_);
  or _76535_ (_26355_, _26354_, _26062_);
  nand _76536_ (_26356_, _26355_, _13012_);
  nor _76537_ (_26357_, _13012_, _05932_);
  nor _76538_ (_26358_, _26357_, _11284_);
  nand _76539_ (_26359_, _26358_, _26356_);
  and _76540_ (_26360_, _11284_, _06028_);
  nor _76541_ (_26362_, _26360_, _06281_);
  and _76542_ (_26363_, _26362_, _26359_);
  and _76543_ (_26364_, _09257_, _06281_);
  or _76544_ (_26365_, _26364_, _26363_);
  nand _76545_ (_26366_, _26365_, _05964_);
  and _76546_ (_26367_, _06452_, _25646_);
  nor _76547_ (_26368_, _26367_, _06362_);
  nand _76548_ (_26369_, _26368_, _26366_);
  nor _76549_ (_26370_, _26076_, _13004_);
  and _76550_ (_26371_, _12243_, _13004_);
  nor _76551_ (_26373_, _26371_, _26370_);
  and _76552_ (_26374_, _26373_, _06362_);
  nor _76553_ (_26375_, _26374_, _13031_);
  nand _76554_ (_26376_, _26375_, _26369_);
  nor _76555_ (_26377_, _13030_, _06028_);
  nor _76556_ (_26378_, _26377_, _06568_);
  and _76557_ (_26379_, _26378_, _26376_);
  or _76558_ (_26380_, _26379_, _26061_);
  nand _76559_ (_26381_, _26380_, _13037_);
  nor _76560_ (_26382_, _13037_, _06027_);
  nor _76561_ (_26384_, _26382_, _07695_);
  nand _76562_ (_26385_, _26384_, _26381_);
  and _76563_ (_26386_, _07695_, _06452_);
  nor _76564_ (_26387_, _26386_, _05927_);
  nand _76565_ (_26388_, _26387_, _26385_);
  and _76566_ (_26389_, _26373_, _05927_);
  nor _76567_ (_26390_, _26389_, _13053_);
  nand _76568_ (_26391_, _26390_, _26388_);
  nor _76569_ (_26392_, _13052_, _06028_);
  nor _76570_ (_26393_, _26392_, _06278_);
  and _76571_ (_26395_, _26393_, _26391_);
  or _76572_ (_26396_, _26395_, _26060_);
  nand _76573_ (_26397_, _26396_, _12141_);
  nor _76574_ (_26398_, _12141_, _06027_);
  nor _76575_ (_26399_, _26398_, _25301_);
  nand _76576_ (_26400_, _26399_, _26397_);
  and _76577_ (_26401_, _25301_, _06452_);
  nor _76578_ (_26402_, _26401_, _13068_);
  and _76579_ (_26403_, _26402_, _26400_);
  or _76580_ (_26404_, _26403_, _26059_);
  or _76581_ (_26406_, _26404_, _01351_);
  or _76582_ (_26407_, _01347_, \oc8051_golden_model_1.PC [3]);
  and _76583_ (_26408_, _26407_, _42618_);
  and _76584_ (_43249_, _26408_, _26406_);
  and _76585_ (_26409_, _08892_, _07695_);
  and _76586_ (_26410_, _12451_, _10558_);
  and _76587_ (_26411_, _12472_, _12469_);
  nor _76588_ (_26412_, _26411_, _12473_);
  and _76589_ (_26413_, _26412_, \oc8051_golden_model_1.PSW [7]);
  or _76590_ (_26414_, _26413_, _26410_);
  and _76591_ (_26416_, _26414_, _12800_);
  nor _76592_ (_26417_, _12452_, _11342_);
  and _76593_ (_26418_, _26412_, _11342_);
  or _76594_ (_26419_, _26418_, _26417_);
  and _76595_ (_26420_, _26419_, _12755_);
  and _76596_ (_26421_, _12451_, _11342_);
  and _76597_ (_26422_, _26412_, _12759_);
  or _76598_ (_26423_, _26422_, _26421_);
  and _76599_ (_26424_, _26423_, _12733_);
  nor _76600_ (_26425_, _12451_, _09030_);
  and _76601_ (_26427_, _12452_, _06257_);
  not _76602_ (_26428_, \oc8051_golden_model_1.PC [4]);
  nor _76603_ (_26429_, _05616_, _26428_);
  and _76604_ (_26430_, _05616_, _26428_);
  nor _76605_ (_26431_, _26430_, _26429_);
  not _76606_ (_26432_, _26431_);
  and _76607_ (_26433_, _26432_, _12174_);
  and _76608_ (_26434_, _12452_, _06268_);
  nor _76609_ (_26435_, _26431_, _12550_);
  nand _76610_ (_26436_, _26412_, _25366_);
  or _76611_ (_26437_, _12393_, _12452_);
  and _76612_ (_26438_, _26437_, _26436_);
  and _76613_ (_26439_, _26438_, _12387_);
  nor _76614_ (_26440_, _26432_, _12512_);
  and _76615_ (_26441_, _08892_, _06758_);
  or _76616_ (_26442_, _07486_, _26428_);
  and _76617_ (_26443_, _26442_, _07142_);
  and _76618_ (_26444_, _12452_, _07141_);
  or _76619_ (_26445_, _26444_, _06781_);
  or _76620_ (_26446_, _26445_, _26443_);
  or _76621_ (_26448_, _26432_, _12513_);
  and _76622_ (_26449_, _26448_, _07504_);
  and _76623_ (_26450_, _26449_, _26446_);
  nor _76624_ (_26451_, _26450_, _12516_);
  not _76625_ (_26452_, _26451_);
  nor _76626_ (_26453_, _26452_, _26441_);
  or _76627_ (_26454_, _26453_, _12387_);
  nor _76628_ (_26455_, _26454_, _26440_);
  or _76629_ (_26456_, _26455_, _26439_);
  nand _76630_ (_26457_, _26456_, _07155_);
  and _76631_ (_26459_, _26432_, _07154_);
  nor _76632_ (_26460_, _26459_, _06341_);
  nand _76633_ (_26461_, _26460_, _26457_);
  or _76634_ (_26462_, _12534_, _12238_);
  and _76635_ (_26463_, _12265_, _12262_);
  nor _76636_ (_26464_, _26463_, _12266_);
  or _76637_ (_26465_, _26464_, _12536_);
  and _76638_ (_26466_, _26465_, _06341_);
  nand _76639_ (_26467_, _26466_, _26462_);
  and _76640_ (_26468_, _26467_, _12541_);
  and _76641_ (_26469_, _26468_, _26461_);
  nor _76642_ (_26470_, _26431_, _12541_);
  or _76643_ (_26471_, _26470_, _26469_);
  nand _76644_ (_26472_, _26471_, _06273_);
  and _76645_ (_26473_, _12452_, _06272_);
  nor _76646_ (_26474_, _26473_, _07611_);
  and _76647_ (_26475_, _26474_, _26472_);
  nor _76648_ (_26476_, _08892_, _06010_);
  or _76649_ (_26477_, _26476_, _06461_);
  nor _76650_ (_26478_, _26477_, _26475_);
  and _76651_ (_26479_, _12452_, _06461_);
  or _76652_ (_26480_, _26479_, _26478_);
  and _76653_ (_26481_, _26480_, _12550_);
  or _76654_ (_26482_, _26481_, _26435_);
  nand _76655_ (_26483_, _26482_, _06465_);
  and _76656_ (_26484_, _12452_, _06464_);
  nor _76657_ (_26485_, _26484_, _25401_);
  nand _76658_ (_26486_, _26485_, _26483_);
  nor _76659_ (_26487_, _26432_, _12560_);
  nor _76660_ (_26488_, _26487_, _06268_);
  and _76661_ (_26489_, _26488_, _26486_);
  or _76662_ (_26490_, _26489_, _26434_);
  nand _76663_ (_26491_, _26490_, _06013_);
  and _76664_ (_26492_, _08892_, _12563_);
  nor _76665_ (_26493_, _26492_, _06267_);
  nand _76666_ (_26494_, _26493_, _26491_);
  and _76667_ (_26495_, _12451_, _06267_);
  nor _76668_ (_26496_, _26495_, _12379_);
  and _76669_ (_26497_, _26496_, _26494_);
  and _76670_ (_26498_, _12371_, _12238_);
  not _76671_ (_26499_, _26464_);
  nor _76672_ (_26500_, _26499_, _12371_);
  or _76673_ (_26501_, _26500_, _12378_);
  nor _76674_ (_26502_, _26501_, _26498_);
  nor _76675_ (_26503_, _26502_, _26497_);
  or _76676_ (_26504_, _26503_, _06347_);
  and _76677_ (_26505_, _26464_, _12335_);
  and _76678_ (_26506_, _12333_, _12238_);
  or _76679_ (_26507_, _26506_, _12177_);
  or _76680_ (_26508_, _26507_, _26505_);
  nand _76681_ (_26509_, _26508_, _26504_);
  or _76682_ (_26510_, _26509_, _06480_);
  nor _76683_ (_26511_, _26499_, _12587_);
  and _76684_ (_26512_, _12587_, _12238_);
  nor _76685_ (_26513_, _26512_, _26511_);
  or _76686_ (_26514_, _26513_, _06774_);
  and _76687_ (_26515_, _26514_, _26510_);
  or _76688_ (_26516_, _26515_, _06371_);
  and _76689_ (_26517_, _12604_, _12238_);
  not _76690_ (_26518_, _12604_);
  and _76691_ (_26520_, _26464_, _26518_);
  or _76692_ (_26521_, _26520_, _26517_);
  and _76693_ (_26522_, _26521_, _06371_);
  nor _76694_ (_26523_, _26522_, _12174_);
  and _76695_ (_26524_, _26523_, _26516_);
  or _76696_ (_26525_, _26524_, _26433_);
  nand _76697_ (_26526_, _26525_, _06262_);
  and _76698_ (_26527_, _12452_, _06261_);
  nor _76699_ (_26528_, _26527_, _12613_);
  nand _76700_ (_26529_, _26528_, _26526_);
  nor _76701_ (_26531_, _08892_, _06007_);
  nor _76702_ (_26532_, _26531_, _25445_);
  nand _76703_ (_26533_, _26532_, _26529_);
  nor _76704_ (_26534_, _25322_, _12451_);
  nor _76705_ (_26535_, _26534_, _12631_);
  nand _76706_ (_26536_, _26535_, _26533_);
  nor _76707_ (_26537_, _26432_, _12630_);
  nor _76708_ (_26538_, _26537_, _06505_);
  nand _76709_ (_26539_, _26538_, _26536_);
  and _76710_ (_26540_, _12452_, _06505_);
  nor _76711_ (_26541_, _26540_, _25158_);
  and _76712_ (_26542_, _26541_, _26539_);
  nor _76713_ (_26543_, _08892_, _06020_);
  or _76714_ (_26544_, _26543_, _06504_);
  or _76715_ (_26545_, _26544_, _26542_);
  and _76716_ (_26546_, _12452_, _06504_);
  nor _76717_ (_26547_, _26546_, _26197_);
  nand _76718_ (_26548_, _26547_, _26545_);
  nor _76719_ (_26549_, _26432_, _12639_);
  nor _76720_ (_26550_, _26549_, _12644_);
  nand _76721_ (_26552_, _26550_, _26548_);
  nor _76722_ (_26553_, _12451_, _12643_);
  nor _76723_ (_26554_, _26553_, _10515_);
  nand _76724_ (_26555_, _26554_, _26552_);
  nor _76725_ (_26556_, _26432_, _05984_);
  nor _76726_ (_26557_, _26556_, _06257_);
  and _76727_ (_26558_, _26557_, _26555_);
  or _76728_ (_26559_, _26558_, _26427_);
  nand _76729_ (_26560_, _26559_, _05978_);
  and _76730_ (_26561_, _08892_, _06254_);
  nor _76731_ (_26563_, _26561_, _06373_);
  nand _76732_ (_26564_, _26563_, _26560_);
  and _76733_ (_26565_, _12238_, _06373_);
  nor _76734_ (_26566_, _26565_, _12659_);
  nand _76735_ (_26567_, _26566_, _26564_);
  nor _76736_ (_26568_, _12451_, _07216_);
  nor _76737_ (_26569_, _26568_, _10094_);
  and _76738_ (_26570_, _26569_, _26567_);
  nor _76739_ (_26571_, _12239_, _05982_);
  nor _76740_ (_26572_, _26571_, _26570_);
  nand _76741_ (_26574_, _26572_, _12172_);
  nor _76742_ (_26575_, _26431_, _12172_);
  nor _76743_ (_26576_, _26575_, _06323_);
  nand _76744_ (_26577_, _26576_, _26574_);
  and _76745_ (_26578_, _12451_, _06323_);
  nor _76746_ (_26579_, _26578_, _12668_);
  nand _76747_ (_26580_, _26579_, _26577_);
  and _76748_ (_26581_, _08892_, _12668_);
  nor _76749_ (_26582_, _26581_, _12674_);
  nand _76750_ (_26583_, _26582_, _26580_);
  and _76751_ (_26585_, _26412_, _12674_);
  nor _76752_ (_26586_, _26585_, _09031_);
  and _76753_ (_26587_, _26586_, _26583_);
  or _76754_ (_26588_, _26587_, _26425_);
  nand _76755_ (_26589_, _26588_, _06219_);
  and _76756_ (_26590_, _12239_, _06218_);
  nor _76757_ (_26591_, _26590_, _10929_);
  nand _76758_ (_26592_, _26591_, _26589_);
  and _76759_ (_26593_, _12451_, _10929_);
  nor _76760_ (_26594_, _26593_, _12690_);
  nand _76761_ (_26595_, _26594_, _26592_);
  and _76762_ (_26596_, _12709_, _12706_);
  nor _76763_ (_26597_, _26596_, _12710_);
  nor _76764_ (_26598_, _26597_, _12691_);
  nor _76765_ (_26599_, _26598_, _06322_);
  nand _76766_ (_26600_, _26599_, _26595_);
  and _76767_ (_26601_, _12451_, _06322_);
  nor _76768_ (_26602_, _26601_, _06217_);
  nand _76769_ (_26603_, _26602_, _26600_);
  and _76770_ (_26604_, _08892_, _06217_);
  nor _76771_ (_26606_, _26604_, _12733_);
  and _76772_ (_26607_, _26606_, _26603_);
  or _76773_ (_26608_, _26607_, _26424_);
  nand _76774_ (_26609_, _26608_, _12169_);
  not _76775_ (_26610_, _12166_);
  nor _76776_ (_26611_, _26432_, _12169_);
  nor _76777_ (_26612_, _26611_, _26610_);
  nand _76778_ (_26613_, _26612_, _26609_);
  nor _76779_ (_26614_, _12451_, _12166_);
  nor _76780_ (_26615_, _26614_, _06369_);
  nand _76781_ (_26617_, _26615_, _26613_);
  and _76782_ (_26618_, _12238_, _06369_);
  nor _76783_ (_26619_, _26618_, _06536_);
  and _76784_ (_26620_, _26619_, _26617_);
  and _76785_ (_26621_, _12452_, _06536_);
  or _76786_ (_26622_, _26621_, _26620_);
  nand _76787_ (_26623_, _26622_, _05955_);
  and _76788_ (_26624_, _08892_, _12750_);
  nor _76789_ (_26625_, _26624_, _12755_);
  and _76790_ (_26626_, _26625_, _26623_);
  or _76791_ (_26628_, _26626_, _26420_);
  nand _76792_ (_26629_, _26628_, _10979_);
  not _76793_ (_26630_, _12164_);
  nor _76794_ (_26631_, _26432_, _10979_);
  nor _76795_ (_26632_, _26631_, _26630_);
  nand _76796_ (_26633_, _26632_, _26629_);
  nor _76797_ (_26634_, _12164_, _12451_);
  nor _76798_ (_26635_, _26634_, _06375_);
  nand _76799_ (_26636_, _26635_, _26633_);
  and _76800_ (_26637_, _12238_, _06375_);
  nor _76801_ (_26639_, _26637_, _06545_);
  and _76802_ (_26640_, _26639_, _26636_);
  and _76803_ (_26641_, _12452_, _06545_);
  or _76804_ (_26642_, _26641_, _26640_);
  nand _76805_ (_26643_, _26642_, _05961_);
  and _76806_ (_26644_, _08892_, _07233_);
  nor _76807_ (_26645_, _26644_, _12776_);
  and _76808_ (_26646_, _26645_, _26643_);
  and _76809_ (_26647_, _12451_, \oc8051_golden_model_1.PSW [7]);
  and _76810_ (_26648_, _26412_, _10558_);
  or _76811_ (_26650_, _26648_, _26647_);
  and _76812_ (_26651_, _26650_, _12776_);
  or _76813_ (_26652_, _26651_, _26646_);
  nand _76814_ (_26653_, _26652_, _12162_);
  nor _76815_ (_26654_, _26432_, _12162_);
  nor _76816_ (_26655_, _26654_, _11023_);
  nand _76817_ (_26656_, _26655_, _26653_);
  nor _76818_ (_26657_, _12451_, _11022_);
  nor _76819_ (_26658_, _26657_, _06366_);
  nand _76820_ (_26659_, _26658_, _26656_);
  and _76821_ (_26660_, _12238_, _06366_);
  nor _76822_ (_26661_, _26660_, _06528_);
  and _76823_ (_26662_, _26661_, _26659_);
  and _76824_ (_26663_, _12452_, _06528_);
  or _76825_ (_26664_, _26663_, _26662_);
  nand _76826_ (_26665_, _26664_, _05966_);
  and _76827_ (_26666_, _08892_, _12795_);
  nor _76828_ (_26667_, _26666_, _12800_);
  and _76829_ (_26668_, _26667_, _26665_);
  or _76830_ (_26669_, _26668_, _26416_);
  nand _76831_ (_26671_, _26669_, _12154_);
  nor _76832_ (_26672_, _26432_, _12154_);
  nor _76833_ (_26673_, _26672_, _14297_);
  nand _76834_ (_26674_, _26673_, _26671_);
  nor _76835_ (_26675_, _12451_, _12153_);
  nor _76836_ (_26676_, _26675_, _11125_);
  nand _76837_ (_26677_, _26676_, _26674_);
  and _76838_ (_26678_, _26431_, _11125_);
  nor _76839_ (_26679_, _26678_, _06551_);
  and _76840_ (_26680_, _26679_, _26677_);
  and _76841_ (_26682_, _09212_, _06551_);
  or _76842_ (_26683_, _26682_, _26680_);
  nand _76843_ (_26684_, _26683_, _05959_);
  and _76844_ (_26685_, _08892_, _07253_);
  nor _76845_ (_26686_, _26685_, _06365_);
  and _76846_ (_26687_, _26686_, _26684_);
  nor _76847_ (_26688_, _12239_, _13004_);
  and _76848_ (_26689_, _26464_, _13004_);
  nor _76849_ (_26690_, _26689_, _26688_);
  nor _76850_ (_26691_, _26690_, _06558_);
  or _76851_ (_26693_, _26691_, _26687_);
  nand _76852_ (_26694_, _26693_, _12151_);
  nor _76853_ (_26695_, _26432_, _12151_);
  nor _76854_ (_26696_, _26695_, _19056_);
  nand _76855_ (_26697_, _26696_, _26694_);
  nor _76856_ (_26698_, _13012_, _12451_);
  nor _76857_ (_26699_, _26698_, _11284_);
  nand _76858_ (_26700_, _26699_, _26697_);
  and _76859_ (_26701_, _26431_, _11284_);
  nor _76860_ (_26702_, _26701_, _06281_);
  nand _76861_ (_26704_, _26702_, _26700_);
  and _76862_ (_26705_, _09212_, _06281_);
  nor _76863_ (_26706_, _26705_, _25646_);
  nand _76864_ (_26707_, _26706_, _26704_);
  nor _76865_ (_26708_, _08892_, _05964_);
  nor _76866_ (_26709_, _26708_, _06362_);
  nand _76867_ (_26710_, _26709_, _26707_);
  and _76868_ (_26711_, _12239_, _13004_);
  nor _76869_ (_26712_, _26464_, _13004_);
  nor _76870_ (_26713_, _26712_, _26711_);
  nor _76871_ (_26715_, _26713_, _06921_);
  nor _76872_ (_26716_, _26715_, _13031_);
  nand _76873_ (_26717_, _26716_, _26710_);
  nor _76874_ (_26718_, _26432_, _13030_);
  nor _76875_ (_26719_, _26718_, _06568_);
  nand _76876_ (_26720_, _26719_, _26717_);
  and _76877_ (_26721_, _12452_, _06568_);
  nor _76878_ (_26722_, _26721_, _13038_);
  nand _76879_ (_26723_, _26722_, _26720_);
  nor _76880_ (_26724_, _26432_, _13037_);
  nor _76881_ (_26725_, _26724_, _07695_);
  and _76882_ (_26726_, _26725_, _26723_);
  or _76883_ (_26727_, _26726_, _26409_);
  nand _76884_ (_26728_, _26727_, _05928_);
  nor _76885_ (_26729_, _26713_, _05928_);
  nor _76886_ (_26730_, _26729_, _13053_);
  nand _76887_ (_26731_, _26730_, _26728_);
  nor _76888_ (_26732_, _26432_, _13052_);
  nor _76889_ (_26733_, _26732_, _06278_);
  nand _76890_ (_26734_, _26733_, _26731_);
  and _76891_ (_26736_, _12452_, _06278_);
  nor _76892_ (_26737_, _26736_, _13059_);
  nand _76893_ (_26738_, _26737_, _26734_);
  nor _76894_ (_26739_, _26432_, _12141_);
  nor _76895_ (_26740_, _26739_, _25301_);
  nand _76896_ (_26741_, _26740_, _26738_);
  and _76897_ (_26742_, _25301_, _08892_);
  nor _76898_ (_26743_, _26742_, _13068_);
  and _76899_ (_26744_, _26743_, _26741_);
  and _76900_ (_26745_, _26431_, _13068_);
  or _76901_ (_26747_, _26745_, _26744_);
  or _76902_ (_26748_, _26747_, _01351_);
  or _76903_ (_26749_, _01347_, \oc8051_golden_model_1.PC [4]);
  and _76904_ (_26750_, _26749_, _42618_);
  and _76905_ (_43250_, _26750_, _26748_);
  and _76906_ (_26751_, _12446_, _06278_);
  and _76907_ (_26752_, _12446_, _06568_);
  nor _76908_ (_26753_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor _76909_ (_26754_, _12446_, _05630_);
  nor _76910_ (_26755_, _26754_, _26753_);
  nor _76911_ (_26757_, _26755_, _12151_);
  nor _76912_ (_26758_, _26755_, _12154_);
  nor _76913_ (_26759_, _26755_, _12162_);
  nor _76914_ (_26760_, _26755_, _10979_);
  nor _76915_ (_26761_, _26755_, _12169_);
  nor _76916_ (_26762_, _12446_, _09030_);
  nor _76917_ (_26763_, _25322_, _12446_);
  not _76918_ (_26764_, _26755_);
  and _76919_ (_26765_, _26764_, _12174_);
  or _76920_ (_26766_, _12534_, _12233_);
  or _76921_ (_26768_, _12236_, _12235_);
  not _76922_ (_26769_, _26768_);
  nor _76923_ (_26770_, _26769_, _12267_);
  and _76924_ (_26771_, _26769_, _12267_);
  nor _76925_ (_26772_, _26771_, _26770_);
  not _76926_ (_26773_, _26772_);
  or _76927_ (_26774_, _26773_, _12536_);
  and _76928_ (_26775_, _26774_, _26766_);
  or _76929_ (_26776_, _26775_, _07151_);
  and _76930_ (_26777_, _12507_, _12446_);
  or _76931_ (_26779_, _12448_, _12449_);
  and _76932_ (_26780_, _26779_, _12474_);
  nor _76933_ (_26781_, _26779_, _12474_);
  nor _76934_ (_26782_, _26781_, _26780_);
  and _76935_ (_26783_, _26782_, _12393_);
  nor _76936_ (_26784_, _26783_, _26777_);
  nand _76937_ (_26785_, _26784_, _12387_);
  nor _76938_ (_26786_, _07486_, \oc8051_golden_model_1.PC [5]);
  nor _76939_ (_26787_, _26786_, _07141_);
  and _76940_ (_26788_, _12446_, _07141_);
  nor _76941_ (_26789_, _26788_, _06781_);
  not _76942_ (_26790_, _26789_);
  nor _76943_ (_26791_, _26790_, _26787_);
  not _76944_ (_26792_, _26791_);
  nor _76945_ (_26793_, _26755_, _12513_);
  nor _76946_ (_26794_, _26793_, _06758_);
  and _76947_ (_26795_, _26794_, _26792_);
  nor _76948_ (_26796_, _08926_, _07504_);
  or _76949_ (_26797_, _26796_, _12516_);
  nor _76950_ (_26798_, _26797_, _26795_);
  nor _76951_ (_26800_, _26755_, _12512_);
  nor _76952_ (_26801_, _26800_, _26798_);
  nor _76953_ (_26802_, _26801_, _12387_);
  nor _76954_ (_26803_, _26802_, _07154_);
  and _76955_ (_26804_, _26803_, _26785_);
  and _76956_ (_26805_, _26755_, _07154_);
  or _76957_ (_26806_, _26805_, _06341_);
  or _76958_ (_26807_, _26806_, _26804_);
  nand _76959_ (_26808_, _26807_, _26776_);
  nand _76960_ (_26809_, _26808_, _12541_);
  nor _76961_ (_26811_, _26755_, _12541_);
  nor _76962_ (_26812_, _26811_, _06272_);
  nand _76963_ (_26813_, _26812_, _26809_);
  and _76964_ (_26814_, _12446_, _06272_);
  nor _76965_ (_26815_, _26814_, _07611_);
  nand _76966_ (_26816_, _26815_, _26813_);
  and _76967_ (_26817_, _08926_, _07611_);
  nor _76968_ (_26818_, _26817_, _06461_);
  nand _76969_ (_26819_, _26818_, _26816_);
  and _76970_ (_26820_, _12446_, _06461_);
  nor _76971_ (_26822_, _26820_, _12551_);
  nand _76972_ (_26823_, _26822_, _26819_);
  nor _76973_ (_26824_, _26755_, _12550_);
  nor _76974_ (_26825_, _26824_, _06464_);
  nand _76975_ (_26826_, _26825_, _26823_);
  and _76976_ (_26827_, _12446_, _06464_);
  nor _76977_ (_26828_, _26827_, _25401_);
  nand _76978_ (_26829_, _26828_, _26826_);
  nor _76979_ (_26830_, _26755_, _12560_);
  nor _76980_ (_26831_, _26830_, _06268_);
  nand _76981_ (_26833_, _26831_, _26829_);
  and _76982_ (_26834_, _12446_, _06268_);
  nor _76983_ (_26835_, _26834_, _12563_);
  nand _76984_ (_26836_, _26835_, _26833_);
  and _76985_ (_26837_, _08926_, _12563_);
  nor _76986_ (_26838_, _26837_, _06267_);
  nand _76987_ (_26839_, _26838_, _26836_);
  and _76988_ (_26840_, _12446_, _06267_);
  nor _76989_ (_26841_, _26840_, _12379_);
  nand _76990_ (_26842_, _26841_, _26839_);
  and _76991_ (_26844_, _12371_, _12233_);
  nor _76992_ (_26845_, _26772_, _12371_);
  or _76993_ (_26846_, _26845_, _26844_);
  nor _76994_ (_26847_, _26846_, _12378_);
  nor _76995_ (_26848_, _26847_, _06347_);
  nand _76996_ (_26849_, _26848_, _26842_);
  or _76997_ (_26850_, _26772_, _12333_);
  or _76998_ (_26851_, _12335_, _12234_);
  nand _76999_ (_26852_, _26851_, _26850_);
  nand _77000_ (_26853_, _26852_, _06347_);
  and _77001_ (_26854_, _26853_, _06774_);
  nand _77002_ (_26855_, _26854_, _26849_);
  nor _77003_ (_26856_, _26772_, _12587_);
  not _77004_ (_26857_, _26856_);
  and _77005_ (_26858_, _12587_, _12233_);
  nor _77006_ (_26859_, _26858_, _06774_);
  and _77007_ (_26860_, _26859_, _26857_);
  nor _77008_ (_26861_, _26860_, _06371_);
  nand _77009_ (_26862_, _26861_, _26855_);
  and _77010_ (_26863_, _12604_, _12234_);
  and _77011_ (_26865_, _26772_, _26518_);
  or _77012_ (_26866_, _26865_, _12176_);
  nor _77013_ (_26867_, _26866_, _26863_);
  nor _77014_ (_26868_, _26867_, _12174_);
  and _77015_ (_26869_, _26868_, _26862_);
  or _77016_ (_26870_, _26869_, _26765_);
  nand _77017_ (_26871_, _26870_, _06262_);
  and _77018_ (_26872_, _12447_, _06261_);
  nor _77019_ (_26873_, _26872_, _12613_);
  nand _77020_ (_26874_, _26873_, _26871_);
  nor _77021_ (_26876_, _08926_, _06007_);
  nor _77022_ (_26877_, _26876_, _25445_);
  and _77023_ (_26878_, _26877_, _26874_);
  or _77024_ (_26879_, _26878_, _26763_);
  nand _77025_ (_26880_, _26879_, _12630_);
  nor _77026_ (_26881_, _26755_, _12630_);
  nor _77027_ (_26882_, _26881_, _06505_);
  nand _77028_ (_26883_, _26882_, _26880_);
  and _77029_ (_26884_, _12446_, _06505_);
  nor _77030_ (_26885_, _26884_, _25158_);
  nand _77031_ (_26887_, _26885_, _26883_);
  and _77032_ (_26888_, _08926_, _25158_);
  nor _77033_ (_26889_, _26888_, _06504_);
  nand _77034_ (_26890_, _26889_, _26887_);
  and _77035_ (_26891_, _12446_, _06504_);
  nor _77036_ (_26892_, _26891_, _26197_);
  and _77037_ (_26893_, _26892_, _26890_);
  nor _77038_ (_26894_, _26755_, _12639_);
  or _77039_ (_26895_, _26894_, _26893_);
  nand _77040_ (_26896_, _26895_, _12643_);
  nor _77041_ (_26898_, _12446_, _12643_);
  nor _77042_ (_26899_, _26898_, _10515_);
  nand _77043_ (_26900_, _26899_, _26896_);
  nor _77044_ (_26901_, _26764_, _05984_);
  nor _77045_ (_26902_, _26901_, _06257_);
  and _77046_ (_26903_, _26902_, _26900_);
  and _77047_ (_26904_, _12447_, _06257_);
  or _77048_ (_26905_, _26904_, _26903_);
  nand _77049_ (_26906_, _26905_, _05978_);
  and _77050_ (_26907_, _08926_, _06254_);
  nor _77051_ (_26909_, _26907_, _06373_);
  nand _77052_ (_26910_, _26909_, _26906_);
  and _77053_ (_26911_, _12233_, _06373_);
  nor _77054_ (_26912_, _26911_, _12659_);
  nand _77055_ (_26913_, _26912_, _26910_);
  nor _77056_ (_26914_, _12446_, _07216_);
  nor _77057_ (_26915_, _26914_, _10094_);
  nand _77058_ (_26916_, _26915_, _26913_);
  nor _77059_ (_26917_, _12234_, _05982_);
  nor _77060_ (_26918_, _26917_, _25492_);
  nand _77061_ (_26920_, _26918_, _26916_);
  nor _77062_ (_26921_, _26755_, _12172_);
  nor _77063_ (_26922_, _26921_, _06323_);
  nand _77064_ (_26923_, _26922_, _26920_);
  and _77065_ (_26924_, _12446_, _06323_);
  nor _77066_ (_26925_, _26924_, _12668_);
  nand _77067_ (_26926_, _26925_, _26923_);
  and _77068_ (_26927_, _08926_, _12668_);
  nor _77069_ (_26928_, _26927_, _12674_);
  nand _77070_ (_26929_, _26928_, _26926_);
  and _77071_ (_26931_, _26782_, _12674_);
  nor _77072_ (_26932_, _26931_, _09031_);
  and _77073_ (_26933_, _26932_, _26929_);
  or _77074_ (_26934_, _26933_, _26762_);
  nand _77075_ (_26935_, _26934_, _06219_);
  and _77076_ (_26936_, _12234_, _06218_);
  nor _77077_ (_26937_, _26936_, _10929_);
  nand _77078_ (_26938_, _26937_, _26935_);
  and _77079_ (_26939_, _12446_, _10929_);
  nor _77080_ (_26940_, _26939_, _12690_);
  nand _77081_ (_26941_, _26940_, _26938_);
  and _77082_ (_26942_, _12711_, _12704_);
  nor _77083_ (_26943_, _26942_, _12712_);
  nor _77084_ (_26944_, _26943_, _12691_);
  nor _77085_ (_26945_, _26944_, _06322_);
  nand _77086_ (_26946_, _26945_, _26941_);
  and _77087_ (_26947_, _12446_, _06322_);
  nor _77088_ (_26948_, _26947_, _06217_);
  nand _77089_ (_26949_, _26948_, _26946_);
  and _77090_ (_26950_, _08926_, _06217_);
  nor _77091_ (_26952_, _26950_, _12733_);
  nand _77092_ (_26953_, _26952_, _26949_);
  and _77093_ (_26954_, _12446_, _11342_);
  and _77094_ (_26955_, _26782_, _12759_);
  or _77095_ (_26956_, _26955_, _26954_);
  and _77096_ (_26957_, _26956_, _12733_);
  nor _77097_ (_26958_, _26957_, _12737_);
  and _77098_ (_26959_, _26958_, _26953_);
  or _77099_ (_26960_, _26959_, _26761_);
  nand _77100_ (_26961_, _26960_, _12166_);
  nor _77101_ (_26963_, _12446_, _12166_);
  nor _77102_ (_26964_, _26963_, _06369_);
  nand _77103_ (_26965_, _26964_, _26961_);
  and _77104_ (_26966_, _12233_, _06369_);
  nor _77105_ (_26967_, _26966_, _06536_);
  and _77106_ (_26968_, _26967_, _26965_);
  and _77107_ (_26969_, _12447_, _06536_);
  or _77108_ (_26970_, _26969_, _26968_);
  nand _77109_ (_26971_, _26970_, _05955_);
  and _77110_ (_26972_, _08926_, _12750_);
  nor _77111_ (_26974_, _26972_, _12755_);
  nand _77112_ (_26975_, _26974_, _26971_);
  nor _77113_ (_26976_, _12447_, _11342_);
  and _77114_ (_26977_, _26782_, _11342_);
  or _77115_ (_26978_, _26977_, _26976_);
  and _77116_ (_26979_, _26978_, _12755_);
  nor _77117_ (_26980_, _26979_, _10980_);
  and _77118_ (_26981_, _26980_, _26975_);
  or _77119_ (_26982_, _26981_, _26760_);
  nand _77120_ (_26983_, _26982_, _12164_);
  nor _77121_ (_26985_, _12164_, _12446_);
  nor _77122_ (_26986_, _26985_, _06375_);
  nand _77123_ (_26987_, _26986_, _26983_);
  and _77124_ (_26988_, _12233_, _06375_);
  nor _77125_ (_26989_, _26988_, _06545_);
  and _77126_ (_26990_, _26989_, _26987_);
  and _77127_ (_26991_, _12447_, _06545_);
  or _77128_ (_26992_, _26991_, _26990_);
  nand _77129_ (_26993_, _26992_, _05961_);
  and _77130_ (_26994_, _08926_, _07233_);
  nor _77131_ (_26996_, _26994_, _12776_);
  nand _77132_ (_26997_, _26996_, _26993_);
  nor _77133_ (_26998_, _26782_, \oc8051_golden_model_1.PSW [7]);
  nor _77134_ (_26999_, _12446_, _10558_);
  nor _77135_ (_27000_, _26999_, _12782_);
  not _77136_ (_27001_, _27000_);
  nor _77137_ (_27002_, _27001_, _26998_);
  nor _77138_ (_27003_, _27002_, _12780_);
  and _77139_ (_27004_, _27003_, _26997_);
  or _77140_ (_27005_, _27004_, _26759_);
  nand _77141_ (_27006_, _27005_, _11022_);
  nor _77142_ (_27007_, _12446_, _11022_);
  nor _77143_ (_27008_, _27007_, _06366_);
  nand _77144_ (_27009_, _27008_, _27006_);
  and _77145_ (_27010_, _12233_, _06366_);
  nor _77146_ (_27011_, _27010_, _06528_);
  and _77147_ (_27012_, _27011_, _27009_);
  and _77148_ (_27013_, _12447_, _06528_);
  or _77149_ (_27014_, _27013_, _27012_);
  nand _77150_ (_27015_, _27014_, _05966_);
  and _77151_ (_27017_, _08926_, _12795_);
  nor _77152_ (_27018_, _27017_, _12800_);
  nand _77153_ (_27019_, _27018_, _27015_);
  and _77154_ (_27020_, _12446_, _10558_);
  and _77155_ (_27021_, _26782_, \oc8051_golden_model_1.PSW [7]);
  or _77156_ (_27022_, _27021_, _27020_);
  and _77157_ (_27023_, _27022_, _12800_);
  nor _77158_ (_27024_, _27023_, _12804_);
  and _77159_ (_27025_, _27024_, _27019_);
  or _77160_ (_27026_, _27025_, _26758_);
  nand _77161_ (_27028_, _27026_, _12153_);
  nor _77162_ (_27029_, _12446_, _12153_);
  nor _77163_ (_27030_, _27029_, _11125_);
  nand _77164_ (_27031_, _27030_, _27028_);
  and _77165_ (_27032_, _26755_, _11125_);
  nor _77166_ (_27033_, _27032_, _06551_);
  and _77167_ (_27034_, _27033_, _27031_);
  and _77168_ (_27035_, _09167_, _06551_);
  or _77169_ (_27036_, _27035_, _27034_);
  nand _77170_ (_27037_, _27036_, _05959_);
  and _77171_ (_27039_, _08926_, _07253_);
  nor _77172_ (_27040_, _27039_, _06365_);
  nand _77173_ (_27041_, _27040_, _27037_);
  and _77174_ (_27042_, _26772_, _13004_);
  nor _77175_ (_27043_, _12233_, _13004_);
  or _77176_ (_27044_, _27043_, _06558_);
  or _77177_ (_27045_, _27044_, _27042_);
  and _77178_ (_27046_, _27045_, _12151_);
  and _77179_ (_27047_, _27046_, _27041_);
  or _77180_ (_27048_, _27047_, _26757_);
  nand _77181_ (_27050_, _27048_, _13012_);
  nor _77182_ (_27051_, _13012_, _12446_);
  nor _77183_ (_27052_, _27051_, _11284_);
  nand _77184_ (_27053_, _27052_, _27050_);
  and _77185_ (_27054_, _26755_, _11284_);
  nor _77186_ (_27055_, _27054_, _06281_);
  and _77187_ (_27056_, _27055_, _27053_);
  and _77188_ (_27057_, _09167_, _06281_);
  or _77189_ (_27058_, _27057_, _27056_);
  nand _77190_ (_27059_, _27058_, _05964_);
  and _77191_ (_27061_, _08926_, _25646_);
  nor _77192_ (_27062_, _27061_, _06362_);
  nand _77193_ (_27063_, _27062_, _27059_);
  and _77194_ (_27064_, _12234_, _13004_);
  nor _77195_ (_27065_, _26773_, _13004_);
  nor _77196_ (_27066_, _27065_, _27064_);
  and _77197_ (_27067_, _27066_, _06362_);
  nor _77198_ (_27068_, _27067_, _13031_);
  nand _77199_ (_27069_, _27068_, _27063_);
  nor _77200_ (_27070_, _26755_, _13030_);
  nor _77201_ (_27072_, _27070_, _06568_);
  and _77202_ (_27073_, _27072_, _27069_);
  or _77203_ (_27074_, _27073_, _26752_);
  nand _77204_ (_27075_, _27074_, _13037_);
  nor _77205_ (_27076_, _26764_, _13037_);
  nor _77206_ (_27077_, _27076_, _07695_);
  nand _77207_ (_27078_, _27077_, _27075_);
  and _77208_ (_27079_, _08926_, _07695_);
  nor _77209_ (_27080_, _27079_, _05927_);
  nand _77210_ (_27081_, _27080_, _27078_);
  and _77211_ (_27083_, _27066_, _05927_);
  nor _77212_ (_27084_, _27083_, _13053_);
  nand _77213_ (_27085_, _27084_, _27081_);
  nor _77214_ (_27086_, _26755_, _13052_);
  nor _77215_ (_27087_, _27086_, _06278_);
  and _77216_ (_27088_, _27087_, _27085_);
  or _77217_ (_27089_, _27088_, _26751_);
  nand _77218_ (_27090_, _27089_, _12141_);
  nor _77219_ (_27091_, _26764_, _12141_);
  nor _77220_ (_27092_, _27091_, _25301_);
  nand _77221_ (_27094_, _27092_, _27090_);
  and _77222_ (_27095_, _25301_, _08926_);
  nor _77223_ (_27096_, _27095_, _13068_);
  and _77224_ (_27097_, _27096_, _27094_);
  and _77225_ (_27098_, _26755_, _13068_);
  or _77226_ (_27099_, _27098_, _27097_);
  or _77227_ (_27100_, _27099_, _01351_);
  or _77228_ (_27101_, _01347_, \oc8051_golden_model_1.PC [5]);
  and _77229_ (_27102_, _27101_, _42618_);
  and _77230_ (_43251_, _27102_, _27100_);
  and _77231_ (_27104_, _08657_, _12142_);
  and _77232_ (_27105_, _08656_, _12142_);
  nor _77233_ (_27106_, _27105_, \oc8051_golden_model_1.PC [6]);
  nor _77234_ (_27107_, _27106_, _27104_);
  and _77235_ (_27108_, _27107_, _13068_);
  and _77236_ (_27109_, _08857_, _07695_);
  not _77237_ (_27110_, _27107_);
  and _77238_ (_27111_, _27110_, _11284_);
  and _77239_ (_27112_, _12226_, _06366_);
  and _77240_ (_27113_, _12226_, _06375_);
  and _77241_ (_27115_, _12226_, _06369_);
  nor _77242_ (_27116_, _25322_, _12439_);
  and _77243_ (_27117_, _27110_, _12174_);
  and _77244_ (_27118_, _12333_, _12226_);
  and _77245_ (_27119_, _12269_, _12230_);
  nor _77246_ (_27120_, _27119_, _12270_);
  not _77247_ (_27121_, _27120_);
  and _77248_ (_27122_, _27121_, _12335_);
  nor _77249_ (_27123_, _27122_, _27118_);
  nor _77250_ (_27124_, _27123_, _12177_);
  and _77251_ (_27126_, _12440_, _06268_);
  nor _77252_ (_27127_, _27107_, _12550_);
  or _77253_ (_27128_, _27120_, _12536_);
  or _77254_ (_27129_, _12534_, _12225_);
  and _77255_ (_27130_, _27129_, _06341_);
  nand _77256_ (_27131_, _27130_, _27128_);
  and _77257_ (_27132_, _12507_, _12439_);
  nor _77258_ (_27133_, _12476_, _12443_);
  nor _77259_ (_27134_, _27133_, _12477_);
  and _77260_ (_27135_, _27134_, _12393_);
  nor _77261_ (_27137_, _27135_, _27132_);
  nand _77262_ (_27138_, _27137_, _12387_);
  and _77263_ (_27139_, _08857_, _06758_);
  and _77264_ (_27140_, _12440_, _07141_);
  nor _77265_ (_27141_, _27140_, _06781_);
  and _77266_ (_27142_, _07487_, \oc8051_golden_model_1.PC [6]);
  or _77267_ (_27143_, _27142_, _07141_);
  and _77268_ (_27144_, _27143_, _27141_);
  nor _77269_ (_27145_, _27110_, _12513_);
  or _77270_ (_27146_, _27145_, _06758_);
  nor _77271_ (_27148_, _27146_, _27144_);
  nor _77272_ (_27149_, _27148_, _12516_);
  not _77273_ (_27150_, _27149_);
  nor _77274_ (_27151_, _27150_, _27139_);
  nor _77275_ (_27152_, _27110_, _12512_);
  nor _77276_ (_27153_, _27152_, _12387_);
  not _77277_ (_27154_, _27153_);
  nor _77278_ (_27155_, _27154_, _27151_);
  not _77279_ (_27156_, _27155_);
  nor _77280_ (_27157_, _07154_, _06341_);
  and _77281_ (_27159_, _27157_, _27156_);
  nand _77282_ (_27160_, _27159_, _27138_);
  nand _77283_ (_27161_, _27160_, _27131_);
  and _77284_ (_27162_, _27161_, _12541_);
  or _77285_ (_27163_, _12542_, _07154_);
  and _77286_ (_27164_, _27163_, _27107_);
  or _77287_ (_27165_, _27164_, _06272_);
  or _77288_ (_27166_, _27165_, _27162_);
  and _77289_ (_27167_, _12440_, _06272_);
  nor _77290_ (_27168_, _27167_, _07611_);
  and _77291_ (_27170_, _27168_, _27166_);
  nor _77292_ (_27171_, _08857_, _06010_);
  or _77293_ (_27172_, _27171_, _06461_);
  nor _77294_ (_27173_, _27172_, _27170_);
  and _77295_ (_27174_, _12440_, _06461_);
  or _77296_ (_27175_, _27174_, _27173_);
  and _77297_ (_27176_, _27175_, _12550_);
  or _77298_ (_27177_, _27176_, _27127_);
  nand _77299_ (_27178_, _27177_, _06465_);
  and _77300_ (_27179_, _12440_, _06464_);
  nor _77301_ (_27181_, _27179_, _25401_);
  nand _77302_ (_27182_, _27181_, _27178_);
  nor _77303_ (_27183_, _27110_, _12560_);
  nor _77304_ (_27184_, _27183_, _06268_);
  and _77305_ (_27185_, _27184_, _27182_);
  or _77306_ (_27186_, _27185_, _27126_);
  nand _77307_ (_27187_, _27186_, _06013_);
  and _77308_ (_27188_, _08857_, _12563_);
  nor _77309_ (_27189_, _27188_, _06267_);
  nand _77310_ (_27190_, _27189_, _27187_);
  and _77311_ (_27192_, _12439_, _06267_);
  nor _77312_ (_27193_, _27192_, _12379_);
  and _77313_ (_27194_, _27193_, _27190_);
  and _77314_ (_27195_, _12371_, _12225_);
  nor _77315_ (_27196_, _27121_, _12371_);
  or _77316_ (_27197_, _27196_, _12378_);
  nor _77317_ (_27198_, _27197_, _27195_);
  or _77318_ (_27199_, _27198_, _27194_);
  and _77319_ (_27200_, _27199_, _12177_);
  nor _77320_ (_27201_, _27200_, _27124_);
  or _77321_ (_27203_, _27201_, _06480_);
  nor _77322_ (_27204_, _27121_, _12587_);
  and _77323_ (_27205_, _12587_, _12225_);
  or _77324_ (_27206_, _27205_, _06774_);
  or _77325_ (_27207_, _27206_, _27204_);
  and _77326_ (_27208_, _27207_, _12176_);
  nand _77327_ (_27209_, _27208_, _27203_);
  and _77328_ (_27210_, _12604_, _12225_);
  and _77329_ (_27211_, _27120_, _26518_);
  or _77330_ (_27212_, _27211_, _27210_);
  and _77331_ (_27214_, _27212_, _06371_);
  nor _77332_ (_27215_, _27214_, _12174_);
  and _77333_ (_27216_, _27215_, _27209_);
  or _77334_ (_27217_, _27216_, _27117_);
  nand _77335_ (_27218_, _27217_, _06262_);
  and _77336_ (_27219_, _12440_, _06261_);
  nor _77337_ (_27220_, _27219_, _12613_);
  nand _77338_ (_27221_, _27220_, _27218_);
  nor _77339_ (_27222_, _08857_, _06007_);
  nor _77340_ (_27223_, _27222_, _25445_);
  and _77341_ (_27225_, _27223_, _27221_);
  or _77342_ (_27226_, _27225_, _27116_);
  nand _77343_ (_27227_, _27226_, _12630_);
  nor _77344_ (_27228_, _27107_, _12630_);
  nor _77345_ (_27229_, _27228_, _06505_);
  nand _77346_ (_27230_, _27229_, _27227_);
  and _77347_ (_27231_, _12439_, _06505_);
  nor _77348_ (_27232_, _27231_, _25158_);
  nand _77349_ (_27233_, _27232_, _27230_);
  and _77350_ (_27234_, _08857_, _25158_);
  nor _77351_ (_27235_, _27234_, _06504_);
  nand _77352_ (_27236_, _27235_, _27233_);
  and _77353_ (_27237_, _12439_, _06504_);
  nor _77354_ (_27238_, _27237_, _26197_);
  nand _77355_ (_27239_, _27238_, _27236_);
  nor _77356_ (_27240_, _27107_, _12639_);
  nor _77357_ (_27241_, _27240_, _12644_);
  nand _77358_ (_27242_, _27241_, _27239_);
  nor _77359_ (_27243_, _12440_, _12643_);
  nor _77360_ (_27244_, _27243_, _10515_);
  and _77361_ (_27247_, _27244_, _27242_);
  nor _77362_ (_27248_, _27107_, _05984_);
  or _77363_ (_27249_, _27248_, _27247_);
  nand _77364_ (_27250_, _27249_, _06258_);
  and _77365_ (_27251_, _12440_, _06257_);
  nor _77366_ (_27252_, _27251_, _06254_);
  nand _77367_ (_27253_, _27252_, _27250_);
  nor _77368_ (_27254_, _08857_, _05978_);
  nor _77369_ (_27255_, _27254_, _06373_);
  nand _77370_ (_27256_, _27255_, _27253_);
  and _77371_ (_27258_, _12226_, _06373_);
  nor _77372_ (_27259_, _27258_, _12659_);
  nand _77373_ (_27260_, _27259_, _27256_);
  nor _77374_ (_27261_, _12440_, _07216_);
  nor _77375_ (_27262_, _27261_, _10094_);
  nand _77376_ (_27263_, _27262_, _27260_);
  nor _77377_ (_27264_, _12225_, _05982_);
  nor _77378_ (_27265_, _27264_, _25492_);
  nand _77379_ (_27266_, _27265_, _27263_);
  nor _77380_ (_27267_, _27110_, _12172_);
  nor _77381_ (_27269_, _27267_, _06323_);
  nand _77382_ (_27270_, _27269_, _27266_);
  and _77383_ (_27271_, _12440_, _06323_);
  nor _77384_ (_27272_, _27271_, _12668_);
  nand _77385_ (_27273_, _27272_, _27270_);
  nor _77386_ (_27274_, _08857_, _05946_);
  nor _77387_ (_27275_, _27274_, _12674_);
  nand _77388_ (_27276_, _27275_, _27273_);
  nor _77389_ (_27277_, _27134_, _12679_);
  nor _77390_ (_27278_, _27277_, _09031_);
  nand _77391_ (_27280_, _27278_, _27276_);
  nor _77392_ (_27281_, _12440_, _09030_);
  nor _77393_ (_27282_, _27281_, _06218_);
  nand _77394_ (_27283_, _27282_, _27280_);
  and _77395_ (_27284_, _12226_, _06218_);
  nor _77396_ (_27285_, _27284_, _10929_);
  nand _77397_ (_27286_, _27285_, _27283_);
  and _77398_ (_27287_, _12439_, _10929_);
  nor _77399_ (_27288_, _27287_, _12690_);
  nand _77400_ (_27289_, _27288_, _27286_);
  and _77401_ (_27291_, _12713_, _12700_);
  nor _77402_ (_27292_, _27291_, _12714_);
  nor _77403_ (_27293_, _27292_, _12691_);
  nor _77404_ (_27294_, _27293_, _06322_);
  nand _77405_ (_27295_, _27294_, _27289_);
  and _77406_ (_27296_, _12439_, _06322_);
  nor _77407_ (_27297_, _27296_, _06217_);
  nand _77408_ (_27298_, _27297_, _27295_);
  and _77409_ (_27299_, _08857_, _06217_);
  nor _77410_ (_27300_, _27299_, _12733_);
  nand _77411_ (_27302_, _27300_, _27298_);
  and _77412_ (_27303_, _12439_, _11342_);
  and _77413_ (_27304_, _27134_, _12759_);
  or _77414_ (_27305_, _27304_, _27303_);
  and _77415_ (_27306_, _27305_, _12733_);
  nor _77416_ (_27307_, _27306_, _12737_);
  nand _77417_ (_27308_, _27307_, _27302_);
  nor _77418_ (_27309_, _27107_, _12169_);
  nor _77419_ (_27310_, _27309_, _26610_);
  nand _77420_ (_27311_, _27310_, _27308_);
  nor _77421_ (_27313_, _12440_, _12166_);
  nor _77422_ (_27314_, _27313_, _06369_);
  and _77423_ (_27315_, _27314_, _27311_);
  or _77424_ (_27316_, _27315_, _27115_);
  nand _77425_ (_27317_, _27316_, _07240_);
  and _77426_ (_27318_, _12440_, _06536_);
  nor _77427_ (_27319_, _27318_, _12750_);
  and _77428_ (_27320_, _27319_, _27317_);
  nor _77429_ (_27321_, _08857_, _05955_);
  or _77430_ (_27322_, _27321_, _27320_);
  nand _77431_ (_27324_, _27322_, _25061_);
  nor _77432_ (_27325_, _12440_, _11342_);
  and _77433_ (_27326_, _27134_, _11342_);
  or _77434_ (_27327_, _27326_, _27325_);
  and _77435_ (_27328_, _27327_, _12755_);
  nor _77436_ (_27329_, _27328_, _10980_);
  nand _77437_ (_27330_, _27329_, _27324_);
  nor _77438_ (_27331_, _27107_, _10979_);
  nor _77439_ (_27332_, _27331_, _26630_);
  nand _77440_ (_27333_, _27332_, _27330_);
  nor _77441_ (_27335_, _12164_, _12440_);
  nor _77442_ (_27336_, _27335_, _06375_);
  and _77443_ (_27337_, _27336_, _27333_);
  or _77444_ (_27338_, _27337_, _27113_);
  nand _77445_ (_27339_, _27338_, _07234_);
  and _77446_ (_27340_, _12440_, _06545_);
  nor _77447_ (_27341_, _27340_, _07233_);
  and _77448_ (_27342_, _27341_, _27339_);
  nor _77449_ (_27343_, _08857_, _05961_);
  or _77450_ (_27344_, _27343_, _27342_);
  nand _77451_ (_27346_, _27344_, _12782_);
  nor _77452_ (_27347_, _27134_, \oc8051_golden_model_1.PSW [7]);
  nor _77453_ (_27348_, _12439_, _10558_);
  nor _77454_ (_27349_, _27348_, _12782_);
  not _77455_ (_27350_, _27349_);
  nor _77456_ (_27351_, _27350_, _27347_);
  nor _77457_ (_27352_, _27351_, _12780_);
  nand _77458_ (_27353_, _27352_, _27346_);
  nor _77459_ (_27354_, _27107_, _12162_);
  nor _77460_ (_27355_, _27354_, _11023_);
  nand _77461_ (_27357_, _27355_, _27353_);
  nor _77462_ (_27358_, _12440_, _11022_);
  nor _77463_ (_27359_, _27358_, _06366_);
  and _77464_ (_27360_, _27359_, _27357_);
  or _77465_ (_27361_, _27360_, _27112_);
  nand _77466_ (_27362_, _27361_, _09061_);
  and _77467_ (_27363_, _12440_, _06528_);
  nor _77468_ (_27364_, _27363_, _12795_);
  and _77469_ (_27365_, _27364_, _27362_);
  nor _77470_ (_27366_, _08857_, _05966_);
  or _77471_ (_27368_, _27366_, _27365_);
  nand _77472_ (_27369_, _27368_, _25056_);
  and _77473_ (_27370_, _12439_, _10558_);
  and _77474_ (_27371_, _27134_, \oc8051_golden_model_1.PSW [7]);
  or _77475_ (_27372_, _27371_, _27370_);
  and _77476_ (_27373_, _27372_, _12800_);
  nor _77477_ (_27374_, _27373_, _12804_);
  nand _77478_ (_27375_, _27374_, _27369_);
  nor _77479_ (_27376_, _27107_, _12154_);
  nor _77480_ (_27377_, _27376_, _14297_);
  nand _77481_ (_27379_, _27377_, _27375_);
  nor _77482_ (_27380_, _12440_, _12153_);
  nor _77483_ (_27381_, _27380_, _11125_);
  nand _77484_ (_27382_, _27381_, _27379_);
  and _77485_ (_27383_, _27110_, _11125_);
  nor _77486_ (_27384_, _27383_, _06551_);
  nand _77487_ (_27385_, _27384_, _27382_);
  and _77488_ (_27386_, _09446_, _06551_);
  nor _77489_ (_27387_, _27386_, _07253_);
  nand _77490_ (_27388_, _27387_, _27385_);
  and _77491_ (_27390_, _08857_, _07253_);
  nor _77492_ (_27391_, _27390_, _06365_);
  nand _77493_ (_27392_, _27391_, _27388_);
  nor _77494_ (_27393_, _12225_, _13004_);
  and _77495_ (_27394_, _27121_, _13004_);
  or _77496_ (_27395_, _27394_, _06558_);
  or _77497_ (_27396_, _27395_, _27393_);
  and _77498_ (_27397_, _27396_, _12151_);
  nand _77499_ (_27398_, _27397_, _27392_);
  nor _77500_ (_27399_, _27107_, _12151_);
  nor _77501_ (_27401_, _27399_, _19056_);
  nand _77502_ (_27402_, _27401_, _27398_);
  nor _77503_ (_27403_, _13012_, _12440_);
  nor _77504_ (_27404_, _27403_, _11284_);
  and _77505_ (_27405_, _27404_, _27402_);
  or _77506_ (_27406_, _27405_, _27111_);
  nand _77507_ (_27407_, _27406_, _06282_);
  and _77508_ (_27408_, _09122_, _06281_);
  nor _77509_ (_27409_, _27408_, _25646_);
  nand _77510_ (_27410_, _27409_, _27407_);
  nor _77511_ (_27412_, _08857_, _05964_);
  nor _77512_ (_27413_, _27412_, _06362_);
  and _77513_ (_27414_, _27413_, _27410_);
  nor _77514_ (_27415_, _27120_, _13004_);
  and _77515_ (_27416_, _12226_, _13004_);
  nor _77516_ (_27417_, _27416_, _27415_);
  nor _77517_ (_27418_, _27417_, _06921_);
  or _77518_ (_27419_, _27418_, _27414_);
  and _77519_ (_27420_, _27419_, _13030_);
  nor _77520_ (_27421_, _27107_, _13030_);
  or _77521_ (_27423_, _27421_, _27420_);
  nand _77522_ (_27424_, _27423_, _06926_);
  and _77523_ (_27425_, _12440_, _06568_);
  nor _77524_ (_27426_, _27425_, _13038_);
  nand _77525_ (_27427_, _27426_, _27424_);
  nor _77526_ (_27428_, _27110_, _13037_);
  nor _77527_ (_27429_, _27428_, _07695_);
  and _77528_ (_27430_, _27429_, _27427_);
  or _77529_ (_27431_, _27430_, _27109_);
  nand _77530_ (_27432_, _27431_, _05928_);
  nor _77531_ (_27434_, _27417_, _05928_);
  nor _77532_ (_27435_, _27434_, _13053_);
  nand _77533_ (_27436_, _27435_, _27432_);
  nor _77534_ (_27437_, _27110_, _13052_);
  nor _77535_ (_27438_, _27437_, _06278_);
  nand _77536_ (_27439_, _27438_, _27436_);
  and _77537_ (_27440_, _12440_, _06278_);
  nor _77538_ (_27441_, _27440_, _13059_);
  nand _77539_ (_27442_, _27441_, _27439_);
  nor _77540_ (_27443_, _27110_, _12141_);
  nor _77541_ (_27445_, _27443_, _25301_);
  nand _77542_ (_27446_, _27445_, _27442_);
  and _77543_ (_27447_, _25301_, _08857_);
  nor _77544_ (_27448_, _27447_, _13068_);
  and _77545_ (_27449_, _27448_, _27446_);
  or _77546_ (_27450_, _27449_, _27108_);
  or _77547_ (_27451_, _27450_, _01351_);
  or _77548_ (_27452_, _01347_, \oc8051_golden_model_1.PC [6]);
  and _77549_ (_27453_, _27452_, _42618_);
  and _77550_ (_43252_, _27453_, _27451_);
  and _77551_ (_27455_, _08661_, _06278_);
  and _77552_ (_27456_, _27104_, \oc8051_golden_model_1.PC [7]);
  nor _77553_ (_27457_, _27104_, \oc8051_golden_model_1.PC [7]);
  nor _77554_ (_27458_, _27457_, _27456_);
  nor _77555_ (_27459_, _27458_, _12151_);
  nor _77556_ (_27460_, _27458_, _12154_);
  nor _77557_ (_27461_, _27458_, _12162_);
  nor _77558_ (_27462_, _27458_, _10979_);
  nor _77559_ (_27463_, _27458_, _12169_);
  nor _77560_ (_27464_, _09030_, _08661_);
  nor _77561_ (_27466_, _27458_, _12639_);
  nor _77562_ (_27467_, _25322_, _08661_);
  or _77563_ (_27468_, _12534_, _09415_);
  or _77564_ (_27469_, _12221_, _12222_);
  and _77565_ (_27470_, _27469_, _12271_);
  nor _77566_ (_27471_, _27469_, _12271_);
  nor _77567_ (_27472_, _27471_, _27470_);
  or _77568_ (_27473_, _27472_, _12536_);
  and _77569_ (_27474_, _27473_, _27468_);
  or _77570_ (_27475_, _27474_, _07151_);
  and _77571_ (_27477_, _12507_, _08661_);
  and _77572_ (_27478_, _12478_, _12436_);
  nor _77573_ (_27479_, _27478_, _12479_);
  and _77574_ (_27480_, _27479_, _12393_);
  nor _77575_ (_27481_, _27480_, _27477_);
  nand _77576_ (_27482_, _27481_, _12387_);
  nor _77577_ (_27483_, _07486_, \oc8051_golden_model_1.PC [7]);
  nor _77578_ (_27484_, _27483_, _07141_);
  and _77579_ (_27485_, _08661_, _07141_);
  nor _77580_ (_27486_, _27485_, _06781_);
  not _77581_ (_27488_, _27486_);
  nor _77582_ (_27489_, _27488_, _27484_);
  not _77583_ (_27490_, _27489_);
  nor _77584_ (_27491_, _27458_, _12513_);
  nor _77585_ (_27492_, _27491_, _06758_);
  and _77586_ (_27493_, _27492_, _27490_);
  nor _77587_ (_27494_, _08608_, _07504_);
  or _77588_ (_27495_, _27494_, _12516_);
  nor _77589_ (_27496_, _27495_, _27493_);
  nor _77590_ (_27497_, _27458_, _12512_);
  nor _77591_ (_27499_, _27497_, _27496_);
  nor _77592_ (_27500_, _27499_, _12387_);
  nor _77593_ (_27501_, _27500_, _07154_);
  and _77594_ (_27502_, _27501_, _27482_);
  and _77595_ (_27503_, _27458_, _07154_);
  or _77596_ (_27504_, _27503_, _06341_);
  or _77597_ (_27505_, _27504_, _27502_);
  nand _77598_ (_27506_, _27505_, _27475_);
  nand _77599_ (_27507_, _27506_, _12541_);
  nor _77600_ (_27508_, _27458_, _12541_);
  nor _77601_ (_27510_, _27508_, _06272_);
  nand _77602_ (_27511_, _27510_, _27507_);
  and _77603_ (_27512_, _08661_, _06272_);
  nor _77604_ (_27513_, _27512_, _07611_);
  nand _77605_ (_27514_, _27513_, _27511_);
  and _77606_ (_27515_, _08608_, _07611_);
  nor _77607_ (_27516_, _27515_, _06461_);
  nand _77608_ (_27517_, _27516_, _27514_);
  and _77609_ (_27518_, _08661_, _06461_);
  nor _77610_ (_27519_, _27518_, _12551_);
  nand _77611_ (_27521_, _27519_, _27517_);
  nor _77612_ (_27522_, _27458_, _12550_);
  nor _77613_ (_27523_, _27522_, _06464_);
  nand _77614_ (_27524_, _27523_, _27521_);
  and _77615_ (_27525_, _08661_, _06464_);
  nor _77616_ (_27526_, _27525_, _25401_);
  nand _77617_ (_27527_, _27526_, _27524_);
  nor _77618_ (_27528_, _27458_, _12560_);
  nor _77619_ (_27529_, _27528_, _06268_);
  nand _77620_ (_27530_, _27529_, _27527_);
  and _77621_ (_27532_, _08661_, _06268_);
  nor _77622_ (_27533_, _27532_, _12563_);
  nand _77623_ (_27534_, _27533_, _27530_);
  and _77624_ (_27535_, _08608_, _12563_);
  nor _77625_ (_27536_, _27535_, _06267_);
  nand _77626_ (_27537_, _27536_, _27534_);
  and _77627_ (_27538_, _08661_, _06267_);
  nor _77628_ (_27539_, _27538_, _12379_);
  nand _77629_ (_27540_, _27539_, _27537_);
  and _77630_ (_27541_, _12371_, _09415_);
  not _77631_ (_27543_, _27472_);
  nor _77632_ (_27544_, _27543_, _12371_);
  or _77633_ (_27545_, _27544_, _12378_);
  nor _77634_ (_27546_, _27545_, _27541_);
  nor _77635_ (_27547_, _27546_, _06347_);
  nand _77636_ (_27548_, _27547_, _27540_);
  or _77637_ (_27549_, _27543_, _12333_);
  or _77638_ (_27550_, _12335_, _09416_);
  nand _77639_ (_27551_, _27550_, _27549_);
  nand _77640_ (_27552_, _27551_, _06347_);
  and _77641_ (_27554_, _27552_, _06774_);
  and _77642_ (_27555_, _27554_, _27548_);
  and _77643_ (_27556_, _12587_, _09415_);
  nor _77644_ (_27557_, _27543_, _12587_);
  or _77645_ (_27558_, _27557_, _06774_);
  nor _77646_ (_27559_, _27558_, _27556_);
  or _77647_ (_27560_, _27559_, _06371_);
  or _77648_ (_27561_, _27560_, _27555_);
  nand _77649_ (_27562_, _12604_, _09415_);
  nand _77650_ (_27563_, _27472_, _26518_);
  and _77651_ (_27565_, _27563_, _27562_);
  or _77652_ (_27566_, _27565_, _12176_);
  and _77653_ (_27567_, _27566_, _27561_);
  or _77654_ (_27568_, _27567_, _12174_);
  nand _77655_ (_27569_, _27458_, _12174_);
  and _77656_ (_27570_, _27569_, _27568_);
  nand _77657_ (_27571_, _27570_, _06262_);
  and _77658_ (_27572_, _08794_, _06261_);
  nor _77659_ (_27573_, _27572_, _12613_);
  nand _77660_ (_27574_, _27573_, _27571_);
  nor _77661_ (_27576_, _08608_, _06007_);
  nor _77662_ (_27577_, _27576_, _25445_);
  and _77663_ (_27578_, _27577_, _27574_);
  or _77664_ (_27579_, _27578_, _27467_);
  nand _77665_ (_27580_, _27579_, _12630_);
  nor _77666_ (_27581_, _27458_, _12630_);
  nor _77667_ (_27582_, _27581_, _06505_);
  nand _77668_ (_27583_, _27582_, _27580_);
  and _77669_ (_27584_, _08661_, _06505_);
  nor _77670_ (_27585_, _27584_, _25158_);
  nand _77671_ (_27587_, _27585_, _27583_);
  and _77672_ (_27588_, _08608_, _25158_);
  nor _77673_ (_27589_, _27588_, _06504_);
  nand _77674_ (_27590_, _27589_, _27587_);
  and _77675_ (_27591_, _08661_, _06504_);
  nor _77676_ (_27592_, _27591_, _26197_);
  and _77677_ (_27593_, _27592_, _27590_);
  or _77678_ (_27594_, _27593_, _27466_);
  nand _77679_ (_27595_, _27594_, _12643_);
  nor _77680_ (_27596_, _12643_, _08661_);
  nor _77681_ (_27598_, _27596_, _10515_);
  nand _77682_ (_27599_, _27598_, _27595_);
  not _77683_ (_27600_, _27458_);
  nor _77684_ (_27601_, _27600_, _05984_);
  nor _77685_ (_27602_, _27601_, _06257_);
  and _77686_ (_27603_, _27602_, _27599_);
  and _77687_ (_27604_, _08794_, _06257_);
  or _77688_ (_27605_, _27604_, _27603_);
  nand _77689_ (_27606_, _27605_, _05978_);
  and _77690_ (_27607_, _08608_, _06254_);
  nor _77691_ (_27609_, _27607_, _06373_);
  nand _77692_ (_27610_, _27609_, _27606_);
  and _77693_ (_27611_, _09415_, _06373_);
  nor _77694_ (_27612_, _27611_, _12659_);
  nand _77695_ (_27613_, _27612_, _27610_);
  nor _77696_ (_27614_, _08661_, _07216_);
  nor _77697_ (_27615_, _27614_, _10094_);
  nand _77698_ (_27616_, _27615_, _27613_);
  nor _77699_ (_27617_, _09416_, _05982_);
  nor _77700_ (_27618_, _27617_, _25492_);
  nand _77701_ (_27620_, _27618_, _27616_);
  nor _77702_ (_27621_, _27458_, _12172_);
  nor _77703_ (_27622_, _27621_, _06323_);
  nand _77704_ (_27623_, _27622_, _27620_);
  and _77705_ (_27624_, _08661_, _06323_);
  nor _77706_ (_27625_, _27624_, _12668_);
  nand _77707_ (_27626_, _27625_, _27623_);
  and _77708_ (_27627_, _08608_, _12668_);
  nor _77709_ (_27628_, _27627_, _12674_);
  nand _77710_ (_27629_, _27628_, _27626_);
  and _77711_ (_27631_, _27479_, _12674_);
  nor _77712_ (_27632_, _27631_, _09031_);
  and _77713_ (_27633_, _27632_, _27629_);
  or _77714_ (_27634_, _27633_, _27464_);
  nand _77715_ (_27635_, _27634_, _06219_);
  and _77716_ (_27636_, _09416_, _06218_);
  nor _77717_ (_27637_, _27636_, _10929_);
  nand _77718_ (_27638_, _27637_, _27635_);
  and _77719_ (_27639_, _10929_, _08661_);
  nor _77720_ (_27640_, _27639_, _12690_);
  nand _77721_ (_27642_, _27640_, _27638_);
  or _77722_ (_27643_, _12695_, _12694_);
  not _77723_ (_27644_, _27643_);
  and _77724_ (_27645_, _27644_, _12715_);
  nor _77725_ (_27646_, _27644_, _12715_);
  nor _77726_ (_27647_, _27646_, _27645_);
  and _77727_ (_27648_, _27647_, _12690_);
  nor _77728_ (_27649_, _27648_, _06322_);
  nand _77729_ (_27650_, _27649_, _27642_);
  and _77730_ (_27651_, _08661_, _06322_);
  nor _77731_ (_27653_, _27651_, _06217_);
  nand _77732_ (_27654_, _27653_, _27650_);
  and _77733_ (_27655_, _08608_, _06217_);
  nor _77734_ (_27656_, _27655_, _12733_);
  nand _77735_ (_27657_, _27656_, _27654_);
  and _77736_ (_27658_, _11342_, _08661_);
  and _77737_ (_27659_, _27479_, _12759_);
  or _77738_ (_27660_, _27659_, _27658_);
  and _77739_ (_27661_, _27660_, _12733_);
  nor _77740_ (_27662_, _27661_, _12737_);
  and _77741_ (_27664_, _27662_, _27657_);
  or _77742_ (_27665_, _27664_, _27463_);
  nand _77743_ (_27666_, _27665_, _12166_);
  nor _77744_ (_27667_, _12166_, _08661_);
  nor _77745_ (_27668_, _27667_, _06369_);
  nand _77746_ (_27669_, _27668_, _27666_);
  and _77747_ (_27670_, _09415_, _06369_);
  nor _77748_ (_27671_, _27670_, _06536_);
  and _77749_ (_27672_, _27671_, _27669_);
  and _77750_ (_27673_, _08794_, _06536_);
  or _77751_ (_27675_, _27673_, _27672_);
  nand _77752_ (_27676_, _27675_, _05955_);
  and _77753_ (_27677_, _08608_, _12750_);
  nor _77754_ (_27678_, _27677_, _12755_);
  nand _77755_ (_27679_, _27678_, _27676_);
  nor _77756_ (_27680_, _11342_, _08794_);
  and _77757_ (_27681_, _27479_, _11342_);
  or _77758_ (_27682_, _27681_, _27680_);
  and _77759_ (_27683_, _27682_, _12755_);
  nor _77760_ (_27684_, _27683_, _10980_);
  and _77761_ (_27686_, _27684_, _27679_);
  or _77762_ (_27687_, _27686_, _27462_);
  nand _77763_ (_27688_, _27687_, _12164_);
  nor _77764_ (_27689_, _12164_, _08661_);
  nor _77765_ (_27690_, _27689_, _06375_);
  nand _77766_ (_27691_, _27690_, _27688_);
  and _77767_ (_27692_, _09415_, _06375_);
  nor _77768_ (_27693_, _27692_, _06545_);
  and _77769_ (_27694_, _27693_, _27691_);
  and _77770_ (_27695_, _08794_, _06545_);
  or _77771_ (_27697_, _27695_, _27694_);
  nand _77772_ (_27698_, _27697_, _05961_);
  and _77773_ (_27699_, _08608_, _07233_);
  nor _77774_ (_27700_, _27699_, _12776_);
  nand _77775_ (_27701_, _27700_, _27698_);
  nor _77776_ (_27702_, _27479_, \oc8051_golden_model_1.PSW [7]);
  nor _77777_ (_27703_, _08661_, _10558_);
  nor _77778_ (_27704_, _27703_, _12782_);
  not _77779_ (_27705_, _27704_);
  nor _77780_ (_27706_, _27705_, _27702_);
  nor _77781_ (_27708_, _27706_, _12780_);
  and _77782_ (_27709_, _27708_, _27701_);
  or _77783_ (_27710_, _27709_, _27461_);
  nand _77784_ (_27711_, _27710_, _11022_);
  nor _77785_ (_27712_, _11022_, _08661_);
  nor _77786_ (_27713_, _27712_, _06366_);
  nand _77787_ (_27714_, _27713_, _27711_);
  and _77788_ (_27715_, _09415_, _06366_);
  nor _77789_ (_27716_, _27715_, _06528_);
  and _77790_ (_27717_, _27716_, _27714_);
  and _77791_ (_27719_, _08794_, _06528_);
  or _77792_ (_27720_, _27719_, _27717_);
  nand _77793_ (_27721_, _27720_, _05966_);
  and _77794_ (_27722_, _08608_, _12795_);
  nor _77795_ (_27723_, _27722_, _12800_);
  nand _77796_ (_27724_, _27723_, _27721_);
  and _77797_ (_27725_, _08661_, _10558_);
  and _77798_ (_27726_, _27479_, \oc8051_golden_model_1.PSW [7]);
  or _77799_ (_27727_, _27726_, _27725_);
  and _77800_ (_27728_, _27727_, _12800_);
  nor _77801_ (_27730_, _27728_, _12804_);
  and _77802_ (_27731_, _27730_, _27724_);
  or _77803_ (_27732_, _27731_, _27460_);
  nand _77804_ (_27733_, _27732_, _12153_);
  nor _77805_ (_27734_, _12153_, _08661_);
  nor _77806_ (_27735_, _27734_, _11125_);
  nand _77807_ (_27736_, _27735_, _27733_);
  and _77808_ (_27737_, _27458_, _11125_);
  nor _77809_ (_27738_, _27737_, _06551_);
  and _77810_ (_27739_, _27738_, _27736_);
  nor _77811_ (_27741_, _08755_, _06716_);
  or _77812_ (_27742_, _27741_, _27739_);
  nand _77813_ (_27743_, _27742_, _05959_);
  and _77814_ (_27744_, _08608_, _07253_);
  nor _77815_ (_27745_, _27744_, _06365_);
  nand _77816_ (_27746_, _27745_, _27743_);
  and _77817_ (_27747_, _27543_, _13004_);
  nor _77818_ (_27748_, _09415_, _13004_);
  or _77819_ (_27749_, _27748_, _06558_);
  or _77820_ (_27750_, _27749_, _27747_);
  and _77821_ (_27752_, _27750_, _12151_);
  and _77822_ (_27753_, _27752_, _27746_);
  or _77823_ (_27754_, _27753_, _27459_);
  nand _77824_ (_27755_, _27754_, _13012_);
  nor _77825_ (_27756_, _13012_, _08661_);
  nor _77826_ (_27757_, _27756_, _11284_);
  nand _77827_ (_27758_, _27757_, _27755_);
  and _77828_ (_27759_, _27458_, _11284_);
  nor _77829_ (_27760_, _27759_, _06281_);
  and _77830_ (_27761_, _27760_, _27758_);
  nor _77831_ (_27763_, _08755_, _06282_);
  or _77832_ (_27764_, _27763_, _27761_);
  nand _77833_ (_27765_, _27764_, _05964_);
  and _77834_ (_27766_, _08608_, _25646_);
  nor _77835_ (_27767_, _27766_, _06362_);
  nand _77836_ (_27768_, _27767_, _27765_);
  and _77837_ (_27769_, _09416_, _13004_);
  nor _77838_ (_27770_, _27472_, _13004_);
  nor _77839_ (_27771_, _27770_, _27769_);
  and _77840_ (_27772_, _27771_, _06362_);
  nor _77841_ (_27774_, _27772_, _13031_);
  nand _77842_ (_27775_, _27774_, _27768_);
  nor _77843_ (_27776_, _27458_, _13030_);
  nor _77844_ (_27777_, _27776_, _06568_);
  nand _77845_ (_27778_, _27777_, _27775_);
  and _77846_ (_27779_, _08661_, _06568_);
  nor _77847_ (_27780_, _27779_, _13038_);
  and _77848_ (_27781_, _27780_, _27778_);
  nor _77849_ (_27782_, _27458_, _13037_);
  or _77850_ (_27783_, _27782_, _27781_);
  nand _77851_ (_27785_, _27783_, _07271_);
  and _77852_ (_27786_, _08608_, _07695_);
  nor _77853_ (_27787_, _27786_, _05927_);
  nand _77854_ (_27788_, _27787_, _27785_);
  and _77855_ (_27789_, _27771_, _05927_);
  nor _77856_ (_27790_, _27789_, _13053_);
  nand _77857_ (_27791_, _27790_, _27788_);
  nor _77858_ (_27792_, _27458_, _13052_);
  nor _77859_ (_27793_, _27792_, _06278_);
  and _77860_ (_27794_, _27793_, _27791_);
  or _77861_ (_27796_, _27794_, _27455_);
  nand _77862_ (_27797_, _27796_, _12141_);
  nor _77863_ (_27798_, _27600_, _12141_);
  nor _77864_ (_27799_, _27798_, _25301_);
  nand _77865_ (_27800_, _27799_, _27797_);
  and _77866_ (_27801_, _25301_, _08608_);
  nor _77867_ (_27802_, _27801_, _13068_);
  and _77868_ (_27803_, _27802_, _27800_);
  and _77869_ (_27804_, _27458_, _13068_);
  or _77870_ (_27805_, _27804_, _27803_);
  or _77871_ (_27807_, _27805_, _01351_);
  or _77872_ (_27808_, _01347_, \oc8051_golden_model_1.PC [7]);
  and _77873_ (_27809_, _27808_, _42618_);
  and _77874_ (_43253_, _27809_, _27807_);
  nor _77875_ (_27810_, _12140_, _06251_);
  nor _77876_ (_27811_, _14508_, _06251_);
  and _77877_ (_27812_, _27456_, \oc8051_golden_model_1.PC [8]);
  nor _77878_ (_27813_, _27456_, \oc8051_golden_model_1.PC [8]);
  nor _77879_ (_27814_, _27813_, _27812_);
  nor _77880_ (_27815_, _27814_, _12151_);
  nor _77881_ (_27817_, _27814_, _12154_);
  nor _77882_ (_27818_, _27814_, _12162_);
  nor _77883_ (_27819_, _27814_, _10979_);
  and _77884_ (_27820_, _12275_, _06369_);
  nor _77885_ (_27821_, _27814_, _12169_);
  nor _77886_ (_27822_, _12431_, _09030_);
  and _77887_ (_27823_, _12431_, _06323_);
  nor _77888_ (_27824_, _25322_, _12431_);
  and _77889_ (_27825_, _12431_, _06268_);
  or _77890_ (_27826_, _06461_, _07611_);
  nand _77891_ (_27828_, _12431_, _06272_);
  and _77892_ (_27829_, _12536_, _12276_);
  nor _77893_ (_27830_, _12279_, _12273_);
  nor _77894_ (_27831_, _27830_, _12280_);
  not _77895_ (_27832_, _27831_);
  and _77896_ (_27833_, _27832_, _12534_);
  or _77897_ (_27834_, _27833_, _27829_);
  and _77898_ (_27835_, _27834_, _06341_);
  not _77899_ (_27836_, _12431_);
  or _77900_ (_27837_, _12393_, _27836_);
  and _77901_ (_27839_, _12483_, _12480_);
  nor _77902_ (_27840_, _27839_, _12484_);
  nand _77903_ (_27841_, _27840_, _12393_);
  and _77904_ (_27842_, _27841_, _27837_);
  and _77905_ (_27843_, _27842_, _12387_);
  nand _77906_ (_27844_, _12431_, _07141_);
  nand _77907_ (_27845_, _07142_, \oc8051_golden_model_1.PC [8]);
  or _77908_ (_27846_, _27845_, _07486_);
  and _77909_ (_27847_, _27846_, _27844_);
  or _77910_ (_27848_, _27847_, _06781_);
  and _77911_ (_27850_, _27848_, _07504_);
  or _77912_ (_27851_, _27850_, _12516_);
  not _77913_ (_27852_, _27814_);
  or _77914_ (_27853_, _27852_, _12514_);
  and _77915_ (_27854_, _27853_, _08654_);
  and _77916_ (_27855_, _27854_, _27851_);
  or _77917_ (_27856_, _27855_, _07154_);
  or _77918_ (_27857_, _27856_, _27843_);
  nand _77919_ (_27858_, _27814_, _07154_);
  and _77920_ (_27859_, _27858_, _07151_);
  and _77921_ (_27861_, _27859_, _27857_);
  or _77922_ (_27862_, _27861_, _27835_);
  and _77923_ (_27863_, _27862_, _12541_);
  nor _77924_ (_27864_, _27814_, _12541_);
  or _77925_ (_27865_, _27864_, _06272_);
  or _77926_ (_27866_, _27865_, _27863_);
  and _77927_ (_27867_, _27866_, _27828_);
  nor _77928_ (_27868_, _27867_, _27826_);
  and _77929_ (_27869_, _12431_, _06461_);
  nor _77930_ (_27870_, _27869_, _12551_);
  not _77931_ (_27871_, _27870_);
  nor _77932_ (_27872_, _27871_, _27868_);
  nor _77933_ (_27873_, _27814_, _12550_);
  nor _77934_ (_27874_, _27873_, _06464_);
  not _77935_ (_27875_, _27874_);
  nor _77936_ (_27876_, _27875_, _27872_);
  and _77937_ (_27877_, _12431_, _06464_);
  nor _77938_ (_27878_, _27877_, _25401_);
  not _77939_ (_27879_, _27878_);
  or _77940_ (_27880_, _27879_, _27876_);
  nor _77941_ (_27883_, _27814_, _12560_);
  nor _77942_ (_27884_, _27883_, _06268_);
  and _77943_ (_27885_, _27884_, _27880_);
  or _77944_ (_27886_, _27885_, _27825_);
  nand _77945_ (_27887_, _27886_, _12564_);
  and _77946_ (_27888_, _12431_, _06267_);
  nor _77947_ (_27889_, _27888_, _12379_);
  nand _77948_ (_27890_, _27889_, _27887_);
  and _77949_ (_27891_, _12371_, _12275_);
  nor _77950_ (_27892_, _27832_, _12371_);
  or _77951_ (_27894_, _27892_, _27891_);
  nor _77952_ (_27895_, _27894_, _12378_);
  nor _77953_ (_27896_, _27895_, _06347_);
  nand _77954_ (_27897_, _27896_, _27890_);
  and _77955_ (_27898_, _27831_, _12335_);
  and _77956_ (_27899_, _12333_, _12275_);
  nor _77957_ (_27900_, _27899_, _27898_);
  nor _77958_ (_27901_, _27900_, _12177_);
  nor _77959_ (_27902_, _27901_, _06480_);
  nand _77960_ (_27903_, _27902_, _27897_);
  and _77961_ (_27905_, _12587_, _12275_);
  not _77962_ (_27906_, _27905_);
  nor _77963_ (_27907_, _27832_, _12587_);
  nor _77964_ (_27908_, _27907_, _06774_);
  and _77965_ (_27909_, _27908_, _27906_);
  nor _77966_ (_27910_, _27909_, _06371_);
  nand _77967_ (_27911_, _27910_, _27903_);
  and _77968_ (_27912_, _12604_, _12275_);
  and _77969_ (_27913_, _27831_, _26518_);
  or _77970_ (_27914_, _27913_, _27912_);
  and _77971_ (_27916_, _27914_, _06371_);
  nor _77972_ (_27917_, _27916_, _12174_);
  nand _77973_ (_27918_, _27917_, _27911_);
  and _77974_ (_27919_, _27852_, _12174_);
  nor _77975_ (_27920_, _27919_, _06261_);
  nand _77976_ (_27921_, _27920_, _27918_);
  and _77977_ (_27922_, _12431_, _06261_);
  not _77978_ (_27923_, _27922_);
  and _77979_ (_27924_, _25322_, _06007_);
  and _77980_ (_27925_, _27924_, _27923_);
  and _77981_ (_27927_, _27925_, _27921_);
  or _77982_ (_27928_, _27927_, _27824_);
  nand _77983_ (_27929_, _27928_, _12630_);
  nor _77984_ (_27930_, _27814_, _12630_);
  nor _77985_ (_27931_, _27930_, _06505_);
  nand _77986_ (_27932_, _27931_, _27929_);
  and _77987_ (_27933_, _12431_, _06505_);
  nor _77988_ (_27934_, _27933_, _25158_);
  nand _77989_ (_27935_, _27934_, _27932_);
  nand _77990_ (_27936_, _27935_, _14057_);
  and _77991_ (_27938_, _12431_, _06504_);
  nor _77992_ (_27939_, _27938_, _26197_);
  and _77993_ (_27940_, _27939_, _27936_);
  nor _77994_ (_27941_, _27814_, _12639_);
  or _77995_ (_27942_, _27941_, _27940_);
  nand _77996_ (_27943_, _27942_, _12643_);
  nor _77997_ (_27944_, _12431_, _12643_);
  nor _77998_ (_27945_, _27944_, _10515_);
  nand _77999_ (_27946_, _27945_, _27943_);
  nor _78000_ (_27947_, _27852_, _05984_);
  nor _78001_ (_27949_, _27947_, _06257_);
  nand _78002_ (_27950_, _27949_, _27946_);
  nor _78003_ (_27951_, _06373_, _06254_);
  not _78004_ (_27952_, _27951_);
  and _78005_ (_27953_, _27836_, _06257_);
  nor _78006_ (_27954_, _27953_, _27952_);
  nand _78007_ (_27955_, _27954_, _27950_);
  and _78008_ (_27956_, _12275_, _06373_);
  nor _78009_ (_27957_, _27956_, _12659_);
  nand _78010_ (_27958_, _27957_, _27955_);
  nor _78011_ (_27960_, _12431_, _07216_);
  nor _78012_ (_27961_, _27960_, _10094_);
  nand _78013_ (_27962_, _27961_, _27958_);
  nor _78014_ (_27963_, _12276_, _05982_);
  nor _78015_ (_27964_, _27963_, _25492_);
  nand _78016_ (_27965_, _27964_, _27962_);
  nor _78017_ (_27966_, _27814_, _12172_);
  nor _78018_ (_27967_, _27966_, _06323_);
  and _78019_ (_27968_, _27967_, _27965_);
  or _78020_ (_27969_, _27968_, _27823_);
  nor _78021_ (_27971_, _12674_, _12668_);
  nand _78022_ (_27972_, _27971_, _27969_);
  and _78023_ (_27973_, _27840_, _12674_);
  nor _78024_ (_27974_, _27973_, _09031_);
  and _78025_ (_27975_, _27974_, _27972_);
  or _78026_ (_27976_, _27975_, _27822_);
  nand _78027_ (_27977_, _27976_, _06219_);
  and _78028_ (_27978_, _12276_, _06218_);
  nor _78029_ (_27979_, _27978_, _10929_);
  nand _78030_ (_27980_, _27979_, _27977_);
  and _78031_ (_27982_, _12431_, _10929_);
  nor _78032_ (_27983_, _27982_, _12690_);
  nand _78033_ (_27984_, _27983_, _27980_);
  and _78034_ (_27985_, _12717_, _12693_);
  nor _78035_ (_27986_, _27985_, _12718_);
  nor _78036_ (_27987_, _27986_, _12691_);
  nor _78037_ (_27988_, _27987_, _06322_);
  nand _78038_ (_27989_, _27988_, _27984_);
  and _78039_ (_27990_, _12431_, _06322_);
  nor _78040_ (_27991_, _27990_, _06217_);
  nand _78041_ (_27993_, _27991_, _27989_);
  nand _78042_ (_27994_, _27993_, _25064_);
  and _78043_ (_27995_, _12431_, _11342_);
  and _78044_ (_27996_, _27840_, _12759_);
  or _78045_ (_27997_, _27996_, _27995_);
  and _78046_ (_27998_, _27997_, _12733_);
  nor _78047_ (_27999_, _27998_, _12737_);
  and _78048_ (_28000_, _27999_, _27994_);
  or _78049_ (_28001_, _28000_, _27821_);
  nand _78050_ (_28002_, _28001_, _12166_);
  nor _78051_ (_28004_, _12431_, _12166_);
  nor _78052_ (_28005_, _28004_, _06369_);
  and _78053_ (_28006_, _28005_, _28002_);
  or _78054_ (_28007_, _28006_, _27820_);
  nand _78055_ (_28008_, _28007_, _07240_);
  and _78056_ (_28009_, _12431_, _06536_);
  nor _78057_ (_28010_, _28009_, _12750_);
  nand _78058_ (_28011_, _28010_, _28008_);
  nand _78059_ (_28012_, _28011_, _25061_);
  nor _78060_ (_28013_, _27836_, _11342_);
  and _78061_ (_28015_, _27840_, _11342_);
  or _78062_ (_28016_, _28015_, _28013_);
  and _78063_ (_28017_, _28016_, _12755_);
  nor _78064_ (_28018_, _28017_, _10980_);
  and _78065_ (_28019_, _28018_, _28012_);
  or _78066_ (_28020_, _28019_, _27819_);
  nand _78067_ (_28021_, _28020_, _12164_);
  nor _78068_ (_28022_, _12164_, _12431_);
  nor _78069_ (_28023_, _28022_, _06375_);
  nand _78070_ (_28024_, _28023_, _28021_);
  and _78071_ (_28026_, _12275_, _06375_);
  nor _78072_ (_28027_, _28026_, _06545_);
  nand _78073_ (_28028_, _28027_, _28024_);
  nor _78074_ (_28029_, _12776_, _07233_);
  and _78075_ (_28030_, _27836_, _06545_);
  not _78076_ (_28031_, _28030_);
  and _78077_ (_28032_, _28031_, _28029_);
  nand _78078_ (_28033_, _28032_, _28028_);
  nor _78079_ (_28034_, _27840_, \oc8051_golden_model_1.PSW [7]);
  nor _78080_ (_28035_, _12431_, _10558_);
  nor _78081_ (_28037_, _28035_, _12782_);
  not _78082_ (_28038_, _28037_);
  nor _78083_ (_28039_, _28038_, _28034_);
  nor _78084_ (_28040_, _28039_, _12780_);
  and _78085_ (_28041_, _28040_, _28033_);
  or _78086_ (_28042_, _28041_, _27818_);
  nand _78087_ (_28043_, _28042_, _11022_);
  nor _78088_ (_28044_, _12431_, _11022_);
  nor _78089_ (_28045_, _28044_, _06366_);
  nand _78090_ (_28046_, _28045_, _28043_);
  and _78091_ (_28048_, _12275_, _06366_);
  nor _78092_ (_28049_, _28048_, _06528_);
  nand _78093_ (_28050_, _28049_, _28046_);
  nor _78094_ (_28051_, _12800_, _12795_);
  and _78095_ (_28052_, _27836_, _06528_);
  not _78096_ (_28053_, _28052_);
  and _78097_ (_28054_, _28053_, _28051_);
  nand _78098_ (_28055_, _28054_, _28050_);
  and _78099_ (_28056_, _12431_, _10558_);
  and _78100_ (_28057_, _27840_, \oc8051_golden_model_1.PSW [7]);
  or _78101_ (_28059_, _28057_, _28056_);
  and _78102_ (_28060_, _28059_, _12800_);
  nor _78103_ (_28061_, _28060_, _12804_);
  and _78104_ (_28062_, _28061_, _28055_);
  or _78105_ (_28063_, _28062_, _27817_);
  nand _78106_ (_28064_, _28063_, _12153_);
  nor _78107_ (_28065_, _12431_, _12153_);
  nor _78108_ (_28066_, _28065_, _11125_);
  and _78109_ (_28067_, _28066_, _28064_);
  and _78110_ (_28068_, _27814_, _11125_);
  or _78111_ (_28070_, _28068_, _28067_);
  nand _78112_ (_28071_, _28070_, _06716_);
  and _78113_ (_28072_, _07133_, _06551_);
  nor _78114_ (_28073_, _28072_, _07253_);
  nand _78115_ (_28074_, _28073_, _28071_);
  nand _78116_ (_28075_, _28074_, _06558_);
  and _78117_ (_28076_, _27832_, _13004_);
  nor _78118_ (_28077_, _12275_, _13004_);
  or _78119_ (_28078_, _28077_, _06558_);
  or _78120_ (_28079_, _28078_, _28076_);
  and _78121_ (_28081_, _28079_, _12151_);
  and _78122_ (_28082_, _28081_, _28075_);
  or _78123_ (_28083_, _28082_, _27815_);
  nand _78124_ (_28084_, _28083_, _13012_);
  nor _78125_ (_28085_, _13012_, _12431_);
  nor _78126_ (_28086_, _28085_, _11284_);
  and _78127_ (_28087_, _28086_, _28084_);
  and _78128_ (_28088_, _27814_, _11284_);
  or _78129_ (_28089_, _28088_, _28087_);
  nand _78130_ (_28090_, _28089_, _06282_);
  and _78131_ (_28092_, _07133_, _06281_);
  nor _78132_ (_28093_, _28092_, _25646_);
  nand _78133_ (_28094_, _28093_, _28090_);
  nand _78134_ (_28095_, _28094_, _06921_);
  and _78135_ (_28096_, _12276_, _13004_);
  nor _78136_ (_28097_, _27831_, _13004_);
  nor _78137_ (_28098_, _28097_, _28096_);
  and _78138_ (_28099_, _28098_, _06362_);
  nor _78139_ (_28100_, _28099_, _13031_);
  nand _78140_ (_28101_, _28100_, _28095_);
  nor _78141_ (_28103_, _27814_, _13030_);
  nor _78142_ (_28104_, _28103_, _06568_);
  nand _78143_ (_28105_, _28104_, _28101_);
  and _78144_ (_28106_, _12431_, _06568_);
  nor _78145_ (_28107_, _28106_, _13038_);
  nand _78146_ (_28108_, _28107_, _28105_);
  nor _78147_ (_28109_, _27814_, _13037_);
  nor _78148_ (_28110_, _28109_, _06361_);
  and _78149_ (_28111_, _28110_, _28108_);
  or _78150_ (_28112_, _28111_, _27811_);
  nor _78151_ (_28114_, _05940_, _05927_);
  nand _78152_ (_28115_, _28114_, _28112_);
  and _78153_ (_28116_, _28098_, _05927_);
  nor _78154_ (_28117_, _28116_, _13053_);
  nand _78155_ (_28118_, _28117_, _28115_);
  nor _78156_ (_28119_, _27814_, _13052_);
  nor _78157_ (_28120_, _28119_, _06278_);
  nand _78158_ (_28121_, _28120_, _28118_);
  and _78159_ (_28122_, _12431_, _06278_);
  nor _78160_ (_28123_, _28122_, _13059_);
  nand _78161_ (_28125_, _28123_, _28121_);
  nor _78162_ (_28126_, _27814_, _12141_);
  nor _78163_ (_28127_, _28126_, _06379_);
  and _78164_ (_28128_, _28127_, _28125_);
  or _78165_ (_28129_, _28128_, _27810_);
  nor _78166_ (_28130_, _13068_, _05939_);
  and _78167_ (_28131_, _28130_, _28129_);
  and _78168_ (_28132_, _27814_, _13068_);
  or _78169_ (_28133_, _28132_, _28131_);
  or _78170_ (_28134_, _28133_, _01351_);
  or _78171_ (_28136_, _01347_, \oc8051_golden_model_1.PC [8]);
  and _78172_ (_28137_, _28136_, _42618_);
  and _78173_ (_43254_, _28137_, _28134_);
  nor _78174_ (_28138_, _07004_, _12140_);
  nor _78175_ (_28139_, _07004_, _14508_);
  and _78176_ (_28140_, _27812_, \oc8051_golden_model_1.PC [9]);
  nor _78177_ (_28141_, _27812_, \oc8051_golden_model_1.PC [9]);
  nor _78178_ (_28142_, _28141_, _28140_);
  nor _78179_ (_28143_, _28142_, _12151_);
  nor _78180_ (_28144_, _28142_, _12154_);
  and _78181_ (_28146_, _12216_, _06366_);
  nor _78182_ (_28147_, _28142_, _12162_);
  and _78183_ (_28148_, _12216_, _06375_);
  nor _78184_ (_28149_, _28142_, _10979_);
  and _78185_ (_28150_, _12216_, _06369_);
  nor _78186_ (_28151_, _28142_, _12169_);
  nor _78187_ (_28152_, _12426_, _09030_);
  and _78188_ (_28153_, _12426_, _06323_);
  and _78189_ (_28154_, _12426_, _06504_);
  nor _78190_ (_28155_, _06504_, _25158_);
  not _78191_ (_28157_, _28142_);
  and _78192_ (_28158_, _28157_, _12174_);
  nor _78193_ (_28159_, _12280_, _12277_);
  and _78194_ (_28160_, _28159_, _12220_);
  nor _78195_ (_28161_, _28159_, _12220_);
  nor _78196_ (_28162_, _28161_, _28160_);
  and _78197_ (_28163_, _28162_, _12335_);
  and _78198_ (_28164_, _12333_, _12217_);
  nor _78199_ (_28165_, _28164_, _28163_);
  nor _78200_ (_28166_, _28165_, _12177_);
  nand _78201_ (_28168_, _12426_, _07141_);
  nand _78202_ (_28169_, _07142_, \oc8051_golden_model_1.PC [9]);
  or _78203_ (_28170_, _28169_, _07486_);
  and _78204_ (_28171_, _28170_, _28168_);
  or _78205_ (_28172_, _28171_, _06781_);
  and _78206_ (_28173_, _28172_, _07504_);
  or _78207_ (_28174_, _28173_, _12516_);
  or _78208_ (_28175_, _28157_, _12514_);
  and _78209_ (_28176_, _28175_, _08654_);
  and _78210_ (_28177_, _28176_, _28174_);
  and _78211_ (_28178_, _12507_, _12426_);
  or _78212_ (_28179_, _12427_, _12428_);
  not _78213_ (_28180_, _28179_);
  nor _78214_ (_28181_, _28180_, _12485_);
  and _78215_ (_28182_, _28180_, _12485_);
  nor _78216_ (_28183_, _28182_, _28181_);
  nor _78217_ (_28184_, _28183_, _12507_);
  nor _78218_ (_28185_, _28184_, _28178_);
  and _78219_ (_28186_, _28185_, _12387_);
  or _78220_ (_28187_, _28186_, _28177_);
  nand _78221_ (_28190_, _28187_, _07155_);
  and _78222_ (_28191_, _28157_, _07154_);
  nor _78223_ (_28192_, _28191_, _06341_);
  and _78224_ (_28193_, _28192_, _28190_);
  and _78225_ (_28194_, _28162_, _12534_);
  and _78226_ (_28195_, _12536_, _12217_);
  or _78227_ (_28196_, _28195_, _07151_);
  nor _78228_ (_28197_, _28196_, _28194_);
  or _78229_ (_28198_, _28197_, _12542_);
  or _78230_ (_28199_, _28198_, _28193_);
  nor _78231_ (_28201_, _28142_, _12541_);
  nor _78232_ (_28202_, _28201_, _06272_);
  nand _78233_ (_28203_, _28202_, _28199_);
  and _78234_ (_28204_, _12426_, _06272_);
  nor _78235_ (_28205_, _28204_, _07611_);
  nand _78236_ (_28206_, _28205_, _28203_);
  nand _78237_ (_28207_, _28206_, _07166_);
  and _78238_ (_28208_, _12426_, _06461_);
  nor _78239_ (_28209_, _28208_, _12551_);
  nand _78240_ (_28210_, _28209_, _28207_);
  nor _78241_ (_28212_, _28142_, _12550_);
  nor _78242_ (_28213_, _28212_, _06464_);
  nand _78243_ (_28214_, _28213_, _28210_);
  and _78244_ (_28215_, _12426_, _06464_);
  nor _78245_ (_28216_, _28215_, _25401_);
  nand _78246_ (_28217_, _28216_, _28214_);
  nor _78247_ (_28218_, _28142_, _12560_);
  nor _78248_ (_28219_, _28218_, _06268_);
  nand _78249_ (_28220_, _28219_, _28217_);
  and _78250_ (_28221_, _12426_, _06268_);
  nor _78251_ (_28223_, _28221_, _12563_);
  nand _78252_ (_28224_, _28223_, _28220_);
  nand _78253_ (_28225_, _28224_, _07303_);
  and _78254_ (_28226_, _12426_, _06267_);
  nor _78255_ (_28227_, _28226_, _12379_);
  and _78256_ (_28228_, _28227_, _28225_);
  and _78257_ (_28229_, _12371_, _12216_);
  nor _78258_ (_28230_, _28162_, _12371_);
  or _78259_ (_28231_, _28230_, _12378_);
  nor _78260_ (_28232_, _28231_, _28229_);
  or _78261_ (_28234_, _28232_, _28228_);
  and _78262_ (_28235_, _28234_, _12177_);
  or _78263_ (_28236_, _28235_, _28166_);
  or _78264_ (_28237_, _28236_, _06480_);
  nor _78265_ (_28238_, _28162_, _12587_);
  and _78266_ (_28239_, _12587_, _12216_);
  nor _78267_ (_28240_, _28239_, _28238_);
  or _78268_ (_28241_, _28240_, _06774_);
  and _78269_ (_28242_, _28241_, _28237_);
  or _78270_ (_28243_, _28242_, _06371_);
  and _78271_ (_28245_, _12604_, _12216_);
  nor _78272_ (_28246_, _28162_, _12604_);
  or _78273_ (_28247_, _28246_, _28245_);
  and _78274_ (_28248_, _28247_, _06371_);
  nor _78275_ (_28249_, _28248_, _12174_);
  and _78276_ (_28250_, _28249_, _28243_);
  or _78277_ (_28251_, _28250_, _28158_);
  nand _78278_ (_28252_, _28251_, _06262_);
  not _78279_ (_28253_, _12426_);
  and _78280_ (_28254_, _28253_, _06261_);
  not _78281_ (_28256_, _28254_);
  and _78282_ (_28257_, _28256_, _27924_);
  nand _78283_ (_28258_, _28257_, _28252_);
  nor _78284_ (_28259_, _25322_, _28253_);
  nor _78285_ (_28260_, _28259_, _12631_);
  nand _78286_ (_28261_, _28260_, _28258_);
  nor _78287_ (_28262_, _28142_, _12630_);
  nor _78288_ (_28263_, _28262_, _06505_);
  and _78289_ (_28264_, _28263_, _28261_);
  and _78290_ (_28265_, _12426_, _06505_);
  or _78291_ (_28267_, _28265_, _28264_);
  and _78292_ (_28268_, _28267_, _28155_);
  or _78293_ (_28269_, _28268_, _28154_);
  nand _78294_ (_28270_, _28269_, _12639_);
  nor _78295_ (_28271_, _28157_, _12639_);
  nor _78296_ (_28272_, _28271_, _12644_);
  nand _78297_ (_28273_, _28272_, _28270_);
  nor _78298_ (_28274_, _12426_, _12643_);
  nor _78299_ (_28275_, _28274_, _10515_);
  nand _78300_ (_28276_, _28275_, _28273_);
  nor _78301_ (_28278_, _28157_, _05984_);
  nor _78302_ (_28279_, _28278_, _06257_);
  nand _78303_ (_28280_, _28279_, _28276_);
  and _78304_ (_28281_, _28253_, _06257_);
  nor _78305_ (_28282_, _28281_, _27952_);
  nand _78306_ (_28283_, _28282_, _28280_);
  and _78307_ (_28284_, _12216_, _06373_);
  nor _78308_ (_28285_, _28284_, _12659_);
  nand _78309_ (_28286_, _28285_, _28283_);
  nor _78310_ (_28287_, _12426_, _07216_);
  nor _78311_ (_28289_, _28287_, _10094_);
  nand _78312_ (_28290_, _28289_, _28286_);
  nor _78313_ (_28291_, _12217_, _05982_);
  nor _78314_ (_28292_, _28291_, _25492_);
  nand _78315_ (_28293_, _28292_, _28290_);
  nor _78316_ (_28294_, _28142_, _12172_);
  nor _78317_ (_28295_, _28294_, _06323_);
  and _78318_ (_28296_, _28295_, _28293_);
  or _78319_ (_28297_, _28296_, _28153_);
  nand _78320_ (_28298_, _28297_, _27971_);
  nor _78321_ (_28300_, _28183_, _12679_);
  nor _78322_ (_28301_, _28300_, _09031_);
  and _78323_ (_28302_, _28301_, _28298_);
  or _78324_ (_28303_, _28302_, _28152_);
  nand _78325_ (_28304_, _28303_, _06219_);
  and _78326_ (_28305_, _12217_, _06218_);
  nor _78327_ (_28306_, _28305_, _10929_);
  nand _78328_ (_28307_, _28306_, _28304_);
  and _78329_ (_28308_, _12426_, _10929_);
  nor _78330_ (_28309_, _28308_, _12690_);
  nand _78331_ (_28311_, _28309_, _28307_);
  nor _78332_ (_28312_, _12718_, \oc8051_golden_model_1.DPH [1]);
  nor _78333_ (_28313_, _28312_, _12719_);
  nor _78334_ (_28314_, _28313_, _12691_);
  nor _78335_ (_28315_, _28314_, _06322_);
  nand _78336_ (_28316_, _28315_, _28311_);
  and _78337_ (_28317_, _12426_, _06322_);
  nor _78338_ (_28318_, _28317_, _06217_);
  nand _78339_ (_28319_, _28318_, _28316_);
  nand _78340_ (_28320_, _28319_, _25064_);
  and _78341_ (_28322_, _12426_, _11342_);
  nor _78342_ (_28323_, _28183_, _11342_);
  or _78343_ (_28324_, _28323_, _28322_);
  and _78344_ (_28325_, _28324_, _12733_);
  nor _78345_ (_28326_, _28325_, _12737_);
  and _78346_ (_28327_, _28326_, _28320_);
  or _78347_ (_28328_, _28327_, _28151_);
  nand _78348_ (_28329_, _28328_, _12166_);
  nor _78349_ (_28330_, _12426_, _12166_);
  nor _78350_ (_28331_, _28330_, _06369_);
  and _78351_ (_28333_, _28331_, _28329_);
  or _78352_ (_28334_, _28333_, _28150_);
  nand _78353_ (_28335_, _28334_, _07240_);
  and _78354_ (_28336_, _12426_, _06536_);
  nor _78355_ (_28337_, _28336_, _12750_);
  nand _78356_ (_28338_, _28337_, _28335_);
  nand _78357_ (_28339_, _28338_, _25061_);
  and _78358_ (_28340_, _28183_, _11342_);
  nor _78359_ (_28341_, _12426_, _11342_);
  nor _78360_ (_28342_, _28341_, _25061_);
  not _78361_ (_28344_, _28342_);
  nor _78362_ (_28345_, _28344_, _28340_);
  nor _78363_ (_28346_, _28345_, _10980_);
  and _78364_ (_28347_, _28346_, _28339_);
  or _78365_ (_28348_, _28347_, _28149_);
  nand _78366_ (_28349_, _28348_, _12164_);
  nor _78367_ (_28350_, _12164_, _12426_);
  nor _78368_ (_28351_, _28350_, _06375_);
  and _78369_ (_28352_, _28351_, _28349_);
  or _78370_ (_28353_, _28352_, _28148_);
  nand _78371_ (_28355_, _28353_, _07234_);
  and _78372_ (_28356_, _12426_, _06545_);
  nor _78373_ (_28357_, _28356_, _07233_);
  nand _78374_ (_28358_, _28357_, _28355_);
  nand _78375_ (_28359_, _28358_, _12782_);
  and _78376_ (_28360_, _12426_, \oc8051_golden_model_1.PSW [7]);
  nor _78377_ (_28361_, _28183_, \oc8051_golden_model_1.PSW [7]);
  or _78378_ (_28362_, _28361_, _28360_);
  and _78379_ (_28363_, _28362_, _12776_);
  nor _78380_ (_28364_, _28363_, _12780_);
  and _78381_ (_28366_, _28364_, _28359_);
  or _78382_ (_28367_, _28366_, _28147_);
  nand _78383_ (_28368_, _28367_, _11022_);
  nor _78384_ (_28369_, _12426_, _11022_);
  nor _78385_ (_28370_, _28369_, _06366_);
  and _78386_ (_28371_, _28370_, _28368_);
  or _78387_ (_28372_, _28371_, _28146_);
  nand _78388_ (_28373_, _28372_, _09061_);
  and _78389_ (_28374_, _12426_, _06528_);
  nor _78390_ (_28375_, _28374_, _12795_);
  nand _78391_ (_28377_, _28375_, _28373_);
  nand _78392_ (_28378_, _28377_, _25056_);
  and _78393_ (_28379_, _12426_, _10558_);
  nor _78394_ (_28380_, _28183_, _10558_);
  or _78395_ (_28381_, _28380_, _28379_);
  and _78396_ (_28382_, _28381_, _12800_);
  nor _78397_ (_28383_, _28382_, _12804_);
  and _78398_ (_28384_, _28383_, _28378_);
  or _78399_ (_28385_, _28384_, _28144_);
  nand _78400_ (_28386_, _28385_, _12153_);
  nor _78401_ (_28388_, _12426_, _12153_);
  nor _78402_ (_28389_, _28388_, _11125_);
  nand _78403_ (_28390_, _28389_, _28386_);
  and _78404_ (_28391_, _28142_, _11125_);
  nor _78405_ (_28392_, _28391_, _06551_);
  nand _78406_ (_28393_, _28392_, _28390_);
  nor _78407_ (_28394_, _06365_, _07253_);
  not _78408_ (_28395_, _28394_);
  and _78409_ (_28396_, _07357_, _06551_);
  nor _78410_ (_28397_, _28396_, _28395_);
  nand _78411_ (_28399_, _28397_, _28393_);
  nor _78412_ (_28400_, _12216_, _13004_);
  and _78413_ (_28401_, _28162_, _13004_);
  or _78414_ (_28402_, _28401_, _06558_);
  or _78415_ (_28403_, _28402_, _28400_);
  and _78416_ (_28404_, _28403_, _12151_);
  and _78417_ (_28405_, _28404_, _28399_);
  or _78418_ (_28406_, _28405_, _28143_);
  nand _78419_ (_28407_, _28406_, _13012_);
  nor _78420_ (_28408_, _13012_, _12426_);
  nor _78421_ (_28410_, _28408_, _11284_);
  nand _78422_ (_28411_, _28410_, _28407_);
  and _78423_ (_28412_, _28142_, _11284_);
  nor _78424_ (_28413_, _28412_, _06281_);
  nand _78425_ (_28414_, _28413_, _28411_);
  nor _78426_ (_28415_, _06362_, _25646_);
  not _78427_ (_28416_, _28415_);
  and _78428_ (_28417_, _07357_, _06281_);
  nor _78429_ (_28418_, _28417_, _28416_);
  nand _78430_ (_28419_, _28418_, _28414_);
  and _78431_ (_28421_, _12216_, _13004_);
  nor _78432_ (_28422_, _28162_, _13004_);
  or _78433_ (_28423_, _28422_, _28421_);
  and _78434_ (_28424_, _28423_, _06362_);
  nor _78435_ (_28425_, _28424_, _13031_);
  nand _78436_ (_28426_, _28425_, _28419_);
  nor _78437_ (_28427_, _28142_, _13030_);
  nor _78438_ (_28428_, _28427_, _06568_);
  nand _78439_ (_28429_, _28428_, _28426_);
  and _78440_ (_28430_, _12426_, _06568_);
  nor _78441_ (_28432_, _28430_, _13038_);
  nand _78442_ (_28433_, _28432_, _28429_);
  nor _78443_ (_28434_, _28142_, _13037_);
  nor _78444_ (_28435_, _28434_, _06361_);
  and _78445_ (_28436_, _28435_, _28433_);
  or _78446_ (_28437_, _28436_, _28139_);
  nand _78447_ (_28438_, _28437_, _28114_);
  and _78448_ (_28439_, _28423_, _05927_);
  nor _78449_ (_28440_, _28439_, _13053_);
  nand _78450_ (_28441_, _28440_, _28438_);
  nor _78451_ (_28443_, _28142_, _13052_);
  nor _78452_ (_28444_, _28443_, _06278_);
  nand _78453_ (_28445_, _28444_, _28441_);
  and _78454_ (_28446_, _12426_, _06278_);
  nor _78455_ (_28447_, _28446_, _13059_);
  nand _78456_ (_28448_, _28447_, _28445_);
  nor _78457_ (_28449_, _28142_, _12141_);
  nor _78458_ (_28450_, _28449_, _06379_);
  and _78459_ (_28451_, _28450_, _28448_);
  or _78460_ (_28452_, _28451_, _28138_);
  and _78461_ (_28454_, _28452_, _28130_);
  and _78462_ (_28455_, _28142_, _13068_);
  or _78463_ (_28456_, _28455_, _28454_);
  or _78464_ (_28457_, _28456_, _01351_);
  or _78465_ (_28458_, _01347_, \oc8051_golden_model_1.PC [9]);
  and _78466_ (_28459_, _28458_, _42618_);
  and _78467_ (_43255_, _28459_, _28457_);
  nand _78468_ (_28460_, _12203_, _06366_);
  nand _78469_ (_28461_, _12203_, _06375_);
  nand _78470_ (_28462_, _12203_, _06369_);
  nand _78471_ (_28464_, _07412_, _05925_);
  and _78472_ (_28465_, _28140_, \oc8051_golden_model_1.PC [10]);
  nor _78473_ (_28466_, _28140_, \oc8051_golden_model_1.PC [10]);
  nor _78474_ (_28467_, _28466_, _28465_);
  and _78475_ (_28468_, _28467_, _25492_);
  and _78476_ (_28469_, _28467_, _25401_);
  or _78477_ (_28470_, _28467_, _12550_);
  and _78478_ (_28471_, _28467_, _27163_);
  nor _78479_ (_28472_, _12284_, _12281_);
  not _78480_ (_28473_, _28472_);
  and _78481_ (_28475_, _28473_, _12213_);
  nor _78482_ (_28476_, _28473_, _12213_);
  nor _78483_ (_28477_, _28476_, _28475_);
  or _78484_ (_28478_, _28477_, _12536_);
  or _78485_ (_28479_, _12534_, _12202_);
  and _78486_ (_28480_, _28479_, _06341_);
  and _78487_ (_28481_, _28480_, _28478_);
  and _78488_ (_28482_, _12507_, _12421_);
  nor _78489_ (_28483_, _12488_, _12424_);
  nor _78490_ (_28484_, _28483_, _12489_);
  and _78491_ (_28486_, _28484_, _12393_);
  or _78492_ (_28487_, _28486_, _28482_);
  or _78493_ (_28488_, _28487_, _08654_);
  and _78494_ (_28489_, _12421_, _07141_);
  nand _78495_ (_28490_, _07142_, \oc8051_golden_model_1.PC [10]);
  nor _78496_ (_28491_, _28490_, _07486_);
  or _78497_ (_28492_, _28491_, _28489_);
  and _78498_ (_28493_, _28492_, _06782_);
  or _78499_ (_28494_, _28493_, _06758_);
  and _78500_ (_28495_, _28494_, _12512_);
  not _78501_ (_28497_, _12514_);
  and _78502_ (_28498_, _28467_, _28497_);
  or _78503_ (_28499_, _28498_, _12387_);
  or _78504_ (_28500_, _28499_, _28495_);
  and _78505_ (_28501_, _28500_, _27157_);
  and _78506_ (_28502_, _28501_, _28488_);
  or _78507_ (_28503_, _28502_, _28481_);
  and _78508_ (_28504_, _28503_, _12541_);
  or _78509_ (_28505_, _28504_, _28471_);
  and _78510_ (_28506_, _28505_, _06466_);
  and _78511_ (_28508_, _12421_, _06467_);
  nor _78512_ (_28509_, _28508_, _07611_);
  nand _78513_ (_28510_, _28509_, _12550_);
  or _78514_ (_28511_, _28510_, _28506_);
  and _78515_ (_28512_, _28511_, _28470_);
  or _78516_ (_28513_, _28512_, _06464_);
  or _78517_ (_28514_, _12421_, _06465_);
  and _78518_ (_28515_, _28514_, _12560_);
  and _78519_ (_28516_, _28515_, _28513_);
  or _78520_ (_28517_, _28516_, _28469_);
  and _78521_ (_28519_, _28517_, _06269_);
  and _78522_ (_28520_, _12421_, _06268_);
  or _78523_ (_28521_, _28520_, _12563_);
  or _78524_ (_28522_, _28521_, _28519_);
  and _78525_ (_28523_, _28522_, _07303_);
  nand _78526_ (_28524_, _12421_, _06267_);
  nand _78527_ (_28525_, _28524_, _12378_);
  or _78528_ (_28526_, _28525_, _28523_);
  or _78529_ (_28527_, _28477_, _12371_);
  nand _78530_ (_28528_, _12371_, _12203_);
  and _78531_ (_28529_, _28528_, _28527_);
  or _78532_ (_28530_, _28529_, _12378_);
  and _78533_ (_28531_, _28530_, _12177_);
  and _78534_ (_28532_, _28531_, _28526_);
  and _78535_ (_28533_, _28477_, _12335_);
  and _78536_ (_28534_, _12333_, _12202_);
  or _78537_ (_28535_, _28534_, _28533_);
  and _78538_ (_28536_, _28535_, _06347_);
  or _78539_ (_28537_, _28536_, _06480_);
  or _78540_ (_28538_, _28537_, _28532_);
  and _78541_ (_28541_, _12587_, _12202_);
  not _78542_ (_28542_, _12587_);
  and _78543_ (_28543_, _28477_, _28542_);
  or _78544_ (_28544_, _28543_, _06774_);
  or _78545_ (_28545_, _28544_, _28541_);
  and _78546_ (_28546_, _28545_, _12176_);
  and _78547_ (_28547_, _28546_, _28538_);
  or _78548_ (_28548_, _28477_, _12604_);
  nand _78549_ (_28549_, _12604_, _12203_);
  and _78550_ (_28550_, _28549_, _06371_);
  and _78551_ (_28552_, _28550_, _28548_);
  or _78552_ (_28553_, _28552_, _12174_);
  or _78553_ (_28554_, _28553_, _28547_);
  or _78554_ (_28555_, _28467_, _12175_);
  and _78555_ (_28556_, _25322_, _06262_);
  and _78556_ (_28557_, _28556_, _28555_);
  and _78557_ (_28558_, _28557_, _28554_);
  not _78558_ (_28559_, _12421_);
  nor _78559_ (_28560_, _28556_, _28559_);
  nand _78560_ (_28561_, _12630_, _06007_);
  or _78561_ (_28563_, _28561_, _28560_);
  or _78562_ (_28564_, _28563_, _28558_);
  or _78563_ (_28565_, _28467_, _12630_);
  and _78564_ (_28566_, _28565_, _14058_);
  and _78565_ (_28567_, _28566_, _28564_);
  or _78566_ (_28568_, _28567_, _25158_);
  and _78567_ (_28569_, _28568_, _14057_);
  or _78568_ (_28570_, _28559_, _06506_);
  nand _78569_ (_28571_, _28570_, _12639_);
  or _78570_ (_28572_, _28571_, _28569_);
  or _78571_ (_28574_, _28467_, _12639_);
  and _78572_ (_28575_, _28574_, _12643_);
  and _78573_ (_28576_, _28575_, _28572_);
  nor _78574_ (_28577_, _28559_, _12643_);
  or _78575_ (_28578_, _28577_, _10515_);
  or _78576_ (_28579_, _28578_, _28576_);
  or _78577_ (_28580_, _28467_, _05984_);
  and _78578_ (_28581_, _28580_, _06258_);
  and _78579_ (_28582_, _28581_, _28579_);
  nand _78580_ (_28583_, _12421_, _06257_);
  nand _78581_ (_28585_, _28583_, _27951_);
  or _78582_ (_28586_, _28585_, _28582_);
  nand _78583_ (_28587_, _12203_, _06373_);
  and _78584_ (_28588_, _28587_, _07216_);
  and _78585_ (_28589_, _28588_, _28586_);
  nor _78586_ (_28590_, _28559_, _07216_);
  or _78587_ (_28591_, _28590_, _10094_);
  or _78588_ (_28592_, _28591_, _28589_);
  or _78589_ (_28593_, _12202_, _05982_);
  and _78590_ (_28594_, _28593_, _12172_);
  and _78591_ (_28596_, _28594_, _28592_);
  nor _78592_ (_28597_, _28596_, _28468_);
  nor _78593_ (_28598_, _28597_, _06323_);
  nand _78594_ (_28599_, _12421_, _06323_);
  nand _78595_ (_28600_, _28599_, _27971_);
  or _78596_ (_28601_, _28600_, _28598_);
  or _78597_ (_28602_, _28484_, _12679_);
  and _78598_ (_28603_, _28602_, _09030_);
  and _78599_ (_28604_, _28603_, _28601_);
  nor _78600_ (_28605_, _28559_, _09030_);
  or _78601_ (_28607_, _28605_, _06218_);
  or _78602_ (_28608_, _28607_, _28604_);
  and _78603_ (_28609_, _12203_, _06218_);
  nor _78604_ (_28610_, _28609_, _10929_);
  and _78605_ (_28611_, _28610_, _28608_);
  and _78606_ (_28612_, _12421_, _10929_);
  or _78607_ (_28613_, _28612_, _12690_);
  or _78608_ (_28614_, _28613_, _28611_);
  nor _78609_ (_28615_, _12719_, \oc8051_golden_model_1.DPH [2]);
  nor _78610_ (_28616_, _28615_, _12720_);
  or _78611_ (_28618_, _28616_, _12691_);
  and _78612_ (_28619_, _28618_, _06881_);
  and _78613_ (_28620_, _28619_, _28614_);
  and _78614_ (_28621_, _12421_, _06322_);
  or _78615_ (_28622_, _28621_, _28620_);
  and _78616_ (_28623_, _28622_, _28464_);
  or _78617_ (_28624_, _28484_, _11342_);
  or _78618_ (_28625_, _12421_, _12759_);
  and _78619_ (_28626_, _28625_, _12733_);
  and _78620_ (_28627_, _28626_, _28624_);
  or _78621_ (_28629_, _28627_, _12737_);
  or _78622_ (_28630_, _28629_, _28623_);
  or _78623_ (_28631_, _28467_, _12169_);
  and _78624_ (_28632_, _28631_, _12166_);
  and _78625_ (_28633_, _28632_, _28630_);
  nor _78626_ (_28634_, _28559_, _12166_);
  or _78627_ (_28635_, _28634_, _06369_);
  or _78628_ (_28636_, _28635_, _28633_);
  and _78629_ (_28637_, _28636_, _28462_);
  or _78630_ (_28638_, _28637_, _06536_);
  nand _78631_ (_28640_, _28559_, _06536_);
  nor _78632_ (_28641_, _12755_, _12750_);
  and _78633_ (_28642_, _28641_, _28640_);
  and _78634_ (_28643_, _28642_, _28638_);
  or _78635_ (_28644_, _28484_, _12759_);
  or _78636_ (_28645_, _12421_, _11342_);
  and _78637_ (_28646_, _28645_, _12755_);
  and _78638_ (_28647_, _28646_, _28644_);
  or _78639_ (_28648_, _28647_, _10980_);
  or _78640_ (_28649_, _28648_, _28643_);
  or _78641_ (_28651_, _28467_, _10979_);
  and _78642_ (_28652_, _28651_, _12164_);
  and _78643_ (_28653_, _28652_, _28649_);
  nor _78644_ (_28654_, _12164_, _28559_);
  or _78645_ (_28655_, _28654_, _06375_);
  or _78646_ (_28656_, _28655_, _28653_);
  and _78647_ (_28657_, _28656_, _28461_);
  or _78648_ (_28658_, _28657_, _06545_);
  nand _78649_ (_28659_, _28559_, _06545_);
  and _78650_ (_28660_, _28659_, _28029_);
  and _78651_ (_28662_, _28660_, _28658_);
  or _78652_ (_28663_, _28484_, \oc8051_golden_model_1.PSW [7]);
  or _78653_ (_28664_, _12421_, _10558_);
  and _78654_ (_28665_, _28664_, _12776_);
  and _78655_ (_28666_, _28665_, _28663_);
  or _78656_ (_28667_, _28666_, _12780_);
  or _78657_ (_28668_, _28667_, _28662_);
  or _78658_ (_28669_, _28467_, _12162_);
  and _78659_ (_28670_, _28669_, _11022_);
  and _78660_ (_28671_, _28670_, _28668_);
  nor _78661_ (_28673_, _28559_, _11022_);
  or _78662_ (_28674_, _28673_, _06366_);
  or _78663_ (_28675_, _28674_, _28671_);
  and _78664_ (_28676_, _28675_, _28460_);
  or _78665_ (_28677_, _28676_, _06528_);
  nand _78666_ (_28678_, _28559_, _06528_);
  and _78667_ (_28679_, _28678_, _28051_);
  and _78668_ (_28680_, _28679_, _28677_);
  or _78669_ (_28681_, _28484_, _10558_);
  or _78670_ (_28682_, _12421_, \oc8051_golden_model_1.PSW [7]);
  and _78671_ (_28684_, _28682_, _12800_);
  and _78672_ (_28685_, _28684_, _28681_);
  or _78673_ (_28686_, _28685_, _12804_);
  or _78674_ (_28687_, _28686_, _28680_);
  or _78675_ (_28688_, _28467_, _12154_);
  and _78676_ (_28689_, _28688_, _12153_);
  and _78677_ (_28690_, _28689_, _28687_);
  nor _78678_ (_28691_, _28559_, _12153_);
  or _78679_ (_28692_, _28691_, _11125_);
  or _78680_ (_28693_, _28692_, _28690_);
  or _78681_ (_28695_, _28467_, _11126_);
  and _78682_ (_28696_, _28695_, _28693_);
  or _78683_ (_28697_, _28696_, _06551_);
  nand _78684_ (_28698_, _07776_, _06551_);
  and _78685_ (_28699_, _28698_, _28394_);
  and _78686_ (_28700_, _28699_, _28697_);
  not _78687_ (_28701_, _13004_);
  or _78688_ (_28702_, _28477_, _28701_);
  or _78689_ (_28703_, _12202_, _13004_);
  and _78690_ (_28704_, _28703_, _06365_);
  and _78691_ (_28706_, _28704_, _28702_);
  or _78692_ (_28707_, _28706_, _25625_);
  or _78693_ (_28708_, _28707_, _28700_);
  or _78694_ (_28709_, _28467_, _12151_);
  and _78695_ (_28710_, _28709_, _13012_);
  and _78696_ (_28711_, _28710_, _28708_);
  nor _78697_ (_28712_, _13012_, _28559_);
  or _78698_ (_28713_, _28712_, _11284_);
  or _78699_ (_28714_, _28713_, _28711_);
  or _78700_ (_28715_, _28467_, _11285_);
  and _78701_ (_28717_, _28715_, _28714_);
  or _78702_ (_28718_, _28717_, _06281_);
  nand _78703_ (_28719_, _07776_, _06281_);
  and _78704_ (_28720_, _28719_, _28415_);
  and _78705_ (_28721_, _28720_, _28718_);
  or _78706_ (_28722_, _28477_, _13004_);
  nand _78707_ (_28723_, _12203_, _13004_);
  and _78708_ (_28724_, _28723_, _28722_);
  and _78709_ (_28725_, _28724_, _06362_);
  or _78710_ (_28726_, _28725_, _13031_);
  or _78711_ (_28728_, _28726_, _28721_);
  or _78712_ (_28729_, _28467_, _13030_);
  and _78713_ (_28730_, _28729_, _28728_);
  or _78714_ (_28731_, _28730_, _06568_);
  nand _78715_ (_28732_, _28559_, _06568_);
  and _78716_ (_28733_, _28732_, _13037_);
  and _78717_ (_28734_, _28733_, _28731_);
  and _78718_ (_28735_, _28467_, _13038_);
  or _78719_ (_28736_, _28735_, _06361_);
  or _78720_ (_28737_, _28736_, _28734_);
  nand _78721_ (_28739_, _06656_, _06361_);
  and _78722_ (_28740_, _28739_, _28114_);
  and _78723_ (_28741_, _28740_, _28737_);
  and _78724_ (_28742_, _28724_, _05927_);
  or _78725_ (_28743_, _28742_, _13053_);
  or _78726_ (_28744_, _28743_, _28741_);
  or _78727_ (_28745_, _28467_, _13052_);
  and _78728_ (_28746_, _28745_, _28744_);
  or _78729_ (_28747_, _28746_, _06278_);
  nand _78730_ (_28748_, _28559_, _06278_);
  and _78731_ (_28750_, _28748_, _12141_);
  and _78732_ (_28751_, _28750_, _28747_);
  and _78733_ (_28752_, _28467_, _13059_);
  or _78734_ (_28753_, _28752_, _06379_);
  or _78735_ (_28754_, _28753_, _28751_);
  nand _78736_ (_28755_, _06656_, _06379_);
  and _78737_ (_28756_, _28755_, _28130_);
  and _78738_ (_28757_, _28756_, _28754_);
  and _78739_ (_28758_, _28467_, _13068_);
  or _78740_ (_28759_, _28758_, _28757_);
  or _78741_ (_28761_, _28759_, _01351_);
  or _78742_ (_28762_, _01347_, \oc8051_golden_model_1.PC [10]);
  and _78743_ (_28763_, _28762_, _42618_);
  and _78744_ (_43256_, _28763_, _28761_);
  and _78745_ (_28764_, _28465_, \oc8051_golden_model_1.PC [11]);
  nor _78746_ (_28765_, _28465_, \oc8051_golden_model_1.PC [11]);
  nor _78747_ (_28766_, _28765_, _28764_);
  or _78748_ (_28767_, _28766_, _12151_);
  or _78749_ (_28768_, _28766_, _12162_);
  or _78750_ (_28769_, _28766_, _10979_);
  or _78751_ (_28771_, _28766_, _12169_);
  or _78752_ (_28772_, _12417_, _09030_);
  nor _78753_ (_28773_, _12208_, _05982_);
  and _78754_ (_28774_, _12333_, _12207_);
  nor _78755_ (_28775_, _28475_, _12204_);
  and _78756_ (_28776_, _28775_, _12211_);
  nor _78757_ (_28777_, _28775_, _12211_);
  or _78758_ (_28778_, _28777_, _28776_);
  and _78759_ (_28779_, _28778_, _12335_);
  or _78760_ (_28780_, _28779_, _12177_);
  or _78761_ (_28782_, _28780_, _28774_);
  nand _78762_ (_28783_, _12371_, _12208_);
  or _78763_ (_28784_, _28778_, _12371_);
  and _78764_ (_28785_, _28784_, _12379_);
  and _78765_ (_28786_, _28785_, _28783_);
  and _78766_ (_28787_, _12417_, _06464_);
  or _78767_ (_28788_, _12545_, _12417_);
  or _78768_ (_28789_, _12534_, _12207_);
  or _78769_ (_28790_, _28778_, _12536_);
  and _78770_ (_28791_, _28790_, _06341_);
  and _78771_ (_28793_, _28791_, _28789_);
  or _78772_ (_28794_, _12418_, _12419_);
  nand _78773_ (_28795_, _28794_, _12490_);
  or _78774_ (_28796_, _28794_, _12490_);
  and _78775_ (_28797_, _28796_, _28795_);
  and _78776_ (_28798_, _28797_, _25366_);
  or _78777_ (_28799_, _28798_, _08654_);
  and _78778_ (_28800_, _12507_, _12417_);
  or _78779_ (_28801_, _28800_, _28799_);
  or _78780_ (_28802_, _12517_, _12417_);
  nor _78781_ (_28804_, _06781_, _07141_);
  nor _78782_ (_28805_, _06758_, \oc8051_golden_model_1.PC [11]);
  nand _78783_ (_28806_, _28805_, _28804_);
  or _78784_ (_28807_, _28806_, _07486_);
  nand _78785_ (_28808_, _28807_, _28802_);
  nand _78786_ (_28809_, _28808_, _12512_);
  or _78787_ (_28810_, _28766_, _12514_);
  and _78788_ (_28811_, _28810_, _28809_);
  or _78789_ (_28812_, _28811_, _12387_);
  and _78790_ (_28813_, _28812_, _27157_);
  and _78791_ (_28815_, _28813_, _28801_);
  or _78792_ (_28816_, _28815_, _28793_);
  and _78793_ (_28817_, _28816_, _12541_);
  and _78794_ (_28818_, _28766_, _27163_);
  or _78795_ (_28819_, _28818_, _12546_);
  or _78796_ (_28820_, _28819_, _28817_);
  and _78797_ (_28821_, _28820_, _28788_);
  or _78798_ (_28822_, _28821_, _12551_);
  or _78799_ (_28823_, _28766_, _12550_);
  and _78800_ (_28824_, _28823_, _06465_);
  and _78801_ (_28826_, _28824_, _28822_);
  or _78802_ (_28827_, _28826_, _28787_);
  and _78803_ (_28828_, _28827_, _12560_);
  and _78804_ (_28829_, _28766_, _25401_);
  or _78805_ (_28830_, _28829_, _12566_);
  or _78806_ (_28831_, _28830_, _28828_);
  or _78807_ (_28832_, _12565_, _12417_);
  and _78808_ (_28833_, _28832_, _12378_);
  and _78809_ (_28834_, _28833_, _28831_);
  or _78810_ (_28835_, _28834_, _28786_);
  or _78811_ (_28837_, _28835_, _06347_);
  and _78812_ (_28838_, _28837_, _06774_);
  and _78813_ (_28839_, _28838_, _28782_);
  and _78814_ (_28840_, _28778_, _28542_);
  and _78815_ (_28841_, _12587_, _12207_);
  or _78816_ (_28842_, _28841_, _28840_);
  and _78817_ (_28843_, _28842_, _06480_);
  or _78818_ (_28844_, _28843_, _28839_);
  and _78819_ (_28845_, _28844_, _12176_);
  or _78820_ (_28846_, _28778_, _12604_);
  nand _78821_ (_28848_, _12604_, _12208_);
  and _78822_ (_28849_, _28848_, _06371_);
  and _78823_ (_28850_, _28849_, _28846_);
  or _78824_ (_28851_, _28850_, _28845_);
  and _78825_ (_28852_, _28851_, _12175_);
  nand _78826_ (_28853_, _28766_, _12174_);
  nand _78827_ (_28854_, _28853_, _12623_);
  or _78828_ (_28855_, _28854_, _28852_);
  or _78829_ (_28856_, _12623_, _12417_);
  and _78830_ (_28857_, _28856_, _12630_);
  and _78831_ (_28859_, _28857_, _28855_);
  and _78832_ (_28860_, _28766_, _12631_);
  or _78833_ (_28861_, _28860_, _12636_);
  or _78834_ (_28862_, _28861_, _28859_);
  or _78835_ (_28863_, _12635_, _12417_);
  and _78836_ (_28864_, _28863_, _12639_);
  and _78837_ (_28865_, _28864_, _28862_);
  and _78838_ (_28866_, _28766_, _26197_);
  or _78839_ (_28867_, _28866_, _12644_);
  or _78840_ (_28868_, _28867_, _28865_);
  or _78841_ (_28870_, _12417_, _12643_);
  and _78842_ (_28871_, _28870_, _05984_);
  and _78843_ (_28872_, _28871_, _28868_);
  nand _78844_ (_28873_, _28766_, _10515_);
  nand _78845_ (_28874_, _28873_, _12652_);
  or _78846_ (_28875_, _28874_, _28872_);
  or _78847_ (_28876_, _12652_, _12417_);
  and _78848_ (_28877_, _28876_, _06374_);
  and _78849_ (_28878_, _28877_, _28875_);
  nand _78850_ (_28879_, _12207_, _06373_);
  nand _78851_ (_28881_, _28879_, _07216_);
  or _78852_ (_28882_, _28881_, _28878_);
  or _78853_ (_28883_, _12417_, _07216_);
  and _78854_ (_28884_, _28883_, _05982_);
  and _78855_ (_28885_, _28884_, _28882_);
  or _78856_ (_28886_, _28885_, _28773_);
  and _78857_ (_28887_, _28886_, _12172_);
  and _78858_ (_28888_, _28766_, _25492_);
  or _78859_ (_28889_, _28888_, _12670_);
  or _78860_ (_28890_, _28889_, _28887_);
  or _78861_ (_28892_, _12669_, _12417_);
  and _78862_ (_28893_, _28892_, _12679_);
  and _78863_ (_28894_, _28893_, _28890_);
  and _78864_ (_28895_, _28797_, _12674_);
  or _78865_ (_28896_, _28895_, _09031_);
  or _78866_ (_28897_, _28896_, _28894_);
  and _78867_ (_28898_, _28897_, _28772_);
  or _78868_ (_28899_, _28898_, _06218_);
  and _78869_ (_28900_, _12208_, _06218_);
  nor _78870_ (_28901_, _28900_, _10929_);
  and _78871_ (_28902_, _28901_, _28899_);
  and _78872_ (_28903_, _12417_, _10929_);
  or _78873_ (_28904_, _28903_, _28902_);
  and _78874_ (_28905_, _28904_, _12691_);
  or _78875_ (_28906_, _12720_, \oc8051_golden_model_1.DPH [3]);
  nor _78876_ (_28907_, _12721_, _12691_);
  and _78877_ (_28908_, _28907_, _28906_);
  or _78878_ (_28909_, _28908_, _12730_);
  or _78879_ (_28910_, _28909_, _28905_);
  or _78880_ (_28911_, _12729_, _12417_);
  and _78881_ (_28914_, _28911_, _25064_);
  and _78882_ (_28915_, _28914_, _28910_);
  or _78883_ (_28916_, _28797_, _11342_);
  or _78884_ (_28917_, _12417_, _12759_);
  and _78885_ (_28918_, _28917_, _12733_);
  and _78886_ (_28919_, _28918_, _28916_);
  or _78887_ (_28920_, _28919_, _12737_);
  or _78888_ (_28921_, _28920_, _28915_);
  and _78889_ (_28922_, _28921_, _28771_);
  or _78890_ (_28923_, _28922_, _26610_);
  or _78891_ (_28925_, _12417_, _12166_);
  and _78892_ (_28926_, _28925_, _07237_);
  and _78893_ (_28927_, _28926_, _28923_);
  nand _78894_ (_28928_, _12207_, _06369_);
  nand _78895_ (_28929_, _28928_, _12751_);
  or _78896_ (_28930_, _28929_, _28927_);
  or _78897_ (_28931_, _12751_, _12417_);
  and _78898_ (_28932_, _28931_, _25061_);
  and _78899_ (_28933_, _28932_, _28930_);
  or _78900_ (_28934_, _28797_, _12759_);
  or _78901_ (_28936_, _12417_, _11342_);
  and _78902_ (_28937_, _28936_, _12755_);
  and _78903_ (_28938_, _28937_, _28934_);
  or _78904_ (_28939_, _28938_, _10980_);
  or _78905_ (_28940_, _28939_, _28933_);
  and _78906_ (_28941_, _28940_, _28769_);
  or _78907_ (_28942_, _28941_, _26630_);
  or _78908_ (_28943_, _12164_, _12417_);
  and _78909_ (_28944_, _28943_, _07242_);
  and _78910_ (_28945_, _28944_, _28942_);
  nand _78911_ (_28947_, _12207_, _06375_);
  nand _78912_ (_28948_, _28947_, _12772_);
  or _78913_ (_28949_, _28948_, _28945_);
  or _78914_ (_28950_, _12772_, _12417_);
  and _78915_ (_28951_, _28950_, _12782_);
  and _78916_ (_28952_, _28951_, _28949_);
  or _78917_ (_28953_, _28797_, \oc8051_golden_model_1.PSW [7]);
  or _78918_ (_28954_, _12417_, _10558_);
  and _78919_ (_28955_, _28954_, _12776_);
  and _78920_ (_28956_, _28955_, _28953_);
  or _78921_ (_28958_, _28956_, _12780_);
  or _78922_ (_28959_, _28958_, _28952_);
  and _78923_ (_28960_, _28959_, _28768_);
  or _78924_ (_28961_, _28960_, _11023_);
  or _78925_ (_28962_, _12417_, _11022_);
  and _78926_ (_28963_, _28962_, _09056_);
  and _78927_ (_28964_, _28963_, _28961_);
  nand _78928_ (_28965_, _12207_, _06366_);
  nand _78929_ (_28966_, _28965_, _12796_);
  or _78930_ (_28967_, _28966_, _28964_);
  or _78931_ (_28969_, _12796_, _12417_);
  and _78932_ (_28970_, _28969_, _25056_);
  and _78933_ (_28971_, _28970_, _28967_);
  or _78934_ (_28972_, _28797_, _10558_);
  or _78935_ (_28973_, _12417_, \oc8051_golden_model_1.PSW [7]);
  and _78936_ (_28974_, _28973_, _12800_);
  and _78937_ (_28975_, _28974_, _28972_);
  or _78938_ (_28976_, _28975_, _28971_);
  and _78939_ (_28977_, _28976_, _12154_);
  and _78940_ (_28978_, _28766_, _12804_);
  or _78941_ (_28980_, _28978_, _14297_);
  or _78942_ (_28981_, _28980_, _28977_);
  or _78943_ (_28982_, _12417_, _12153_);
  and _78944_ (_28983_, _28982_, _11126_);
  and _78945_ (_28984_, _28983_, _28981_);
  and _78946_ (_28985_, _28766_, _11125_);
  or _78947_ (_28986_, _28985_, _06551_);
  or _78948_ (_28987_, _28986_, _28984_);
  nand _78949_ (_28988_, _07594_, _06551_);
  and _78950_ (_28989_, _28988_, _28987_);
  or _78951_ (_28991_, _28989_, _07253_);
  nor _78952_ (_28992_, _12417_, _05959_);
  nor _78953_ (_28993_, _28992_, _06365_);
  and _78954_ (_28994_, _28993_, _28991_);
  or _78955_ (_28995_, _28778_, _28701_);
  or _78956_ (_28996_, _12207_, _13004_);
  and _78957_ (_28997_, _28996_, _06365_);
  and _78958_ (_28998_, _28997_, _28995_);
  or _78959_ (_28999_, _28998_, _25625_);
  or _78960_ (_29000_, _28999_, _28994_);
  and _78961_ (_29002_, _29000_, _28767_);
  or _78962_ (_29003_, _29002_, _19056_);
  or _78963_ (_29004_, _13012_, _12417_);
  and _78964_ (_29005_, _29004_, _11285_);
  and _78965_ (_29006_, _29005_, _29003_);
  and _78966_ (_29007_, _28766_, _11284_);
  or _78967_ (_29008_, _29007_, _06281_);
  or _78968_ (_29009_, _29008_, _29006_);
  nand _78969_ (_29010_, _07594_, _06281_);
  and _78970_ (_29011_, _29010_, _29009_);
  or _78971_ (_29013_, _29011_, _25646_);
  nor _78972_ (_29014_, _12417_, _05964_);
  nor _78973_ (_29015_, _29014_, _06362_);
  and _78974_ (_29016_, _29015_, _29013_);
  or _78975_ (_29017_, _28778_, _13004_);
  nand _78976_ (_29018_, _12208_, _13004_);
  and _78977_ (_29019_, _29018_, _29017_);
  and _78978_ (_29020_, _29019_, _06362_);
  or _78979_ (_29021_, _29020_, _13031_);
  or _78980_ (_29022_, _29021_, _29016_);
  or _78981_ (_29024_, _28766_, _13030_);
  and _78982_ (_29025_, _29024_, _06926_);
  and _78983_ (_29026_, _29025_, _29022_);
  nand _78984_ (_29027_, _12417_, _06568_);
  nand _78985_ (_29028_, _29027_, _13037_);
  or _78986_ (_29029_, _29028_, _29026_);
  or _78987_ (_29030_, _28766_, _13037_);
  and _78988_ (_29031_, _29030_, _14508_);
  and _78989_ (_29032_, _29031_, _29029_);
  nor _78990_ (_29033_, _14508_, _06213_);
  or _78991_ (_29035_, _29033_, _05940_);
  or _78992_ (_29036_, _29035_, _29032_);
  or _78993_ (_29037_, _12417_, _14710_);
  and _78994_ (_29038_, _29037_, _05928_);
  and _78995_ (_29039_, _29038_, _29036_);
  and _78996_ (_29040_, _29019_, _05927_);
  or _78997_ (_29041_, _29040_, _13053_);
  or _78998_ (_29042_, _29041_, _29039_);
  or _78999_ (_29043_, _28766_, _13052_);
  and _79000_ (_29044_, _29043_, _06279_);
  and _79001_ (_29046_, _29044_, _29042_);
  nand _79002_ (_29047_, _12417_, _06278_);
  nand _79003_ (_29048_, _29047_, _12141_);
  or _79004_ (_29049_, _29048_, _29046_);
  or _79005_ (_29050_, _28766_, _12141_);
  and _79006_ (_29051_, _29050_, _12140_);
  and _79007_ (_29052_, _29051_, _29049_);
  nor _79008_ (_29053_, _12140_, _06213_);
  or _79009_ (_29054_, _29053_, _05939_);
  or _79010_ (_29055_, _29054_, _29052_);
  not _79011_ (_29057_, _13068_);
  not _79012_ (_29058_, _05939_);
  or _79013_ (_29059_, _12417_, _29058_);
  and _79014_ (_29060_, _29059_, _29057_);
  and _79015_ (_29061_, _29060_, _29055_);
  and _79016_ (_29062_, _28766_, _13068_);
  or _79017_ (_29063_, _29062_, _29061_);
  or _79018_ (_29064_, _29063_, _01351_);
  or _79019_ (_29065_, _01347_, \oc8051_golden_model_1.PC [11]);
  and _79020_ (_29066_, _29065_, _42618_);
  and _79021_ (_43257_, _29066_, _29064_);
  and _79022_ (_29068_, _06968_, _06379_);
  or _79023_ (_29069_, _29068_, _05939_);
  and _79024_ (_29070_, _28764_, \oc8051_golden_model_1.PC [12]);
  nor _79025_ (_29071_, _28764_, \oc8051_golden_model_1.PC [12]);
  nor _79026_ (_29072_, _29071_, _29070_);
  not _79027_ (_29073_, _29072_);
  and _79028_ (_29074_, _29073_, _11284_);
  not _79029_ (_29075_, _12414_);
  nor _79030_ (_29076_, _12796_, _29075_);
  nor _79031_ (_29078_, _12772_, _29075_);
  nor _79032_ (_29079_, _12751_, _29075_);
  and _79033_ (_29080_, _12291_, _12288_);
  nor _79034_ (_29081_, _29080_, _12292_);
  or _79035_ (_29082_, _29081_, _12333_);
  or _79036_ (_29083_, _12335_, _12198_);
  and _79037_ (_29084_, _29083_, _06347_);
  nand _79038_ (_29085_, _29084_, _29082_);
  nand _79039_ (_29086_, _12371_, _12198_);
  not _79040_ (_29087_, _29081_);
  or _79041_ (_29089_, _29087_, _12371_);
  and _79042_ (_29090_, _29089_, _12379_);
  and _79043_ (_29091_, _29090_, _29086_);
  or _79044_ (_29092_, _29087_, _12536_);
  or _79045_ (_29093_, _12534_, _12199_);
  nand _79046_ (_29094_, _29093_, _29092_);
  nand _79047_ (_29095_, _29094_, _06341_);
  and _79048_ (_29096_, _12507_, _12414_);
  nor _79049_ (_29097_, _12494_, _12492_);
  nor _79050_ (_29098_, _29097_, _12495_);
  and _79051_ (_29100_, _29098_, _12393_);
  nor _79052_ (_29101_, _29100_, _29096_);
  nand _79053_ (_29102_, _29101_, _12387_);
  nor _79054_ (_29103_, _29073_, _12514_);
  not _79055_ (_29104_, _29103_);
  nor _79056_ (_29105_, _12517_, _29075_);
  and _79057_ (_29106_, _28804_, _07504_);
  and _79058_ (_29107_, _07487_, \oc8051_golden_model_1.PC [12]);
  and _79059_ (_29108_, _29107_, _29106_);
  nor _79060_ (_29109_, _29108_, _29105_);
  nor _79061_ (_29111_, _29109_, _12516_);
  nor _79062_ (_29112_, _29111_, _12387_);
  and _79063_ (_29113_, _29112_, _29104_);
  not _79064_ (_29114_, _29113_);
  and _79065_ (_29115_, _29114_, _27157_);
  nand _79066_ (_29116_, _29115_, _29102_);
  nand _79067_ (_29117_, _29116_, _29095_);
  and _79068_ (_29118_, _29117_, _12541_);
  and _79069_ (_29119_, _29072_, _27163_);
  or _79070_ (_29120_, _29119_, _12546_);
  or _79071_ (_29122_, _29120_, _29118_);
  nor _79072_ (_29123_, _12545_, _12414_);
  nor _79073_ (_29124_, _29123_, _12551_);
  and _79074_ (_29125_, _29124_, _29122_);
  nor _79075_ (_29126_, _29073_, _12550_);
  or _79076_ (_29127_, _29126_, _06464_);
  nor _79077_ (_29128_, _29127_, _29125_);
  and _79078_ (_29129_, _29075_, _06464_);
  or _79079_ (_29130_, _29129_, _29128_);
  nand _79080_ (_29131_, _29130_, _12560_);
  nor _79081_ (_29133_, _29072_, _12560_);
  nor _79082_ (_29134_, _29133_, _12566_);
  and _79083_ (_29135_, _29134_, _29131_);
  nor _79084_ (_29136_, _12565_, _29075_);
  or _79085_ (_29137_, _29136_, _12379_);
  nor _79086_ (_29138_, _29137_, _29135_);
  or _79087_ (_29139_, _29138_, _06347_);
  or _79088_ (_29140_, _29139_, _29091_);
  and _79089_ (_29141_, _29140_, _29085_);
  nand _79090_ (_29142_, _29141_, _06774_);
  nor _79091_ (_29144_, _29087_, _12587_);
  and _79092_ (_29145_, _12587_, _12198_);
  or _79093_ (_29146_, _29145_, _29144_);
  nor _79094_ (_29147_, _29146_, _06774_);
  nor _79095_ (_29148_, _29147_, _06371_);
  nand _79096_ (_29149_, _29148_, _29142_);
  and _79097_ (_29150_, _12604_, _12198_);
  and _79098_ (_29151_, _29081_, _26518_);
  or _79099_ (_29152_, _29151_, _29150_);
  and _79100_ (_29153_, _29152_, _06371_);
  nor _79101_ (_29155_, _29153_, _12174_);
  and _79102_ (_29156_, _29155_, _29149_);
  and _79103_ (_29157_, _29073_, _12174_);
  or _79104_ (_29158_, _29157_, _29156_);
  and _79105_ (_29159_, _29158_, _12623_);
  nor _79106_ (_29160_, _12623_, _12414_);
  or _79107_ (_29161_, _29160_, _29159_);
  nand _79108_ (_29162_, _29161_, _12630_);
  nor _79109_ (_29163_, _29072_, _12630_);
  nor _79110_ (_29164_, _29163_, _12636_);
  nand _79111_ (_29166_, _29164_, _29162_);
  nor _79112_ (_29167_, _12635_, _29075_);
  nor _79113_ (_29168_, _29167_, _26197_);
  nand _79114_ (_29169_, _29168_, _29166_);
  nor _79115_ (_29170_, _29072_, _12639_);
  nor _79116_ (_29171_, _29170_, _12644_);
  nand _79117_ (_29172_, _29171_, _29169_);
  nor _79118_ (_29173_, _29075_, _12643_);
  nor _79119_ (_29174_, _29173_, _10515_);
  nand _79120_ (_29175_, _29174_, _29172_);
  nor _79121_ (_29177_, _29072_, _05984_);
  nor _79122_ (_29178_, _29177_, _12653_);
  nand _79123_ (_29179_, _29178_, _29175_);
  nor _79124_ (_29180_, _12652_, _29075_);
  nor _79125_ (_29181_, _29180_, _06373_);
  nand _79126_ (_29182_, _29181_, _29179_);
  and _79127_ (_29183_, _12199_, _06373_);
  nor _79128_ (_29184_, _29183_, _12659_);
  nand _79129_ (_29185_, _29184_, _29182_);
  nor _79130_ (_29186_, _29075_, _07216_);
  nor _79131_ (_29188_, _29186_, _10094_);
  nand _79132_ (_29189_, _29188_, _29185_);
  nor _79133_ (_29190_, _12198_, _05982_);
  nor _79134_ (_29191_, _29190_, _25492_);
  nand _79135_ (_29192_, _29191_, _29189_);
  nor _79136_ (_29193_, _29073_, _12172_);
  nor _79137_ (_29194_, _29193_, _12670_);
  nand _79138_ (_29195_, _29194_, _29192_);
  nor _79139_ (_29196_, _12669_, _12414_);
  nor _79140_ (_29197_, _29196_, _12674_);
  and _79141_ (_29199_, _29197_, _29195_);
  and _79142_ (_29200_, _29098_, _12674_);
  nor _79143_ (_29201_, _29200_, _29199_);
  or _79144_ (_29202_, _29201_, _09031_);
  or _79145_ (_29203_, _29075_, _09030_);
  and _79146_ (_29204_, _29203_, _06219_);
  nand _79147_ (_29205_, _29204_, _29202_);
  and _79148_ (_29206_, _12199_, _06218_);
  nor _79149_ (_29207_, _29206_, _10929_);
  nand _79150_ (_29208_, _29207_, _29205_);
  and _79151_ (_29210_, _12414_, _10929_);
  nor _79152_ (_29211_, _29210_, _12690_);
  and _79153_ (_29212_, _29211_, _29208_);
  nor _79154_ (_29213_, _12721_, \oc8051_golden_model_1.DPH [4]);
  nor _79155_ (_29214_, _29213_, _12722_);
  nor _79156_ (_29215_, _29214_, _12691_);
  or _79157_ (_29216_, _29215_, _29212_);
  nand _79158_ (_29217_, _29216_, _12729_);
  nor _79159_ (_29218_, _12729_, _12414_);
  nor _79160_ (_29219_, _29218_, _12733_);
  nand _79161_ (_29221_, _29219_, _29217_);
  nor _79162_ (_29222_, _29098_, _11342_);
  nor _79163_ (_29223_, _12414_, _12759_);
  nor _79164_ (_29224_, _29223_, _25064_);
  not _79165_ (_29225_, _29224_);
  nor _79166_ (_29226_, _29225_, _29222_);
  nor _79167_ (_29227_, _29226_, _12737_);
  nand _79168_ (_29228_, _29227_, _29221_);
  nor _79169_ (_29229_, _29072_, _12169_);
  nor _79170_ (_29230_, _29229_, _26610_);
  nand _79171_ (_29232_, _29230_, _29228_);
  nor _79172_ (_29233_, _29075_, _12166_);
  nor _79173_ (_29234_, _29233_, _06369_);
  nand _79174_ (_29235_, _29234_, _29232_);
  and _79175_ (_29236_, _12199_, _06369_);
  nor _79176_ (_29237_, _29236_, _12752_);
  and _79177_ (_29238_, _29237_, _29235_);
  or _79178_ (_29239_, _29238_, _29079_);
  nand _79179_ (_29240_, _29239_, _25061_);
  and _79180_ (_29241_, _12414_, _12759_);
  and _79181_ (_29243_, _29098_, _11342_);
  or _79182_ (_29244_, _29243_, _29241_);
  and _79183_ (_29245_, _29244_, _12755_);
  nor _79184_ (_29246_, _29245_, _10980_);
  nand _79185_ (_29247_, _29246_, _29240_);
  nor _79186_ (_29248_, _29072_, _10979_);
  nor _79187_ (_29249_, _29248_, _26630_);
  nand _79188_ (_29250_, _29249_, _29247_);
  nor _79189_ (_29251_, _12164_, _29075_);
  nor _79190_ (_29252_, _29251_, _06375_);
  nand _79191_ (_29254_, _29252_, _29250_);
  and _79192_ (_29255_, _12199_, _06375_);
  nor _79193_ (_29256_, _29255_, _12773_);
  and _79194_ (_29257_, _29256_, _29254_);
  or _79195_ (_29258_, _29257_, _29078_);
  nand _79196_ (_29259_, _29258_, _12782_);
  and _79197_ (_29260_, _12414_, \oc8051_golden_model_1.PSW [7]);
  and _79198_ (_29261_, _29098_, _10558_);
  or _79199_ (_29262_, _29261_, _29260_);
  and _79200_ (_29263_, _29262_, _12776_);
  nor _79201_ (_29265_, _29263_, _12780_);
  nand _79202_ (_29266_, _29265_, _29259_);
  nor _79203_ (_29267_, _29072_, _12162_);
  nor _79204_ (_29268_, _29267_, _11023_);
  nand _79205_ (_29269_, _29268_, _29266_);
  nor _79206_ (_29270_, _29075_, _11022_);
  nor _79207_ (_29271_, _29270_, _06366_);
  nand _79208_ (_29272_, _29271_, _29269_);
  and _79209_ (_29273_, _12199_, _06366_);
  nor _79210_ (_29274_, _29273_, _12797_);
  and _79211_ (_29276_, _29274_, _29272_);
  or _79212_ (_29277_, _29276_, _29076_);
  nand _79213_ (_29278_, _29277_, _25056_);
  and _79214_ (_29279_, _12414_, _10558_);
  and _79215_ (_29280_, _29098_, \oc8051_golden_model_1.PSW [7]);
  or _79216_ (_29281_, _29280_, _29279_);
  and _79217_ (_29282_, _29281_, _12800_);
  nor _79218_ (_29283_, _29282_, _12804_);
  nand _79219_ (_29284_, _29283_, _29278_);
  nor _79220_ (_29285_, _29072_, _12154_);
  nor _79221_ (_29287_, _29285_, _14297_);
  nand _79222_ (_29288_, _29287_, _29284_);
  nor _79223_ (_29289_, _29075_, _12153_);
  nor _79224_ (_29290_, _29289_, _11125_);
  nand _79225_ (_29291_, _29290_, _29288_);
  and _79226_ (_29292_, _29073_, _11125_);
  nor _79227_ (_29293_, _29292_, _06551_);
  and _79228_ (_29294_, _29293_, _29291_);
  nor _79229_ (_29295_, _08541_, _06716_);
  or _79230_ (_29296_, _29295_, _07253_);
  or _79231_ (_29298_, _29296_, _29294_);
  nor _79232_ (_29299_, _12414_, _05959_);
  nor _79233_ (_29300_, _29299_, _06365_);
  nand _79234_ (_29301_, _29300_, _29298_);
  and _79235_ (_29302_, _29087_, _13004_);
  nor _79236_ (_29303_, _12198_, _13004_);
  or _79237_ (_29304_, _29303_, _06558_);
  or _79238_ (_29305_, _29304_, _29302_);
  and _79239_ (_29306_, _29305_, _12151_);
  nand _79240_ (_29307_, _29306_, _29301_);
  nor _79241_ (_29309_, _29072_, _12151_);
  nor _79242_ (_29310_, _29309_, _19056_);
  nand _79243_ (_29311_, _29310_, _29307_);
  nor _79244_ (_29312_, _13012_, _29075_);
  nor _79245_ (_29313_, _29312_, _11284_);
  and _79246_ (_29314_, _29313_, _29311_);
  or _79247_ (_29315_, _29314_, _29074_);
  nand _79248_ (_29316_, _29315_, _06282_);
  and _79249_ (_29317_, _08541_, _06281_);
  nor _79250_ (_29318_, _29317_, _25646_);
  and _79251_ (_29320_, _29318_, _29316_);
  nor _79252_ (_29321_, _29075_, _05964_);
  or _79253_ (_29322_, _29321_, _06362_);
  nor _79254_ (_29323_, _29322_, _29320_);
  nor _79255_ (_29324_, _29081_, _13004_);
  and _79256_ (_29325_, _12199_, _13004_);
  nor _79257_ (_29326_, _29325_, _29324_);
  nor _79258_ (_29327_, _29326_, _06921_);
  or _79259_ (_29328_, _29327_, _29323_);
  and _79260_ (_29329_, _29328_, _13030_);
  nor _79261_ (_29331_, _29072_, _13030_);
  or _79262_ (_29332_, _29331_, _29329_);
  nand _79263_ (_29333_, _29332_, _06926_);
  and _79264_ (_29334_, _29075_, _06568_);
  nor _79265_ (_29335_, _29334_, _13038_);
  nand _79266_ (_29336_, _29335_, _29333_);
  nor _79267_ (_29337_, _29073_, _13037_);
  nor _79268_ (_29338_, _29337_, _06361_);
  nand _79269_ (_29339_, _29338_, _29336_);
  and _79270_ (_29340_, _06968_, _06361_);
  nor _79271_ (_29342_, _29340_, _05940_);
  nand _79272_ (_29343_, _29342_, _29339_);
  and _79273_ (_29344_, _12414_, _05940_);
  nor _79274_ (_29345_, _29344_, _05927_);
  nand _79275_ (_29346_, _29345_, _29343_);
  nor _79276_ (_29347_, _29326_, _05928_);
  nor _79277_ (_29348_, _29347_, _13053_);
  nand _79278_ (_29349_, _29348_, _29346_);
  nor _79279_ (_29350_, _29073_, _13052_);
  nor _79280_ (_29351_, _29350_, _06278_);
  nand _79281_ (_29353_, _29351_, _29349_);
  and _79282_ (_29354_, _29075_, _06278_);
  nor _79283_ (_29355_, _29354_, _13059_);
  nand _79284_ (_29356_, _29355_, _29353_);
  nor _79285_ (_29357_, _29073_, _12141_);
  nor _79286_ (_29358_, _29357_, _06379_);
  and _79287_ (_29359_, _29358_, _29356_);
  or _79288_ (_29360_, _29359_, _29069_);
  and _79289_ (_29361_, _12414_, _05939_);
  nor _79290_ (_29362_, _29361_, _13068_);
  and _79291_ (_29364_, _29362_, _29360_);
  and _79292_ (_29365_, _29073_, _13068_);
  nor _79293_ (_29366_, _29365_, _29364_);
  or _79294_ (_29367_, _29366_, _01351_);
  or _79295_ (_29368_, _01347_, \oc8051_golden_model_1.PC [12]);
  and _79296_ (_29369_, _29368_, _42618_);
  and _79297_ (_43258_, _29369_, _29367_);
  and _79298_ (_29370_, _29070_, \oc8051_golden_model_1.PC [13]);
  nor _79299_ (_29371_, _29070_, \oc8051_golden_model_1.PC [13]);
  nor _79300_ (_29372_, _29371_, _29370_);
  or _79301_ (_29374_, _29372_, _12151_);
  or _79302_ (_29375_, _29372_, _12154_);
  or _79303_ (_29376_, _29372_, _12162_);
  or _79304_ (_29377_, _29372_, _10979_);
  or _79305_ (_29378_, _29372_, _12169_);
  or _79306_ (_29379_, _12409_, _09030_);
  nor _79307_ (_29380_, _12194_, _05982_);
  or _79308_ (_29381_, _12196_, _12195_);
  not _79309_ (_29382_, _29381_);
  nor _79310_ (_29383_, _29382_, _12293_);
  and _79311_ (_29385_, _29382_, _12293_);
  or _79312_ (_29386_, _29385_, _29383_);
  or _79313_ (_29387_, _29386_, _12587_);
  nand _79314_ (_29388_, _12587_, _12194_);
  and _79315_ (_29389_, _29388_, _06480_);
  and _79316_ (_29390_, _29389_, _29387_);
  and _79317_ (_29391_, _12333_, _12193_);
  and _79318_ (_29392_, _29386_, _12335_);
  or _79319_ (_29393_, _29392_, _12177_);
  or _79320_ (_29394_, _29393_, _29391_);
  nand _79321_ (_29396_, _12371_, _12194_);
  or _79322_ (_29397_, _29386_, _12371_);
  and _79323_ (_29398_, _29397_, _12379_);
  and _79324_ (_29399_, _29398_, _29396_);
  and _79325_ (_29400_, _12409_, _06464_);
  or _79326_ (_29401_, _12545_, _12409_);
  or _79327_ (_29402_, _29386_, _12536_);
  or _79328_ (_29403_, _12534_, _12193_);
  and _79329_ (_29404_, _29403_, _06341_);
  and _79330_ (_29405_, _29404_, _29402_);
  or _79331_ (_29407_, _12410_, _12411_);
  not _79332_ (_29408_, _29407_);
  nor _79333_ (_29409_, _29408_, _12496_);
  and _79334_ (_29410_, _29408_, _12496_);
  or _79335_ (_29411_, _29410_, _29409_);
  and _79336_ (_29412_, _29411_, _25366_);
  or _79337_ (_29413_, _29412_, _08654_);
  and _79338_ (_29414_, _12507_, _12409_);
  or _79339_ (_29415_, _29414_, _29413_);
  or _79340_ (_29416_, _29372_, _12514_);
  or _79341_ (_29418_, _12517_, _12409_);
  nor _79342_ (_29419_, _07486_, \oc8051_golden_model_1.PC [13]);
  nand _79343_ (_29420_, _29419_, _29106_);
  and _79344_ (_29421_, _29420_, _29418_);
  or _79345_ (_29422_, _29421_, _12516_);
  and _79346_ (_29423_, _29422_, _29416_);
  or _79347_ (_29424_, _29423_, _12387_);
  and _79348_ (_29425_, _29424_, _27157_);
  and _79349_ (_29426_, _29425_, _29415_);
  or _79350_ (_29427_, _29426_, _29405_);
  and _79351_ (_29428_, _29427_, _12541_);
  and _79352_ (_29429_, _29372_, _27163_);
  or _79353_ (_29430_, _29429_, _12546_);
  or _79354_ (_29431_, _29430_, _29428_);
  and _79355_ (_29432_, _29431_, _29401_);
  or _79356_ (_29433_, _29432_, _12551_);
  or _79357_ (_29434_, _29372_, _12550_);
  and _79358_ (_29435_, _29434_, _06465_);
  and _79359_ (_29436_, _29435_, _29433_);
  or _79360_ (_29437_, _29436_, _29400_);
  and _79361_ (_29440_, _29437_, _12560_);
  and _79362_ (_29441_, _29372_, _25401_);
  or _79363_ (_29442_, _29441_, _12566_);
  or _79364_ (_29443_, _29442_, _29440_);
  or _79365_ (_29444_, _12565_, _12409_);
  and _79366_ (_29445_, _29444_, _12378_);
  and _79367_ (_29446_, _29445_, _29443_);
  or _79368_ (_29447_, _29446_, _29399_);
  or _79369_ (_29448_, _29447_, _06347_);
  and _79370_ (_29449_, _29448_, _06774_);
  and _79371_ (_29451_, _29449_, _29394_);
  or _79372_ (_29452_, _29451_, _29390_);
  and _79373_ (_29453_, _29452_, _12176_);
  or _79374_ (_29454_, _29386_, _12604_);
  nand _79375_ (_29455_, _12604_, _12194_);
  and _79376_ (_29456_, _29455_, _06371_);
  and _79377_ (_29457_, _29456_, _29454_);
  or _79378_ (_29458_, _29457_, _29453_);
  and _79379_ (_29459_, _29458_, _12175_);
  nand _79380_ (_29460_, _29372_, _12174_);
  nand _79381_ (_29462_, _29460_, _12623_);
  or _79382_ (_29463_, _29462_, _29459_);
  or _79383_ (_29464_, _12623_, _12409_);
  and _79384_ (_29465_, _29464_, _12630_);
  and _79385_ (_29466_, _29465_, _29463_);
  and _79386_ (_29467_, _29372_, _12631_);
  or _79387_ (_29468_, _29467_, _12636_);
  or _79388_ (_29469_, _29468_, _29466_);
  or _79389_ (_29470_, _12635_, _12409_);
  and _79390_ (_29471_, _29470_, _12639_);
  and _79391_ (_29473_, _29471_, _29469_);
  and _79392_ (_29474_, _29372_, _26197_);
  or _79393_ (_29475_, _29474_, _12644_);
  or _79394_ (_29476_, _29475_, _29473_);
  or _79395_ (_29477_, _12409_, _12643_);
  and _79396_ (_29478_, _29477_, _05984_);
  and _79397_ (_29479_, _29478_, _29476_);
  nand _79398_ (_29480_, _29372_, _10515_);
  nand _79399_ (_29481_, _29480_, _12652_);
  or _79400_ (_29482_, _29481_, _29479_);
  or _79401_ (_29484_, _12652_, _12409_);
  and _79402_ (_29485_, _29484_, _06374_);
  and _79403_ (_29486_, _29485_, _29482_);
  nand _79404_ (_29487_, _12193_, _06373_);
  nand _79405_ (_29488_, _29487_, _07216_);
  or _79406_ (_29489_, _29488_, _29486_);
  or _79407_ (_29490_, _12409_, _07216_);
  and _79408_ (_29491_, _29490_, _05982_);
  and _79409_ (_29492_, _29491_, _29489_);
  or _79410_ (_29493_, _29492_, _29380_);
  and _79411_ (_29495_, _29493_, _12172_);
  and _79412_ (_29496_, _29372_, _25492_);
  or _79413_ (_29497_, _29496_, _12670_);
  or _79414_ (_29498_, _29497_, _29495_);
  or _79415_ (_29499_, _12669_, _12409_);
  and _79416_ (_29500_, _29499_, _12679_);
  and _79417_ (_29501_, _29500_, _29498_);
  and _79418_ (_29502_, _29411_, _12674_);
  or _79419_ (_29503_, _29502_, _09031_);
  or _79420_ (_29504_, _29503_, _29501_);
  and _79421_ (_29506_, _29504_, _29379_);
  or _79422_ (_29507_, _29506_, _06218_);
  and _79423_ (_29508_, _12194_, _06218_);
  nor _79424_ (_29509_, _29508_, _10929_);
  and _79425_ (_29510_, _29509_, _29507_);
  and _79426_ (_29511_, _12409_, _10929_);
  or _79427_ (_29512_, _29511_, _29510_);
  and _79428_ (_29513_, _29512_, _12691_);
  or _79429_ (_29514_, _12722_, \oc8051_golden_model_1.DPH [5]);
  nor _79430_ (_29515_, _12723_, _12691_);
  and _79431_ (_29517_, _29515_, _29514_);
  or _79432_ (_29518_, _29517_, _12730_);
  or _79433_ (_29519_, _29518_, _29513_);
  or _79434_ (_29520_, _12729_, _12409_);
  and _79435_ (_29521_, _29520_, _25064_);
  and _79436_ (_29522_, _29521_, _29519_);
  or _79437_ (_29523_, _29411_, _11342_);
  or _79438_ (_29524_, _12409_, _12759_);
  and _79439_ (_29525_, _29524_, _12733_);
  and _79440_ (_29526_, _29525_, _29523_);
  or _79441_ (_29528_, _29526_, _12737_);
  or _79442_ (_29529_, _29528_, _29522_);
  and _79443_ (_29530_, _29529_, _29378_);
  or _79444_ (_29531_, _29530_, _26610_);
  or _79445_ (_29532_, _12409_, _12166_);
  and _79446_ (_29533_, _29532_, _07237_);
  and _79447_ (_29534_, _29533_, _29531_);
  nand _79448_ (_29535_, _12193_, _06369_);
  nand _79449_ (_29536_, _29535_, _12751_);
  or _79450_ (_29537_, _29536_, _29534_);
  or _79451_ (_29539_, _12751_, _12409_);
  and _79452_ (_29540_, _29539_, _25061_);
  and _79453_ (_29541_, _29540_, _29537_);
  or _79454_ (_29542_, _29411_, _12759_);
  or _79455_ (_29543_, _12409_, _11342_);
  and _79456_ (_29544_, _29543_, _12755_);
  and _79457_ (_29545_, _29544_, _29542_);
  or _79458_ (_29546_, _29545_, _10980_);
  or _79459_ (_29547_, _29546_, _29541_);
  and _79460_ (_29548_, _29547_, _29377_);
  or _79461_ (_29550_, _29548_, _26630_);
  or _79462_ (_29551_, _12164_, _12409_);
  and _79463_ (_29552_, _29551_, _07242_);
  and _79464_ (_29553_, _29552_, _29550_);
  nand _79465_ (_29554_, _12193_, _06375_);
  nand _79466_ (_29555_, _29554_, _12772_);
  or _79467_ (_29556_, _29555_, _29553_);
  or _79468_ (_29557_, _12772_, _12409_);
  and _79469_ (_29558_, _29557_, _12782_);
  and _79470_ (_29559_, _29558_, _29556_);
  or _79471_ (_29561_, _29411_, \oc8051_golden_model_1.PSW [7]);
  or _79472_ (_29562_, _12409_, _10558_);
  and _79473_ (_29563_, _29562_, _12776_);
  and _79474_ (_29564_, _29563_, _29561_);
  or _79475_ (_29565_, _29564_, _12780_);
  or _79476_ (_29566_, _29565_, _29559_);
  and _79477_ (_29567_, _29566_, _29376_);
  or _79478_ (_29568_, _29567_, _11023_);
  or _79479_ (_29569_, _12409_, _11022_);
  and _79480_ (_29570_, _29569_, _09056_);
  and _79481_ (_29572_, _29570_, _29568_);
  nand _79482_ (_29573_, _12193_, _06366_);
  nand _79483_ (_29574_, _29573_, _12796_);
  or _79484_ (_29575_, _29574_, _29572_);
  or _79485_ (_29576_, _12796_, _12409_);
  and _79486_ (_29577_, _29576_, _25056_);
  and _79487_ (_29578_, _29577_, _29575_);
  or _79488_ (_29579_, _29411_, _10558_);
  or _79489_ (_29580_, _12409_, \oc8051_golden_model_1.PSW [7]);
  and _79490_ (_29581_, _29580_, _12800_);
  and _79491_ (_29583_, _29581_, _29579_);
  or _79492_ (_29584_, _29583_, _12804_);
  or _79493_ (_29585_, _29584_, _29578_);
  and _79494_ (_29586_, _29585_, _29375_);
  or _79495_ (_29587_, _29586_, _14297_);
  or _79496_ (_29588_, _12409_, _12153_);
  and _79497_ (_29589_, _29588_, _11126_);
  and _79498_ (_29590_, _29589_, _29587_);
  and _79499_ (_29591_, _29372_, _11125_);
  or _79500_ (_29592_, _29591_, _06551_);
  or _79501_ (_29594_, _29592_, _29590_);
  nand _79502_ (_29595_, _08244_, _06551_);
  and _79503_ (_29596_, _29595_, _29594_);
  or _79504_ (_29597_, _29596_, _07253_);
  nor _79505_ (_29598_, _12409_, _05959_);
  nor _79506_ (_29599_, _29598_, _06365_);
  and _79507_ (_29600_, _29599_, _29597_);
  or _79508_ (_29601_, _29386_, _28701_);
  or _79509_ (_29602_, _12193_, _13004_);
  and _79510_ (_29603_, _29602_, _06365_);
  and _79511_ (_29605_, _29603_, _29601_);
  or _79512_ (_29606_, _29605_, _25625_);
  or _79513_ (_29607_, _29606_, _29600_);
  and _79514_ (_29608_, _29607_, _29374_);
  or _79515_ (_29609_, _29608_, _19056_);
  or _79516_ (_29610_, _13012_, _12409_);
  and _79517_ (_29611_, _29610_, _11285_);
  and _79518_ (_29612_, _29611_, _29609_);
  and _79519_ (_29613_, _29372_, _11284_);
  or _79520_ (_29614_, _29613_, _06281_);
  or _79521_ (_29616_, _29614_, _29612_);
  nand _79522_ (_29617_, _08244_, _06281_);
  and _79523_ (_29618_, _29617_, _29616_);
  or _79524_ (_29619_, _29618_, _25646_);
  nor _79525_ (_29620_, _12409_, _05964_);
  nor _79526_ (_29621_, _29620_, _06362_);
  and _79527_ (_29622_, _29621_, _29619_);
  or _79528_ (_29623_, _29386_, _13004_);
  nand _79529_ (_29624_, _12194_, _13004_);
  and _79530_ (_29625_, _29624_, _29623_);
  and _79531_ (_29627_, _29625_, _06362_);
  or _79532_ (_29628_, _29627_, _13031_);
  or _79533_ (_29629_, _29628_, _29622_);
  or _79534_ (_29630_, _29372_, _13030_);
  and _79535_ (_29631_, _29630_, _06926_);
  and _79536_ (_29632_, _29631_, _29629_);
  nand _79537_ (_29633_, _12409_, _06568_);
  nand _79538_ (_29634_, _29633_, _13037_);
  or _79539_ (_29635_, _29634_, _29632_);
  or _79540_ (_29636_, _29372_, _13037_);
  and _79541_ (_29638_, _29636_, _14508_);
  and _79542_ (_29639_, _29638_, _29635_);
  nor _79543_ (_29640_, _06611_, _14508_);
  or _79544_ (_29641_, _29640_, _05940_);
  or _79545_ (_29642_, _29641_, _29639_);
  or _79546_ (_29643_, _12409_, _14710_);
  and _79547_ (_29644_, _29643_, _05928_);
  and _79548_ (_29645_, _29644_, _29642_);
  and _79549_ (_29646_, _29625_, _05927_);
  or _79550_ (_29647_, _29646_, _13053_);
  or _79551_ (_29649_, _29647_, _29645_);
  or _79552_ (_29650_, _29372_, _13052_);
  and _79553_ (_29651_, _29650_, _06279_);
  and _79554_ (_29652_, _29651_, _29649_);
  nand _79555_ (_29653_, _12409_, _06278_);
  nand _79556_ (_29654_, _29653_, _12141_);
  or _79557_ (_29655_, _29654_, _29652_);
  or _79558_ (_29656_, _29372_, _12141_);
  and _79559_ (_29657_, _29656_, _12140_);
  and _79560_ (_29658_, _29657_, _29655_);
  nor _79561_ (_29660_, _06611_, _12140_);
  or _79562_ (_29661_, _29660_, _05939_);
  or _79563_ (_29662_, _29661_, _29658_);
  or _79564_ (_29663_, _12409_, _29058_);
  and _79565_ (_29664_, _29663_, _29057_);
  and _79566_ (_29665_, _29664_, _29662_);
  and _79567_ (_29666_, _29372_, _13068_);
  or _79568_ (_29667_, _29666_, _29665_);
  or _79569_ (_29668_, _29667_, _01351_);
  or _79570_ (_29669_, _01347_, \oc8051_golden_model_1.PC [13]);
  and _79571_ (_29671_, _29669_, _42618_);
  and _79572_ (_43260_, _29671_, _29668_);
  and _79573_ (_29672_, _29370_, \oc8051_golden_model_1.PC [14]);
  nor _79574_ (_29673_, _29370_, \oc8051_golden_model_1.PC [14]);
  nor _79575_ (_29674_, _29673_, _29672_);
  nor _79576_ (_29675_, _29674_, _11285_);
  not _79577_ (_29676_, _12403_);
  nor _79578_ (_29677_, _12796_, _29676_);
  nor _79579_ (_29678_, _12772_, _29676_);
  nor _79580_ (_29679_, _12751_, _29676_);
  nor _79581_ (_29681_, _12729_, _29676_);
  and _79582_ (_29682_, _12295_, _12191_);
  nor _79583_ (_29683_, _29682_, _12296_);
  not _79584_ (_29684_, _29683_);
  nand _79585_ (_29685_, _29684_, _12335_);
  or _79586_ (_29686_, _12335_, _12186_);
  and _79587_ (_29687_, _29686_, _06347_);
  nand _79588_ (_29688_, _29687_, _29685_);
  not _79589_ (_29689_, _29674_);
  nor _79590_ (_29690_, _29689_, _12560_);
  nor _79591_ (_29692_, _29674_, _12550_);
  or _79592_ (_29693_, _29683_, _12536_);
  or _79593_ (_29694_, _12534_, _12186_);
  and _79594_ (_29695_, _29694_, _29693_);
  nor _79595_ (_29696_, _29695_, _07151_);
  or _79596_ (_29697_, _12393_, _29676_);
  and _79597_ (_29698_, _12498_, _12407_);
  nor _79598_ (_29699_, _29698_, _12499_);
  nand _79599_ (_29700_, _29699_, _25366_);
  and _79600_ (_29701_, _29700_, _12387_);
  nand _79601_ (_29702_, _29701_, _29697_);
  nor _79602_ (_29703_, _29689_, _12514_);
  not _79603_ (_29704_, _29703_);
  nor _79604_ (_29705_, _12517_, _29676_);
  and _79605_ (_29706_, _07487_, \oc8051_golden_model_1.PC [14]);
  and _79606_ (_29707_, _29706_, _29106_);
  nor _79607_ (_29708_, _29707_, _29705_);
  nor _79608_ (_29709_, _29708_, _12516_);
  nor _79609_ (_29710_, _29709_, _12387_);
  and _79610_ (_29711_, _29710_, _29704_);
  nor _79611_ (_29714_, _29711_, _07154_);
  nand _79612_ (_29715_, _29714_, _29702_);
  and _79613_ (_29716_, _29674_, _07154_);
  nor _79614_ (_29717_, _29716_, _06341_);
  and _79615_ (_29718_, _29717_, _29715_);
  or _79616_ (_29719_, _29718_, _29696_);
  nand _79617_ (_29720_, _29719_, _12541_);
  nor _79618_ (_29721_, _29674_, _12541_);
  nor _79619_ (_29722_, _29721_, _12546_);
  and _79620_ (_29723_, _29722_, _29720_);
  nor _79621_ (_29725_, _12545_, _29676_);
  nor _79622_ (_29726_, _29725_, _29723_);
  and _79623_ (_29727_, _29726_, _12550_);
  or _79624_ (_29728_, _29727_, _29692_);
  nand _79625_ (_29729_, _29728_, _06465_);
  nor _79626_ (_29730_, _12403_, _06465_);
  nor _79627_ (_29731_, _29730_, _25401_);
  and _79628_ (_29732_, _29731_, _29729_);
  or _79629_ (_29733_, _29732_, _29690_);
  nand _79630_ (_29734_, _29733_, _12565_);
  nor _79631_ (_29736_, _12565_, _29676_);
  nor _79632_ (_29737_, _29736_, _12379_);
  and _79633_ (_29738_, _29737_, _29734_);
  and _79634_ (_29739_, _12371_, _12186_);
  nor _79635_ (_29740_, _29684_, _12371_);
  or _79636_ (_29741_, _29740_, _12378_);
  nor _79637_ (_29742_, _29741_, _29739_);
  or _79638_ (_29743_, _29742_, _06347_);
  or _79639_ (_29744_, _29743_, _29738_);
  and _79640_ (_29745_, _29744_, _29688_);
  nand _79641_ (_29747_, _29745_, _06774_);
  and _79642_ (_29748_, _12587_, _12186_);
  nor _79643_ (_29749_, _29684_, _12587_);
  or _79644_ (_29750_, _29749_, _29748_);
  nor _79645_ (_29751_, _29750_, _06774_);
  nor _79646_ (_29752_, _29751_, _06371_);
  nand _79647_ (_29753_, _29752_, _29747_);
  and _79648_ (_29754_, _12604_, _12186_);
  and _79649_ (_29755_, _29683_, _26518_);
  or _79650_ (_29756_, _29755_, _29754_);
  and _79651_ (_29758_, _29756_, _06371_);
  nor _79652_ (_29759_, _29758_, _12174_);
  and _79653_ (_29760_, _29759_, _29753_);
  nor _79654_ (_29761_, _29674_, _12175_);
  or _79655_ (_29762_, _29761_, _29760_);
  and _79656_ (_29763_, _29762_, _12623_);
  nor _79657_ (_29764_, _12623_, _12403_);
  or _79658_ (_29765_, _29764_, _29763_);
  nand _79659_ (_29766_, _29765_, _12630_);
  nor _79660_ (_29767_, _29674_, _12630_);
  nor _79661_ (_29769_, _29767_, _12636_);
  nand _79662_ (_29770_, _29769_, _29766_);
  nor _79663_ (_29771_, _12635_, _29676_);
  nor _79664_ (_29772_, _29771_, _26197_);
  nand _79665_ (_29773_, _29772_, _29770_);
  nor _79666_ (_29774_, _29674_, _12639_);
  nor _79667_ (_29775_, _29774_, _12644_);
  nand _79668_ (_29776_, _29775_, _29773_);
  nor _79669_ (_29777_, _29676_, _12643_);
  nor _79670_ (_29778_, _29777_, _10515_);
  nand _79671_ (_29780_, _29778_, _29776_);
  nor _79672_ (_29781_, _29674_, _05984_);
  nor _79673_ (_29782_, _29781_, _12653_);
  nand _79674_ (_29783_, _29782_, _29780_);
  nor _79675_ (_29784_, _12652_, _29676_);
  nor _79676_ (_29785_, _29784_, _06373_);
  nand _79677_ (_29786_, _29785_, _29783_);
  nor _79678_ (_29787_, _12186_, _06374_);
  nor _79679_ (_29788_, _29787_, _12659_);
  nand _79680_ (_29789_, _29788_, _29786_);
  nor _79681_ (_29791_, _29676_, _07216_);
  nor _79682_ (_29792_, _29791_, _10094_);
  nand _79683_ (_29793_, _29792_, _29789_);
  nor _79684_ (_29794_, _12186_, _05982_);
  nor _79685_ (_29795_, _29794_, _25492_);
  nand _79686_ (_29796_, _29795_, _29793_);
  nor _79687_ (_29797_, _29689_, _12172_);
  nor _79688_ (_29798_, _29797_, _12670_);
  nand _79689_ (_29799_, _29798_, _29796_);
  nor _79690_ (_29800_, _12669_, _12403_);
  nor _79691_ (_29802_, _29800_, _12674_);
  and _79692_ (_29803_, _29802_, _29799_);
  and _79693_ (_29804_, _29699_, _12674_);
  nor _79694_ (_29805_, _29804_, _29803_);
  or _79695_ (_29806_, _29805_, _09031_);
  or _79696_ (_29807_, _29676_, _09030_);
  and _79697_ (_29808_, _29807_, _06219_);
  nand _79698_ (_29809_, _29808_, _29806_);
  nor _79699_ (_29810_, _12186_, _06219_);
  nor _79700_ (_29811_, _29810_, _10929_);
  nand _79701_ (_29813_, _29811_, _29809_);
  and _79702_ (_29814_, _12403_, _10929_);
  nor _79703_ (_29815_, _29814_, _12690_);
  nand _79704_ (_29816_, _29815_, _29813_);
  nor _79705_ (_29817_, _12723_, \oc8051_golden_model_1.DPH [6]);
  nor _79706_ (_29818_, _29817_, _12724_);
  nor _79707_ (_29819_, _29818_, _12691_);
  nor _79708_ (_29820_, _29819_, _12730_);
  and _79709_ (_29821_, _29820_, _29816_);
  or _79710_ (_29822_, _29821_, _29681_);
  nand _79711_ (_29824_, _29822_, _25064_);
  and _79712_ (_29825_, _12403_, _11342_);
  and _79713_ (_29826_, _29699_, _12759_);
  or _79714_ (_29827_, _29826_, _29825_);
  and _79715_ (_29828_, _29827_, _12733_);
  nor _79716_ (_29829_, _29828_, _12737_);
  nand _79717_ (_29830_, _29829_, _29824_);
  nor _79718_ (_29831_, _29674_, _12169_);
  nor _79719_ (_29832_, _29831_, _26610_);
  nand _79720_ (_29833_, _29832_, _29830_);
  nor _79721_ (_29835_, _29676_, _12166_);
  nor _79722_ (_29836_, _29835_, _06369_);
  nand _79723_ (_29837_, _29836_, _29833_);
  nor _79724_ (_29838_, _12186_, _07237_);
  nor _79725_ (_29839_, _29838_, _12752_);
  and _79726_ (_29840_, _29839_, _29837_);
  or _79727_ (_29841_, _29840_, _29679_);
  nand _79728_ (_29842_, _29841_, _25061_);
  and _79729_ (_29843_, _12403_, _12759_);
  and _79730_ (_29844_, _29699_, _11342_);
  or _79731_ (_29846_, _29844_, _29843_);
  and _79732_ (_29847_, _29846_, _12755_);
  nor _79733_ (_29848_, _29847_, _10980_);
  nand _79734_ (_29849_, _29848_, _29842_);
  nor _79735_ (_29850_, _29674_, _10979_);
  nor _79736_ (_29851_, _29850_, _26630_);
  nand _79737_ (_29852_, _29851_, _29849_);
  nor _79738_ (_29853_, _12164_, _29676_);
  nor _79739_ (_29854_, _29853_, _06375_);
  nand _79740_ (_29855_, _29854_, _29852_);
  nor _79741_ (_29857_, _12186_, _07242_);
  nor _79742_ (_29858_, _29857_, _12773_);
  and _79743_ (_29859_, _29858_, _29855_);
  or _79744_ (_29860_, _29859_, _29678_);
  nand _79745_ (_29861_, _29860_, _12782_);
  and _79746_ (_29862_, _12403_, \oc8051_golden_model_1.PSW [7]);
  and _79747_ (_29863_, _29699_, _10558_);
  or _79748_ (_29864_, _29863_, _29862_);
  and _79749_ (_29865_, _29864_, _12776_);
  nor _79750_ (_29866_, _29865_, _12780_);
  nand _79751_ (_29868_, _29866_, _29861_);
  nor _79752_ (_29869_, _29674_, _12162_);
  nor _79753_ (_29870_, _29869_, _11023_);
  nand _79754_ (_29871_, _29870_, _29868_);
  nor _79755_ (_29872_, _29676_, _11022_);
  nor _79756_ (_29873_, _29872_, _06366_);
  nand _79757_ (_29874_, _29873_, _29871_);
  nor _79758_ (_29875_, _12186_, _09056_);
  nor _79759_ (_29876_, _29875_, _12797_);
  and _79760_ (_29877_, _29876_, _29874_);
  or _79761_ (_29879_, _29877_, _29677_);
  nand _79762_ (_29880_, _29879_, _25056_);
  and _79763_ (_29881_, _12403_, _10558_);
  and _79764_ (_29882_, _29699_, \oc8051_golden_model_1.PSW [7]);
  or _79765_ (_29883_, _29882_, _29881_);
  and _79766_ (_29884_, _29883_, _12800_);
  nor _79767_ (_29885_, _29884_, _12804_);
  nand _79768_ (_29886_, _29885_, _29880_);
  nor _79769_ (_29887_, _29674_, _12154_);
  nor _79770_ (_29888_, _29887_, _14297_);
  nand _79771_ (_29890_, _29888_, _29886_);
  nor _79772_ (_29891_, _29676_, _12153_);
  nor _79773_ (_29892_, _29891_, _11125_);
  nand _79774_ (_29893_, _29892_, _29890_);
  nor _79775_ (_29894_, _29674_, _11126_);
  nor _79776_ (_29895_, _29894_, _06551_);
  nand _79777_ (_29896_, _29895_, _29893_);
  nor _79778_ (_29897_, _08142_, _06716_);
  nor _79779_ (_29898_, _29897_, _07253_);
  nand _79780_ (_29899_, _29898_, _29896_);
  nor _79781_ (_29901_, _12403_, _05959_);
  nor _79782_ (_29902_, _29901_, _06365_);
  nand _79783_ (_29903_, _29902_, _29899_);
  and _79784_ (_29904_, _29684_, _13004_);
  nor _79785_ (_29905_, _12186_, _13004_);
  or _79786_ (_29906_, _29905_, _06558_);
  or _79787_ (_29907_, _29906_, _29904_);
  and _79788_ (_29908_, _29907_, _12151_);
  nand _79789_ (_29909_, _29908_, _29903_);
  nor _79790_ (_29910_, _29674_, _12151_);
  nor _79791_ (_29912_, _29910_, _19056_);
  nand _79792_ (_29913_, _29912_, _29909_);
  nor _79793_ (_29914_, _13012_, _29676_);
  nor _79794_ (_29915_, _29914_, _11284_);
  and _79795_ (_29916_, _29915_, _29913_);
  or _79796_ (_29917_, _29916_, _29675_);
  nand _79797_ (_29918_, _29917_, _06282_);
  and _79798_ (_29919_, _08142_, _06281_);
  nor _79799_ (_29920_, _29919_, _25646_);
  nand _79800_ (_29921_, _29920_, _29918_);
  and _79801_ (_29923_, _12403_, _25646_);
  nor _79802_ (_29924_, _29923_, _06362_);
  and _79803_ (_29925_, _29924_, _29921_);
  and _79804_ (_29926_, _12187_, _13004_);
  nor _79805_ (_29927_, _29683_, _13004_);
  nor _79806_ (_29928_, _29927_, _29926_);
  nor _79807_ (_29929_, _29928_, _06921_);
  or _79808_ (_29930_, _29929_, _29925_);
  and _79809_ (_29931_, _29930_, _13030_);
  nor _79810_ (_29932_, _29674_, _13030_);
  or _79811_ (_29934_, _29932_, _29931_);
  nand _79812_ (_29935_, _29934_, _06926_);
  nor _79813_ (_29936_, _12403_, _06926_);
  nor _79814_ (_29937_, _29936_, _13038_);
  nand _79815_ (_29938_, _29937_, _29935_);
  nor _79816_ (_29939_, _29689_, _13037_);
  nor _79817_ (_29940_, _29939_, _06361_);
  nand _79818_ (_29941_, _29940_, _29938_);
  and _79819_ (_29942_, _06361_, _06317_);
  nor _79820_ (_29943_, _29942_, _05940_);
  nand _79821_ (_29945_, _29943_, _29941_);
  and _79822_ (_29946_, _12403_, _05940_);
  nor _79823_ (_29947_, _29946_, _05927_);
  nand _79824_ (_29948_, _29947_, _29945_);
  nor _79825_ (_29949_, _29928_, _05928_);
  nor _79826_ (_29950_, _29949_, _13053_);
  nand _79827_ (_29951_, _29950_, _29948_);
  nor _79828_ (_29952_, _29689_, _13052_);
  nor _79829_ (_29953_, _29952_, _06278_);
  nand _79830_ (_29954_, _29953_, _29951_);
  nor _79831_ (_29956_, _12403_, _06279_);
  nor _79832_ (_29957_, _29956_, _13059_);
  nand _79833_ (_29958_, _29957_, _29954_);
  nor _79834_ (_29959_, _29689_, _12141_);
  nor _79835_ (_29960_, _29959_, _06379_);
  and _79836_ (_29961_, _29960_, _29958_);
  and _79837_ (_29962_, _06379_, _06317_);
  or _79838_ (_29963_, _29962_, _29961_);
  nand _79839_ (_29964_, _29963_, _29058_);
  nor _79840_ (_29965_, _12403_, _29058_);
  nor _79841_ (_29967_, _29965_, _13068_);
  and _79842_ (_29968_, _29967_, _29964_);
  and _79843_ (_29969_, _29674_, _13068_);
  or _79844_ (_29970_, _29969_, _29968_);
  or _79845_ (_29971_, _29970_, _01351_);
  or _79846_ (_29972_, _01347_, \oc8051_golden_model_1.PC [14]);
  and _79847_ (_29973_, _29972_, _42618_);
  and _79848_ (_43261_, _29973_, _29971_);
  nand _79849_ (_29974_, _11263_, _07904_);
  and _79850_ (_29975_, _13077_, \oc8051_golden_model_1.P2 [0]);
  nor _79851_ (_29977_, _29975_, _07234_);
  nand _79852_ (_29978_, _29977_, _29974_);
  and _79853_ (_29979_, _07904_, _07133_);
  or _79854_ (_29980_, _29979_, _29975_);
  or _79855_ (_29981_, _29980_, _07215_);
  nor _79856_ (_29982_, _08390_, _13077_);
  or _79857_ (_29983_, _29982_, _29975_);
  or _79858_ (_29984_, _29983_, _07151_);
  and _79859_ (_29985_, _07904_, \oc8051_golden_model_1.ACC [0]);
  or _79860_ (_29986_, _29985_, _29975_);
  and _79861_ (_29988_, _29986_, _07141_);
  and _79862_ (_29989_, _07142_, \oc8051_golden_model_1.P2 [0]);
  or _79863_ (_29990_, _29989_, _06341_);
  or _79864_ (_29991_, _29990_, _29988_);
  and _79865_ (_29992_, _29991_, _06273_);
  and _79866_ (_29993_, _29992_, _29984_);
  and _79867_ (_29994_, _13085_, \oc8051_golden_model_1.P2 [0]);
  and _79868_ (_29995_, _14382_, _08624_);
  or _79869_ (_29996_, _29995_, _29994_);
  and _79870_ (_29997_, _29996_, _06272_);
  or _79871_ (_29999_, _29997_, _29993_);
  and _79872_ (_30000_, _29999_, _07166_);
  and _79873_ (_30001_, _29980_, _06461_);
  or _79874_ (_30002_, _30001_, _06464_);
  or _79875_ (_30003_, _30002_, _30000_);
  or _79876_ (_30004_, _29986_, _06465_);
  and _79877_ (_30005_, _30004_, _06269_);
  and _79878_ (_30006_, _30005_, _30003_);
  and _79879_ (_30007_, _29975_, _06268_);
  or _79880_ (_30008_, _30007_, _06261_);
  or _79881_ (_30010_, _30008_, _30006_);
  or _79882_ (_30011_, _29983_, _06262_);
  and _79883_ (_30012_, _30011_, _06258_);
  and _79884_ (_30013_, _30012_, _30010_);
  and _79885_ (_30014_, _14413_, _08624_);
  or _79886_ (_30015_, _30014_, _29994_);
  and _79887_ (_30016_, _30015_, _06257_);
  or _79888_ (_30017_, _30016_, _10080_);
  or _79889_ (_30018_, _30017_, _30013_);
  and _79890_ (_30019_, _30018_, _29981_);
  or _79891_ (_30021_, _30019_, _07460_);
  and _79892_ (_30022_, _09392_, _07904_);
  or _79893_ (_30023_, _29975_, _07208_);
  or _79894_ (_30024_, _30023_, _30022_);
  and _79895_ (_30025_, _30024_, _30021_);
  or _79896_ (_30026_, _30025_, _10094_);
  and _79897_ (_30027_, _14467_, _07904_);
  or _79898_ (_30028_, _29975_, _05982_);
  or _79899_ (_30029_, _30028_, _30027_);
  and _79900_ (_30030_, _30029_, _06219_);
  and _79901_ (_30032_, _30030_, _30026_);
  and _79902_ (_30033_, _07904_, _08954_);
  or _79903_ (_30034_, _30033_, _29975_);
  and _79904_ (_30035_, _30034_, _06218_);
  or _79905_ (_30036_, _30035_, _06369_);
  or _79906_ (_30037_, _30036_, _30032_);
  and _79907_ (_30038_, _14366_, _07904_);
  or _79908_ (_30039_, _30038_, _29975_);
  or _79909_ (_30040_, _30039_, _07237_);
  and _79910_ (_30041_, _30040_, _07240_);
  and _79911_ (_30043_, _30041_, _30037_);
  nor _79912_ (_30044_, _12580_, _13077_);
  or _79913_ (_30045_, _30044_, _29975_);
  and _79914_ (_30046_, _29974_, _06536_);
  and _79915_ (_30047_, _30046_, _30045_);
  or _79916_ (_30048_, _30047_, _30043_);
  and _79917_ (_30049_, _30048_, _07242_);
  nand _79918_ (_30050_, _30034_, _06375_);
  nor _79919_ (_30051_, _30050_, _29982_);
  or _79920_ (_30052_, _30051_, _06545_);
  or _79921_ (_30054_, _30052_, _30049_);
  and _79922_ (_30055_, _30054_, _29978_);
  or _79923_ (_30056_, _30055_, _06366_);
  and _79924_ (_30057_, _14363_, _07904_);
  or _79925_ (_30058_, _29975_, _09056_);
  or _79926_ (_30059_, _30058_, _30057_);
  and _79927_ (_30060_, _30059_, _09061_);
  and _79928_ (_30061_, _30060_, _30056_);
  and _79929_ (_30062_, _30045_, _06528_);
  or _79930_ (_30063_, _30062_, _06568_);
  or _79931_ (_30065_, _30063_, _30061_);
  or _79932_ (_30066_, _29983_, _06926_);
  and _79933_ (_30067_, _30066_, _30065_);
  or _79934_ (_30068_, _30067_, _05927_);
  or _79935_ (_30069_, _29975_, _05928_);
  and _79936_ (_30070_, _30069_, _30068_);
  or _79937_ (_30071_, _30070_, _06278_);
  or _79938_ (_30072_, _29983_, _06279_);
  and _79939_ (_30073_, _30072_, _01347_);
  and _79940_ (_30074_, _30073_, _30071_);
  nor _79941_ (_30076_, \oc8051_golden_model_1.P2 [0], rst);
  nor _79942_ (_30077_, _30076_, _01354_);
  or _79943_ (_43262_, _30077_, _30074_);
  nor _79944_ (_30078_, \oc8051_golden_model_1.P2 [1], rst);
  nor _79945_ (_30079_, _30078_, _01354_);
  and _79946_ (_30080_, _13077_, \oc8051_golden_model_1.P2 [1]);
  nor _79947_ (_30081_, _11261_, _13077_);
  or _79948_ (_30082_, _30081_, _30080_);
  or _79949_ (_30083_, _30082_, _09061_);
  nand _79950_ (_30084_, _07904_, _07038_);
  or _79951_ (_30086_, _07904_, \oc8051_golden_model_1.P2 [1]);
  and _79952_ (_30087_, _30086_, _06218_);
  and _79953_ (_30088_, _30087_, _30084_);
  nor _79954_ (_30089_, _13077_, _07357_);
  or _79955_ (_30090_, _30089_, _30080_);
  and _79956_ (_30091_, _30090_, _06461_);
  and _79957_ (_30092_, _13085_, \oc8051_golden_model_1.P2 [1]);
  and _79958_ (_30093_, _14557_, _08624_);
  or _79959_ (_30094_, _30093_, _30092_);
  or _79960_ (_30095_, _30094_, _06273_);
  and _79961_ (_30097_, _14562_, _07904_);
  not _79962_ (_30098_, _30097_);
  and _79963_ (_30099_, _30098_, _30086_);
  and _79964_ (_30100_, _30099_, _06341_);
  and _79965_ (_30101_, _07142_, \oc8051_golden_model_1.P2 [1]);
  and _79966_ (_30102_, _07904_, \oc8051_golden_model_1.ACC [1]);
  or _79967_ (_30103_, _30102_, _30080_);
  and _79968_ (_30104_, _30103_, _07141_);
  or _79969_ (_30105_, _30104_, _30101_);
  and _79970_ (_30106_, _30105_, _07151_);
  or _79971_ (_30108_, _30106_, _06272_);
  or _79972_ (_30109_, _30108_, _30100_);
  and _79973_ (_30110_, _30109_, _30095_);
  and _79974_ (_30111_, _30110_, _07166_);
  or _79975_ (_30112_, _30111_, _30091_);
  or _79976_ (_30113_, _30112_, _06464_);
  or _79977_ (_30114_, _30103_, _06465_);
  and _79978_ (_30115_, _30114_, _06269_);
  and _79979_ (_30116_, _30115_, _30113_);
  and _79980_ (_30117_, _14560_, _08624_);
  or _79981_ (_30119_, _30117_, _30092_);
  and _79982_ (_30120_, _30119_, _06268_);
  or _79983_ (_30121_, _30120_, _06261_);
  or _79984_ (_30122_, _30121_, _30116_);
  or _79985_ (_30123_, _30092_, _14556_);
  and _79986_ (_30124_, _30123_, _30094_);
  or _79987_ (_30125_, _30124_, _06262_);
  and _79988_ (_30126_, _30125_, _06258_);
  and _79989_ (_30127_, _30126_, _30122_);
  or _79990_ (_30128_, _30092_, _14597_);
  and _79991_ (_30130_, _30128_, _06257_);
  and _79992_ (_30131_, _30130_, _30094_);
  or _79993_ (_30132_, _30131_, _10080_);
  or _79994_ (_30133_, _30132_, _30127_);
  or _79995_ (_30134_, _30090_, _07215_);
  and _79996_ (_30135_, _30134_, _30133_);
  or _79997_ (_30136_, _30135_, _07460_);
  and _79998_ (_30137_, _09451_, _07904_);
  or _79999_ (_30138_, _30080_, _07208_);
  or _80000_ (_30139_, _30138_, _30137_);
  and _80001_ (_30141_, _30139_, _05982_);
  and _80002_ (_30142_, _30141_, _30136_);
  and _80003_ (_30143_, _14653_, _07904_);
  or _80004_ (_30144_, _30143_, _30080_);
  and _80005_ (_30145_, _30144_, _10094_);
  or _80006_ (_30146_, _30145_, _30142_);
  and _80007_ (_30147_, _30146_, _06219_);
  or _80008_ (_30148_, _30147_, _30088_);
  and _80009_ (_30149_, _30148_, _07237_);
  or _80010_ (_30150_, _14668_, _13077_);
  and _80011_ (_30152_, _30086_, _06369_);
  and _80012_ (_30153_, _30152_, _30150_);
  or _80013_ (_30154_, _30153_, _06536_);
  or _80014_ (_30155_, _30154_, _30149_);
  nand _80015_ (_30156_, _11260_, _07904_);
  and _80016_ (_30157_, _30156_, _30082_);
  or _80017_ (_30158_, _30157_, _07240_);
  and _80018_ (_30159_, _30158_, _07242_);
  and _80019_ (_30160_, _30159_, _30155_);
  or _80020_ (_30161_, _14666_, _13077_);
  and _80021_ (_30163_, _30086_, _06375_);
  and _80022_ (_30164_, _30163_, _30161_);
  or _80023_ (_30165_, _30164_, _06545_);
  or _80024_ (_30166_, _30165_, _30160_);
  nor _80025_ (_30167_, _30080_, _07234_);
  nand _80026_ (_30168_, _30167_, _30156_);
  and _80027_ (_30169_, _30168_, _09056_);
  and _80028_ (_30170_, _30169_, _30166_);
  or _80029_ (_30171_, _30084_, _08341_);
  and _80030_ (_30172_, _30086_, _06366_);
  and _80031_ (_30174_, _30172_, _30171_);
  or _80032_ (_30175_, _30174_, _06528_);
  or _80033_ (_30176_, _30175_, _30170_);
  and _80034_ (_30177_, _30176_, _30083_);
  or _80035_ (_30178_, _30177_, _06568_);
  or _80036_ (_30179_, _30099_, _06926_);
  and _80037_ (_30180_, _30179_, _05928_);
  and _80038_ (_30181_, _30180_, _30178_);
  and _80039_ (_30182_, _30119_, _05927_);
  or _80040_ (_30183_, _30182_, _06278_);
  or _80041_ (_30185_, _30183_, _30181_);
  or _80042_ (_30186_, _30080_, _06279_);
  or _80043_ (_30187_, _30186_, _30097_);
  and _80044_ (_30188_, _30187_, _01347_);
  and _80045_ (_30189_, _30188_, _30185_);
  or _80046_ (_43264_, _30189_, _30079_);
  and _80047_ (_30190_, _13077_, \oc8051_golden_model_1.P2 [2]);
  nor _80048_ (_30191_, _13077_, _07776_);
  or _80049_ (_30192_, _30191_, _30190_);
  or _80050_ (_30193_, _30192_, _07215_);
  or _80051_ (_30195_, _30192_, _07166_);
  and _80052_ (_30196_, _14770_, _07904_);
  or _80053_ (_30197_, _30196_, _30190_);
  or _80054_ (_30198_, _30197_, _07151_);
  and _80055_ (_30199_, _07904_, \oc8051_golden_model_1.ACC [2]);
  or _80056_ (_30200_, _30199_, _30190_);
  and _80057_ (_30201_, _30200_, _07141_);
  and _80058_ (_30202_, _07142_, \oc8051_golden_model_1.P2 [2]);
  or _80059_ (_30203_, _30202_, _06341_);
  or _80060_ (_30204_, _30203_, _30201_);
  and _80061_ (_30206_, _30204_, _06273_);
  and _80062_ (_30207_, _30206_, _30198_);
  and _80063_ (_30208_, _13085_, \oc8051_golden_model_1.P2 [2]);
  and _80064_ (_30209_, _14774_, _08624_);
  or _80065_ (_30210_, _30209_, _30208_);
  and _80066_ (_30211_, _30210_, _06272_);
  or _80067_ (_30212_, _30211_, _06461_);
  or _80068_ (_30213_, _30212_, _30207_);
  and _80069_ (_30214_, _30213_, _30195_);
  or _80070_ (_30215_, _30214_, _06464_);
  or _80071_ (_30217_, _30200_, _06465_);
  and _80072_ (_30218_, _30217_, _06269_);
  and _80073_ (_30219_, _30218_, _30215_);
  and _80074_ (_30220_, _14756_, _08624_);
  or _80075_ (_30221_, _30220_, _30208_);
  and _80076_ (_30222_, _30221_, _06268_);
  or _80077_ (_30223_, _30222_, _06261_);
  or _80078_ (_30224_, _30223_, _30219_);
  and _80079_ (_30225_, _30209_, _14789_);
  or _80080_ (_30226_, _30208_, _06262_);
  or _80081_ (_30228_, _30226_, _30225_);
  and _80082_ (_30229_, _30228_, _06258_);
  and _80083_ (_30230_, _30229_, _30224_);
  and _80084_ (_30231_, _14804_, _08624_);
  or _80085_ (_30232_, _30231_, _30208_);
  and _80086_ (_30233_, _30232_, _06257_);
  or _80087_ (_30234_, _30233_, _10080_);
  or _80088_ (_30235_, _30234_, _30230_);
  and _80089_ (_30236_, _30235_, _30193_);
  or _80090_ (_30237_, _30236_, _07460_);
  and _80091_ (_30239_, _09450_, _07904_);
  or _80092_ (_30240_, _30190_, _07208_);
  or _80093_ (_30241_, _30240_, _30239_);
  and _80094_ (_30242_, _30241_, _05982_);
  and _80095_ (_30243_, _30242_, _30237_);
  and _80096_ (_30244_, _14859_, _07904_);
  or _80097_ (_30245_, _30244_, _30190_);
  and _80098_ (_30246_, _30245_, _10094_);
  or _80099_ (_30247_, _30246_, _06218_);
  or _80100_ (_30248_, _30247_, _30243_);
  and _80101_ (_30250_, _07904_, _08973_);
  or _80102_ (_30251_, _30250_, _30190_);
  or _80103_ (_30252_, _30251_, _06219_);
  and _80104_ (_30253_, _30252_, _30248_);
  or _80105_ (_30254_, _30253_, _06369_);
  and _80106_ (_30255_, _14751_, _07904_);
  or _80107_ (_30256_, _30255_, _30190_);
  or _80108_ (_30257_, _30256_, _07237_);
  and _80109_ (_30258_, _30257_, _07240_);
  and _80110_ (_30259_, _30258_, _30254_);
  and _80111_ (_30261_, _11259_, _07904_);
  or _80112_ (_30262_, _30261_, _30190_);
  and _80113_ (_30263_, _30262_, _06536_);
  or _80114_ (_30264_, _30263_, _30259_);
  and _80115_ (_30265_, _30264_, _07242_);
  or _80116_ (_30266_, _30190_, _08440_);
  and _80117_ (_30267_, _30251_, _06375_);
  and _80118_ (_30268_, _30267_, _30266_);
  or _80119_ (_30269_, _30268_, _30265_);
  and _80120_ (_30270_, _30269_, _07234_);
  and _80121_ (_30272_, _30200_, _06545_);
  and _80122_ (_30273_, _30272_, _30266_);
  or _80123_ (_30274_, _30273_, _06366_);
  or _80124_ (_30275_, _30274_, _30270_);
  and _80125_ (_30276_, _14748_, _07904_);
  or _80126_ (_30277_, _30190_, _09056_);
  or _80127_ (_30278_, _30277_, _30276_);
  and _80128_ (_30279_, _30278_, _09061_);
  and _80129_ (_30280_, _30279_, _30275_);
  nor _80130_ (_30281_, _11258_, _13077_);
  or _80131_ (_30283_, _30281_, _30190_);
  and _80132_ (_30284_, _30283_, _06528_);
  or _80133_ (_30285_, _30284_, _06568_);
  or _80134_ (_30286_, _30285_, _30280_);
  or _80135_ (_30287_, _30197_, _06926_);
  and _80136_ (_30288_, _30287_, _05928_);
  and _80137_ (_30289_, _30288_, _30286_);
  and _80138_ (_30290_, _30221_, _05927_);
  or _80139_ (_30291_, _30290_, _06278_);
  or _80140_ (_30292_, _30291_, _30289_);
  and _80141_ (_30294_, _14926_, _07904_);
  or _80142_ (_30295_, _30190_, _06279_);
  or _80143_ (_30296_, _30295_, _30294_);
  and _80144_ (_30297_, _30296_, _01347_);
  and _80145_ (_30298_, _30297_, _30292_);
  nor _80146_ (_30299_, \oc8051_golden_model_1.P2 [2], rst);
  nor _80147_ (_30300_, _30299_, _01354_);
  or _80148_ (_43265_, _30300_, _30298_);
  and _80149_ (_30301_, _13077_, \oc8051_golden_model_1.P2 [3]);
  nor _80150_ (_30302_, _13077_, _07594_);
  or _80151_ (_30304_, _30302_, _30301_);
  or _80152_ (_30305_, _30304_, _07215_);
  and _80153_ (_30306_, _14953_, _07904_);
  or _80154_ (_30307_, _30306_, _30301_);
  or _80155_ (_30308_, _30307_, _07151_);
  and _80156_ (_30309_, _07904_, \oc8051_golden_model_1.ACC [3]);
  or _80157_ (_30310_, _30309_, _30301_);
  and _80158_ (_30311_, _30310_, _07141_);
  and _80159_ (_30312_, _07142_, \oc8051_golden_model_1.P2 [3]);
  or _80160_ (_30313_, _30312_, _06341_);
  or _80161_ (_30315_, _30313_, _30311_);
  and _80162_ (_30316_, _30315_, _06273_);
  and _80163_ (_30317_, _30316_, _30308_);
  and _80164_ (_30318_, _13085_, \oc8051_golden_model_1.P2 [3]);
  and _80165_ (_30319_, _14950_, _08624_);
  or _80166_ (_30320_, _30319_, _30318_);
  and _80167_ (_30321_, _30320_, _06272_);
  or _80168_ (_30322_, _30321_, _06461_);
  or _80169_ (_30323_, _30322_, _30317_);
  or _80170_ (_30324_, _30304_, _07166_);
  and _80171_ (_30325_, _30324_, _30323_);
  or _80172_ (_30326_, _30325_, _06464_);
  or _80173_ (_30327_, _30310_, _06465_);
  and _80174_ (_30328_, _30327_, _06269_);
  and _80175_ (_30329_, _30328_, _30326_);
  and _80176_ (_30330_, _14948_, _08624_);
  or _80177_ (_30331_, _30330_, _30318_);
  and _80178_ (_30332_, _30331_, _06268_);
  or _80179_ (_30333_, _30332_, _06261_);
  or _80180_ (_30334_, _30333_, _30329_);
  or _80181_ (_30337_, _30318_, _14979_);
  and _80182_ (_30338_, _30337_, _30320_);
  or _80183_ (_30339_, _30338_, _06262_);
  and _80184_ (_30340_, _30339_, _06258_);
  and _80185_ (_30341_, _30340_, _30334_);
  or _80186_ (_30342_, _30318_, _14992_);
  and _80187_ (_30343_, _30342_, _06257_);
  and _80188_ (_30344_, _30343_, _30320_);
  or _80189_ (_30345_, _30344_, _10080_);
  or _80190_ (_30346_, _30345_, _30341_);
  and _80191_ (_30348_, _30346_, _30305_);
  or _80192_ (_30349_, _30348_, _07460_);
  and _80193_ (_30350_, _09449_, _07904_);
  or _80194_ (_30351_, _30301_, _07208_);
  or _80195_ (_30352_, _30351_, _30350_);
  and _80196_ (_30353_, _30352_, _05982_);
  and _80197_ (_30354_, _30353_, _30349_);
  and _80198_ (_30355_, _15048_, _07904_);
  or _80199_ (_30356_, _30355_, _30301_);
  and _80200_ (_30357_, _30356_, _10094_);
  or _80201_ (_30359_, _30357_, _06218_);
  or _80202_ (_30360_, _30359_, _30354_);
  and _80203_ (_30361_, _07904_, _08930_);
  or _80204_ (_30362_, _30361_, _30301_);
  or _80205_ (_30363_, _30362_, _06219_);
  and _80206_ (_30364_, _30363_, _30360_);
  or _80207_ (_30365_, _30364_, _06369_);
  and _80208_ (_30366_, _14943_, _07904_);
  or _80209_ (_30367_, _30366_, _30301_);
  or _80210_ (_30368_, _30367_, _07237_);
  and _80211_ (_30370_, _30368_, _07240_);
  and _80212_ (_30371_, _30370_, _30365_);
  and _80213_ (_30372_, _12577_, _07904_);
  or _80214_ (_30373_, _30372_, _30301_);
  and _80215_ (_30374_, _30373_, _06536_);
  or _80216_ (_30375_, _30374_, _30371_);
  and _80217_ (_30376_, _30375_, _07242_);
  or _80218_ (_30377_, _30301_, _08292_);
  and _80219_ (_30378_, _30362_, _06375_);
  and _80220_ (_30379_, _30378_, _30377_);
  or _80221_ (_30381_, _30379_, _30376_);
  and _80222_ (_30382_, _30381_, _07234_);
  and _80223_ (_30383_, _30310_, _06545_);
  and _80224_ (_30384_, _30383_, _30377_);
  or _80225_ (_30385_, _30384_, _06366_);
  or _80226_ (_30386_, _30385_, _30382_);
  and _80227_ (_30387_, _14940_, _07904_);
  or _80228_ (_30388_, _30301_, _09056_);
  or _80229_ (_30389_, _30388_, _30387_);
  and _80230_ (_30390_, _30389_, _09061_);
  and _80231_ (_30392_, _30390_, _30386_);
  nor _80232_ (_30393_, _11256_, _13077_);
  or _80233_ (_30394_, _30393_, _30301_);
  and _80234_ (_30395_, _30394_, _06528_);
  or _80235_ (_30396_, _30395_, _06568_);
  or _80236_ (_30397_, _30396_, _30392_);
  or _80237_ (_30398_, _30307_, _06926_);
  and _80238_ (_30399_, _30398_, _05928_);
  and _80239_ (_30400_, _30399_, _30397_);
  and _80240_ (_30401_, _30331_, _05927_);
  or _80241_ (_30403_, _30401_, _06278_);
  or _80242_ (_30404_, _30403_, _30400_);
  and _80243_ (_30405_, _15128_, _07904_);
  or _80244_ (_30406_, _30301_, _06279_);
  or _80245_ (_30407_, _30406_, _30405_);
  and _80246_ (_30408_, _30407_, _01347_);
  and _80247_ (_30409_, _30408_, _30404_);
  nor _80248_ (_30410_, \oc8051_golden_model_1.P2 [3], rst);
  nor _80249_ (_30411_, _30410_, _01354_);
  or _80250_ (_43266_, _30411_, _30409_);
  nor _80251_ (_30413_, \oc8051_golden_model_1.P2 [4], rst);
  nor _80252_ (_30414_, _30413_, _01354_);
  and _80253_ (_30415_, _13077_, \oc8051_golden_model_1.P2 [4]);
  nor _80254_ (_30416_, _08541_, _13077_);
  or _80255_ (_30417_, _30416_, _30415_);
  or _80256_ (_30418_, _30417_, _07215_);
  and _80257_ (_30419_, _13085_, \oc8051_golden_model_1.P2 [4]);
  and _80258_ (_30420_, _15176_, _08624_);
  or _80259_ (_30421_, _30420_, _30419_);
  and _80260_ (_30422_, _30421_, _06268_);
  and _80261_ (_30424_, _15162_, _07904_);
  or _80262_ (_30425_, _30424_, _30415_);
  or _80263_ (_30426_, _30425_, _07151_);
  and _80264_ (_30427_, _07904_, \oc8051_golden_model_1.ACC [4]);
  or _80265_ (_30428_, _30427_, _30415_);
  and _80266_ (_30429_, _30428_, _07141_);
  and _80267_ (_30430_, _07142_, \oc8051_golden_model_1.P2 [4]);
  or _80268_ (_30431_, _30430_, _06341_);
  or _80269_ (_30432_, _30431_, _30429_);
  and _80270_ (_30433_, _30432_, _06273_);
  and _80271_ (_30435_, _30433_, _30426_);
  and _80272_ (_30436_, _15166_, _08624_);
  or _80273_ (_30437_, _30436_, _30419_);
  and _80274_ (_30438_, _30437_, _06272_);
  or _80275_ (_30439_, _30438_, _06461_);
  or _80276_ (_30440_, _30439_, _30435_);
  or _80277_ (_30441_, _30417_, _07166_);
  and _80278_ (_30442_, _30441_, _30440_);
  or _80279_ (_30443_, _30442_, _06464_);
  or _80280_ (_30444_, _30428_, _06465_);
  and _80281_ (_30446_, _30444_, _06269_);
  and _80282_ (_30447_, _30446_, _30443_);
  or _80283_ (_30448_, _30447_, _30422_);
  and _80284_ (_30449_, _30448_, _06262_);
  and _80285_ (_30450_, _15184_, _08624_);
  or _80286_ (_30451_, _30450_, _30419_);
  and _80287_ (_30452_, _30451_, _06261_);
  or _80288_ (_30453_, _30452_, _30449_);
  and _80289_ (_30454_, _30453_, _06258_);
  and _80290_ (_30455_, _15200_, _08624_);
  or _80291_ (_30457_, _30455_, _30419_);
  and _80292_ (_30458_, _30457_, _06257_);
  or _80293_ (_30459_, _30458_, _10080_);
  or _80294_ (_30460_, _30459_, _30454_);
  and _80295_ (_30461_, _30460_, _30418_);
  or _80296_ (_30462_, _30461_, _07460_);
  and _80297_ (_30463_, _09448_, _07904_);
  or _80298_ (_30464_, _30415_, _07208_);
  or _80299_ (_30465_, _30464_, _30463_);
  and _80300_ (_30466_, _30465_, _05982_);
  and _80301_ (_30468_, _30466_, _30462_);
  and _80302_ (_30469_, _15254_, _07904_);
  or _80303_ (_30470_, _30469_, _30415_);
  and _80304_ (_30471_, _30470_, _10094_);
  or _80305_ (_30472_, _30471_, _06218_);
  or _80306_ (_30473_, _30472_, _30468_);
  and _80307_ (_30474_, _08959_, _07904_);
  or _80308_ (_30475_, _30474_, _30415_);
  or _80309_ (_30476_, _30475_, _06219_);
  and _80310_ (_30477_, _30476_, _30473_);
  or _80311_ (_30479_, _30477_, _06369_);
  and _80312_ (_30480_, _15269_, _07904_);
  or _80313_ (_30481_, _30480_, _30415_);
  or _80314_ (_30482_, _30481_, _07237_);
  and _80315_ (_30483_, _30482_, _07240_);
  and _80316_ (_30484_, _30483_, _30479_);
  and _80317_ (_30485_, _11254_, _07904_);
  or _80318_ (_30486_, _30485_, _30415_);
  and _80319_ (_30487_, _30486_, _06536_);
  or _80320_ (_30488_, _30487_, _30484_);
  and _80321_ (_30490_, _30488_, _07242_);
  or _80322_ (_30491_, _30415_, _08544_);
  and _80323_ (_30492_, _30475_, _06375_);
  and _80324_ (_30493_, _30492_, _30491_);
  or _80325_ (_30494_, _30493_, _30490_);
  and _80326_ (_30495_, _30494_, _07234_);
  and _80327_ (_30496_, _30428_, _06545_);
  and _80328_ (_30497_, _30496_, _30491_);
  or _80329_ (_30498_, _30497_, _06366_);
  or _80330_ (_30499_, _30498_, _30495_);
  and _80331_ (_30501_, _15266_, _07904_);
  or _80332_ (_30502_, _30415_, _09056_);
  or _80333_ (_30503_, _30502_, _30501_);
  and _80334_ (_30504_, _30503_, _09061_);
  and _80335_ (_30505_, _30504_, _30499_);
  nor _80336_ (_30506_, _11253_, _13077_);
  or _80337_ (_30507_, _30506_, _30415_);
  and _80338_ (_30508_, _30507_, _06528_);
  or _80339_ (_30509_, _30508_, _06568_);
  or _80340_ (_30510_, _30509_, _30505_);
  or _80341_ (_30512_, _30425_, _06926_);
  and _80342_ (_30513_, _30512_, _05928_);
  and _80343_ (_30514_, _30513_, _30510_);
  and _80344_ (_30515_, _30421_, _05927_);
  or _80345_ (_30516_, _30515_, _06278_);
  or _80346_ (_30517_, _30516_, _30514_);
  and _80347_ (_30518_, _15329_, _07904_);
  or _80348_ (_30519_, _30415_, _06279_);
  or _80349_ (_30520_, _30519_, _30518_);
  and _80350_ (_30521_, _30520_, _01347_);
  and _80351_ (_30523_, _30521_, _30517_);
  or _80352_ (_43267_, _30523_, _30414_);
  and _80353_ (_30524_, _13077_, \oc8051_golden_model_1.P2 [5]);
  and _80354_ (_30525_, _15358_, _07904_);
  or _80355_ (_30526_, _30525_, _30524_);
  or _80356_ (_30527_, _30526_, _07151_);
  and _80357_ (_30528_, _07904_, \oc8051_golden_model_1.ACC [5]);
  or _80358_ (_30529_, _30528_, _30524_);
  and _80359_ (_30530_, _30529_, _07141_);
  and _80360_ (_30531_, _07142_, \oc8051_golden_model_1.P2 [5]);
  or _80361_ (_30533_, _30531_, _06341_);
  or _80362_ (_30534_, _30533_, _30530_);
  and _80363_ (_30535_, _30534_, _06273_);
  and _80364_ (_30536_, _30535_, _30527_);
  and _80365_ (_30537_, _13085_, \oc8051_golden_model_1.P2 [5]);
  and _80366_ (_30538_, _15372_, _08624_);
  or _80367_ (_30539_, _30538_, _30537_);
  and _80368_ (_30540_, _30539_, _06272_);
  or _80369_ (_30541_, _30540_, _06461_);
  or _80370_ (_30542_, _30541_, _30536_);
  nor _80371_ (_30544_, _08244_, _13077_);
  or _80372_ (_30545_, _30544_, _30524_);
  or _80373_ (_30546_, _30545_, _07166_);
  and _80374_ (_30547_, _30546_, _30542_);
  or _80375_ (_30548_, _30547_, _06464_);
  or _80376_ (_30549_, _30529_, _06465_);
  and _80377_ (_30550_, _30549_, _06269_);
  and _80378_ (_30551_, _30550_, _30548_);
  and _80379_ (_30552_, _15355_, _08624_);
  or _80380_ (_30553_, _30552_, _30537_);
  and _80381_ (_30555_, _30553_, _06268_);
  or _80382_ (_30556_, _30555_, _06261_);
  or _80383_ (_30557_, _30556_, _30551_);
  or _80384_ (_30558_, _30537_, _15387_);
  and _80385_ (_30559_, _30558_, _30539_);
  or _80386_ (_30560_, _30559_, _06262_);
  and _80387_ (_30561_, _30560_, _06258_);
  and _80388_ (_30562_, _30561_, _30557_);
  or _80389_ (_30563_, _30537_, _15403_);
  and _80390_ (_30564_, _30563_, _06257_);
  and _80391_ (_30566_, _30564_, _30539_);
  or _80392_ (_30567_, _30566_, _10080_);
  or _80393_ (_30568_, _30567_, _30562_);
  or _80394_ (_30569_, _30545_, _07215_);
  and _80395_ (_30570_, _30569_, _30568_);
  or _80396_ (_30571_, _30570_, _07460_);
  and _80397_ (_30572_, _09447_, _07904_);
  or _80398_ (_30573_, _30524_, _07208_);
  or _80399_ (_30574_, _30573_, _30572_);
  and _80400_ (_30575_, _30574_, _05982_);
  and _80401_ (_30577_, _30575_, _30571_);
  and _80402_ (_30578_, _15459_, _07904_);
  or _80403_ (_30579_, _30578_, _30524_);
  and _80404_ (_30580_, _30579_, _10094_);
  or _80405_ (_30581_, _30580_, _06218_);
  or _80406_ (_30582_, _30581_, _30577_);
  and _80407_ (_30583_, _08946_, _07904_);
  or _80408_ (_30584_, _30583_, _30524_);
  or _80409_ (_30585_, _30584_, _06219_);
  and _80410_ (_30586_, _30585_, _30582_);
  or _80411_ (_30588_, _30586_, _06369_);
  and _80412_ (_30589_, _15353_, _07904_);
  or _80413_ (_30590_, _30589_, _30524_);
  or _80414_ (_30591_, _30590_, _07237_);
  and _80415_ (_30592_, _30591_, _07240_);
  and _80416_ (_30593_, _30592_, _30588_);
  and _80417_ (_30594_, _11250_, _07904_);
  or _80418_ (_30595_, _30594_, _30524_);
  and _80419_ (_30596_, _30595_, _06536_);
  or _80420_ (_30597_, _30596_, _30593_);
  and _80421_ (_30599_, _30597_, _07242_);
  or _80422_ (_30600_, _30524_, _08247_);
  and _80423_ (_30601_, _30584_, _06375_);
  and _80424_ (_30602_, _30601_, _30600_);
  or _80425_ (_30603_, _30602_, _30599_);
  and _80426_ (_30604_, _30603_, _07234_);
  and _80427_ (_30605_, _30529_, _06545_);
  and _80428_ (_30606_, _30605_, _30600_);
  or _80429_ (_30607_, _30606_, _06366_);
  or _80430_ (_30608_, _30607_, _30604_);
  and _80431_ (_30610_, _15350_, _07904_);
  or _80432_ (_30611_, _30524_, _09056_);
  or _80433_ (_30612_, _30611_, _30610_);
  and _80434_ (_30613_, _30612_, _09061_);
  and _80435_ (_30614_, _30613_, _30608_);
  nor _80436_ (_30615_, _11249_, _13077_);
  or _80437_ (_30616_, _30615_, _30524_);
  and _80438_ (_30617_, _30616_, _06528_);
  or _80439_ (_30618_, _30617_, _06568_);
  or _80440_ (_30619_, _30618_, _30614_);
  or _80441_ (_30621_, _30526_, _06926_);
  and _80442_ (_30622_, _30621_, _05928_);
  and _80443_ (_30623_, _30622_, _30619_);
  and _80444_ (_30624_, _30553_, _05927_);
  or _80445_ (_30625_, _30624_, _06278_);
  or _80446_ (_30626_, _30625_, _30623_);
  and _80447_ (_30627_, _15532_, _07904_);
  or _80448_ (_30628_, _30524_, _06279_);
  or _80449_ (_30629_, _30628_, _30627_);
  and _80450_ (_30630_, _30629_, _01347_);
  and _80451_ (_30632_, _30630_, _30626_);
  nor _80452_ (_30633_, \oc8051_golden_model_1.P2 [5], rst);
  nor _80453_ (_30634_, _30633_, _01354_);
  or _80454_ (_43268_, _30634_, _30632_);
  nor _80455_ (_30635_, \oc8051_golden_model_1.P2 [6], rst);
  nor _80456_ (_30636_, _30635_, _01354_);
  and _80457_ (_30637_, _13077_, \oc8051_golden_model_1.P2 [6]);
  and _80458_ (_30638_, _15554_, _07904_);
  or _80459_ (_30639_, _30638_, _30637_);
  or _80460_ (_30640_, _30639_, _07151_);
  and _80461_ (_30642_, _07904_, \oc8051_golden_model_1.ACC [6]);
  or _80462_ (_30643_, _30642_, _30637_);
  and _80463_ (_30644_, _30643_, _07141_);
  and _80464_ (_30645_, _07142_, \oc8051_golden_model_1.P2 [6]);
  or _80465_ (_30646_, _30645_, _06341_);
  or _80466_ (_30647_, _30646_, _30644_);
  and _80467_ (_30648_, _30647_, _06273_);
  and _80468_ (_30649_, _30648_, _30640_);
  and _80469_ (_30650_, _13085_, \oc8051_golden_model_1.P2 [6]);
  and _80470_ (_30651_, _15570_, _08624_);
  or _80471_ (_30653_, _30651_, _30650_);
  and _80472_ (_30654_, _30653_, _06272_);
  or _80473_ (_30655_, _30654_, _06461_);
  or _80474_ (_30656_, _30655_, _30649_);
  nor _80475_ (_30657_, _08142_, _13077_);
  or _80476_ (_30658_, _30657_, _30637_);
  or _80477_ (_30659_, _30658_, _07166_);
  and _80478_ (_30660_, _30659_, _30656_);
  or _80479_ (_30661_, _30660_, _06464_);
  or _80480_ (_30662_, _30643_, _06465_);
  and _80481_ (_30664_, _30662_, _06269_);
  and _80482_ (_30665_, _30664_, _30661_);
  and _80483_ (_30666_, _15551_, _08624_);
  or _80484_ (_30667_, _30666_, _30650_);
  and _80485_ (_30668_, _30667_, _06268_);
  or _80486_ (_30669_, _30668_, _06261_);
  or _80487_ (_30670_, _30669_, _30665_);
  or _80488_ (_30671_, _30650_, _15585_);
  and _80489_ (_30672_, _30671_, _30653_);
  or _80490_ (_30673_, _30672_, _06262_);
  and _80491_ (_30675_, _30673_, _06258_);
  and _80492_ (_30676_, _30675_, _30670_);
  and _80493_ (_30677_, _15602_, _08624_);
  or _80494_ (_30678_, _30677_, _30650_);
  and _80495_ (_30679_, _30678_, _06257_);
  or _80496_ (_30680_, _30679_, _10080_);
  or _80497_ (_30681_, _30680_, _30676_);
  or _80498_ (_30682_, _30658_, _07215_);
  and _80499_ (_30683_, _30682_, _30681_);
  or _80500_ (_30684_, _30683_, _07460_);
  and _80501_ (_30686_, _09446_, _07904_);
  or _80502_ (_30687_, _30637_, _07208_);
  or _80503_ (_30688_, _30687_, _30686_);
  and _80504_ (_30689_, _30688_, _05982_);
  and _80505_ (_30690_, _30689_, _30684_);
  and _80506_ (_30691_, _15657_, _07904_);
  or _80507_ (_30692_, _30691_, _30637_);
  and _80508_ (_30693_, _30692_, _10094_);
  or _80509_ (_30694_, _30693_, _06218_);
  or _80510_ (_30695_, _30694_, _30690_);
  and _80511_ (_30697_, _15664_, _07904_);
  or _80512_ (_30698_, _30697_, _30637_);
  or _80513_ (_30699_, _30698_, _06219_);
  and _80514_ (_30700_, _30699_, _30695_);
  or _80515_ (_30701_, _30700_, _06369_);
  and _80516_ (_30702_, _15549_, _07904_);
  or _80517_ (_30703_, _30702_, _30637_);
  or _80518_ (_30704_, _30703_, _07237_);
  and _80519_ (_30705_, _30704_, _07240_);
  and _80520_ (_30706_, _30705_, _30701_);
  and _80521_ (_30708_, _11247_, _07904_);
  or _80522_ (_30709_, _30708_, _30637_);
  and _80523_ (_30710_, _30709_, _06536_);
  or _80524_ (_30711_, _30710_, _30706_);
  and _80525_ (_30712_, _30711_, _07242_);
  or _80526_ (_30713_, _30637_, _08145_);
  and _80527_ (_30714_, _30698_, _06375_);
  and _80528_ (_30715_, _30714_, _30713_);
  or _80529_ (_30716_, _30715_, _30712_);
  and _80530_ (_30717_, _30716_, _07234_);
  and _80531_ (_30719_, _30643_, _06545_);
  and _80532_ (_30720_, _30719_, _30713_);
  or _80533_ (_30721_, _30720_, _06366_);
  or _80534_ (_30722_, _30721_, _30717_);
  and _80535_ (_30723_, _15546_, _07904_);
  or _80536_ (_30724_, _30637_, _09056_);
  or _80537_ (_30725_, _30724_, _30723_);
  and _80538_ (_30726_, _30725_, _09061_);
  and _80539_ (_30727_, _30726_, _30722_);
  nor _80540_ (_30728_, _11246_, _13077_);
  or _80541_ (_30730_, _30728_, _30637_);
  and _80542_ (_30731_, _30730_, _06528_);
  or _80543_ (_30732_, _30731_, _06568_);
  or _80544_ (_30733_, _30732_, _30727_);
  or _80545_ (_30734_, _30639_, _06926_);
  and _80546_ (_30735_, _30734_, _05928_);
  and _80547_ (_30736_, _30735_, _30733_);
  and _80548_ (_30737_, _30667_, _05927_);
  or _80549_ (_30738_, _30737_, _06278_);
  or _80550_ (_30739_, _30738_, _30736_);
  and _80551_ (_30741_, _15734_, _07904_);
  or _80552_ (_30742_, _30637_, _06279_);
  or _80553_ (_30743_, _30742_, _30741_);
  and _80554_ (_30744_, _30743_, _01347_);
  and _80555_ (_30745_, _30744_, _30739_);
  or _80556_ (_43269_, _30745_, _30636_);
  and _80557_ (_30746_, _07894_, \oc8051_golden_model_1.ACC [0]);
  and _80558_ (_30747_, _30746_, _08390_);
  and _80559_ (_30748_, _13180_, \oc8051_golden_model_1.P3 [0]);
  or _80560_ (_30749_, _30748_, _07234_);
  or _80561_ (_30751_, _30749_, _30747_);
  and _80562_ (_30752_, _07894_, _07133_);
  or _80563_ (_30753_, _30752_, _30748_);
  or _80564_ (_30754_, _30753_, _07215_);
  nor _80565_ (_30755_, _08390_, _13180_);
  or _80566_ (_30756_, _30755_, _30748_);
  and _80567_ (_30757_, _30756_, _06341_);
  and _80568_ (_30758_, _07142_, \oc8051_golden_model_1.P3 [0]);
  or _80569_ (_30759_, _30746_, _30748_);
  and _80570_ (_30760_, _30759_, _07141_);
  or _80571_ (_30762_, _30760_, _30758_);
  and _80572_ (_30763_, _30762_, _07151_);
  or _80573_ (_30764_, _30763_, _06272_);
  or _80574_ (_30765_, _30764_, _30757_);
  and _80575_ (_30766_, _14382_, _08628_);
  and _80576_ (_30767_, _13188_, \oc8051_golden_model_1.P3 [0]);
  or _80577_ (_30768_, _30767_, _06273_);
  or _80578_ (_30769_, _30768_, _30766_);
  and _80579_ (_30770_, _30769_, _07166_);
  and _80580_ (_30771_, _30770_, _30765_);
  and _80581_ (_30773_, _30753_, _06461_);
  or _80582_ (_30774_, _30773_, _06464_);
  or _80583_ (_30775_, _30774_, _30771_);
  or _80584_ (_30776_, _30759_, _06465_);
  and _80585_ (_30777_, _30776_, _06269_);
  and _80586_ (_30778_, _30777_, _30775_);
  and _80587_ (_30779_, _30748_, _06268_);
  or _80588_ (_30780_, _30779_, _06261_);
  or _80589_ (_30781_, _30780_, _30778_);
  or _80590_ (_30782_, _30756_, _06262_);
  and _80591_ (_30784_, _30782_, _06258_);
  and _80592_ (_30785_, _30784_, _30781_);
  and _80593_ (_30786_, _14413_, _08628_);
  or _80594_ (_30787_, _30786_, _30767_);
  and _80595_ (_30788_, _30787_, _06257_);
  or _80596_ (_30789_, _30788_, _10080_);
  or _80597_ (_30790_, _30789_, _30785_);
  and _80598_ (_30791_, _30790_, _30754_);
  or _80599_ (_30792_, _30791_, _07460_);
  and _80600_ (_30793_, _09392_, _07894_);
  or _80601_ (_30795_, _30748_, _07208_);
  or _80602_ (_30796_, _30795_, _30793_);
  and _80603_ (_30797_, _30796_, _30792_);
  or _80604_ (_30798_, _30797_, _10094_);
  and _80605_ (_30799_, _14467_, _07894_);
  or _80606_ (_30800_, _30748_, _05982_);
  or _80607_ (_30801_, _30800_, _30799_);
  and _80608_ (_30802_, _30801_, _06219_);
  and _80609_ (_30803_, _30802_, _30798_);
  and _80610_ (_30804_, _07894_, _08954_);
  or _80611_ (_30806_, _30804_, _30748_);
  and _80612_ (_30807_, _30806_, _06218_);
  or _80613_ (_30808_, _30807_, _06369_);
  or _80614_ (_30809_, _30808_, _30803_);
  and _80615_ (_30810_, _14366_, _07894_);
  or _80616_ (_30811_, _30810_, _30748_);
  or _80617_ (_30812_, _30811_, _07237_);
  and _80618_ (_30813_, _30812_, _07240_);
  and _80619_ (_30814_, _30813_, _30809_);
  nor _80620_ (_30815_, _12580_, _13180_);
  or _80621_ (_30817_, _30815_, _30748_);
  nor _80622_ (_30818_, _30747_, _07240_);
  and _80623_ (_30819_, _30818_, _30817_);
  or _80624_ (_30820_, _30819_, _30814_);
  and _80625_ (_30821_, _30820_, _07242_);
  nand _80626_ (_30822_, _30806_, _06375_);
  nor _80627_ (_30823_, _30822_, _30755_);
  or _80628_ (_30824_, _30823_, _06545_);
  or _80629_ (_30825_, _30824_, _30821_);
  and _80630_ (_30826_, _30825_, _30751_);
  or _80631_ (_30828_, _30826_, _06366_);
  and _80632_ (_30829_, _14363_, _07894_);
  or _80633_ (_30830_, _30748_, _09056_);
  or _80634_ (_30831_, _30830_, _30829_);
  and _80635_ (_30832_, _30831_, _09061_);
  and _80636_ (_30833_, _30832_, _30828_);
  and _80637_ (_30834_, _30817_, _06528_);
  or _80638_ (_30835_, _30834_, _06568_);
  or _80639_ (_30836_, _30835_, _30833_);
  or _80640_ (_30837_, _30756_, _06926_);
  and _80641_ (_30839_, _30837_, _30836_);
  or _80642_ (_30840_, _30839_, _05927_);
  or _80643_ (_30841_, _30748_, _05928_);
  and _80644_ (_30842_, _30841_, _30840_);
  or _80645_ (_30843_, _30842_, _06278_);
  or _80646_ (_30844_, _30756_, _06279_);
  and _80647_ (_30845_, _30844_, _01347_);
  and _80648_ (_30846_, _30845_, _30843_);
  nor _80649_ (_30847_, \oc8051_golden_model_1.P3 [0], rst);
  nor _80650_ (_30848_, _30847_, _01354_);
  or _80651_ (_43271_, _30848_, _30846_);
  and _80652_ (_30850_, _13180_, \oc8051_golden_model_1.P3 [1]);
  nor _80653_ (_30851_, _11261_, _13180_);
  or _80654_ (_30852_, _30851_, _30850_);
  or _80655_ (_30853_, _30852_, _09061_);
  nand _80656_ (_30854_, _07894_, _07038_);
  or _80657_ (_30855_, _07894_, \oc8051_golden_model_1.P3 [1]);
  and _80658_ (_30856_, _30855_, _06218_);
  and _80659_ (_30857_, _30856_, _30854_);
  nor _80660_ (_30858_, _13180_, _07357_);
  or _80661_ (_30860_, _30858_, _30850_);
  or _80662_ (_30861_, _30860_, _07166_);
  and _80663_ (_30862_, _14562_, _07894_);
  not _80664_ (_30863_, _30862_);
  and _80665_ (_30864_, _30863_, _30855_);
  or _80666_ (_30865_, _30864_, _07151_);
  and _80667_ (_30866_, _07894_, \oc8051_golden_model_1.ACC [1]);
  or _80668_ (_30867_, _30866_, _30850_);
  and _80669_ (_30868_, _30867_, _07141_);
  and _80670_ (_30869_, _07142_, \oc8051_golden_model_1.P3 [1]);
  or _80671_ (_30871_, _30869_, _06341_);
  or _80672_ (_30872_, _30871_, _30868_);
  and _80673_ (_30873_, _30872_, _06273_);
  and _80674_ (_30874_, _30873_, _30865_);
  and _80675_ (_30875_, _13188_, \oc8051_golden_model_1.P3 [1]);
  and _80676_ (_30876_, _14557_, _08628_);
  or _80677_ (_30877_, _30876_, _30875_);
  and _80678_ (_30878_, _30877_, _06272_);
  or _80679_ (_30879_, _30878_, _06461_);
  or _80680_ (_30880_, _30879_, _30874_);
  and _80681_ (_30882_, _30880_, _30861_);
  or _80682_ (_30883_, _30882_, _06464_);
  or _80683_ (_30884_, _30867_, _06465_);
  and _80684_ (_30885_, _30884_, _06269_);
  and _80685_ (_30886_, _30885_, _30883_);
  and _80686_ (_30887_, _14560_, _08628_);
  or _80687_ (_30888_, _30887_, _30875_);
  and _80688_ (_30889_, _30888_, _06268_);
  or _80689_ (_30890_, _30889_, _06261_);
  or _80690_ (_30891_, _30890_, _30886_);
  and _80691_ (_30893_, _30876_, _14556_);
  or _80692_ (_30894_, _30875_, _06262_);
  or _80693_ (_30895_, _30894_, _30893_);
  and _80694_ (_30896_, _30895_, _06258_);
  and _80695_ (_30897_, _30896_, _30891_);
  or _80696_ (_30898_, _30875_, _14597_);
  and _80697_ (_30899_, _30898_, _06257_);
  and _80698_ (_30900_, _30899_, _30877_);
  or _80699_ (_30901_, _30900_, _10080_);
  or _80700_ (_30902_, _30901_, _30897_);
  or _80701_ (_30904_, _30860_, _07215_);
  and _80702_ (_30905_, _30904_, _30902_);
  or _80703_ (_30906_, _30905_, _07460_);
  and _80704_ (_30907_, _09451_, _07894_);
  or _80705_ (_30908_, _30850_, _07208_);
  or _80706_ (_30909_, _30908_, _30907_);
  and _80707_ (_30910_, _30909_, _05982_);
  and _80708_ (_30911_, _30910_, _30906_);
  and _80709_ (_30912_, _14653_, _07894_);
  or _80710_ (_30913_, _30912_, _30850_);
  and _80711_ (_30915_, _30913_, _10094_);
  or _80712_ (_30916_, _30915_, _30911_);
  and _80713_ (_30917_, _30916_, _06219_);
  or _80714_ (_30918_, _30917_, _30857_);
  and _80715_ (_30919_, _30918_, _07237_);
  or _80716_ (_30920_, _14668_, _13180_);
  and _80717_ (_30921_, _30855_, _06369_);
  and _80718_ (_30922_, _30921_, _30920_);
  or _80719_ (_30923_, _30922_, _06536_);
  or _80720_ (_30924_, _30923_, _30919_);
  and _80721_ (_30926_, _11262_, _07894_);
  or _80722_ (_30927_, _30926_, _30850_);
  or _80723_ (_30928_, _30927_, _07240_);
  and _80724_ (_30929_, _30928_, _07242_);
  and _80725_ (_30930_, _30929_, _30924_);
  or _80726_ (_30931_, _14666_, _13180_);
  and _80727_ (_30932_, _30855_, _06375_);
  and _80728_ (_30933_, _30932_, _30931_);
  or _80729_ (_30934_, _30933_, _06545_);
  or _80730_ (_30935_, _30934_, _30930_);
  and _80731_ (_30937_, _30866_, _08341_);
  or _80732_ (_30938_, _30850_, _07234_);
  or _80733_ (_30939_, _30938_, _30937_);
  and _80734_ (_30940_, _30939_, _09056_);
  and _80735_ (_30941_, _30940_, _30935_);
  or _80736_ (_30942_, _30854_, _08341_);
  and _80737_ (_30943_, _30855_, _06366_);
  and _80738_ (_30944_, _30943_, _30942_);
  or _80739_ (_30945_, _30944_, _06528_);
  or _80740_ (_30946_, _30945_, _30941_);
  and _80741_ (_30948_, _30946_, _30853_);
  or _80742_ (_30949_, _30948_, _06568_);
  or _80743_ (_30950_, _30864_, _06926_);
  and _80744_ (_30951_, _30950_, _05928_);
  and _80745_ (_30952_, _30951_, _30949_);
  and _80746_ (_30953_, _30888_, _05927_);
  or _80747_ (_30954_, _30953_, _06278_);
  or _80748_ (_30955_, _30954_, _30952_);
  or _80749_ (_30956_, _30850_, _06279_);
  or _80750_ (_30957_, _30956_, _30862_);
  and _80751_ (_30959_, _30957_, _01347_);
  and _80752_ (_30960_, _30959_, _30955_);
  nor _80753_ (_30961_, \oc8051_golden_model_1.P3 [1], rst);
  nor _80754_ (_30962_, _30961_, _01354_);
  or _80755_ (_43272_, _30962_, _30960_);
  and _80756_ (_30963_, _13180_, \oc8051_golden_model_1.P3 [2]);
  nor _80757_ (_30964_, _13180_, _07776_);
  or _80758_ (_30965_, _30964_, _30963_);
  or _80759_ (_30966_, _30965_, _07215_);
  or _80760_ (_30967_, _30965_, _07166_);
  and _80761_ (_30969_, _14770_, _07894_);
  or _80762_ (_30970_, _30969_, _30963_);
  or _80763_ (_30971_, _30970_, _07151_);
  and _80764_ (_30972_, _07894_, \oc8051_golden_model_1.ACC [2]);
  or _80765_ (_30973_, _30972_, _30963_);
  and _80766_ (_30974_, _30973_, _07141_);
  and _80767_ (_30975_, _07142_, \oc8051_golden_model_1.P3 [2]);
  or _80768_ (_30976_, _30975_, _06341_);
  or _80769_ (_30977_, _30976_, _30974_);
  and _80770_ (_30978_, _30977_, _06273_);
  and _80771_ (_30980_, _30978_, _30971_);
  and _80772_ (_30981_, _13188_, \oc8051_golden_model_1.P3 [2]);
  and _80773_ (_30982_, _14774_, _08628_);
  or _80774_ (_30983_, _30982_, _30981_);
  and _80775_ (_30984_, _30983_, _06272_);
  or _80776_ (_30985_, _30984_, _06461_);
  or _80777_ (_30986_, _30985_, _30980_);
  and _80778_ (_30987_, _30986_, _30967_);
  or _80779_ (_30988_, _30987_, _06464_);
  or _80780_ (_30989_, _30973_, _06465_);
  and _80781_ (_30991_, _30989_, _06269_);
  and _80782_ (_30992_, _30991_, _30988_);
  and _80783_ (_30993_, _14756_, _08628_);
  or _80784_ (_30994_, _30993_, _30981_);
  and _80785_ (_30995_, _30994_, _06268_);
  or _80786_ (_30996_, _30995_, _06261_);
  or _80787_ (_30997_, _30996_, _30992_);
  and _80788_ (_30998_, _30982_, _14789_);
  or _80789_ (_30999_, _30981_, _06262_);
  or _80790_ (_31000_, _30999_, _30998_);
  and _80791_ (_31002_, _31000_, _06258_);
  and _80792_ (_31003_, _31002_, _30997_);
  and _80793_ (_31004_, _14804_, _08628_);
  or _80794_ (_31005_, _31004_, _30981_);
  and _80795_ (_31006_, _31005_, _06257_);
  or _80796_ (_31007_, _31006_, _10080_);
  or _80797_ (_31008_, _31007_, _31003_);
  and _80798_ (_31009_, _31008_, _30966_);
  or _80799_ (_31010_, _31009_, _07460_);
  and _80800_ (_31011_, _09450_, _07894_);
  or _80801_ (_31013_, _30963_, _07208_);
  or _80802_ (_31014_, _31013_, _31011_);
  and _80803_ (_31015_, _31014_, _05982_);
  and _80804_ (_31016_, _31015_, _31010_);
  and _80805_ (_31017_, _14859_, _07894_);
  or _80806_ (_31018_, _31017_, _30963_);
  and _80807_ (_31019_, _31018_, _10094_);
  or _80808_ (_31020_, _31019_, _06218_);
  or _80809_ (_31021_, _31020_, _31016_);
  and _80810_ (_31022_, _07894_, _08973_);
  or _80811_ (_31024_, _31022_, _30963_);
  or _80812_ (_31025_, _31024_, _06219_);
  and _80813_ (_31026_, _31025_, _31021_);
  or _80814_ (_31027_, _31026_, _06369_);
  and _80815_ (_31028_, _14751_, _07894_);
  or _80816_ (_31029_, _31028_, _30963_);
  or _80817_ (_31030_, _31029_, _07237_);
  and _80818_ (_31031_, _31030_, _07240_);
  and _80819_ (_31032_, _31031_, _31027_);
  and _80820_ (_31033_, _11259_, _07894_);
  or _80821_ (_31035_, _31033_, _30963_);
  and _80822_ (_31036_, _31035_, _06536_);
  or _80823_ (_31037_, _31036_, _31032_);
  and _80824_ (_31038_, _31037_, _07242_);
  or _80825_ (_31039_, _30963_, _08440_);
  and _80826_ (_31040_, _31024_, _06375_);
  and _80827_ (_31041_, _31040_, _31039_);
  or _80828_ (_31042_, _31041_, _31038_);
  and _80829_ (_31043_, _31042_, _07234_);
  and _80830_ (_31044_, _30973_, _06545_);
  and _80831_ (_31047_, _31044_, _31039_);
  or _80832_ (_31048_, _31047_, _06366_);
  or _80833_ (_31049_, _31048_, _31043_);
  and _80834_ (_31050_, _14748_, _07894_);
  or _80835_ (_31051_, _30963_, _09056_);
  or _80836_ (_31052_, _31051_, _31050_);
  and _80837_ (_31053_, _31052_, _09061_);
  and _80838_ (_31054_, _31053_, _31049_);
  nor _80839_ (_31055_, _11258_, _13180_);
  or _80840_ (_31056_, _31055_, _30963_);
  and _80841_ (_31058_, _31056_, _06528_);
  or _80842_ (_31059_, _31058_, _06568_);
  or _80843_ (_31060_, _31059_, _31054_);
  or _80844_ (_31061_, _30970_, _06926_);
  and _80845_ (_31062_, _31061_, _05928_);
  and _80846_ (_31063_, _31062_, _31060_);
  and _80847_ (_31064_, _30994_, _05927_);
  or _80848_ (_31065_, _31064_, _06278_);
  or _80849_ (_31066_, _31065_, _31063_);
  and _80850_ (_31067_, _14926_, _07894_);
  or _80851_ (_31070_, _30963_, _06279_);
  or _80852_ (_31071_, _31070_, _31067_);
  and _80853_ (_31072_, _31071_, _01347_);
  and _80854_ (_31073_, _31072_, _31066_);
  nor _80855_ (_31074_, \oc8051_golden_model_1.P3 [2], rst);
  nor _80856_ (_31075_, _31074_, _01354_);
  or _80857_ (_43273_, _31075_, _31073_);
  nor _80858_ (_31076_, \oc8051_golden_model_1.P3 [3], rst);
  nor _80859_ (_31077_, _31076_, _01354_);
  and _80860_ (_31078_, _13180_, \oc8051_golden_model_1.P3 [3]);
  nor _80861_ (_31080_, _13180_, _07594_);
  or _80862_ (_31081_, _31080_, _31078_);
  or _80863_ (_31082_, _31081_, _07215_);
  and _80864_ (_31083_, _14953_, _07894_);
  or _80865_ (_31084_, _31083_, _31078_);
  or _80866_ (_31085_, _31084_, _07151_);
  and _80867_ (_31086_, _07894_, \oc8051_golden_model_1.ACC [3]);
  or _80868_ (_31087_, _31086_, _31078_);
  and _80869_ (_31088_, _31087_, _07141_);
  and _80870_ (_31089_, _07142_, \oc8051_golden_model_1.P3 [3]);
  or _80871_ (_31092_, _31089_, _06341_);
  or _80872_ (_31093_, _31092_, _31088_);
  and _80873_ (_31094_, _31093_, _06273_);
  and _80874_ (_31095_, _31094_, _31085_);
  and _80875_ (_31096_, _13188_, \oc8051_golden_model_1.P3 [3]);
  and _80876_ (_31097_, _14950_, _08628_);
  or _80877_ (_31098_, _31097_, _31096_);
  and _80878_ (_31099_, _31098_, _06272_);
  or _80879_ (_31100_, _31099_, _06461_);
  or _80880_ (_31101_, _31100_, _31095_);
  or _80881_ (_31103_, _31081_, _07166_);
  and _80882_ (_31104_, _31103_, _31101_);
  or _80883_ (_31105_, _31104_, _06464_);
  or _80884_ (_31106_, _31087_, _06465_);
  and _80885_ (_31107_, _31106_, _06269_);
  and _80886_ (_31108_, _31107_, _31105_);
  and _80887_ (_31109_, _14948_, _08628_);
  or _80888_ (_31110_, _31109_, _31096_);
  and _80889_ (_31111_, _31110_, _06268_);
  or _80890_ (_31112_, _31111_, _06261_);
  or _80891_ (_31115_, _31112_, _31108_);
  or _80892_ (_31116_, _31096_, _14979_);
  and _80893_ (_31117_, _31116_, _31098_);
  or _80894_ (_31118_, _31117_, _06262_);
  and _80895_ (_31119_, _31118_, _06258_);
  and _80896_ (_31120_, _31119_, _31115_);
  or _80897_ (_31121_, _31096_, _14992_);
  and _80898_ (_31122_, _31121_, _06257_);
  and _80899_ (_31123_, _31122_, _31098_);
  or _80900_ (_31124_, _31123_, _10080_);
  or _80901_ (_31126_, _31124_, _31120_);
  and _80902_ (_31127_, _31126_, _31082_);
  or _80903_ (_31128_, _31127_, _07460_);
  and _80904_ (_31129_, _09449_, _07894_);
  or _80905_ (_31130_, _31078_, _07208_);
  or _80906_ (_31131_, _31130_, _31129_);
  and _80907_ (_31132_, _31131_, _05982_);
  and _80908_ (_31133_, _31132_, _31128_);
  and _80909_ (_31134_, _15048_, _07894_);
  or _80910_ (_31135_, _31134_, _31078_);
  and _80911_ (_31137_, _31135_, _10094_);
  or _80912_ (_31138_, _31137_, _06218_);
  or _80913_ (_31139_, _31138_, _31133_);
  and _80914_ (_31140_, _07894_, _08930_);
  or _80915_ (_31141_, _31140_, _31078_);
  or _80916_ (_31142_, _31141_, _06219_);
  and _80917_ (_31143_, _31142_, _31139_);
  or _80918_ (_31144_, _31143_, _06369_);
  and _80919_ (_31145_, _14943_, _07894_);
  or _80920_ (_31146_, _31145_, _31078_);
  or _80921_ (_31148_, _31146_, _07237_);
  and _80922_ (_31149_, _31148_, _07240_);
  and _80923_ (_31150_, _31149_, _31144_);
  and _80924_ (_31151_, _12577_, _07894_);
  or _80925_ (_31152_, _31151_, _31078_);
  and _80926_ (_31153_, _31152_, _06536_);
  or _80927_ (_31154_, _31153_, _31150_);
  and _80928_ (_31155_, _31154_, _07242_);
  or _80929_ (_31156_, _31078_, _08292_);
  and _80930_ (_31157_, _31141_, _06375_);
  and _80931_ (_31158_, _31157_, _31156_);
  or _80932_ (_31159_, _31158_, _31155_);
  and _80933_ (_31160_, _31159_, _07234_);
  and _80934_ (_31161_, _31087_, _06545_);
  and _80935_ (_31162_, _31161_, _31156_);
  or _80936_ (_31163_, _31162_, _06366_);
  or _80937_ (_31164_, _31163_, _31160_);
  and _80938_ (_31165_, _14940_, _07894_);
  or _80939_ (_31166_, _31078_, _09056_);
  or _80940_ (_31167_, _31166_, _31165_);
  and _80941_ (_31170_, _31167_, _09061_);
  and _80942_ (_31171_, _31170_, _31164_);
  nor _80943_ (_31172_, _11256_, _13180_);
  or _80944_ (_31173_, _31172_, _31078_);
  and _80945_ (_31174_, _31173_, _06528_);
  or _80946_ (_31175_, _31174_, _06568_);
  or _80947_ (_31176_, _31175_, _31171_);
  or _80948_ (_31177_, _31084_, _06926_);
  and _80949_ (_31178_, _31177_, _05928_);
  and _80950_ (_31179_, _31178_, _31176_);
  and _80951_ (_31180_, _31110_, _05927_);
  or _80952_ (_31181_, _31180_, _06278_);
  or _80953_ (_31182_, _31181_, _31179_);
  and _80954_ (_31183_, _15128_, _07894_);
  or _80955_ (_31184_, _31078_, _06279_);
  or _80956_ (_31185_, _31184_, _31183_);
  and _80957_ (_31186_, _31185_, _01347_);
  and _80958_ (_31187_, _31186_, _31182_);
  or _80959_ (_43274_, _31187_, _31077_);
  and _80960_ (_31188_, _13180_, \oc8051_golden_model_1.P3 [4]);
  nor _80961_ (_31191_, _08541_, _13180_);
  or _80962_ (_31192_, _31191_, _31188_);
  or _80963_ (_31193_, _31192_, _07215_);
  and _80964_ (_31194_, _13188_, \oc8051_golden_model_1.P3 [4]);
  and _80965_ (_31195_, _15176_, _08628_);
  or _80966_ (_31196_, _31195_, _31194_);
  and _80967_ (_31197_, _31196_, _06268_);
  and _80968_ (_31198_, _15162_, _07894_);
  or _80969_ (_31199_, _31198_, _31188_);
  or _80970_ (_31200_, _31199_, _07151_);
  and _80971_ (_31201_, _07894_, \oc8051_golden_model_1.ACC [4]);
  or _80972_ (_31202_, _31201_, _31188_);
  and _80973_ (_31203_, _31202_, _07141_);
  and _80974_ (_31204_, _07142_, \oc8051_golden_model_1.P3 [4]);
  or _80975_ (_31205_, _31204_, _06341_);
  or _80976_ (_31206_, _31205_, _31203_);
  and _80977_ (_31207_, _31206_, _06273_);
  and _80978_ (_31208_, _31207_, _31200_);
  and _80979_ (_31209_, _15166_, _08628_);
  or _80980_ (_31210_, _31209_, _31194_);
  and _80981_ (_31213_, _31210_, _06272_);
  or _80982_ (_31214_, _31213_, _06461_);
  or _80983_ (_31215_, _31214_, _31208_);
  or _80984_ (_31216_, _31192_, _07166_);
  and _80985_ (_31217_, _31216_, _31215_);
  or _80986_ (_31218_, _31217_, _06464_);
  or _80987_ (_31219_, _31202_, _06465_);
  and _80988_ (_31220_, _31219_, _06269_);
  and _80989_ (_31221_, _31220_, _31218_);
  or _80990_ (_31222_, _31221_, _31197_);
  and _80991_ (_31223_, _31222_, _06262_);
  and _80992_ (_31224_, _15184_, _08628_);
  or _80993_ (_31225_, _31224_, _31194_);
  and _80994_ (_31226_, _31225_, _06261_);
  or _80995_ (_31227_, _31226_, _31223_);
  and _80996_ (_31228_, _31227_, _06258_);
  and _80997_ (_31229_, _15200_, _08628_);
  or _80998_ (_31230_, _31229_, _31194_);
  and _80999_ (_31231_, _31230_, _06257_);
  or _81000_ (_31232_, _31231_, _10080_);
  or _81001_ (_31235_, _31232_, _31228_);
  and _81002_ (_31236_, _31235_, _31193_);
  or _81003_ (_31237_, _31236_, _07460_);
  and _81004_ (_31238_, _09448_, _07894_);
  or _81005_ (_31239_, _31188_, _07208_);
  or _81006_ (_31240_, _31239_, _31238_);
  and _81007_ (_31241_, _31240_, _05982_);
  and _81008_ (_31242_, _31241_, _31237_);
  and _81009_ (_31243_, _15254_, _07894_);
  or _81010_ (_31244_, _31243_, _31188_);
  and _81011_ (_31245_, _31244_, _10094_);
  or _81012_ (_31246_, _31245_, _06218_);
  or _81013_ (_31247_, _31246_, _31242_);
  and _81014_ (_31248_, _08959_, _07894_);
  or _81015_ (_31249_, _31248_, _31188_);
  or _81016_ (_31250_, _31249_, _06219_);
  and _81017_ (_31251_, _31250_, _31247_);
  or _81018_ (_31252_, _31251_, _06369_);
  and _81019_ (_31253_, _15269_, _07894_);
  or _81020_ (_31254_, _31253_, _31188_);
  or _81021_ (_31257_, _31254_, _07237_);
  and _81022_ (_31258_, _31257_, _07240_);
  and _81023_ (_31259_, _31258_, _31252_);
  and _81024_ (_31260_, _11254_, _07894_);
  or _81025_ (_31261_, _31260_, _31188_);
  and _81026_ (_31262_, _31261_, _06536_);
  or _81027_ (_31263_, _31262_, _31259_);
  and _81028_ (_31264_, _31263_, _07242_);
  or _81029_ (_31265_, _31188_, _08544_);
  and _81030_ (_31266_, _31249_, _06375_);
  and _81031_ (_31267_, _31266_, _31265_);
  or _81032_ (_31268_, _31267_, _31264_);
  and _81033_ (_31269_, _31268_, _07234_);
  and _81034_ (_31270_, _31202_, _06545_);
  and _81035_ (_31271_, _31270_, _31265_);
  or _81036_ (_31272_, _31271_, _06366_);
  or _81037_ (_31273_, _31272_, _31269_);
  and _81038_ (_31274_, _15266_, _07894_);
  or _81039_ (_31275_, _31188_, _09056_);
  or _81040_ (_31276_, _31275_, _31274_);
  and _81041_ (_31279_, _31276_, _09061_);
  and _81042_ (_31280_, _31279_, _31273_);
  nor _81043_ (_31281_, _11253_, _13180_);
  or _81044_ (_31282_, _31281_, _31188_);
  and _81045_ (_31283_, _31282_, _06528_);
  or _81046_ (_31284_, _31283_, _06568_);
  or _81047_ (_31285_, _31284_, _31280_);
  or _81048_ (_31286_, _31199_, _06926_);
  and _81049_ (_31287_, _31286_, _05928_);
  and _81050_ (_31288_, _31287_, _31285_);
  and _81051_ (_31289_, _31196_, _05927_);
  or _81052_ (_31290_, _31289_, _06278_);
  or _81053_ (_31291_, _31290_, _31288_);
  and _81054_ (_31292_, _15329_, _07894_);
  or _81055_ (_31293_, _31188_, _06279_);
  or _81056_ (_31294_, _31293_, _31292_);
  and _81057_ (_31295_, _31294_, _01347_);
  and _81058_ (_31296_, _31295_, _31291_);
  nor _81059_ (_31297_, \oc8051_golden_model_1.P3 [4], rst);
  nor _81060_ (_31298_, _31297_, _01354_);
  or _81061_ (_43275_, _31298_, _31296_);
  nor _81062_ (_31301_, \oc8051_golden_model_1.P3 [5], rst);
  nor _81063_ (_31302_, _31301_, _01354_);
  and _81064_ (_31303_, _13180_, \oc8051_golden_model_1.P3 [5]);
  and _81065_ (_31304_, _15358_, _07894_);
  or _81066_ (_31305_, _31304_, _31303_);
  or _81067_ (_31306_, _31305_, _07151_);
  and _81068_ (_31307_, _07894_, \oc8051_golden_model_1.ACC [5]);
  or _81069_ (_31308_, _31307_, _31303_);
  and _81070_ (_31309_, _31308_, _07141_);
  and _81071_ (_31310_, _07142_, \oc8051_golden_model_1.P3 [5]);
  or _81072_ (_31311_, _31310_, _06341_);
  or _81073_ (_31312_, _31311_, _31309_);
  and _81074_ (_31313_, _31312_, _06273_);
  and _81075_ (_31314_, _31313_, _31306_);
  and _81076_ (_31315_, _13188_, \oc8051_golden_model_1.P3 [5]);
  and _81077_ (_31316_, _15372_, _08628_);
  or _81078_ (_31317_, _31316_, _31315_);
  and _81079_ (_31318_, _31317_, _06272_);
  or _81080_ (_31319_, _31318_, _06461_);
  or _81081_ (_31322_, _31319_, _31314_);
  nor _81082_ (_31323_, _08244_, _13180_);
  or _81083_ (_31324_, _31323_, _31303_);
  or _81084_ (_31325_, _31324_, _07166_);
  and _81085_ (_31326_, _31325_, _31322_);
  or _81086_ (_31327_, _31326_, _06464_);
  or _81087_ (_31328_, _31308_, _06465_);
  and _81088_ (_31329_, _31328_, _06269_);
  and _81089_ (_31330_, _31329_, _31327_);
  and _81090_ (_31331_, _15355_, _08628_);
  or _81091_ (_31332_, _31331_, _31315_);
  and _81092_ (_31333_, _31332_, _06268_);
  or _81093_ (_31334_, _31333_, _06261_);
  or _81094_ (_31335_, _31334_, _31330_);
  or _81095_ (_31336_, _31315_, _15387_);
  and _81096_ (_31337_, _31336_, _31317_);
  or _81097_ (_31338_, _31337_, _06262_);
  and _81098_ (_31339_, _31338_, _06258_);
  and _81099_ (_31340_, _31339_, _31335_);
  or _81100_ (_31341_, _31315_, _15403_);
  and _81101_ (_31344_, _31341_, _06257_);
  and _81102_ (_31345_, _31344_, _31317_);
  or _81103_ (_31346_, _31345_, _10080_);
  or _81104_ (_31347_, _31346_, _31340_);
  or _81105_ (_31348_, _31324_, _07215_);
  and _81106_ (_31349_, _31348_, _31347_);
  or _81107_ (_31350_, _31349_, _07460_);
  and _81108_ (_31351_, _09447_, _07894_);
  or _81109_ (_31352_, _31303_, _07208_);
  or _81110_ (_31353_, _31352_, _31351_);
  and _81111_ (_31354_, _31353_, _05982_);
  and _81112_ (_31355_, _31354_, _31350_);
  and _81113_ (_31356_, _15459_, _07894_);
  or _81114_ (_31357_, _31356_, _31303_);
  and _81115_ (_31358_, _31357_, _10094_);
  or _81116_ (_31359_, _31358_, _06218_);
  or _81117_ (_31360_, _31359_, _31355_);
  and _81118_ (_31361_, _08946_, _07894_);
  or _81119_ (_31362_, _31361_, _31303_);
  or _81120_ (_31363_, _31362_, _06219_);
  and _81121_ (_31366_, _31363_, _31360_);
  or _81122_ (_31367_, _31366_, _06369_);
  and _81123_ (_31368_, _15353_, _07894_);
  or _81124_ (_31369_, _31368_, _31303_);
  or _81125_ (_31370_, _31369_, _07237_);
  and _81126_ (_31371_, _31370_, _07240_);
  and _81127_ (_31372_, _31371_, _31367_);
  and _81128_ (_31373_, _11250_, _07894_);
  or _81129_ (_31374_, _31373_, _31303_);
  and _81130_ (_31375_, _31374_, _06536_);
  or _81131_ (_31376_, _31375_, _31372_);
  and _81132_ (_31377_, _31376_, _07242_);
  or _81133_ (_31378_, _31303_, _08247_);
  and _81134_ (_31379_, _31362_, _06375_);
  and _81135_ (_31380_, _31379_, _31378_);
  or _81136_ (_31381_, _31380_, _31377_);
  and _81137_ (_31382_, _31381_, _07234_);
  and _81138_ (_31383_, _31308_, _06545_);
  and _81139_ (_31384_, _31383_, _31378_);
  or _81140_ (_31385_, _31384_, _06366_);
  or _81141_ (_31388_, _31385_, _31382_);
  and _81142_ (_31389_, _15350_, _07894_);
  or _81143_ (_31390_, _31303_, _09056_);
  or _81144_ (_31391_, _31390_, _31389_);
  and _81145_ (_31392_, _31391_, _09061_);
  and _81146_ (_31393_, _31392_, _31388_);
  nor _81147_ (_31394_, _11249_, _13180_);
  or _81148_ (_31395_, _31394_, _31303_);
  and _81149_ (_31396_, _31395_, _06528_);
  or _81150_ (_31397_, _31396_, _06568_);
  or _81151_ (_31398_, _31397_, _31393_);
  or _81152_ (_31399_, _31305_, _06926_);
  and _81153_ (_31400_, _31399_, _05928_);
  and _81154_ (_31401_, _31400_, _31398_);
  and _81155_ (_31402_, _31332_, _05927_);
  or _81156_ (_31403_, _31402_, _06278_);
  or _81157_ (_31404_, _31403_, _31401_);
  and _81158_ (_31405_, _15532_, _07894_);
  or _81159_ (_31406_, _31303_, _06279_);
  or _81160_ (_31407_, _31406_, _31405_);
  and _81161_ (_31410_, _31407_, _01347_);
  and _81162_ (_31411_, _31410_, _31404_);
  or _81163_ (_43276_, _31411_, _31302_);
  and _81164_ (_31412_, _13180_, \oc8051_golden_model_1.P3 [6]);
  and _81165_ (_31413_, _15554_, _07894_);
  or _81166_ (_31414_, _31413_, _31412_);
  or _81167_ (_31415_, _31414_, _07151_);
  and _81168_ (_31416_, _07894_, \oc8051_golden_model_1.ACC [6]);
  or _81169_ (_31417_, _31416_, _31412_);
  and _81170_ (_31418_, _31417_, _07141_);
  and _81171_ (_31419_, _07142_, \oc8051_golden_model_1.P3 [6]);
  or _81172_ (_31420_, _31419_, _06341_);
  or _81173_ (_31421_, _31420_, _31418_);
  and _81174_ (_31422_, _31421_, _06273_);
  and _81175_ (_31423_, _31422_, _31415_);
  and _81176_ (_31424_, _13188_, \oc8051_golden_model_1.P3 [6]);
  and _81177_ (_31425_, _15570_, _08628_);
  or _81178_ (_31426_, _31425_, _31424_);
  and _81179_ (_31427_, _31426_, _06272_);
  or _81180_ (_31428_, _31427_, _06461_);
  or _81181_ (_31431_, _31428_, _31423_);
  nor _81182_ (_31432_, _08142_, _13180_);
  or _81183_ (_31433_, _31432_, _31412_);
  or _81184_ (_31434_, _31433_, _07166_);
  and _81185_ (_31435_, _31434_, _31431_);
  or _81186_ (_31436_, _31435_, _06464_);
  or _81187_ (_31437_, _31417_, _06465_);
  and _81188_ (_31438_, _31437_, _06269_);
  and _81189_ (_31439_, _31438_, _31436_);
  and _81190_ (_31440_, _15551_, _08628_);
  or _81191_ (_31441_, _31440_, _31424_);
  and _81192_ (_31442_, _31441_, _06268_);
  or _81193_ (_31443_, _31442_, _06261_);
  or _81194_ (_31444_, _31443_, _31439_);
  or _81195_ (_31445_, _31424_, _15585_);
  and _81196_ (_31446_, _31445_, _31426_);
  or _81197_ (_31447_, _31446_, _06262_);
  and _81198_ (_31448_, _31447_, _06258_);
  and _81199_ (_31449_, _31448_, _31444_);
  and _81200_ (_31450_, _15602_, _08628_);
  or _81201_ (_31453_, _31450_, _31424_);
  and _81202_ (_31454_, _31453_, _06257_);
  or _81203_ (_31455_, _31454_, _10080_);
  or _81204_ (_31456_, _31455_, _31449_);
  or _81205_ (_31457_, _31433_, _07215_);
  and _81206_ (_31458_, _31457_, _31456_);
  or _81207_ (_31459_, _31458_, _07460_);
  and _81208_ (_31460_, _09446_, _07894_);
  or _81209_ (_31461_, _31412_, _07208_);
  or _81210_ (_31462_, _31461_, _31460_);
  and _81211_ (_31463_, _31462_, _05982_);
  and _81212_ (_31464_, _31463_, _31459_);
  and _81213_ (_31465_, _15657_, _07894_);
  or _81214_ (_31466_, _31465_, _31412_);
  and _81215_ (_31467_, _31466_, _10094_);
  or _81216_ (_31468_, _31467_, _06218_);
  or _81217_ (_31469_, _31468_, _31464_);
  and _81218_ (_31470_, _15664_, _07894_);
  or _81219_ (_31471_, _31470_, _31412_);
  or _81220_ (_31472_, _31471_, _06219_);
  and _81221_ (_31475_, _31472_, _31469_);
  or _81222_ (_31476_, _31475_, _06369_);
  and _81223_ (_31477_, _15549_, _07894_);
  or _81224_ (_31478_, _31477_, _31412_);
  or _81225_ (_31479_, _31478_, _07237_);
  and _81226_ (_31480_, _31479_, _07240_);
  and _81227_ (_31481_, _31480_, _31476_);
  and _81228_ (_31482_, _11247_, _07894_);
  or _81229_ (_31483_, _31482_, _31412_);
  and _81230_ (_31484_, _31483_, _06536_);
  or _81231_ (_31485_, _31484_, _31481_);
  and _81232_ (_31486_, _31485_, _07242_);
  or _81233_ (_31487_, _31412_, _08145_);
  and _81234_ (_31488_, _31471_, _06375_);
  and _81235_ (_31489_, _31488_, _31487_);
  or _81236_ (_31490_, _31489_, _31486_);
  and _81237_ (_31491_, _31490_, _07234_);
  and _81238_ (_31492_, _31417_, _06545_);
  and _81239_ (_31493_, _31492_, _31487_);
  or _81240_ (_31494_, _31493_, _06366_);
  or _81241_ (_31497_, _31494_, _31491_);
  and _81242_ (_31498_, _15546_, _07894_);
  or _81243_ (_31499_, _31412_, _09056_);
  or _81244_ (_31500_, _31499_, _31498_);
  and _81245_ (_31501_, _31500_, _09061_);
  and _81246_ (_31502_, _31501_, _31497_);
  nor _81247_ (_31503_, _11246_, _13180_);
  or _81248_ (_31504_, _31503_, _31412_);
  and _81249_ (_31505_, _31504_, _06528_);
  or _81250_ (_31506_, _31505_, _06568_);
  or _81251_ (_31507_, _31506_, _31502_);
  or _81252_ (_31508_, _31414_, _06926_);
  and _81253_ (_31509_, _31508_, _05928_);
  and _81254_ (_31510_, _31509_, _31507_);
  and _81255_ (_31511_, _31441_, _05927_);
  or _81256_ (_31512_, _31511_, _06278_);
  or _81257_ (_31513_, _31512_, _31510_);
  and _81258_ (_31514_, _15734_, _07894_);
  or _81259_ (_31515_, _31412_, _06279_);
  or _81260_ (_31516_, _31515_, _31514_);
  and _81261_ (_31519_, _31516_, _01347_);
  and _81262_ (_31520_, _31519_, _31513_);
  nor _81263_ (_31521_, \oc8051_golden_model_1.P3 [6], rst);
  nor _81264_ (_31522_, _31521_, _01354_);
  or _81265_ (_43277_, _31522_, _31520_);
  nand _81266_ (_31523_, _11263_, _07926_);
  not _81267_ (_31524_, \oc8051_golden_model_1.P0 [0]);
  nor _81268_ (_31525_, _07926_, _31524_);
  nor _81269_ (_31526_, _31525_, _07234_);
  nand _81270_ (_31527_, _31526_, _31523_);
  and _81271_ (_31528_, _07926_, _07133_);
  or _81272_ (_31529_, _31528_, _31525_);
  or _81273_ (_31530_, _31529_, _07215_);
  nor _81274_ (_31531_, _08390_, _13283_);
  or _81275_ (_31532_, _31531_, _31525_);
  or _81276_ (_31533_, _31532_, _07151_);
  and _81277_ (_31534_, _07926_, \oc8051_golden_model_1.ACC [0]);
  or _81278_ (_31535_, _31534_, _31525_);
  and _81279_ (_31536_, _31535_, _07141_);
  nor _81280_ (_31537_, _07141_, _31524_);
  or _81281_ (_31540_, _31537_, _06341_);
  or _81282_ (_31541_, _31540_, _31536_);
  and _81283_ (_31542_, _31541_, _06273_);
  and _81284_ (_31543_, _31542_, _31533_);
  nor _81285_ (_31544_, _07948_, _31524_);
  and _81286_ (_31545_, _14382_, _07948_);
  or _81287_ (_31546_, _31545_, _31544_);
  and _81288_ (_31547_, _31546_, _06272_);
  or _81289_ (_31548_, _31547_, _31543_);
  and _81290_ (_31549_, _31548_, _07166_);
  and _81291_ (_31550_, _31529_, _06461_);
  or _81292_ (_31551_, _31550_, _06464_);
  or _81293_ (_31552_, _31551_, _31549_);
  or _81294_ (_31553_, _31535_, _06465_);
  and _81295_ (_31554_, _31553_, _06269_);
  and _81296_ (_31555_, _31554_, _31552_);
  and _81297_ (_31556_, _31525_, _06268_);
  or _81298_ (_31557_, _31556_, _06261_);
  or _81299_ (_31558_, _31557_, _31555_);
  or _81300_ (_31559_, _31532_, _06262_);
  and _81301_ (_31562_, _31559_, _06258_);
  and _81302_ (_31563_, _31562_, _31558_);
  and _81303_ (_31564_, _14413_, _07948_);
  or _81304_ (_31565_, _31564_, _31544_);
  and _81305_ (_31566_, _31565_, _06257_);
  or _81306_ (_31567_, _31566_, _10080_);
  or _81307_ (_31568_, _31567_, _31563_);
  and _81308_ (_31569_, _31568_, _31530_);
  or _81309_ (_31570_, _31569_, _07460_);
  and _81310_ (_31571_, _09392_, _07926_);
  or _81311_ (_31572_, _31525_, _07208_);
  or _81312_ (_31573_, _31572_, _31571_);
  and _81313_ (_31574_, _31573_, _31570_);
  or _81314_ (_31575_, _31574_, _10094_);
  and _81315_ (_31576_, _14467_, _07926_);
  or _81316_ (_31577_, _31525_, _05982_);
  or _81317_ (_31578_, _31577_, _31576_);
  and _81318_ (_31579_, _31578_, _06219_);
  and _81319_ (_31580_, _31579_, _31575_);
  and _81320_ (_31581_, _07926_, _08954_);
  or _81321_ (_31584_, _31581_, _31525_);
  and _81322_ (_31585_, _31584_, _06218_);
  or _81323_ (_31586_, _31585_, _06369_);
  or _81324_ (_31587_, _31586_, _31580_);
  and _81325_ (_31588_, _14366_, _07926_);
  or _81326_ (_31589_, _31588_, _31525_);
  or _81327_ (_31590_, _31589_, _07237_);
  and _81328_ (_31591_, _31590_, _07240_);
  and _81329_ (_31592_, _31591_, _31587_);
  nor _81330_ (_31593_, _12580_, _13283_);
  or _81331_ (_31594_, _31593_, _31525_);
  and _81332_ (_31595_, _31523_, _06536_);
  and _81333_ (_31596_, _31595_, _31594_);
  or _81334_ (_31597_, _31596_, _31592_);
  and _81335_ (_31598_, _31597_, _07242_);
  nand _81336_ (_31599_, _31584_, _06375_);
  nor _81337_ (_31600_, _31599_, _31531_);
  or _81338_ (_31601_, _31600_, _06545_);
  or _81339_ (_31602_, _31601_, _31598_);
  and _81340_ (_31603_, _31602_, _31527_);
  or _81341_ (_31606_, _31603_, _06366_);
  and _81342_ (_31607_, _14363_, _07926_);
  or _81343_ (_31608_, _31607_, _31525_);
  or _81344_ (_31609_, _31608_, _09056_);
  and _81345_ (_31610_, _31609_, _09061_);
  and _81346_ (_31611_, _31610_, _31606_);
  and _81347_ (_31612_, _31594_, _06528_);
  or _81348_ (_31613_, _31612_, _06568_);
  or _81349_ (_31614_, _31613_, _31611_);
  or _81350_ (_31615_, _31532_, _06926_);
  and _81351_ (_31616_, _31615_, _31614_);
  or _81352_ (_31617_, _31616_, _05927_);
  or _81353_ (_31618_, _31525_, _05928_);
  and _81354_ (_31619_, _31618_, _31617_);
  or _81355_ (_31620_, _31619_, _06278_);
  or _81356_ (_31621_, _31532_, _06279_);
  and _81357_ (_31622_, _31621_, _01347_);
  and _81358_ (_31623_, _31622_, _31620_);
  nor _81359_ (_31624_, \oc8051_golden_model_1.P0 [0], rst);
  nor _81360_ (_31625_, _31624_, _01354_);
  or _81361_ (_43279_, _31625_, _31623_);
  nor _81362_ (_31628_, \oc8051_golden_model_1.P0 [1], rst);
  nor _81363_ (_31629_, _31628_, _01354_);
  not _81364_ (_31630_, \oc8051_golden_model_1.P0 [1]);
  nor _81365_ (_31631_, _07926_, _31630_);
  nor _81366_ (_31632_, _11261_, _13283_);
  or _81367_ (_31633_, _31632_, _31631_);
  or _81368_ (_31634_, _31633_, _09061_);
  nor _81369_ (_31635_, _13283_, _07357_);
  or _81370_ (_31636_, _31635_, _31631_);
  or _81371_ (_31637_, _31636_, _07166_);
  or _81372_ (_31638_, _07926_, \oc8051_golden_model_1.P0 [1]);
  and _81373_ (_31639_, _14562_, _07926_);
  not _81374_ (_31640_, _31639_);
  and _81375_ (_31641_, _31640_, _31638_);
  or _81376_ (_31642_, _31641_, _07151_);
  and _81377_ (_31643_, _07926_, \oc8051_golden_model_1.ACC [1]);
  or _81378_ (_31644_, _31643_, _31631_);
  and _81379_ (_31645_, _31644_, _07141_);
  nor _81380_ (_31646_, _07141_, _31630_);
  or _81381_ (_31649_, _31646_, _06341_);
  or _81382_ (_31650_, _31649_, _31645_);
  and _81383_ (_31651_, _31650_, _06273_);
  and _81384_ (_31652_, _31651_, _31642_);
  nor _81385_ (_31653_, _07948_, _31630_);
  and _81386_ (_31654_, _14557_, _07948_);
  or _81387_ (_31655_, _31654_, _31653_);
  and _81388_ (_31656_, _31655_, _06272_);
  or _81389_ (_31657_, _31656_, _06461_);
  or _81390_ (_31658_, _31657_, _31652_);
  and _81391_ (_31659_, _31658_, _31637_);
  or _81392_ (_31660_, _31659_, _06464_);
  or _81393_ (_31661_, _31644_, _06465_);
  and _81394_ (_31662_, _31661_, _06269_);
  and _81395_ (_31663_, _31662_, _31660_);
  and _81396_ (_31664_, _14560_, _07948_);
  or _81397_ (_31665_, _31664_, _31653_);
  and _81398_ (_31666_, _31665_, _06268_);
  or _81399_ (_31667_, _31666_, _06261_);
  or _81400_ (_31668_, _31667_, _31663_);
  and _81401_ (_31671_, _31654_, _14556_);
  or _81402_ (_31672_, _31653_, _06262_);
  or _81403_ (_31673_, _31672_, _31671_);
  and _81404_ (_31674_, _31673_, _06258_);
  and _81405_ (_31675_, _31674_, _31668_);
  or _81406_ (_31676_, _31653_, _14597_);
  and _81407_ (_31677_, _31676_, _06257_);
  and _81408_ (_31678_, _31677_, _31655_);
  or _81409_ (_31679_, _31678_, _10080_);
  or _81410_ (_31680_, _31679_, _31675_);
  or _81411_ (_31681_, _31636_, _07215_);
  and _81412_ (_31682_, _31681_, _31680_);
  or _81413_ (_31683_, _31682_, _07460_);
  and _81414_ (_31684_, _09451_, _07926_);
  or _81415_ (_31685_, _31631_, _07208_);
  or _81416_ (_31686_, _31685_, _31684_);
  and _81417_ (_31687_, _31686_, _05982_);
  and _81418_ (_31688_, _31687_, _31683_);
  and _81419_ (_31689_, _14653_, _07926_);
  or _81420_ (_31690_, _31689_, _31631_);
  and _81421_ (_31693_, _31690_, _10094_);
  or _81422_ (_31694_, _31693_, _31688_);
  and _81423_ (_31695_, _31694_, _06219_);
  nand _81424_ (_31696_, _07926_, _07038_);
  and _81425_ (_31697_, _31638_, _06218_);
  and _81426_ (_31698_, _31697_, _31696_);
  or _81427_ (_31699_, _31698_, _31695_);
  and _81428_ (_31700_, _31699_, _07237_);
  or _81429_ (_31701_, _14668_, _13283_);
  and _81430_ (_31702_, _31638_, _06369_);
  and _81431_ (_31703_, _31702_, _31701_);
  or _81432_ (_31704_, _31703_, _06536_);
  or _81433_ (_31705_, _31704_, _31700_);
  nand _81434_ (_31706_, _11260_, _07926_);
  and _81435_ (_31707_, _31706_, _31633_);
  or _81436_ (_31708_, _31707_, _07240_);
  and _81437_ (_31709_, _31708_, _07242_);
  and _81438_ (_31710_, _31709_, _31705_);
  or _81439_ (_31711_, _14666_, _13283_);
  and _81440_ (_31712_, _31638_, _06375_);
  and _81441_ (_31715_, _31712_, _31711_);
  or _81442_ (_31716_, _31715_, _06545_);
  or _81443_ (_31717_, _31716_, _31710_);
  nor _81444_ (_31718_, _31631_, _07234_);
  nand _81445_ (_31719_, _31718_, _31706_);
  and _81446_ (_31720_, _31719_, _09056_);
  and _81447_ (_31721_, _31720_, _31717_);
  or _81448_ (_31722_, _31696_, _08341_);
  and _81449_ (_31723_, _31638_, _06366_);
  and _81450_ (_31724_, _31723_, _31722_);
  or _81451_ (_31725_, _31724_, _06528_);
  or _81452_ (_31726_, _31725_, _31721_);
  and _81453_ (_31727_, _31726_, _31634_);
  or _81454_ (_31728_, _31727_, _06568_);
  or _81455_ (_31729_, _31641_, _06926_);
  and _81456_ (_31730_, _31729_, _05928_);
  and _81457_ (_31731_, _31730_, _31728_);
  and _81458_ (_31732_, _31665_, _05927_);
  or _81459_ (_31733_, _31732_, _06278_);
  or _81460_ (_31734_, _31733_, _31731_);
  or _81461_ (_31737_, _31631_, _06279_);
  or _81462_ (_31738_, _31737_, _31639_);
  and _81463_ (_31739_, _31738_, _01347_);
  and _81464_ (_31740_, _31739_, _31734_);
  or _81465_ (_43280_, _31740_, _31629_);
  and _81466_ (_31741_, _13283_, \oc8051_golden_model_1.P0 [2]);
  nor _81467_ (_31742_, _13283_, _07776_);
  or _81468_ (_31743_, _31742_, _31741_);
  or _81469_ (_31744_, _31743_, _07215_);
  or _81470_ (_31745_, _31743_, _07166_);
  and _81471_ (_31746_, _14770_, _07926_);
  or _81472_ (_31747_, _31746_, _31741_);
  or _81473_ (_31748_, _31747_, _07151_);
  and _81474_ (_31749_, _07926_, \oc8051_golden_model_1.ACC [2]);
  or _81475_ (_31750_, _31749_, _31741_);
  and _81476_ (_31751_, _31750_, _07141_);
  and _81477_ (_31752_, _07142_, \oc8051_golden_model_1.P0 [2]);
  or _81478_ (_31753_, _31752_, _06341_);
  or _81479_ (_31754_, _31753_, _31751_);
  and _81480_ (_31755_, _31754_, _06273_);
  and _81481_ (_31758_, _31755_, _31748_);
  and _81482_ (_31759_, _13291_, \oc8051_golden_model_1.P0 [2]);
  and _81483_ (_31760_, _14774_, _07948_);
  or _81484_ (_31761_, _31760_, _31759_);
  and _81485_ (_31762_, _31761_, _06272_);
  or _81486_ (_31763_, _31762_, _06461_);
  or _81487_ (_31764_, _31763_, _31758_);
  and _81488_ (_31765_, _31764_, _31745_);
  or _81489_ (_31766_, _31765_, _06464_);
  or _81490_ (_31767_, _31750_, _06465_);
  and _81491_ (_31769_, _31767_, _06269_);
  and _81492_ (_31770_, _31769_, _31766_);
  and _81493_ (_31771_, _14756_, _07948_);
  or _81494_ (_31772_, _31771_, _31759_);
  and _81495_ (_31773_, _31772_, _06268_);
  or _81496_ (_31774_, _31773_, _06261_);
  or _81497_ (_31775_, _31774_, _31770_);
  and _81498_ (_31776_, _31760_, _14789_);
  or _81499_ (_31777_, _31759_, _06262_);
  or _81500_ (_31778_, _31777_, _31776_);
  and _81501_ (_31780_, _31778_, _06258_);
  and _81502_ (_31781_, _31780_, _31775_);
  and _81503_ (_31782_, _14804_, _07948_);
  or _81504_ (_31783_, _31782_, _31759_);
  and _81505_ (_31784_, _31783_, _06257_);
  or _81506_ (_31785_, _31784_, _10080_);
  or _81507_ (_31786_, _31785_, _31781_);
  and _81508_ (_31787_, _31786_, _31744_);
  or _81509_ (_31788_, _31787_, _07460_);
  and _81510_ (_31789_, _09450_, _07926_);
  or _81511_ (_31791_, _31741_, _07208_);
  or _81512_ (_31792_, _31791_, _31789_);
  and _81513_ (_31793_, _31792_, _05982_);
  and _81514_ (_31794_, _31793_, _31788_);
  and _81515_ (_31795_, _14859_, _07926_);
  or _81516_ (_31796_, _31795_, _31741_);
  and _81517_ (_31797_, _31796_, _10094_);
  or _81518_ (_31798_, _31797_, _06218_);
  or _81519_ (_31799_, _31798_, _31794_);
  and _81520_ (_31800_, _07926_, _08973_);
  or _81521_ (_31802_, _31800_, _31741_);
  or _81522_ (_31803_, _31802_, _06219_);
  and _81523_ (_31804_, _31803_, _31799_);
  or _81524_ (_31805_, _31804_, _06369_);
  and _81525_ (_31806_, _14751_, _07926_);
  or _81526_ (_31807_, _31806_, _31741_);
  or _81527_ (_31808_, _31807_, _07237_);
  and _81528_ (_31809_, _31808_, _07240_);
  and _81529_ (_31810_, _31809_, _31805_);
  and _81530_ (_31811_, _11259_, _07926_);
  or _81531_ (_31813_, _31811_, _31741_);
  and _81532_ (_31814_, _31813_, _06536_);
  or _81533_ (_31815_, _31814_, _31810_);
  and _81534_ (_31816_, _31815_, _07242_);
  or _81535_ (_31817_, _31741_, _08440_);
  and _81536_ (_31818_, _31802_, _06375_);
  and _81537_ (_31819_, _31818_, _31817_);
  or _81538_ (_31820_, _31819_, _31816_);
  and _81539_ (_31821_, _31820_, _07234_);
  and _81540_ (_31822_, _31750_, _06545_);
  and _81541_ (_31824_, _31822_, _31817_);
  or _81542_ (_31825_, _31824_, _06366_);
  or _81543_ (_31826_, _31825_, _31821_);
  and _81544_ (_31827_, _14748_, _07926_);
  or _81545_ (_31828_, _31741_, _09056_);
  or _81546_ (_31829_, _31828_, _31827_);
  and _81547_ (_31830_, _31829_, _09061_);
  and _81548_ (_31831_, _31830_, _31826_);
  nor _81549_ (_31832_, _11258_, _13283_);
  or _81550_ (_31833_, _31832_, _31741_);
  and _81551_ (_31835_, _31833_, _06528_);
  or _81552_ (_31836_, _31835_, _06568_);
  or _81553_ (_31837_, _31836_, _31831_);
  or _81554_ (_31838_, _31747_, _06926_);
  and _81555_ (_31839_, _31838_, _05928_);
  and _81556_ (_31840_, _31839_, _31837_);
  and _81557_ (_31841_, _31772_, _05927_);
  or _81558_ (_31842_, _31841_, _06278_);
  or _81559_ (_31843_, _31842_, _31840_);
  and _81560_ (_31844_, _14926_, _07926_);
  or _81561_ (_31846_, _31741_, _06279_);
  or _81562_ (_31847_, _31846_, _31844_);
  and _81563_ (_31848_, _31847_, _01347_);
  and _81564_ (_31849_, _31848_, _31843_);
  nor _81565_ (_31850_, \oc8051_golden_model_1.P0 [2], rst);
  nor _81566_ (_31851_, _31850_, _01354_);
  or _81567_ (_43281_, _31851_, _31849_);
  and _81568_ (_31852_, _13283_, \oc8051_golden_model_1.P0 [3]);
  nor _81569_ (_31853_, _13283_, _07594_);
  or _81570_ (_31854_, _31853_, _31852_);
  or _81571_ (_31856_, _31854_, _07215_);
  and _81572_ (_31857_, _14953_, _07926_);
  or _81573_ (_31858_, _31857_, _31852_);
  or _81574_ (_31859_, _31858_, _07151_);
  and _81575_ (_31860_, _07926_, \oc8051_golden_model_1.ACC [3]);
  or _81576_ (_31861_, _31860_, _31852_);
  and _81577_ (_31862_, _31861_, _07141_);
  and _81578_ (_31863_, _07142_, \oc8051_golden_model_1.P0 [3]);
  or _81579_ (_31864_, _31863_, _06341_);
  or _81580_ (_31865_, _31864_, _31862_);
  and _81581_ (_31867_, _31865_, _06273_);
  and _81582_ (_31868_, _31867_, _31859_);
  and _81583_ (_31869_, _13291_, \oc8051_golden_model_1.P0 [3]);
  and _81584_ (_31870_, _14950_, _07948_);
  or _81585_ (_31871_, _31870_, _31869_);
  and _81586_ (_31872_, _31871_, _06272_);
  or _81587_ (_31873_, _31872_, _06461_);
  or _81588_ (_31874_, _31873_, _31868_);
  or _81589_ (_31875_, _31854_, _07166_);
  and _81590_ (_31876_, _31875_, _31874_);
  or _81591_ (_31878_, _31876_, _06464_);
  or _81592_ (_31879_, _31861_, _06465_);
  and _81593_ (_31880_, _31879_, _06269_);
  and _81594_ (_31881_, _31880_, _31878_);
  and _81595_ (_31882_, _14948_, _07948_);
  or _81596_ (_31883_, _31882_, _31869_);
  and _81597_ (_31884_, _31883_, _06268_);
  or _81598_ (_31885_, _31884_, _06261_);
  or _81599_ (_31886_, _31885_, _31881_);
  or _81600_ (_31887_, _31869_, _14979_);
  and _81601_ (_31889_, _31887_, _31871_);
  or _81602_ (_31890_, _31889_, _06262_);
  and _81603_ (_31891_, _31890_, _06258_);
  and _81604_ (_31892_, _31891_, _31886_);
  or _81605_ (_31893_, _31869_, _14992_);
  and _81606_ (_31894_, _31893_, _06257_);
  and _81607_ (_31895_, _31894_, _31871_);
  or _81608_ (_31896_, _31895_, _10080_);
  or _81609_ (_31897_, _31896_, _31892_);
  and _81610_ (_31898_, _31897_, _31856_);
  or _81611_ (_31900_, _31898_, _07460_);
  and _81612_ (_31901_, _09449_, _07926_);
  or _81613_ (_31902_, _31852_, _07208_);
  or _81614_ (_31903_, _31902_, _31901_);
  and _81615_ (_31904_, _31903_, _05982_);
  and _81616_ (_31905_, _31904_, _31900_);
  and _81617_ (_31906_, _15048_, _07926_);
  or _81618_ (_31907_, _31906_, _31852_);
  and _81619_ (_31908_, _31907_, _10094_);
  or _81620_ (_31909_, _31908_, _06218_);
  or _81621_ (_31911_, _31909_, _31905_);
  and _81622_ (_31912_, _07926_, _08930_);
  or _81623_ (_31913_, _31912_, _31852_);
  or _81624_ (_31914_, _31913_, _06219_);
  and _81625_ (_31915_, _31914_, _31911_);
  or _81626_ (_31916_, _31915_, _06369_);
  and _81627_ (_31917_, _14943_, _07926_);
  or _81628_ (_31918_, _31917_, _31852_);
  or _81629_ (_31919_, _31918_, _07237_);
  and _81630_ (_31920_, _31919_, _07240_);
  and _81631_ (_31922_, _31920_, _31916_);
  and _81632_ (_31923_, _12577_, _07926_);
  or _81633_ (_31924_, _31923_, _31852_);
  and _81634_ (_31925_, _31924_, _06536_);
  or _81635_ (_31926_, _31925_, _31922_);
  and _81636_ (_31927_, _31926_, _07242_);
  or _81637_ (_31928_, _31852_, _08292_);
  and _81638_ (_31929_, _31913_, _06375_);
  and _81639_ (_31930_, _31929_, _31928_);
  or _81640_ (_31931_, _31930_, _31927_);
  and _81641_ (_31933_, _31931_, _07234_);
  and _81642_ (_31934_, _31861_, _06545_);
  and _81643_ (_31935_, _31934_, _31928_);
  or _81644_ (_31936_, _31935_, _06366_);
  or _81645_ (_31937_, _31936_, _31933_);
  and _81646_ (_31938_, _14940_, _07926_);
  or _81647_ (_31939_, _31852_, _09056_);
  or _81648_ (_31940_, _31939_, _31938_);
  and _81649_ (_31941_, _31940_, _09061_);
  and _81650_ (_31942_, _31941_, _31937_);
  nor _81651_ (_31944_, _11256_, _13283_);
  or _81652_ (_31945_, _31944_, _31852_);
  and _81653_ (_31946_, _31945_, _06528_);
  or _81654_ (_31947_, _31946_, _06568_);
  or _81655_ (_31948_, _31947_, _31942_);
  or _81656_ (_31949_, _31858_, _06926_);
  and _81657_ (_31950_, _31949_, _05928_);
  and _81658_ (_31951_, _31950_, _31948_);
  and _81659_ (_31952_, _31883_, _05927_);
  or _81660_ (_31953_, _31952_, _06278_);
  or _81661_ (_31954_, _31953_, _31951_);
  and _81662_ (_31955_, _15128_, _07926_);
  or _81663_ (_31956_, _31852_, _06279_);
  or _81664_ (_31957_, _31956_, _31955_);
  and _81665_ (_31958_, _31957_, _01347_);
  and _81666_ (_31959_, _31958_, _31954_);
  nor _81667_ (_31960_, \oc8051_golden_model_1.P0 [3], rst);
  nor _81668_ (_31961_, _31960_, _01354_);
  or _81669_ (_43283_, _31961_, _31959_);
  nor _81670_ (_31962_, \oc8051_golden_model_1.P0 [4], rst);
  nor _81671_ (_31964_, _31962_, _01354_);
  and _81672_ (_31965_, _13283_, \oc8051_golden_model_1.P0 [4]);
  nor _81673_ (_31966_, _08541_, _13283_);
  or _81674_ (_31967_, _31966_, _31965_);
  or _81675_ (_31968_, _31967_, _07215_);
  and _81676_ (_31969_, _13291_, \oc8051_golden_model_1.P0 [4]);
  and _81677_ (_31970_, _15176_, _07948_);
  or _81678_ (_31971_, _31970_, _31969_);
  and _81679_ (_31972_, _31971_, _06268_);
  and _81680_ (_31973_, _15162_, _07926_);
  or _81681_ (_31975_, _31973_, _31965_);
  or _81682_ (_31976_, _31975_, _07151_);
  and _81683_ (_31977_, _07926_, \oc8051_golden_model_1.ACC [4]);
  or _81684_ (_31978_, _31977_, _31965_);
  and _81685_ (_31979_, _31978_, _07141_);
  and _81686_ (_31980_, _07142_, \oc8051_golden_model_1.P0 [4]);
  or _81687_ (_31981_, _31980_, _06341_);
  or _81688_ (_31982_, _31981_, _31979_);
  and _81689_ (_31983_, _31982_, _06273_);
  and _81690_ (_31984_, _31983_, _31976_);
  and _81691_ (_31986_, _15166_, _07948_);
  or _81692_ (_31987_, _31986_, _31969_);
  and _81693_ (_31988_, _31987_, _06272_);
  or _81694_ (_31989_, _31988_, _06461_);
  or _81695_ (_31990_, _31989_, _31984_);
  or _81696_ (_31991_, _31967_, _07166_);
  and _81697_ (_31992_, _31991_, _31990_);
  or _81698_ (_31993_, _31992_, _06464_);
  or _81699_ (_31994_, _31978_, _06465_);
  and _81700_ (_31995_, _31994_, _06269_);
  and _81701_ (_31997_, _31995_, _31993_);
  or _81702_ (_31998_, _31997_, _31972_);
  and _81703_ (_31999_, _31998_, _06262_);
  and _81704_ (_32000_, _15184_, _07948_);
  or _81705_ (_32001_, _32000_, _31969_);
  and _81706_ (_32002_, _32001_, _06261_);
  or _81707_ (_32003_, _32002_, _31999_);
  and _81708_ (_32004_, _32003_, _06258_);
  and _81709_ (_32005_, _15200_, _07948_);
  or _81710_ (_32006_, _32005_, _31969_);
  and _81711_ (_32008_, _32006_, _06257_);
  or _81712_ (_32009_, _32008_, _10080_);
  or _81713_ (_32010_, _32009_, _32004_);
  and _81714_ (_32011_, _32010_, _31968_);
  or _81715_ (_32012_, _32011_, _07460_);
  and _81716_ (_32013_, _09448_, _07926_);
  or _81717_ (_32014_, _31965_, _07208_);
  or _81718_ (_32015_, _32014_, _32013_);
  and _81719_ (_32016_, _32015_, _05982_);
  and _81720_ (_32017_, _32016_, _32012_);
  and _81721_ (_32019_, _15254_, _07926_);
  or _81722_ (_32020_, _32019_, _31965_);
  and _81723_ (_32021_, _32020_, _10094_);
  or _81724_ (_32022_, _32021_, _06218_);
  or _81725_ (_32023_, _32022_, _32017_);
  and _81726_ (_32024_, _08959_, _07926_);
  or _81727_ (_32025_, _32024_, _31965_);
  or _81728_ (_32026_, _32025_, _06219_);
  and _81729_ (_32027_, _32026_, _32023_);
  or _81730_ (_32028_, _32027_, _06369_);
  and _81731_ (_32030_, _15269_, _07926_);
  or _81732_ (_32031_, _32030_, _31965_);
  or _81733_ (_32032_, _32031_, _07237_);
  and _81734_ (_32033_, _32032_, _07240_);
  and _81735_ (_32034_, _32033_, _32028_);
  and _81736_ (_32035_, _11254_, _07926_);
  or _81737_ (_32036_, _32035_, _31965_);
  and _81738_ (_32037_, _32036_, _06536_);
  or _81739_ (_32038_, _32037_, _32034_);
  and _81740_ (_32039_, _32038_, _07242_);
  or _81741_ (_32041_, _31965_, _08544_);
  and _81742_ (_32042_, _32025_, _06375_);
  and _81743_ (_32043_, _32042_, _32041_);
  or _81744_ (_32044_, _32043_, _32039_);
  and _81745_ (_32045_, _32044_, _07234_);
  and _81746_ (_32046_, _31978_, _06545_);
  and _81747_ (_32047_, _32046_, _32041_);
  or _81748_ (_32048_, _32047_, _06366_);
  or _81749_ (_32049_, _32048_, _32045_);
  and _81750_ (_32050_, _15266_, _07926_);
  or _81751_ (_32052_, _31965_, _09056_);
  or _81752_ (_32053_, _32052_, _32050_);
  and _81753_ (_32054_, _32053_, _09061_);
  and _81754_ (_32055_, _32054_, _32049_);
  nor _81755_ (_32056_, _11253_, _13283_);
  or _81756_ (_32057_, _32056_, _31965_);
  and _81757_ (_32058_, _32057_, _06528_);
  or _81758_ (_32059_, _32058_, _06568_);
  or _81759_ (_32060_, _32059_, _32055_);
  or _81760_ (_32061_, _31975_, _06926_);
  and _81761_ (_32063_, _32061_, _05928_);
  and _81762_ (_32064_, _32063_, _32060_);
  and _81763_ (_32065_, _31971_, _05927_);
  or _81764_ (_32066_, _32065_, _06278_);
  or _81765_ (_32067_, _32066_, _32064_);
  and _81766_ (_32068_, _15329_, _07926_);
  or _81767_ (_32069_, _31965_, _06279_);
  or _81768_ (_32070_, _32069_, _32068_);
  and _81769_ (_32071_, _32070_, _01347_);
  and _81770_ (_32072_, _32071_, _32067_);
  or _81771_ (_43284_, _32072_, _31964_);
  and _81772_ (_32074_, _13283_, \oc8051_golden_model_1.P0 [5]);
  and _81773_ (_32075_, _15358_, _07926_);
  or _81774_ (_32076_, _32075_, _32074_);
  or _81775_ (_32077_, _32076_, _07151_);
  and _81776_ (_32078_, _07926_, \oc8051_golden_model_1.ACC [5]);
  or _81777_ (_32079_, _32078_, _32074_);
  and _81778_ (_32080_, _32079_, _07141_);
  and _81779_ (_32081_, _07142_, \oc8051_golden_model_1.P0 [5]);
  or _81780_ (_32082_, _32081_, _06341_);
  or _81781_ (_32084_, _32082_, _32080_);
  and _81782_ (_32085_, _32084_, _06273_);
  and _81783_ (_32086_, _32085_, _32077_);
  and _81784_ (_32087_, _13291_, \oc8051_golden_model_1.P0 [5]);
  and _81785_ (_32088_, _15372_, _07948_);
  or _81786_ (_32089_, _32088_, _32087_);
  and _81787_ (_32090_, _32089_, _06272_);
  or _81788_ (_32091_, _32090_, _06461_);
  or _81789_ (_32092_, _32091_, _32086_);
  nor _81790_ (_32093_, _08244_, _13283_);
  or _81791_ (_32095_, _32093_, _32074_);
  or _81792_ (_32096_, _32095_, _07166_);
  and _81793_ (_32097_, _32096_, _32092_);
  or _81794_ (_32098_, _32097_, _06464_);
  or _81795_ (_32099_, _32079_, _06465_);
  and _81796_ (_32100_, _32099_, _06269_);
  and _81797_ (_32101_, _32100_, _32098_);
  and _81798_ (_32102_, _15355_, _07948_);
  or _81799_ (_32103_, _32102_, _32087_);
  and _81800_ (_32104_, _32103_, _06268_);
  or _81801_ (_32106_, _32104_, _06261_);
  or _81802_ (_32107_, _32106_, _32101_);
  or _81803_ (_32108_, _32087_, _15387_);
  and _81804_ (_32109_, _32108_, _32089_);
  or _81805_ (_32110_, _32109_, _06262_);
  and _81806_ (_32111_, _32110_, _06258_);
  and _81807_ (_32112_, _32111_, _32107_);
  or _81808_ (_32113_, _32087_, _15403_);
  and _81809_ (_32114_, _32113_, _06257_);
  and _81810_ (_32115_, _32114_, _32089_);
  or _81811_ (_32117_, _32115_, _10080_);
  or _81812_ (_32118_, _32117_, _32112_);
  or _81813_ (_32119_, _32095_, _07215_);
  and _81814_ (_32120_, _32119_, _32118_);
  or _81815_ (_32121_, _32120_, _07460_);
  and _81816_ (_32122_, _09447_, _07926_);
  or _81817_ (_32123_, _32074_, _07208_);
  or _81818_ (_32124_, _32123_, _32122_);
  and _81819_ (_32125_, _32124_, _05982_);
  and _81820_ (_32126_, _32125_, _32121_);
  and _81821_ (_32128_, _15459_, _07926_);
  or _81822_ (_32129_, _32128_, _32074_);
  and _81823_ (_32130_, _32129_, _10094_);
  or _81824_ (_32131_, _32130_, _06218_);
  or _81825_ (_32132_, _32131_, _32126_);
  and _81826_ (_32133_, _08946_, _07926_);
  or _81827_ (_32134_, _32133_, _32074_);
  or _81828_ (_32135_, _32134_, _06219_);
  and _81829_ (_32136_, _32135_, _32132_);
  or _81830_ (_32137_, _32136_, _06369_);
  and _81831_ (_32139_, _15353_, _07926_);
  or _81832_ (_32140_, _32139_, _32074_);
  or _81833_ (_32141_, _32140_, _07237_);
  and _81834_ (_32142_, _32141_, _07240_);
  and _81835_ (_32143_, _32142_, _32137_);
  and _81836_ (_32144_, _11250_, _07926_);
  or _81837_ (_32145_, _32144_, _32074_);
  and _81838_ (_32146_, _32145_, _06536_);
  or _81839_ (_32147_, _32146_, _32143_);
  and _81840_ (_32148_, _32147_, _07242_);
  or _81841_ (_32150_, _32074_, _08247_);
  and _81842_ (_32151_, _32134_, _06375_);
  and _81843_ (_32152_, _32151_, _32150_);
  or _81844_ (_32153_, _32152_, _32148_);
  and _81845_ (_32154_, _32153_, _07234_);
  and _81846_ (_32155_, _32079_, _06545_);
  and _81847_ (_32156_, _32155_, _32150_);
  or _81848_ (_32157_, _32156_, _06366_);
  or _81849_ (_32158_, _32157_, _32154_);
  and _81850_ (_32159_, _15350_, _07926_);
  or _81851_ (_32161_, _32074_, _09056_);
  or _81852_ (_32162_, _32161_, _32159_);
  and _81853_ (_32163_, _32162_, _09061_);
  and _81854_ (_32164_, _32163_, _32158_);
  nor _81855_ (_32165_, _11249_, _13283_);
  or _81856_ (_32166_, _32165_, _32074_);
  and _81857_ (_32167_, _32166_, _06528_);
  or _81858_ (_32168_, _32167_, _06568_);
  or _81859_ (_32169_, _32168_, _32164_);
  or _81860_ (_32170_, _32076_, _06926_);
  and _81861_ (_32172_, _32170_, _05928_);
  and _81862_ (_32173_, _32172_, _32169_);
  and _81863_ (_32174_, _32103_, _05927_);
  or _81864_ (_32175_, _32174_, _06278_);
  or _81865_ (_32176_, _32175_, _32173_);
  and _81866_ (_32177_, _15532_, _07926_);
  or _81867_ (_32178_, _32074_, _06279_);
  or _81868_ (_32179_, _32178_, _32177_);
  and _81869_ (_32180_, _32179_, _01347_);
  and _81870_ (_32181_, _32180_, _32176_);
  nor _81871_ (_32183_, \oc8051_golden_model_1.P0 [5], rst);
  nor _81872_ (_32184_, _32183_, _01354_);
  or _81873_ (_43285_, _32184_, _32181_);
  and _81874_ (_32185_, _13283_, \oc8051_golden_model_1.P0 [6]);
  and _81875_ (_32186_, _15554_, _07926_);
  or _81876_ (_32187_, _32186_, _32185_);
  or _81877_ (_32188_, _32187_, _07151_);
  and _81878_ (_32189_, _07926_, \oc8051_golden_model_1.ACC [6]);
  or _81879_ (_32190_, _32189_, _32185_);
  and _81880_ (_32191_, _32190_, _07141_);
  and _81881_ (_32193_, _07142_, \oc8051_golden_model_1.P0 [6]);
  or _81882_ (_32194_, _32193_, _06341_);
  or _81883_ (_32195_, _32194_, _32191_);
  and _81884_ (_32196_, _32195_, _06273_);
  and _81885_ (_32197_, _32196_, _32188_);
  and _81886_ (_32198_, _13291_, \oc8051_golden_model_1.P0 [6]);
  and _81887_ (_32199_, _15570_, _07948_);
  or _81888_ (_32200_, _32199_, _32198_);
  and _81889_ (_32201_, _32200_, _06272_);
  or _81890_ (_32202_, _32201_, _06461_);
  or _81891_ (_32204_, _32202_, _32197_);
  nor _81892_ (_32205_, _08142_, _13283_);
  or _81893_ (_32206_, _32205_, _32185_);
  or _81894_ (_32207_, _32206_, _07166_);
  and _81895_ (_32208_, _32207_, _32204_);
  or _81896_ (_32209_, _32208_, _06464_);
  or _81897_ (_32210_, _32190_, _06465_);
  and _81898_ (_32211_, _32210_, _06269_);
  and _81899_ (_32212_, _32211_, _32209_);
  and _81900_ (_32213_, _15551_, _07948_);
  or _81901_ (_32215_, _32213_, _32198_);
  and _81902_ (_32216_, _32215_, _06268_);
  or _81903_ (_32217_, _32216_, _06261_);
  or _81904_ (_32218_, _32217_, _32212_);
  or _81905_ (_32219_, _32198_, _15585_);
  and _81906_ (_32220_, _32219_, _32200_);
  or _81907_ (_32221_, _32220_, _06262_);
  and _81908_ (_32222_, _32221_, _06258_);
  and _81909_ (_32223_, _32222_, _32218_);
  and _81910_ (_32224_, _15602_, _07948_);
  or _81911_ (_32226_, _32224_, _32198_);
  and _81912_ (_32227_, _32226_, _06257_);
  or _81913_ (_32228_, _32227_, _10080_);
  or _81914_ (_32229_, _32228_, _32223_);
  or _81915_ (_32230_, _32206_, _07215_);
  and _81916_ (_32231_, _32230_, _32229_);
  or _81917_ (_32232_, _32231_, _07460_);
  and _81918_ (_32233_, _09446_, _07926_);
  or _81919_ (_32234_, _32185_, _07208_);
  or _81920_ (_32235_, _32234_, _32233_);
  and _81921_ (_32237_, _32235_, _05982_);
  and _81922_ (_32238_, _32237_, _32232_);
  and _81923_ (_32239_, _15657_, _07926_);
  or _81924_ (_32240_, _32239_, _32185_);
  and _81925_ (_32241_, _32240_, _10094_);
  or _81926_ (_32242_, _32241_, _06218_);
  or _81927_ (_32243_, _32242_, _32238_);
  and _81928_ (_32244_, _15664_, _07926_);
  or _81929_ (_32245_, _32244_, _32185_);
  or _81930_ (_32246_, _32245_, _06219_);
  and _81931_ (_32248_, _32246_, _32243_);
  or _81932_ (_32249_, _32248_, _06369_);
  and _81933_ (_32250_, _15549_, _07926_);
  or _81934_ (_32251_, _32250_, _32185_);
  or _81935_ (_32252_, _32251_, _07237_);
  and _81936_ (_32253_, _32252_, _07240_);
  and _81937_ (_32254_, _32253_, _32249_);
  and _81938_ (_32255_, _11247_, _07926_);
  or _81939_ (_32256_, _32255_, _32185_);
  and _81940_ (_32257_, _32256_, _06536_);
  or _81941_ (_32259_, _32257_, _32254_);
  and _81942_ (_32260_, _32259_, _07242_);
  or _81943_ (_32261_, _32185_, _08145_);
  and _81944_ (_32262_, _32245_, _06375_);
  and _81945_ (_32263_, _32262_, _32261_);
  or _81946_ (_32264_, _32263_, _32260_);
  and _81947_ (_32265_, _32264_, _07234_);
  and _81948_ (_32266_, _32190_, _06545_);
  and _81949_ (_32267_, _32266_, _32261_);
  or _81950_ (_32268_, _32267_, _06366_);
  or _81951_ (_32270_, _32268_, _32265_);
  and _81952_ (_32271_, _15546_, _07926_);
  or _81953_ (_32272_, _32185_, _09056_);
  or _81954_ (_32273_, _32272_, _32271_);
  and _81955_ (_32274_, _32273_, _09061_);
  and _81956_ (_32275_, _32274_, _32270_);
  nor _81957_ (_32276_, _11246_, _13283_);
  or _81958_ (_32277_, _32276_, _32185_);
  and _81959_ (_32278_, _32277_, _06528_);
  or _81960_ (_32279_, _32278_, _06568_);
  or _81961_ (_32281_, _32279_, _32275_);
  or _81962_ (_32282_, _32187_, _06926_);
  and _81963_ (_32283_, _32282_, _05928_);
  and _81964_ (_32284_, _32283_, _32281_);
  and _81965_ (_32285_, _32215_, _05927_);
  or _81966_ (_32286_, _32285_, _06278_);
  or _81967_ (_32287_, _32286_, _32284_);
  and _81968_ (_32288_, _15734_, _07926_);
  or _81969_ (_32289_, _32185_, _06279_);
  or _81970_ (_32290_, _32289_, _32288_);
  and _81971_ (_32292_, _32290_, _01347_);
  and _81972_ (_32293_, _32292_, _32287_);
  nor _81973_ (_32294_, \oc8051_golden_model_1.P0 [6], rst);
  nor _81974_ (_32295_, _32294_, _01354_);
  or _81975_ (_43286_, _32295_, _32293_);
  nor _81976_ (_32296_, \oc8051_golden_model_1.P1 [0], rst);
  nor _81977_ (_32297_, _32296_, _01354_);
  nand _81978_ (_32298_, _11263_, _07971_);
  and _81979_ (_32299_, _13388_, \oc8051_golden_model_1.P1 [0]);
  nor _81980_ (_32300_, _32299_, _07234_);
  nand _81981_ (_32302_, _32300_, _32298_);
  and _81982_ (_32303_, _07971_, _07133_);
  or _81983_ (_32304_, _32303_, _32299_);
  or _81984_ (_32305_, _32304_, _07215_);
  nor _81985_ (_32306_, _08390_, _13388_);
  or _81986_ (_32307_, _32306_, _32299_);
  and _81987_ (_32308_, _32307_, _06341_);
  and _81988_ (_32309_, _07142_, \oc8051_golden_model_1.P1 [0]);
  and _81989_ (_32310_, _07971_, \oc8051_golden_model_1.ACC [0]);
  or _81990_ (_32311_, _32310_, _32299_);
  and _81991_ (_32313_, _32311_, _07141_);
  or _81992_ (_32314_, _32313_, _32309_);
  and _81993_ (_32315_, _32314_, _07151_);
  or _81994_ (_32316_, _32315_, _06272_);
  or _81995_ (_32317_, _32316_, _32308_);
  and _81996_ (_32318_, _14382_, _08620_);
  and _81997_ (_32319_, _13396_, \oc8051_golden_model_1.P1 [0]);
  or _81998_ (_32320_, _32319_, _06273_);
  or _81999_ (_32321_, _32320_, _32318_);
  and _82000_ (_32322_, _32321_, _07166_);
  and _82001_ (_32324_, _32322_, _32317_);
  and _82002_ (_32325_, _32304_, _06461_);
  or _82003_ (_32326_, _32325_, _06464_);
  or _82004_ (_32327_, _32326_, _32324_);
  or _82005_ (_32328_, _32311_, _06465_);
  and _82006_ (_32329_, _32328_, _06269_);
  and _82007_ (_32330_, _32329_, _32327_);
  and _82008_ (_32331_, _32299_, _06268_);
  or _82009_ (_32332_, _32331_, _06261_);
  or _82010_ (_32333_, _32332_, _32330_);
  or _82011_ (_32335_, _32307_, _06262_);
  and _82012_ (_32336_, _32335_, _06258_);
  and _82013_ (_32337_, _32336_, _32333_);
  and _82014_ (_32338_, _14413_, _08620_);
  or _82015_ (_32339_, _32338_, _32319_);
  and _82016_ (_32340_, _32339_, _06257_);
  or _82017_ (_32341_, _32340_, _10080_);
  or _82018_ (_32342_, _32341_, _32337_);
  and _82019_ (_32343_, _32342_, _32305_);
  or _82020_ (_32344_, _32343_, _07460_);
  and _82021_ (_32346_, _09392_, _07971_);
  or _82022_ (_32347_, _32299_, _07208_);
  or _82023_ (_32348_, _32347_, _32346_);
  and _82024_ (_32349_, _32348_, _32344_);
  or _82025_ (_32350_, _32349_, _10094_);
  and _82026_ (_32351_, _14467_, _07971_);
  or _82027_ (_32352_, _32299_, _05982_);
  or _82028_ (_32353_, _32352_, _32351_);
  and _82029_ (_32354_, _32353_, _06219_);
  and _82030_ (_32355_, _32354_, _32350_);
  and _82031_ (_32357_, _07971_, _08954_);
  or _82032_ (_32358_, _32357_, _32299_);
  and _82033_ (_32359_, _32358_, _06218_);
  or _82034_ (_32360_, _32359_, _06369_);
  or _82035_ (_32361_, _32360_, _32355_);
  and _82036_ (_32362_, _14366_, _07971_);
  or _82037_ (_32363_, _32362_, _32299_);
  or _82038_ (_32364_, _32363_, _07237_);
  and _82039_ (_32365_, _32364_, _07240_);
  and _82040_ (_32366_, _32365_, _32361_);
  nor _82041_ (_32368_, _12580_, _13388_);
  or _82042_ (_32369_, _32368_, _32299_);
  and _82043_ (_32370_, _32298_, _06536_);
  and _82044_ (_32371_, _32370_, _32369_);
  or _82045_ (_32372_, _32371_, _32366_);
  and _82046_ (_32373_, _32372_, _07242_);
  nand _82047_ (_32374_, _32358_, _06375_);
  nor _82048_ (_32375_, _32374_, _32306_);
  or _82049_ (_32376_, _32375_, _06545_);
  or _82050_ (_32377_, _32376_, _32373_);
  and _82051_ (_32379_, _32377_, _32302_);
  or _82052_ (_32380_, _32379_, _06366_);
  and _82053_ (_32381_, _14363_, _07971_);
  or _82054_ (_32382_, _32299_, _09056_);
  or _82055_ (_32383_, _32382_, _32381_);
  and _82056_ (_32384_, _32383_, _09061_);
  and _82057_ (_32385_, _32384_, _32380_);
  and _82058_ (_32386_, _32369_, _06528_);
  or _82059_ (_32387_, _32386_, _06568_);
  or _82060_ (_32388_, _32387_, _32385_);
  or _82061_ (_32390_, _32307_, _06926_);
  and _82062_ (_32391_, _32390_, _32388_);
  or _82063_ (_32392_, _32391_, _05927_);
  or _82064_ (_32393_, _32299_, _05928_);
  and _82065_ (_32394_, _32393_, _32392_);
  or _82066_ (_32395_, _32394_, _06278_);
  or _82067_ (_32396_, _32307_, _06279_);
  and _82068_ (_32397_, _32396_, _01347_);
  and _82069_ (_32398_, _32397_, _32395_);
  or _82070_ (_43288_, _32398_, _32297_);
  and _82071_ (_32400_, _13388_, \oc8051_golden_model_1.P1 [1]);
  nor _82072_ (_32401_, _11261_, _13388_);
  or _82073_ (_32402_, _32401_, _32400_);
  or _82074_ (_32403_, _32402_, _09061_);
  nand _82075_ (_32404_, _07971_, _07038_);
  or _82076_ (_32405_, _07971_, \oc8051_golden_model_1.P1 [1]);
  and _82077_ (_32406_, _32405_, _06218_);
  and _82078_ (_32407_, _32406_, _32404_);
  nor _82079_ (_32408_, _13388_, _07357_);
  or _82080_ (_32409_, _32408_, _32400_);
  or _82081_ (_32411_, _32409_, _07166_);
  and _82082_ (_32412_, _14562_, _07971_);
  not _82083_ (_32413_, _32412_);
  and _82084_ (_32414_, _32413_, _32405_);
  or _82085_ (_32415_, _32414_, _07151_);
  and _82086_ (_32416_, _07971_, \oc8051_golden_model_1.ACC [1]);
  or _82087_ (_32417_, _32416_, _32400_);
  and _82088_ (_32418_, _32417_, _07141_);
  and _82089_ (_32419_, _07142_, \oc8051_golden_model_1.P1 [1]);
  or _82090_ (_32420_, _32419_, _06341_);
  or _82091_ (_32422_, _32420_, _32418_);
  and _82092_ (_32423_, _32422_, _06273_);
  and _82093_ (_32424_, _32423_, _32415_);
  and _82094_ (_32425_, _13396_, \oc8051_golden_model_1.P1 [1]);
  and _82095_ (_32426_, _14557_, _08620_);
  or _82096_ (_32427_, _32426_, _32425_);
  and _82097_ (_32428_, _32427_, _06272_);
  or _82098_ (_32429_, _32428_, _06461_);
  or _82099_ (_32430_, _32429_, _32424_);
  and _82100_ (_32431_, _32430_, _32411_);
  or _82101_ (_32433_, _32431_, _06464_);
  or _82102_ (_32434_, _32417_, _06465_);
  and _82103_ (_32435_, _32434_, _06269_);
  and _82104_ (_32436_, _32435_, _32433_);
  and _82105_ (_32437_, _14560_, _08620_);
  or _82106_ (_32438_, _32437_, _32425_);
  and _82107_ (_32439_, _32438_, _06268_);
  or _82108_ (_32440_, _32439_, _06261_);
  or _82109_ (_32441_, _32440_, _32436_);
  and _82110_ (_32442_, _32426_, _14556_);
  or _82111_ (_32444_, _32425_, _06262_);
  or _82112_ (_32445_, _32444_, _32442_);
  and _82113_ (_32446_, _32445_, _06258_);
  and _82114_ (_32447_, _32446_, _32441_);
  or _82115_ (_32448_, _32425_, _14597_);
  and _82116_ (_32449_, _32448_, _06257_);
  and _82117_ (_32450_, _32449_, _32427_);
  or _82118_ (_32451_, _32450_, _10080_);
  or _82119_ (_32452_, _32451_, _32447_);
  or _82120_ (_32453_, _32409_, _07215_);
  and _82121_ (_32455_, _32453_, _32452_);
  or _82122_ (_32456_, _32455_, _07460_);
  and _82123_ (_32457_, _09451_, _07971_);
  or _82124_ (_32458_, _32400_, _07208_);
  or _82125_ (_32459_, _32458_, _32457_);
  and _82126_ (_32460_, _32459_, _05982_);
  and _82127_ (_32461_, _32460_, _32456_);
  and _82128_ (_32462_, _14653_, _07971_);
  or _82129_ (_32463_, _32462_, _32400_);
  and _82130_ (_32464_, _32463_, _10094_);
  or _82131_ (_32466_, _32464_, _32461_);
  and _82132_ (_32467_, _32466_, _06219_);
  or _82133_ (_32468_, _32467_, _32407_);
  and _82134_ (_32469_, _32468_, _07237_);
  or _82135_ (_32470_, _14668_, _13388_);
  and _82136_ (_32471_, _32405_, _06369_);
  and _82137_ (_32472_, _32471_, _32470_);
  or _82138_ (_32473_, _32472_, _06536_);
  or _82139_ (_32474_, _32473_, _32469_);
  and _82140_ (_32475_, _11262_, _07971_);
  or _82141_ (_32476_, _32475_, _32400_);
  or _82142_ (_32477_, _32476_, _07240_);
  and _82143_ (_32478_, _32477_, _07242_);
  and _82144_ (_32479_, _32478_, _32474_);
  or _82145_ (_32480_, _14666_, _13388_);
  and _82146_ (_32481_, _32405_, _06375_);
  and _82147_ (_32482_, _32481_, _32480_);
  or _82148_ (_32483_, _32482_, _06545_);
  or _82149_ (_32484_, _32483_, _32479_);
  and _82150_ (_32485_, _32416_, _08341_);
  or _82151_ (_32487_, _32400_, _07234_);
  or _82152_ (_32488_, _32487_, _32485_);
  and _82153_ (_32489_, _32488_, _09056_);
  and _82154_ (_32490_, _32489_, _32484_);
  or _82155_ (_32491_, _32404_, _08341_);
  and _82156_ (_32492_, _32405_, _06366_);
  and _82157_ (_32493_, _32492_, _32491_);
  or _82158_ (_32494_, _32493_, _06528_);
  or _82159_ (_32495_, _32494_, _32490_);
  and _82160_ (_32496_, _32495_, _32403_);
  or _82161_ (_32498_, _32496_, _06568_);
  or _82162_ (_32499_, _32414_, _06926_);
  and _82163_ (_32500_, _32499_, _05928_);
  and _82164_ (_32501_, _32500_, _32498_);
  and _82165_ (_32502_, _32438_, _05927_);
  or _82166_ (_32503_, _32502_, _06278_);
  or _82167_ (_32504_, _32503_, _32501_);
  or _82168_ (_32505_, _32400_, _06279_);
  or _82169_ (_32506_, _32505_, _32412_);
  and _82170_ (_32507_, _32506_, _01347_);
  and _82171_ (_32509_, _32507_, _32504_);
  nor _82172_ (_32510_, \oc8051_golden_model_1.P1 [1], rst);
  nor _82173_ (_32511_, _32510_, _01354_);
  or _82174_ (_43289_, _32511_, _32509_);
  nor _82175_ (_32512_, \oc8051_golden_model_1.P1 [2], rst);
  nor _82176_ (_32513_, _32512_, _01354_);
  and _82177_ (_32514_, _13388_, \oc8051_golden_model_1.P1 [2]);
  nor _82178_ (_32515_, _13388_, _07776_);
  or _82179_ (_32516_, _32515_, _32514_);
  or _82180_ (_32517_, _32516_, _07215_);
  or _82181_ (_32519_, _32516_, _07166_);
  and _82182_ (_32520_, _14770_, _07971_);
  or _82183_ (_32521_, _32520_, _32514_);
  or _82184_ (_32522_, _32521_, _07151_);
  and _82185_ (_32523_, _07971_, \oc8051_golden_model_1.ACC [2]);
  or _82186_ (_32524_, _32523_, _32514_);
  and _82187_ (_32525_, _32524_, _07141_);
  and _82188_ (_32526_, _07142_, \oc8051_golden_model_1.P1 [2]);
  or _82189_ (_32527_, _32526_, _06341_);
  or _82190_ (_32528_, _32527_, _32525_);
  and _82191_ (_32530_, _32528_, _06273_);
  and _82192_ (_32531_, _32530_, _32522_);
  and _82193_ (_32532_, _13396_, \oc8051_golden_model_1.P1 [2]);
  and _82194_ (_32533_, _14774_, _08620_);
  or _82195_ (_32534_, _32533_, _32532_);
  and _82196_ (_32535_, _32534_, _06272_);
  or _82197_ (_32536_, _32535_, _06461_);
  or _82198_ (_32537_, _32536_, _32531_);
  and _82199_ (_32538_, _32537_, _32519_);
  or _82200_ (_32539_, _32538_, _06464_);
  or _82201_ (_32541_, _32524_, _06465_);
  and _82202_ (_32542_, _32541_, _06269_);
  and _82203_ (_32543_, _32542_, _32539_);
  and _82204_ (_32544_, _14756_, _08620_);
  or _82205_ (_32545_, _32544_, _32532_);
  and _82206_ (_32546_, _32545_, _06268_);
  or _82207_ (_32547_, _32546_, _06261_);
  or _82208_ (_32548_, _32547_, _32543_);
  and _82209_ (_32549_, _32533_, _14789_);
  or _82210_ (_32550_, _32532_, _06262_);
  or _82211_ (_32552_, _32550_, _32549_);
  and _82212_ (_32553_, _32552_, _06258_);
  and _82213_ (_32554_, _32553_, _32548_);
  and _82214_ (_32555_, _14804_, _08620_);
  or _82215_ (_32556_, _32555_, _32532_);
  and _82216_ (_32557_, _32556_, _06257_);
  or _82217_ (_32558_, _32557_, _10080_);
  or _82218_ (_32559_, _32558_, _32554_);
  and _82219_ (_32560_, _32559_, _32517_);
  or _82220_ (_32561_, _32560_, _07460_);
  and _82221_ (_32563_, _09450_, _07971_);
  or _82222_ (_32564_, _32514_, _07208_);
  or _82223_ (_32565_, _32564_, _32563_);
  and _82224_ (_32566_, _32565_, _05982_);
  and _82225_ (_32567_, _32566_, _32561_);
  and _82226_ (_32568_, _14859_, _07971_);
  or _82227_ (_32569_, _32568_, _32514_);
  and _82228_ (_32570_, _32569_, _10094_);
  or _82229_ (_32571_, _32570_, _06218_);
  or _82230_ (_32572_, _32571_, _32567_);
  and _82231_ (_32574_, _07971_, _08973_);
  or _82232_ (_32575_, _32574_, _32514_);
  or _82233_ (_32576_, _32575_, _06219_);
  and _82234_ (_32577_, _32576_, _32572_);
  or _82235_ (_32578_, _32577_, _06369_);
  and _82236_ (_32579_, _14751_, _07971_);
  or _82237_ (_32580_, _32579_, _32514_);
  or _82238_ (_32581_, _32580_, _07237_);
  and _82239_ (_32582_, _32581_, _07240_);
  and _82240_ (_32583_, _32582_, _32578_);
  and _82241_ (_32585_, _11259_, _07971_);
  or _82242_ (_32586_, _32585_, _32514_);
  and _82243_ (_32587_, _32586_, _06536_);
  or _82244_ (_32588_, _32587_, _32583_);
  and _82245_ (_32589_, _32588_, _07242_);
  or _82246_ (_32590_, _32514_, _08440_);
  and _82247_ (_32591_, _32575_, _06375_);
  and _82248_ (_32592_, _32591_, _32590_);
  or _82249_ (_32593_, _32592_, _32589_);
  and _82250_ (_32594_, _32593_, _07234_);
  and _82251_ (_32596_, _32524_, _06545_);
  and _82252_ (_32597_, _32596_, _32590_);
  or _82253_ (_32598_, _32597_, _06366_);
  or _82254_ (_32599_, _32598_, _32594_);
  and _82255_ (_32600_, _14748_, _07971_);
  or _82256_ (_32601_, _32514_, _09056_);
  or _82257_ (_32602_, _32601_, _32600_);
  and _82258_ (_32603_, _32602_, _09061_);
  and _82259_ (_32604_, _32603_, _32599_);
  nor _82260_ (_32605_, _11258_, _13388_);
  or _82261_ (_32607_, _32605_, _32514_);
  and _82262_ (_32608_, _32607_, _06528_);
  or _82263_ (_32609_, _32608_, _06568_);
  or _82264_ (_32610_, _32609_, _32604_);
  or _82265_ (_32611_, _32521_, _06926_);
  and _82266_ (_32612_, _32611_, _05928_);
  and _82267_ (_32613_, _32612_, _32610_);
  and _82268_ (_32614_, _32545_, _05927_);
  or _82269_ (_32615_, _32614_, _06278_);
  or _82270_ (_32616_, _32615_, _32613_);
  and _82271_ (_32618_, _14926_, _07971_);
  or _82272_ (_32619_, _32514_, _06279_);
  or _82273_ (_32620_, _32619_, _32618_);
  and _82274_ (_32621_, _32620_, _01347_);
  and _82275_ (_32622_, _32621_, _32616_);
  or _82276_ (_43290_, _32622_, _32513_);
  and _82277_ (_32623_, _13388_, \oc8051_golden_model_1.P1 [3]);
  nor _82278_ (_32624_, _13388_, _07594_);
  or _82279_ (_32625_, _32624_, _32623_);
  or _82280_ (_32626_, _32625_, _07215_);
  and _82281_ (_32628_, _14953_, _07971_);
  or _82282_ (_32629_, _32628_, _32623_);
  or _82283_ (_32630_, _32629_, _07151_);
  and _82284_ (_32631_, _07971_, \oc8051_golden_model_1.ACC [3]);
  or _82285_ (_32632_, _32631_, _32623_);
  and _82286_ (_32633_, _32632_, _07141_);
  and _82287_ (_32634_, _07142_, \oc8051_golden_model_1.P1 [3]);
  or _82288_ (_32635_, _32634_, _06341_);
  or _82289_ (_32636_, _32635_, _32633_);
  and _82290_ (_32637_, _32636_, _06273_);
  and _82291_ (_32639_, _32637_, _32630_);
  and _82292_ (_32640_, _13396_, \oc8051_golden_model_1.P1 [3]);
  and _82293_ (_32641_, _14950_, _08620_);
  or _82294_ (_32642_, _32641_, _32640_);
  and _82295_ (_32643_, _32642_, _06272_);
  or _82296_ (_32644_, _32643_, _06461_);
  or _82297_ (_32645_, _32644_, _32639_);
  or _82298_ (_32646_, _32625_, _07166_);
  and _82299_ (_32647_, _32646_, _32645_);
  or _82300_ (_32648_, _32647_, _06464_);
  or _82301_ (_32650_, _32632_, _06465_);
  and _82302_ (_32651_, _32650_, _06269_);
  and _82303_ (_32652_, _32651_, _32648_);
  and _82304_ (_32653_, _14948_, _08620_);
  or _82305_ (_32654_, _32653_, _32640_);
  and _82306_ (_32655_, _32654_, _06268_);
  or _82307_ (_32656_, _32655_, _06261_);
  or _82308_ (_32657_, _32656_, _32652_);
  or _82309_ (_32658_, _32640_, _14979_);
  and _82310_ (_32659_, _32658_, _32642_);
  or _82311_ (_32661_, _32659_, _06262_);
  and _82312_ (_32662_, _32661_, _06258_);
  and _82313_ (_32663_, _32662_, _32657_);
  or _82314_ (_32664_, _32640_, _14992_);
  and _82315_ (_32665_, _32664_, _06257_);
  and _82316_ (_32666_, _32665_, _32642_);
  or _82317_ (_32667_, _32666_, _10080_);
  or _82318_ (_32668_, _32667_, _32663_);
  and _82319_ (_32669_, _32668_, _32626_);
  or _82320_ (_32670_, _32669_, _07460_);
  and _82321_ (_32672_, _09449_, _07971_);
  or _82322_ (_32673_, _32623_, _07208_);
  or _82323_ (_32674_, _32673_, _32672_);
  and _82324_ (_32675_, _32674_, _05982_);
  and _82325_ (_32676_, _32675_, _32670_);
  and _82326_ (_32677_, _15048_, _07971_);
  or _82327_ (_32678_, _32677_, _32623_);
  and _82328_ (_32679_, _32678_, _10094_);
  or _82329_ (_32680_, _32679_, _06218_);
  or _82330_ (_32681_, _32680_, _32676_);
  and _82331_ (_32683_, _07971_, _08930_);
  or _82332_ (_32684_, _32683_, _32623_);
  or _82333_ (_32685_, _32684_, _06219_);
  and _82334_ (_32686_, _32685_, _32681_);
  or _82335_ (_32687_, _32686_, _06369_);
  and _82336_ (_32688_, _14943_, _07971_);
  or _82337_ (_32689_, _32688_, _32623_);
  or _82338_ (_32690_, _32689_, _07237_);
  and _82339_ (_32691_, _32690_, _07240_);
  and _82340_ (_32692_, _32691_, _32687_);
  and _82341_ (_32694_, _12577_, _07971_);
  or _82342_ (_32695_, _32694_, _32623_);
  and _82343_ (_32696_, _32695_, _06536_);
  or _82344_ (_32697_, _32696_, _32692_);
  and _82345_ (_32698_, _32697_, _07242_);
  or _82346_ (_32699_, _32623_, _08292_);
  and _82347_ (_32700_, _32684_, _06375_);
  and _82348_ (_32701_, _32700_, _32699_);
  or _82349_ (_32702_, _32701_, _32698_);
  and _82350_ (_32703_, _32702_, _07234_);
  and _82351_ (_32705_, _32632_, _06545_);
  and _82352_ (_32706_, _32705_, _32699_);
  or _82353_ (_32707_, _32706_, _06366_);
  or _82354_ (_32708_, _32707_, _32703_);
  and _82355_ (_32709_, _14940_, _07971_);
  or _82356_ (_32710_, _32623_, _09056_);
  or _82357_ (_32711_, _32710_, _32709_);
  and _82358_ (_32712_, _32711_, _09061_);
  and _82359_ (_32713_, _32712_, _32708_);
  nor _82360_ (_32714_, _11256_, _13388_);
  or _82361_ (_32716_, _32714_, _32623_);
  and _82362_ (_32717_, _32716_, _06528_);
  or _82363_ (_32718_, _32717_, _06568_);
  or _82364_ (_32719_, _32718_, _32713_);
  or _82365_ (_32720_, _32629_, _06926_);
  and _82366_ (_32721_, _32720_, _05928_);
  and _82367_ (_32722_, _32721_, _32719_);
  and _82368_ (_32723_, _32654_, _05927_);
  or _82369_ (_32724_, _32723_, _06278_);
  or _82370_ (_32725_, _32724_, _32722_);
  and _82371_ (_32727_, _15128_, _07971_);
  or _82372_ (_32728_, _32623_, _06279_);
  or _82373_ (_32729_, _32728_, _32727_);
  and _82374_ (_32730_, _32729_, _01347_);
  and _82375_ (_32731_, _32730_, _32725_);
  nor _82376_ (_32732_, \oc8051_golden_model_1.P1 [3], rst);
  nor _82377_ (_32733_, _32732_, _01354_);
  or _82378_ (_43291_, _32733_, _32731_);
  nor _82379_ (_32734_, \oc8051_golden_model_1.P1 [4], rst);
  nor _82380_ (_32735_, _32734_, _01354_);
  and _82381_ (_32737_, _13388_, \oc8051_golden_model_1.P1 [4]);
  nor _82382_ (_32738_, _08541_, _13388_);
  or _82383_ (_32739_, _32738_, _32737_);
  or _82384_ (_32740_, _32739_, _07215_);
  and _82385_ (_32741_, _13396_, \oc8051_golden_model_1.P1 [4]);
  and _82386_ (_32742_, _15176_, _08620_);
  or _82387_ (_32743_, _32742_, _32741_);
  and _82388_ (_32744_, _32743_, _06268_);
  and _82389_ (_32745_, _15162_, _07971_);
  or _82390_ (_32746_, _32745_, _32737_);
  or _82391_ (_32748_, _32746_, _07151_);
  and _82392_ (_32749_, _07971_, \oc8051_golden_model_1.ACC [4]);
  or _82393_ (_32750_, _32749_, _32737_);
  and _82394_ (_32751_, _32750_, _07141_);
  and _82395_ (_32752_, _07142_, \oc8051_golden_model_1.P1 [4]);
  or _82396_ (_32753_, _32752_, _06341_);
  or _82397_ (_32754_, _32753_, _32751_);
  and _82398_ (_32755_, _32754_, _06273_);
  and _82399_ (_32756_, _32755_, _32748_);
  and _82400_ (_32757_, _15166_, _08620_);
  or _82401_ (_32759_, _32757_, _32741_);
  and _82402_ (_32760_, _32759_, _06272_);
  or _82403_ (_32761_, _32760_, _06461_);
  or _82404_ (_32762_, _32761_, _32756_);
  or _82405_ (_32763_, _32739_, _07166_);
  and _82406_ (_32764_, _32763_, _32762_);
  or _82407_ (_32765_, _32764_, _06464_);
  or _82408_ (_32766_, _32750_, _06465_);
  and _82409_ (_32767_, _32766_, _06269_);
  and _82410_ (_32768_, _32767_, _32765_);
  or _82411_ (_32770_, _32768_, _32744_);
  and _82412_ (_32771_, _32770_, _06262_);
  and _82413_ (_32772_, _15184_, _08620_);
  or _82414_ (_32773_, _32772_, _32741_);
  and _82415_ (_32774_, _32773_, _06261_);
  or _82416_ (_32775_, _32774_, _32771_);
  and _82417_ (_32776_, _32775_, _06258_);
  and _82418_ (_32777_, _15200_, _08620_);
  or _82419_ (_32778_, _32777_, _32741_);
  and _82420_ (_32779_, _32778_, _06257_);
  or _82421_ (_32781_, _32779_, _10080_);
  or _82422_ (_32782_, _32781_, _32776_);
  and _82423_ (_32783_, _32782_, _32740_);
  or _82424_ (_32784_, _32783_, _07460_);
  and _82425_ (_32785_, _09448_, _07971_);
  or _82426_ (_32786_, _32737_, _07208_);
  or _82427_ (_32787_, _32786_, _32785_);
  and _82428_ (_32788_, _32787_, _05982_);
  and _82429_ (_32789_, _32788_, _32784_);
  and _82430_ (_32790_, _15254_, _07971_);
  or _82431_ (_32792_, _32790_, _32737_);
  and _82432_ (_32793_, _32792_, _10094_);
  or _82433_ (_32794_, _32793_, _06218_);
  or _82434_ (_32795_, _32794_, _32789_);
  and _82435_ (_32796_, _08959_, _07971_);
  or _82436_ (_32797_, _32796_, _32737_);
  or _82437_ (_32798_, _32797_, _06219_);
  and _82438_ (_32799_, _32798_, _32795_);
  or _82439_ (_32800_, _32799_, _06369_);
  and _82440_ (_32801_, _15269_, _07971_);
  or _82441_ (_32803_, _32801_, _32737_);
  or _82442_ (_32804_, _32803_, _07237_);
  and _82443_ (_32805_, _32804_, _07240_);
  and _82444_ (_32806_, _32805_, _32800_);
  and _82445_ (_32807_, _11254_, _07971_);
  or _82446_ (_32808_, _32807_, _32737_);
  and _82447_ (_32809_, _32808_, _06536_);
  or _82448_ (_32810_, _32809_, _32806_);
  and _82449_ (_32811_, _32810_, _07242_);
  or _82450_ (_32812_, _32737_, _08544_);
  and _82451_ (_32814_, _32797_, _06375_);
  and _82452_ (_32815_, _32814_, _32812_);
  or _82453_ (_32816_, _32815_, _32811_);
  and _82454_ (_32817_, _32816_, _07234_);
  and _82455_ (_32818_, _32750_, _06545_);
  and _82456_ (_32819_, _32818_, _32812_);
  or _82457_ (_32820_, _32819_, _06366_);
  or _82458_ (_32821_, _32820_, _32817_);
  and _82459_ (_32822_, _15266_, _07971_);
  or _82460_ (_32823_, _32737_, _09056_);
  or _82461_ (_32825_, _32823_, _32822_);
  and _82462_ (_32826_, _32825_, _09061_);
  and _82463_ (_32827_, _32826_, _32821_);
  nor _82464_ (_32828_, _11253_, _13388_);
  or _82465_ (_32829_, _32828_, _32737_);
  and _82466_ (_32830_, _32829_, _06528_);
  or _82467_ (_32831_, _32830_, _06568_);
  or _82468_ (_32832_, _32831_, _32827_);
  or _82469_ (_32833_, _32746_, _06926_);
  and _82470_ (_32834_, _32833_, _05928_);
  and _82471_ (_32836_, _32834_, _32832_);
  and _82472_ (_32837_, _32743_, _05927_);
  or _82473_ (_32838_, _32837_, _06278_);
  or _82474_ (_32839_, _32838_, _32836_);
  and _82475_ (_32840_, _15329_, _07971_);
  or _82476_ (_32841_, _32737_, _06279_);
  or _82477_ (_32842_, _32841_, _32840_);
  and _82478_ (_32843_, _32842_, _01347_);
  and _82479_ (_32844_, _32843_, _32839_);
  or _82480_ (_43292_, _32844_, _32735_);
  and _82481_ (_32846_, _13388_, \oc8051_golden_model_1.P1 [5]);
  and _82482_ (_32847_, _15358_, _07971_);
  or _82483_ (_32848_, _32847_, _32846_);
  or _82484_ (_32849_, _32848_, _07151_);
  and _82485_ (_32850_, _07971_, \oc8051_golden_model_1.ACC [5]);
  or _82486_ (_32851_, _32850_, _32846_);
  and _82487_ (_32852_, _32851_, _07141_);
  and _82488_ (_32853_, _07142_, \oc8051_golden_model_1.P1 [5]);
  or _82489_ (_32854_, _32853_, _06341_);
  or _82490_ (_32855_, _32854_, _32852_);
  and _82491_ (_32857_, _32855_, _06273_);
  and _82492_ (_32858_, _32857_, _32849_);
  and _82493_ (_32859_, _13396_, \oc8051_golden_model_1.P1 [5]);
  and _82494_ (_32860_, _15372_, _08620_);
  or _82495_ (_32861_, _32860_, _32859_);
  and _82496_ (_32862_, _32861_, _06272_);
  or _82497_ (_32863_, _32862_, _06461_);
  or _82498_ (_32864_, _32863_, _32858_);
  nor _82499_ (_32865_, _08244_, _13388_);
  or _82500_ (_32866_, _32865_, _32846_);
  or _82501_ (_32868_, _32866_, _07166_);
  and _82502_ (_32869_, _32868_, _32864_);
  or _82503_ (_32870_, _32869_, _06464_);
  or _82504_ (_32871_, _32851_, _06465_);
  and _82505_ (_32872_, _32871_, _06269_);
  and _82506_ (_32873_, _32872_, _32870_);
  and _82507_ (_32874_, _15355_, _08620_);
  or _82508_ (_32875_, _32874_, _32859_);
  and _82509_ (_32876_, _32875_, _06268_);
  or _82510_ (_32877_, _32876_, _06261_);
  or _82511_ (_32879_, _32877_, _32873_);
  or _82512_ (_32880_, _32859_, _15387_);
  and _82513_ (_32881_, _32880_, _32861_);
  or _82514_ (_32882_, _32881_, _06262_);
  and _82515_ (_32883_, _32882_, _06258_);
  and _82516_ (_32884_, _32883_, _32879_);
  or _82517_ (_32885_, _32859_, _15403_);
  and _82518_ (_32886_, _32885_, _06257_);
  and _82519_ (_32887_, _32886_, _32861_);
  or _82520_ (_32888_, _32887_, _10080_);
  or _82521_ (_32890_, _32888_, _32884_);
  or _82522_ (_32891_, _32866_, _07215_);
  and _82523_ (_32892_, _32891_, _32890_);
  or _82524_ (_32893_, _32892_, _07460_);
  and _82525_ (_32894_, _09447_, _07971_);
  or _82526_ (_32895_, _32846_, _07208_);
  or _82527_ (_32896_, _32895_, _32894_);
  and _82528_ (_32897_, _32896_, _05982_);
  and _82529_ (_32898_, _32897_, _32893_);
  and _82530_ (_32899_, _15459_, _07971_);
  or _82531_ (_32901_, _32899_, _32846_);
  and _82532_ (_32902_, _32901_, _10094_);
  or _82533_ (_32903_, _32902_, _06218_);
  or _82534_ (_32904_, _32903_, _32898_);
  and _82535_ (_32905_, _08946_, _07971_);
  or _82536_ (_32906_, _32905_, _32846_);
  or _82537_ (_32907_, _32906_, _06219_);
  and _82538_ (_32908_, _32907_, _32904_);
  or _82539_ (_32909_, _32908_, _06369_);
  and _82540_ (_32910_, _15353_, _07971_);
  or _82541_ (_32912_, _32910_, _32846_);
  or _82542_ (_32913_, _32912_, _07237_);
  and _82543_ (_32914_, _32913_, _07240_);
  and _82544_ (_32915_, _32914_, _32909_);
  and _82545_ (_32916_, _11250_, _07971_);
  or _82546_ (_32917_, _32916_, _32846_);
  and _82547_ (_32918_, _32917_, _06536_);
  or _82548_ (_32919_, _32918_, _32915_);
  and _82549_ (_32920_, _32919_, _07242_);
  or _82550_ (_32921_, _32846_, _08247_);
  and _82551_ (_32923_, _32906_, _06375_);
  and _82552_ (_32924_, _32923_, _32921_);
  or _82553_ (_32925_, _32924_, _32920_);
  and _82554_ (_32926_, _32925_, _07234_);
  and _82555_ (_32927_, _32851_, _06545_);
  and _82556_ (_32928_, _32927_, _32921_);
  or _82557_ (_32929_, _32928_, _06366_);
  or _82558_ (_32930_, _32929_, _32926_);
  and _82559_ (_32931_, _15350_, _07971_);
  or _82560_ (_32932_, _32846_, _09056_);
  or _82561_ (_32934_, _32932_, _32931_);
  and _82562_ (_32935_, _32934_, _09061_);
  and _82563_ (_32936_, _32935_, _32930_);
  nor _82564_ (_32937_, _11249_, _13388_);
  or _82565_ (_32938_, _32937_, _32846_);
  and _82566_ (_32939_, _32938_, _06528_);
  or _82567_ (_32940_, _32939_, _06568_);
  or _82568_ (_32941_, _32940_, _32936_);
  or _82569_ (_32942_, _32848_, _06926_);
  and _82570_ (_32943_, _32942_, _05928_);
  and _82571_ (_32945_, _32943_, _32941_);
  and _82572_ (_32946_, _32875_, _05927_);
  or _82573_ (_32947_, _32946_, _06278_);
  or _82574_ (_32948_, _32947_, _32945_);
  and _82575_ (_32949_, _15532_, _07971_);
  or _82576_ (_32950_, _32846_, _06279_);
  or _82577_ (_32951_, _32950_, _32949_);
  and _82578_ (_32952_, _32951_, _01347_);
  and _82579_ (_32953_, _32952_, _32948_);
  nor _82580_ (_32954_, \oc8051_golden_model_1.P1 [5], rst);
  nor _82581_ (_32956_, _32954_, _01354_);
  or _82582_ (_43293_, _32956_, _32953_);
  and _82583_ (_32957_, _13388_, \oc8051_golden_model_1.P1 [6]);
  and _82584_ (_32958_, _15554_, _07971_);
  or _82585_ (_32959_, _32958_, _32957_);
  or _82586_ (_32960_, _32959_, _07151_);
  and _82587_ (_32961_, _07971_, \oc8051_golden_model_1.ACC [6]);
  or _82588_ (_32962_, _32961_, _32957_);
  and _82589_ (_32963_, _32962_, _07141_);
  and _82590_ (_32964_, _07142_, \oc8051_golden_model_1.P1 [6]);
  or _82591_ (_32966_, _32964_, _06341_);
  or _82592_ (_32967_, _32966_, _32963_);
  and _82593_ (_32968_, _32967_, _06273_);
  and _82594_ (_32969_, _32968_, _32960_);
  and _82595_ (_32970_, _13396_, \oc8051_golden_model_1.P1 [6]);
  and _82596_ (_32971_, _15570_, _08620_);
  or _82597_ (_32972_, _32971_, _32970_);
  and _82598_ (_32973_, _32972_, _06272_);
  or _82599_ (_32974_, _32973_, _06461_);
  or _82600_ (_32975_, _32974_, _32969_);
  nor _82601_ (_32977_, _08142_, _13388_);
  or _82602_ (_32978_, _32977_, _32957_);
  or _82603_ (_32979_, _32978_, _07166_);
  and _82604_ (_32980_, _32979_, _32975_);
  or _82605_ (_32981_, _32980_, _06464_);
  or _82606_ (_32982_, _32962_, _06465_);
  and _82607_ (_32983_, _32982_, _06269_);
  and _82608_ (_32984_, _32983_, _32981_);
  and _82609_ (_32985_, _15551_, _08620_);
  or _82610_ (_32986_, _32985_, _32970_);
  and _82611_ (_32988_, _32986_, _06268_);
  or _82612_ (_32989_, _32988_, _06261_);
  or _82613_ (_32990_, _32989_, _32984_);
  or _82614_ (_32991_, _32970_, _15585_);
  and _82615_ (_32992_, _32991_, _32972_);
  or _82616_ (_32993_, _32992_, _06262_);
  and _82617_ (_32994_, _32993_, _06258_);
  and _82618_ (_32995_, _32994_, _32990_);
  and _82619_ (_32996_, _15602_, _08620_);
  or _82620_ (_32997_, _32996_, _32970_);
  and _82621_ (_32999_, _32997_, _06257_);
  or _82622_ (_33000_, _32999_, _10080_);
  or _82623_ (_33001_, _33000_, _32995_);
  or _82624_ (_33002_, _32978_, _07215_);
  and _82625_ (_33003_, _33002_, _33001_);
  or _82626_ (_33004_, _33003_, _07460_);
  and _82627_ (_33005_, _09446_, _07971_);
  or _82628_ (_33006_, _32957_, _07208_);
  or _82629_ (_33007_, _33006_, _33005_);
  and _82630_ (_33008_, _33007_, _05982_);
  and _82631_ (_33010_, _33008_, _33004_);
  and _82632_ (_33011_, _15657_, _07971_);
  or _82633_ (_33012_, _33011_, _32957_);
  and _82634_ (_33013_, _33012_, _10094_);
  or _82635_ (_33014_, _33013_, _06218_);
  or _82636_ (_33015_, _33014_, _33010_);
  and _82637_ (_33016_, _15664_, _07971_);
  or _82638_ (_33017_, _33016_, _32957_);
  or _82639_ (_33018_, _33017_, _06219_);
  and _82640_ (_33019_, _33018_, _33015_);
  or _82641_ (_33021_, _33019_, _06369_);
  and _82642_ (_33022_, _15549_, _07971_);
  or _82643_ (_33023_, _33022_, _32957_);
  or _82644_ (_33024_, _33023_, _07237_);
  and _82645_ (_33025_, _33024_, _07240_);
  and _82646_ (_33026_, _33025_, _33021_);
  and _82647_ (_33027_, _11247_, _07971_);
  or _82648_ (_33028_, _33027_, _32957_);
  and _82649_ (_33029_, _33028_, _06536_);
  or _82650_ (_33030_, _33029_, _33026_);
  and _82651_ (_33032_, _33030_, _07242_);
  or _82652_ (_33033_, _32957_, _08145_);
  and _82653_ (_33034_, _33017_, _06375_);
  and _82654_ (_33035_, _33034_, _33033_);
  or _82655_ (_33036_, _33035_, _33032_);
  and _82656_ (_33037_, _33036_, _07234_);
  and _82657_ (_33038_, _32962_, _06545_);
  and _82658_ (_33039_, _33038_, _33033_);
  or _82659_ (_33040_, _33039_, _06366_);
  or _82660_ (_33041_, _33040_, _33037_);
  and _82661_ (_33043_, _15546_, _07971_);
  or _82662_ (_33044_, _32957_, _09056_);
  or _82663_ (_33045_, _33044_, _33043_);
  and _82664_ (_33046_, _33045_, _09061_);
  and _82665_ (_33047_, _33046_, _33041_);
  nor _82666_ (_33048_, _11246_, _13388_);
  or _82667_ (_33049_, _33048_, _32957_);
  and _82668_ (_33050_, _33049_, _06528_);
  or _82669_ (_33051_, _33050_, _06568_);
  or _82670_ (_33052_, _33051_, _33047_);
  or _82671_ (_33054_, _32959_, _06926_);
  and _82672_ (_33055_, _33054_, _05928_);
  and _82673_ (_33056_, _33055_, _33052_);
  and _82674_ (_33057_, _32986_, _05927_);
  or _82675_ (_33058_, _33057_, _06278_);
  or _82676_ (_33059_, _33058_, _33056_);
  and _82677_ (_33060_, _15734_, _07971_);
  or _82678_ (_33061_, _32957_, _06279_);
  or _82679_ (_33062_, _33061_, _33060_);
  and _82680_ (_33063_, _33062_, _01347_);
  and _82681_ (_33065_, _33063_, _33059_);
  nor _82682_ (_33066_, \oc8051_golden_model_1.P1 [6], rst);
  nor _82683_ (_33067_, _33066_, _01354_);
  or _82684_ (_43294_, _33067_, _33065_);
  and _82685_ (_33068_, _01351_, \oc8051_golden_model_1.IP [0]);
  and _82686_ (_33069_, _07946_, \oc8051_golden_model_1.ACC [0]);
  and _82687_ (_33070_, _33069_, _08390_);
  and _82688_ (_33071_, _13490_, \oc8051_golden_model_1.IP [0]);
  or _82689_ (_33072_, _33071_, _07234_);
  or _82690_ (_33073_, _33072_, _33070_);
  and _82691_ (_33075_, _07946_, _07133_);
  or _82692_ (_33076_, _33075_, _33071_);
  or _82693_ (_33077_, _33076_, _07215_);
  nor _82694_ (_33078_, _08390_, _13490_);
  or _82695_ (_33079_, _33078_, _33071_);
  and _82696_ (_33080_, _33079_, _06341_);
  and _82697_ (_33081_, _07142_, \oc8051_golden_model_1.IP [0]);
  or _82698_ (_33082_, _33069_, _33071_);
  and _82699_ (_33083_, _33082_, _07141_);
  or _82700_ (_33084_, _33083_, _33081_);
  and _82701_ (_33086_, _33084_, _07151_);
  or _82702_ (_33087_, _33086_, _06272_);
  or _82703_ (_33088_, _33087_, _33080_);
  and _82704_ (_33089_, _14382_, _08632_);
  and _82705_ (_33090_, _13498_, \oc8051_golden_model_1.IP [0]);
  or _82706_ (_33091_, _33090_, _06273_);
  or _82707_ (_33092_, _33091_, _33089_);
  and _82708_ (_33093_, _33092_, _07166_);
  and _82709_ (_33094_, _33093_, _33088_);
  and _82710_ (_33095_, _33076_, _06461_);
  or _82711_ (_33097_, _33095_, _06464_);
  or _82712_ (_33098_, _33097_, _33094_);
  or _82713_ (_33099_, _33082_, _06465_);
  and _82714_ (_33100_, _33099_, _06269_);
  and _82715_ (_33101_, _33100_, _33098_);
  and _82716_ (_33102_, _33071_, _06268_);
  or _82717_ (_33103_, _33102_, _06261_);
  or _82718_ (_33104_, _33103_, _33101_);
  or _82719_ (_33105_, _33079_, _06262_);
  and _82720_ (_33106_, _33105_, _06258_);
  and _82721_ (_33108_, _33106_, _33104_);
  and _82722_ (_33109_, _14413_, _08632_);
  or _82723_ (_33110_, _33109_, _33090_);
  and _82724_ (_33111_, _33110_, _06257_);
  or _82725_ (_33112_, _33111_, _10080_);
  or _82726_ (_33113_, _33112_, _33108_);
  and _82727_ (_33114_, _33113_, _33077_);
  or _82728_ (_33115_, _33114_, _07460_);
  and _82729_ (_33116_, _09392_, _07946_);
  or _82730_ (_33117_, _33071_, _07208_);
  or _82731_ (_33119_, _33117_, _33116_);
  and _82732_ (_33120_, _33119_, _33115_);
  or _82733_ (_33121_, _33120_, _10094_);
  and _82734_ (_33122_, _14467_, _07946_);
  or _82735_ (_33123_, _33071_, _05982_);
  or _82736_ (_33124_, _33123_, _33122_);
  and _82737_ (_33125_, _33124_, _06219_);
  and _82738_ (_33126_, _33125_, _33121_);
  and _82739_ (_33127_, _07946_, _08954_);
  or _82740_ (_33128_, _33127_, _33071_);
  and _82741_ (_33130_, _33128_, _06218_);
  or _82742_ (_33131_, _33130_, _06369_);
  or _82743_ (_33132_, _33131_, _33126_);
  and _82744_ (_33133_, _14366_, _07946_);
  or _82745_ (_33134_, _33133_, _33071_);
  or _82746_ (_33135_, _33134_, _07237_);
  and _82747_ (_33136_, _33135_, _07240_);
  and _82748_ (_33137_, _33136_, _33132_);
  nor _82749_ (_33138_, _12580_, _13490_);
  or _82750_ (_33139_, _33138_, _33071_);
  nor _82751_ (_33141_, _33070_, _07240_);
  and _82752_ (_33142_, _33141_, _33139_);
  or _82753_ (_33143_, _33142_, _33137_);
  and _82754_ (_33144_, _33143_, _07242_);
  nand _82755_ (_33145_, _33128_, _06375_);
  nor _82756_ (_33146_, _33145_, _33078_);
  or _82757_ (_33147_, _33146_, _06545_);
  or _82758_ (_33148_, _33147_, _33144_);
  and _82759_ (_33149_, _33148_, _33073_);
  or _82760_ (_33150_, _33149_, _06366_);
  and _82761_ (_33152_, _14363_, _07946_);
  or _82762_ (_33153_, _33071_, _09056_);
  or _82763_ (_33154_, _33153_, _33152_);
  and _82764_ (_33155_, _33154_, _09061_);
  and _82765_ (_33156_, _33155_, _33150_);
  and _82766_ (_33157_, _33139_, _06528_);
  or _82767_ (_33158_, _33157_, _06568_);
  or _82768_ (_33159_, _33158_, _33156_);
  or _82769_ (_33160_, _33079_, _06926_);
  and _82770_ (_33161_, _33160_, _33159_);
  or _82771_ (_33163_, _33161_, _05927_);
  or _82772_ (_33164_, _33071_, _05928_);
  and _82773_ (_33165_, _33164_, _33163_);
  or _82774_ (_33166_, _33165_, _06278_);
  or _82775_ (_33167_, _33079_, _06279_);
  and _82776_ (_33168_, _33167_, _01347_);
  and _82777_ (_33169_, _33168_, _33166_);
  or _82778_ (_33170_, _33169_, _33068_);
  and _82779_ (_43296_, _33170_, _42618_);
  not _82780_ (_33171_, \oc8051_golden_model_1.IP [1]);
  nor _82781_ (_33173_, _01347_, _33171_);
  nor _82782_ (_33174_, _07946_, _33171_);
  nor _82783_ (_33175_, _11261_, _13490_);
  or _82784_ (_33176_, _33175_, _33174_);
  or _82785_ (_33177_, _33176_, _09061_);
  nand _82786_ (_33178_, _07946_, _07038_);
  or _82787_ (_33179_, _07946_, \oc8051_golden_model_1.IP [1]);
  and _82788_ (_33180_, _33179_, _06218_);
  and _82789_ (_33181_, _33180_, _33178_);
  nor _82790_ (_33182_, _13490_, _07357_);
  or _82791_ (_33184_, _33182_, _33174_);
  or _82792_ (_33185_, _33184_, _07166_);
  and _82793_ (_33186_, _14562_, _07946_);
  not _82794_ (_33187_, _33186_);
  and _82795_ (_33188_, _33187_, _33179_);
  or _82796_ (_33189_, _33188_, _07151_);
  and _82797_ (_33190_, _07946_, \oc8051_golden_model_1.ACC [1]);
  or _82798_ (_33191_, _33190_, _33174_);
  and _82799_ (_33192_, _33191_, _07141_);
  nor _82800_ (_33193_, _07141_, _33171_);
  or _82801_ (_33195_, _33193_, _06341_);
  or _82802_ (_33196_, _33195_, _33192_);
  and _82803_ (_33197_, _33196_, _06273_);
  and _82804_ (_33198_, _33197_, _33189_);
  nor _82805_ (_33199_, _08632_, _33171_);
  and _82806_ (_33200_, _14557_, _08632_);
  or _82807_ (_33201_, _33200_, _33199_);
  and _82808_ (_33202_, _33201_, _06272_);
  or _82809_ (_33203_, _33202_, _06461_);
  or _82810_ (_33204_, _33203_, _33198_);
  and _82811_ (_33206_, _33204_, _33185_);
  or _82812_ (_33207_, _33206_, _06464_);
  or _82813_ (_33208_, _33191_, _06465_);
  and _82814_ (_33209_, _33208_, _06269_);
  and _82815_ (_33210_, _33209_, _33207_);
  and _82816_ (_33211_, _14560_, _08632_);
  or _82817_ (_33212_, _33211_, _33199_);
  and _82818_ (_33213_, _33212_, _06268_);
  or _82819_ (_33214_, _33213_, _06261_);
  or _82820_ (_33215_, _33214_, _33210_);
  and _82821_ (_33216_, _33200_, _14556_);
  or _82822_ (_33217_, _33199_, _06262_);
  or _82823_ (_33218_, _33217_, _33216_);
  and _82824_ (_33219_, _33218_, _06258_);
  and _82825_ (_33220_, _33219_, _33215_);
  or _82826_ (_33221_, _33199_, _14597_);
  and _82827_ (_33222_, _33221_, _06257_);
  and _82828_ (_33223_, _33222_, _33201_);
  or _82829_ (_33224_, _33223_, _10080_);
  or _82830_ (_33225_, _33224_, _33220_);
  or _82831_ (_33227_, _33184_, _07215_);
  and _82832_ (_33228_, _33227_, _33225_);
  or _82833_ (_33229_, _33228_, _07460_);
  and _82834_ (_33230_, _09451_, _07946_);
  or _82835_ (_33231_, _33174_, _07208_);
  or _82836_ (_33232_, _33231_, _33230_);
  and _82837_ (_33233_, _33232_, _05982_);
  and _82838_ (_33234_, _33233_, _33229_);
  and _82839_ (_33235_, _14653_, _07946_);
  or _82840_ (_33236_, _33235_, _33174_);
  and _82841_ (_33238_, _33236_, _10094_);
  or _82842_ (_33239_, _33238_, _33234_);
  and _82843_ (_33240_, _33239_, _06219_);
  or _82844_ (_33241_, _33240_, _33181_);
  and _82845_ (_33242_, _33241_, _07237_);
  or _82846_ (_33243_, _14668_, _13490_);
  and _82847_ (_33244_, _33179_, _06369_);
  and _82848_ (_33245_, _33244_, _33243_);
  or _82849_ (_33246_, _33245_, _06536_);
  or _82850_ (_33247_, _33246_, _33242_);
  nand _82851_ (_33249_, _11260_, _07946_);
  and _82852_ (_33250_, _33249_, _33176_);
  or _82853_ (_33251_, _33250_, _07240_);
  and _82854_ (_33252_, _33251_, _07242_);
  and _82855_ (_33253_, _33252_, _33247_);
  or _82856_ (_33254_, _14666_, _13490_);
  and _82857_ (_33255_, _33179_, _06375_);
  and _82858_ (_33256_, _33255_, _33254_);
  or _82859_ (_33257_, _33256_, _06545_);
  or _82860_ (_33258_, _33257_, _33253_);
  nor _82861_ (_33260_, _33174_, _07234_);
  nand _82862_ (_33261_, _33260_, _33249_);
  and _82863_ (_33262_, _33261_, _09056_);
  and _82864_ (_33263_, _33262_, _33258_);
  or _82865_ (_33264_, _33178_, _08341_);
  and _82866_ (_33265_, _33179_, _06366_);
  and _82867_ (_33266_, _33265_, _33264_);
  or _82868_ (_33267_, _33266_, _06528_);
  or _82869_ (_33268_, _33267_, _33263_);
  and _82870_ (_33269_, _33268_, _33177_);
  or _82871_ (_33271_, _33269_, _06568_);
  or _82872_ (_33272_, _33188_, _06926_);
  and _82873_ (_33273_, _33272_, _05928_);
  and _82874_ (_33274_, _33273_, _33271_);
  and _82875_ (_33275_, _33212_, _05927_);
  or _82876_ (_33276_, _33275_, _06278_);
  or _82877_ (_33277_, _33276_, _33274_);
  or _82878_ (_33278_, _33174_, _06279_);
  or _82879_ (_33279_, _33278_, _33186_);
  and _82880_ (_33280_, _33279_, _01347_);
  and _82881_ (_33282_, _33280_, _33277_);
  or _82882_ (_33283_, _33282_, _33173_);
  and _82883_ (_43297_, _33283_, _42618_);
  and _82884_ (_33284_, _01351_, \oc8051_golden_model_1.IP [2]);
  and _82885_ (_33285_, _13490_, \oc8051_golden_model_1.IP [2]);
  nor _82886_ (_33286_, _13490_, _07776_);
  or _82887_ (_33287_, _33286_, _33285_);
  or _82888_ (_33288_, _33287_, _07215_);
  or _82889_ (_33289_, _33287_, _07166_);
  and _82890_ (_33290_, _14770_, _07946_);
  or _82891_ (_33292_, _33290_, _33285_);
  or _82892_ (_33293_, _33292_, _07151_);
  and _82893_ (_33294_, _07946_, \oc8051_golden_model_1.ACC [2]);
  or _82894_ (_33295_, _33294_, _33285_);
  and _82895_ (_33296_, _33295_, _07141_);
  and _82896_ (_33297_, _07142_, \oc8051_golden_model_1.IP [2]);
  or _82897_ (_33298_, _33297_, _06341_);
  or _82898_ (_33299_, _33298_, _33296_);
  and _82899_ (_33300_, _33299_, _06273_);
  and _82900_ (_33301_, _33300_, _33293_);
  and _82901_ (_33303_, _13498_, \oc8051_golden_model_1.IP [2]);
  and _82902_ (_33304_, _14774_, _08632_);
  or _82903_ (_33305_, _33304_, _33303_);
  and _82904_ (_33306_, _33305_, _06272_);
  or _82905_ (_33307_, _33306_, _06461_);
  or _82906_ (_33308_, _33307_, _33301_);
  and _82907_ (_33309_, _33308_, _33289_);
  or _82908_ (_33310_, _33309_, _06464_);
  or _82909_ (_33311_, _33295_, _06465_);
  and _82910_ (_33312_, _33311_, _06269_);
  and _82911_ (_33314_, _33312_, _33310_);
  and _82912_ (_33315_, _14756_, _08632_);
  or _82913_ (_33316_, _33315_, _33303_);
  and _82914_ (_33317_, _33316_, _06268_);
  or _82915_ (_33318_, _33317_, _06261_);
  or _82916_ (_33319_, _33318_, _33314_);
  and _82917_ (_33320_, _33304_, _14789_);
  or _82918_ (_33321_, _33303_, _06262_);
  or _82919_ (_33322_, _33321_, _33320_);
  and _82920_ (_33323_, _33322_, _06258_);
  and _82921_ (_33325_, _33323_, _33319_);
  and _82922_ (_33326_, _14804_, _08632_);
  or _82923_ (_33327_, _33326_, _33303_);
  and _82924_ (_33328_, _33327_, _06257_);
  or _82925_ (_33329_, _33328_, _10080_);
  or _82926_ (_33330_, _33329_, _33325_);
  and _82927_ (_33331_, _33330_, _33288_);
  or _82928_ (_33332_, _33331_, _07460_);
  and _82929_ (_33333_, _09450_, _07946_);
  or _82930_ (_33334_, _33285_, _07208_);
  or _82931_ (_33336_, _33334_, _33333_);
  and _82932_ (_33337_, _33336_, _05982_);
  and _82933_ (_33338_, _33337_, _33332_);
  and _82934_ (_33339_, _14859_, _07946_);
  or _82935_ (_33340_, _33339_, _33285_);
  and _82936_ (_33341_, _33340_, _10094_);
  or _82937_ (_33342_, _33341_, _06218_);
  or _82938_ (_33343_, _33342_, _33338_);
  and _82939_ (_33344_, _07946_, _08973_);
  or _82940_ (_33345_, _33344_, _33285_);
  or _82941_ (_33347_, _33345_, _06219_);
  and _82942_ (_33348_, _33347_, _33343_);
  or _82943_ (_33349_, _33348_, _06369_);
  and _82944_ (_33350_, _14751_, _07946_);
  or _82945_ (_33351_, _33350_, _33285_);
  or _82946_ (_33352_, _33351_, _07237_);
  and _82947_ (_33353_, _33352_, _07240_);
  and _82948_ (_33354_, _33353_, _33349_);
  and _82949_ (_33355_, _11259_, _07946_);
  or _82950_ (_33356_, _33355_, _33285_);
  and _82951_ (_33358_, _33356_, _06536_);
  or _82952_ (_33359_, _33358_, _33354_);
  and _82953_ (_33360_, _33359_, _07242_);
  or _82954_ (_33361_, _33285_, _08440_);
  and _82955_ (_33362_, _33345_, _06375_);
  and _82956_ (_33363_, _33362_, _33361_);
  or _82957_ (_33364_, _33363_, _33360_);
  and _82958_ (_33365_, _33364_, _07234_);
  and _82959_ (_33366_, _33295_, _06545_);
  and _82960_ (_33367_, _33366_, _33361_);
  or _82961_ (_33369_, _33367_, _06366_);
  or _82962_ (_33370_, _33369_, _33365_);
  and _82963_ (_33371_, _14748_, _07946_);
  or _82964_ (_33372_, _33285_, _09056_);
  or _82965_ (_33373_, _33372_, _33371_);
  and _82966_ (_33374_, _33373_, _09061_);
  and _82967_ (_33375_, _33374_, _33370_);
  nor _82968_ (_33376_, _11258_, _13490_);
  or _82969_ (_33377_, _33376_, _33285_);
  and _82970_ (_33378_, _33377_, _06528_);
  or _82971_ (_33380_, _33378_, _06568_);
  or _82972_ (_33381_, _33380_, _33375_);
  or _82973_ (_33382_, _33292_, _06926_);
  and _82974_ (_33383_, _33382_, _05928_);
  and _82975_ (_33384_, _33383_, _33381_);
  and _82976_ (_33385_, _33316_, _05927_);
  or _82977_ (_33386_, _33385_, _06278_);
  or _82978_ (_33387_, _33386_, _33384_);
  and _82979_ (_33388_, _14926_, _07946_);
  or _82980_ (_33389_, _33285_, _06279_);
  or _82981_ (_33391_, _33389_, _33388_);
  and _82982_ (_33392_, _33391_, _01347_);
  and _82983_ (_33393_, _33392_, _33387_);
  or _82984_ (_33394_, _33393_, _33284_);
  and _82985_ (_43298_, _33394_, _42618_);
  and _82986_ (_33395_, _01351_, \oc8051_golden_model_1.IP [3]);
  and _82987_ (_33396_, _13490_, \oc8051_golden_model_1.IP [3]);
  nor _82988_ (_33397_, _13490_, _07594_);
  or _82989_ (_33398_, _33397_, _33396_);
  or _82990_ (_33399_, _33398_, _07215_);
  and _82991_ (_33401_, _14953_, _07946_);
  or _82992_ (_33402_, _33401_, _33396_);
  or _82993_ (_33403_, _33402_, _07151_);
  and _82994_ (_33404_, _07946_, \oc8051_golden_model_1.ACC [3]);
  or _82995_ (_33405_, _33404_, _33396_);
  and _82996_ (_33406_, _33405_, _07141_);
  and _82997_ (_33407_, _07142_, \oc8051_golden_model_1.IP [3]);
  or _82998_ (_33408_, _33407_, _06341_);
  or _82999_ (_33409_, _33408_, _33406_);
  and _83000_ (_33410_, _33409_, _06273_);
  and _83001_ (_33412_, _33410_, _33403_);
  and _83002_ (_33413_, _13498_, \oc8051_golden_model_1.IP [3]);
  and _83003_ (_33414_, _14950_, _08632_);
  or _83004_ (_33415_, _33414_, _33413_);
  and _83005_ (_33416_, _33415_, _06272_);
  or _83006_ (_33417_, _33416_, _06461_);
  or _83007_ (_33418_, _33417_, _33412_);
  or _83008_ (_33419_, _33398_, _07166_);
  and _83009_ (_33420_, _33419_, _33418_);
  or _83010_ (_33421_, _33420_, _06464_);
  or _83011_ (_33423_, _33405_, _06465_);
  and _83012_ (_33424_, _33423_, _06269_);
  and _83013_ (_33425_, _33424_, _33421_);
  and _83014_ (_33426_, _14948_, _08632_);
  or _83015_ (_33427_, _33426_, _33413_);
  and _83016_ (_33428_, _33427_, _06268_);
  or _83017_ (_33429_, _33428_, _06261_);
  or _83018_ (_33430_, _33429_, _33425_);
  or _83019_ (_33431_, _33413_, _14979_);
  and _83020_ (_33432_, _33431_, _33415_);
  or _83021_ (_33434_, _33432_, _06262_);
  and _83022_ (_33435_, _33434_, _06258_);
  and _83023_ (_33436_, _33435_, _33430_);
  or _83024_ (_33437_, _33413_, _14992_);
  and _83025_ (_33438_, _33437_, _06257_);
  and _83026_ (_33439_, _33438_, _33415_);
  or _83027_ (_33440_, _33439_, _10080_);
  or _83028_ (_33441_, _33440_, _33436_);
  and _83029_ (_33442_, _33441_, _33399_);
  or _83030_ (_33443_, _33442_, _07460_);
  and _83031_ (_33445_, _09449_, _07946_);
  or _83032_ (_33446_, _33396_, _07208_);
  or _83033_ (_33447_, _33446_, _33445_);
  and _83034_ (_33448_, _33447_, _05982_);
  and _83035_ (_33449_, _33448_, _33443_);
  and _83036_ (_33450_, _15048_, _07946_);
  or _83037_ (_33451_, _33450_, _33396_);
  and _83038_ (_33452_, _33451_, _10094_);
  or _83039_ (_33453_, _33452_, _06218_);
  or _83040_ (_33454_, _33453_, _33449_);
  and _83041_ (_33456_, _07946_, _08930_);
  or _83042_ (_33457_, _33456_, _33396_);
  or _83043_ (_33458_, _33457_, _06219_);
  and _83044_ (_33459_, _33458_, _33454_);
  or _83045_ (_33460_, _33459_, _06369_);
  and _83046_ (_33461_, _14943_, _07946_);
  or _83047_ (_33462_, _33461_, _33396_);
  or _83048_ (_33463_, _33462_, _07237_);
  and _83049_ (_33464_, _33463_, _07240_);
  and _83050_ (_33465_, _33464_, _33460_);
  and _83051_ (_33467_, _12577_, _07946_);
  or _83052_ (_33468_, _33467_, _33396_);
  and _83053_ (_33469_, _33468_, _06536_);
  or _83054_ (_33470_, _33469_, _33465_);
  and _83055_ (_33471_, _33470_, _07242_);
  or _83056_ (_33472_, _33396_, _08292_);
  and _83057_ (_33473_, _33457_, _06375_);
  and _83058_ (_33474_, _33473_, _33472_);
  or _83059_ (_33475_, _33474_, _33471_);
  and _83060_ (_33476_, _33475_, _07234_);
  and _83061_ (_33478_, _33405_, _06545_);
  and _83062_ (_33479_, _33478_, _33472_);
  or _83063_ (_33480_, _33479_, _06366_);
  or _83064_ (_33481_, _33480_, _33476_);
  and _83065_ (_33482_, _14940_, _07946_);
  or _83066_ (_33483_, _33396_, _09056_);
  or _83067_ (_33484_, _33483_, _33482_);
  and _83068_ (_33485_, _33484_, _09061_);
  and _83069_ (_33486_, _33485_, _33481_);
  nor _83070_ (_33487_, _11256_, _13490_);
  or _83071_ (_33489_, _33487_, _33396_);
  and _83072_ (_33490_, _33489_, _06528_);
  or _83073_ (_33491_, _33490_, _06568_);
  or _83074_ (_33492_, _33491_, _33486_);
  or _83075_ (_33493_, _33402_, _06926_);
  and _83076_ (_33494_, _33493_, _05928_);
  and _83077_ (_33495_, _33494_, _33492_);
  and _83078_ (_33496_, _33427_, _05927_);
  or _83079_ (_33497_, _33496_, _06278_);
  or _83080_ (_33498_, _33497_, _33495_);
  and _83081_ (_33500_, _15128_, _07946_);
  or _83082_ (_33501_, _33396_, _06279_);
  or _83083_ (_33502_, _33501_, _33500_);
  and _83084_ (_33503_, _33502_, _01347_);
  and _83085_ (_33504_, _33503_, _33498_);
  or _83086_ (_33505_, _33504_, _33395_);
  and _83087_ (_43299_, _33505_, _42618_);
  and _83088_ (_33506_, _01351_, \oc8051_golden_model_1.IP [4]);
  and _83089_ (_33507_, _13490_, \oc8051_golden_model_1.IP [4]);
  nor _83090_ (_33508_, _08541_, _13490_);
  or _83091_ (_33510_, _33508_, _33507_);
  or _83092_ (_33511_, _33510_, _07215_);
  and _83093_ (_33512_, _13498_, \oc8051_golden_model_1.IP [4]);
  and _83094_ (_33513_, _15176_, _08632_);
  or _83095_ (_33514_, _33513_, _33512_);
  and _83096_ (_33515_, _33514_, _06268_);
  and _83097_ (_33516_, _15162_, _07946_);
  or _83098_ (_33517_, _33516_, _33507_);
  or _83099_ (_33518_, _33517_, _07151_);
  and _83100_ (_33519_, _07946_, \oc8051_golden_model_1.ACC [4]);
  or _83101_ (_33521_, _33519_, _33507_);
  and _83102_ (_33522_, _33521_, _07141_);
  and _83103_ (_33523_, _07142_, \oc8051_golden_model_1.IP [4]);
  or _83104_ (_33524_, _33523_, _06341_);
  or _83105_ (_33525_, _33524_, _33522_);
  and _83106_ (_33526_, _33525_, _06273_);
  and _83107_ (_33527_, _33526_, _33518_);
  and _83108_ (_33528_, _15166_, _08632_);
  or _83109_ (_33529_, _33528_, _33512_);
  and _83110_ (_33530_, _33529_, _06272_);
  or _83111_ (_33532_, _33530_, _06461_);
  or _83112_ (_33533_, _33532_, _33527_);
  or _83113_ (_33534_, _33510_, _07166_);
  and _83114_ (_33535_, _33534_, _33533_);
  or _83115_ (_33536_, _33535_, _06464_);
  or _83116_ (_33537_, _33521_, _06465_);
  and _83117_ (_33538_, _33537_, _06269_);
  and _83118_ (_33539_, _33538_, _33536_);
  or _83119_ (_33540_, _33539_, _33515_);
  and _83120_ (_33541_, _33540_, _06262_);
  or _83121_ (_33543_, _33512_, _15183_);
  and _83122_ (_33544_, _33543_, _06261_);
  and _83123_ (_33545_, _33544_, _33529_);
  or _83124_ (_33546_, _33545_, _33541_);
  and _83125_ (_33547_, _33546_, _06258_);
  and _83126_ (_33548_, _15200_, _08632_);
  or _83127_ (_33549_, _33548_, _33512_);
  and _83128_ (_33550_, _33549_, _06257_);
  or _83129_ (_33551_, _33550_, _10080_);
  or _83130_ (_33552_, _33551_, _33547_);
  and _83131_ (_33554_, _33552_, _33511_);
  or _83132_ (_33555_, _33554_, _07460_);
  and _83133_ (_33556_, _09448_, _07946_);
  or _83134_ (_33557_, _33507_, _07208_);
  or _83135_ (_33558_, _33557_, _33556_);
  and _83136_ (_33559_, _33558_, _05982_);
  and _83137_ (_33560_, _33559_, _33555_);
  and _83138_ (_33561_, _15254_, _07946_);
  or _83139_ (_33562_, _33561_, _33507_);
  and _83140_ (_33563_, _33562_, _10094_);
  or _83141_ (_33565_, _33563_, _06218_);
  or _83142_ (_33566_, _33565_, _33560_);
  and _83143_ (_33567_, _08959_, _07946_);
  or _83144_ (_33568_, _33567_, _33507_);
  or _83145_ (_33569_, _33568_, _06219_);
  and _83146_ (_33570_, _33569_, _33566_);
  or _83147_ (_33571_, _33570_, _06369_);
  and _83148_ (_33572_, _15269_, _07946_);
  or _83149_ (_33573_, _33572_, _33507_);
  or _83150_ (_33574_, _33573_, _07237_);
  and _83151_ (_33576_, _33574_, _07240_);
  and _83152_ (_33577_, _33576_, _33571_);
  and _83153_ (_33578_, _11254_, _07946_);
  or _83154_ (_33579_, _33578_, _33507_);
  and _83155_ (_33580_, _33579_, _06536_);
  or _83156_ (_33581_, _33580_, _33577_);
  and _83157_ (_33582_, _33581_, _07242_);
  or _83158_ (_33583_, _33507_, _08544_);
  and _83159_ (_33584_, _33568_, _06375_);
  and _83160_ (_33585_, _33584_, _33583_);
  or _83161_ (_33587_, _33585_, _33582_);
  and _83162_ (_33588_, _33587_, _07234_);
  and _83163_ (_33589_, _33521_, _06545_);
  and _83164_ (_33590_, _33589_, _33583_);
  or _83165_ (_33591_, _33590_, _06366_);
  or _83166_ (_33592_, _33591_, _33588_);
  and _83167_ (_33593_, _15266_, _07946_);
  or _83168_ (_33594_, _33507_, _09056_);
  or _83169_ (_33595_, _33594_, _33593_);
  and _83170_ (_33596_, _33595_, _09061_);
  and _83171_ (_33598_, _33596_, _33592_);
  nor _83172_ (_33599_, _11253_, _13490_);
  or _83173_ (_33600_, _33599_, _33507_);
  and _83174_ (_33601_, _33600_, _06528_);
  or _83175_ (_33602_, _33601_, _06568_);
  or _83176_ (_33603_, _33602_, _33598_);
  or _83177_ (_33604_, _33517_, _06926_);
  and _83178_ (_33605_, _33604_, _05928_);
  and _83179_ (_33606_, _33605_, _33603_);
  and _83180_ (_33607_, _33514_, _05927_);
  or _83181_ (_33609_, _33607_, _06278_);
  or _83182_ (_33610_, _33609_, _33606_);
  and _83183_ (_33611_, _15329_, _07946_);
  or _83184_ (_33612_, _33507_, _06279_);
  or _83185_ (_33613_, _33612_, _33611_);
  and _83186_ (_33614_, _33613_, _01347_);
  and _83187_ (_33615_, _33614_, _33610_);
  or _83188_ (_33616_, _33615_, _33506_);
  and _83189_ (_43300_, _33616_, _42618_);
  and _83190_ (_33617_, _01351_, \oc8051_golden_model_1.IP [5]);
  and _83191_ (_33619_, _13490_, \oc8051_golden_model_1.IP [5]);
  and _83192_ (_33620_, _15358_, _07946_);
  or _83193_ (_33621_, _33620_, _33619_);
  or _83194_ (_33622_, _33621_, _07151_);
  and _83195_ (_33623_, _07946_, \oc8051_golden_model_1.ACC [5]);
  or _83196_ (_33624_, _33623_, _33619_);
  and _83197_ (_33625_, _33624_, _07141_);
  and _83198_ (_33626_, _07142_, \oc8051_golden_model_1.IP [5]);
  or _83199_ (_33627_, _33626_, _06341_);
  or _83200_ (_33628_, _33627_, _33625_);
  and _83201_ (_33630_, _33628_, _06273_);
  and _83202_ (_33631_, _33630_, _33622_);
  and _83203_ (_33632_, _13498_, \oc8051_golden_model_1.IP [5]);
  and _83204_ (_33633_, _15372_, _08632_);
  or _83205_ (_33634_, _33633_, _33632_);
  and _83206_ (_33635_, _33634_, _06272_);
  or _83207_ (_33636_, _33635_, _06461_);
  or _83208_ (_33637_, _33636_, _33631_);
  nor _83209_ (_33638_, _08244_, _13490_);
  or _83210_ (_33639_, _33638_, _33619_);
  or _83211_ (_33641_, _33639_, _07166_);
  and _83212_ (_33642_, _33641_, _33637_);
  or _83213_ (_33643_, _33642_, _06464_);
  or _83214_ (_33644_, _33624_, _06465_);
  and _83215_ (_33645_, _33644_, _06269_);
  and _83216_ (_33646_, _33645_, _33643_);
  and _83217_ (_33647_, _15355_, _08632_);
  or _83218_ (_33648_, _33647_, _33632_);
  and _83219_ (_33649_, _33648_, _06268_);
  or _83220_ (_33650_, _33649_, _06261_);
  or _83221_ (_33652_, _33650_, _33646_);
  or _83222_ (_33653_, _33632_, _15387_);
  and _83223_ (_33654_, _33653_, _33634_);
  or _83224_ (_33655_, _33654_, _06262_);
  and _83225_ (_33656_, _33655_, _06258_);
  and _83226_ (_33657_, _33656_, _33652_);
  or _83227_ (_33658_, _33632_, _15403_);
  and _83228_ (_33659_, _33658_, _06257_);
  and _83229_ (_33660_, _33659_, _33634_);
  or _83230_ (_33661_, _33660_, _10080_);
  or _83231_ (_33663_, _33661_, _33657_);
  or _83232_ (_33664_, _33639_, _07215_);
  and _83233_ (_33665_, _33664_, _33663_);
  or _83234_ (_33666_, _33665_, _07460_);
  and _83235_ (_33667_, _09447_, _07946_);
  or _83236_ (_33668_, _33619_, _07208_);
  or _83237_ (_33669_, _33668_, _33667_);
  and _83238_ (_33670_, _33669_, _05982_);
  and _83239_ (_33671_, _33670_, _33666_);
  and _83240_ (_33672_, _15459_, _07946_);
  or _83241_ (_33674_, _33672_, _33619_);
  and _83242_ (_33675_, _33674_, _10094_);
  or _83243_ (_33676_, _33675_, _06218_);
  or _83244_ (_33677_, _33676_, _33671_);
  and _83245_ (_33678_, _08946_, _07946_);
  or _83246_ (_33679_, _33678_, _33619_);
  or _83247_ (_33680_, _33679_, _06219_);
  and _83248_ (_33681_, _33680_, _33677_);
  or _83249_ (_33682_, _33681_, _06369_);
  and _83250_ (_33683_, _15353_, _07946_);
  or _83251_ (_33685_, _33683_, _33619_);
  or _83252_ (_33686_, _33685_, _07237_);
  and _83253_ (_33687_, _33686_, _07240_);
  and _83254_ (_33688_, _33687_, _33682_);
  and _83255_ (_33689_, _11250_, _07946_);
  or _83256_ (_33690_, _33689_, _33619_);
  and _83257_ (_33691_, _33690_, _06536_);
  or _83258_ (_33692_, _33691_, _33688_);
  and _83259_ (_33693_, _33692_, _07242_);
  or _83260_ (_33694_, _33619_, _08247_);
  and _83261_ (_33696_, _33679_, _06375_);
  and _83262_ (_33697_, _33696_, _33694_);
  or _83263_ (_33698_, _33697_, _33693_);
  and _83264_ (_33699_, _33698_, _07234_);
  and _83265_ (_33700_, _33624_, _06545_);
  and _83266_ (_33701_, _33700_, _33694_);
  or _83267_ (_33702_, _33701_, _06366_);
  or _83268_ (_33703_, _33702_, _33699_);
  and _83269_ (_33704_, _15350_, _07946_);
  or _83270_ (_33705_, _33619_, _09056_);
  or _83271_ (_33707_, _33705_, _33704_);
  and _83272_ (_33708_, _33707_, _09061_);
  and _83273_ (_33709_, _33708_, _33703_);
  nor _83274_ (_33710_, _11249_, _13490_);
  or _83275_ (_33711_, _33710_, _33619_);
  and _83276_ (_33712_, _33711_, _06528_);
  or _83277_ (_33713_, _33712_, _06568_);
  or _83278_ (_33714_, _33713_, _33709_);
  or _83279_ (_33715_, _33621_, _06926_);
  and _83280_ (_33716_, _33715_, _05928_);
  and _83281_ (_33718_, _33716_, _33714_);
  and _83282_ (_33719_, _33648_, _05927_);
  or _83283_ (_33720_, _33719_, _06278_);
  or _83284_ (_33721_, _33720_, _33718_);
  and _83285_ (_33722_, _15532_, _07946_);
  or _83286_ (_33723_, _33619_, _06279_);
  or _83287_ (_33724_, _33723_, _33722_);
  and _83288_ (_33725_, _33724_, _01347_);
  and _83289_ (_33726_, _33725_, _33721_);
  or _83290_ (_33727_, _33726_, _33617_);
  and _83291_ (_43302_, _33727_, _42618_);
  and _83292_ (_33729_, _01351_, \oc8051_golden_model_1.IP [6]);
  and _83293_ (_33730_, _13490_, \oc8051_golden_model_1.IP [6]);
  and _83294_ (_33731_, _15554_, _07946_);
  or _83295_ (_33732_, _33731_, _33730_);
  or _83296_ (_33733_, _33732_, _07151_);
  and _83297_ (_33734_, _07946_, \oc8051_golden_model_1.ACC [6]);
  or _83298_ (_33735_, _33734_, _33730_);
  and _83299_ (_33736_, _33735_, _07141_);
  and _83300_ (_33737_, _07142_, \oc8051_golden_model_1.IP [6]);
  or _83301_ (_33739_, _33737_, _06341_);
  or _83302_ (_33740_, _33739_, _33736_);
  and _83303_ (_33741_, _33740_, _06273_);
  and _83304_ (_33742_, _33741_, _33733_);
  and _83305_ (_33743_, _13498_, \oc8051_golden_model_1.IP [6]);
  and _83306_ (_33744_, _15570_, _08632_);
  or _83307_ (_33745_, _33744_, _33743_);
  and _83308_ (_33746_, _33745_, _06272_);
  or _83309_ (_33747_, _33746_, _06461_);
  or _83310_ (_33748_, _33747_, _33742_);
  nor _83311_ (_33750_, _08142_, _13490_);
  or _83312_ (_33751_, _33750_, _33730_);
  or _83313_ (_33752_, _33751_, _07166_);
  and _83314_ (_33753_, _33752_, _33748_);
  or _83315_ (_33754_, _33753_, _06464_);
  or _83316_ (_33755_, _33735_, _06465_);
  and _83317_ (_33756_, _33755_, _06269_);
  and _83318_ (_33757_, _33756_, _33754_);
  and _83319_ (_33758_, _15551_, _08632_);
  or _83320_ (_33759_, _33758_, _33743_);
  and _83321_ (_33761_, _33759_, _06268_);
  or _83322_ (_33762_, _33761_, _06261_);
  or _83323_ (_33763_, _33762_, _33757_);
  or _83324_ (_33764_, _33743_, _15585_);
  and _83325_ (_33765_, _33764_, _33745_);
  or _83326_ (_33766_, _33765_, _06262_);
  and _83327_ (_33767_, _33766_, _06258_);
  and _83328_ (_33768_, _33767_, _33763_);
  and _83329_ (_33769_, _15602_, _08632_);
  or _83330_ (_33770_, _33769_, _33743_);
  and _83331_ (_33772_, _33770_, _06257_);
  or _83332_ (_33773_, _33772_, _10080_);
  or _83333_ (_33774_, _33773_, _33768_);
  or _83334_ (_33775_, _33751_, _07215_);
  and _83335_ (_33776_, _33775_, _33774_);
  or _83336_ (_33777_, _33776_, _07460_);
  and _83337_ (_33778_, _09446_, _07946_);
  or _83338_ (_33779_, _33730_, _07208_);
  or _83339_ (_33780_, _33779_, _33778_);
  and _83340_ (_33781_, _33780_, _05982_);
  and _83341_ (_33783_, _33781_, _33777_);
  and _83342_ (_33784_, _15657_, _07946_);
  or _83343_ (_33785_, _33784_, _33730_);
  and _83344_ (_33786_, _33785_, _10094_);
  or _83345_ (_33787_, _33786_, _06218_);
  or _83346_ (_33788_, _33787_, _33783_);
  and _83347_ (_33789_, _15664_, _07946_);
  or _83348_ (_33790_, _33789_, _33730_);
  or _83349_ (_33791_, _33790_, _06219_);
  and _83350_ (_33792_, _33791_, _33788_);
  or _83351_ (_33794_, _33792_, _06369_);
  and _83352_ (_33795_, _15549_, _07946_);
  or _83353_ (_33796_, _33795_, _33730_);
  or _83354_ (_33797_, _33796_, _07237_);
  and _83355_ (_33798_, _33797_, _07240_);
  and _83356_ (_33799_, _33798_, _33794_);
  and _83357_ (_33800_, _11247_, _07946_);
  or _83358_ (_33801_, _33800_, _33730_);
  and _83359_ (_33802_, _33801_, _06536_);
  or _83360_ (_33803_, _33802_, _33799_);
  and _83361_ (_33805_, _33803_, _07242_);
  or _83362_ (_33806_, _33730_, _08145_);
  and _83363_ (_33807_, _33790_, _06375_);
  and _83364_ (_33808_, _33807_, _33806_);
  or _83365_ (_33809_, _33808_, _33805_);
  and _83366_ (_33810_, _33809_, _07234_);
  and _83367_ (_33811_, _33735_, _06545_);
  and _83368_ (_33812_, _33811_, _33806_);
  or _83369_ (_33813_, _33812_, _06366_);
  or _83370_ (_33814_, _33813_, _33810_);
  and _83371_ (_33816_, _15546_, _07946_);
  or _83372_ (_33817_, _33730_, _09056_);
  or _83373_ (_33818_, _33817_, _33816_);
  and _83374_ (_33819_, _33818_, _09061_);
  and _83375_ (_33820_, _33819_, _33814_);
  nor _83376_ (_33821_, _11246_, _13490_);
  or _83377_ (_33822_, _33821_, _33730_);
  and _83378_ (_33823_, _33822_, _06528_);
  or _83379_ (_33824_, _33823_, _06568_);
  or _83380_ (_33825_, _33824_, _33820_);
  or _83381_ (_33827_, _33732_, _06926_);
  and _83382_ (_33828_, _33827_, _05928_);
  and _83383_ (_33829_, _33828_, _33825_);
  and _83384_ (_33830_, _33759_, _05927_);
  or _83385_ (_33831_, _33830_, _06278_);
  or _83386_ (_33832_, _33831_, _33829_);
  and _83387_ (_33833_, _15734_, _07946_);
  or _83388_ (_33834_, _33730_, _06279_);
  or _83389_ (_33835_, _33834_, _33833_);
  and _83390_ (_33836_, _33835_, _01347_);
  and _83391_ (_33838_, _33836_, _33832_);
  or _83392_ (_33839_, _33838_, _33729_);
  and _83393_ (_43303_, _33839_, _42618_);
  and _83394_ (_33840_, _01351_, \oc8051_golden_model_1.IE [0]);
  and _83395_ (_33841_, _07900_, \oc8051_golden_model_1.ACC [0]);
  and _83396_ (_33842_, _33841_, _08390_);
  and _83397_ (_33843_, _13593_, \oc8051_golden_model_1.IE [0]);
  or _83398_ (_33844_, _33843_, _07234_);
  or _83399_ (_33845_, _33844_, _33842_);
  and _83400_ (_33846_, _07900_, _07133_);
  or _83401_ (_33848_, _33846_, _33843_);
  or _83402_ (_33849_, _33848_, _07215_);
  nor _83403_ (_33850_, _08390_, _13593_);
  or _83404_ (_33851_, _33850_, _33843_);
  and _83405_ (_33852_, _33851_, _06341_);
  and _83406_ (_33853_, _07142_, \oc8051_golden_model_1.IE [0]);
  or _83407_ (_33854_, _33841_, _33843_);
  and _83408_ (_33855_, _33854_, _07141_);
  or _83409_ (_33856_, _33855_, _33853_);
  and _83410_ (_33857_, _33856_, _07151_);
  or _83411_ (_33859_, _33857_, _06272_);
  or _83412_ (_33860_, _33859_, _33852_);
  and _83413_ (_33861_, _14382_, _08626_);
  and _83414_ (_33862_, _13601_, \oc8051_golden_model_1.IE [0]);
  or _83415_ (_33863_, _33862_, _06273_);
  or _83416_ (_33864_, _33863_, _33861_);
  and _83417_ (_33865_, _33864_, _07166_);
  and _83418_ (_33866_, _33865_, _33860_);
  and _83419_ (_33867_, _33848_, _06461_);
  or _83420_ (_33868_, _33867_, _06464_);
  or _83421_ (_33870_, _33868_, _33866_);
  or _83422_ (_33871_, _33854_, _06465_);
  and _83423_ (_33872_, _33871_, _06269_);
  and _83424_ (_33873_, _33872_, _33870_);
  and _83425_ (_33874_, _33843_, _06268_);
  or _83426_ (_33875_, _33874_, _06261_);
  or _83427_ (_33876_, _33875_, _33873_);
  or _83428_ (_33877_, _33851_, _06262_);
  and _83429_ (_33878_, _33877_, _06258_);
  and _83430_ (_33879_, _33878_, _33876_);
  and _83431_ (_33881_, _14413_, _08626_);
  or _83432_ (_33882_, _33881_, _33862_);
  and _83433_ (_33883_, _33882_, _06257_);
  or _83434_ (_33884_, _33883_, _10080_);
  or _83435_ (_33885_, _33884_, _33879_);
  and _83436_ (_33886_, _33885_, _33849_);
  or _83437_ (_33887_, _33886_, _07460_);
  and _83438_ (_33888_, _09392_, _07900_);
  or _83439_ (_33889_, _33843_, _07208_);
  or _83440_ (_33890_, _33889_, _33888_);
  and _83441_ (_33892_, _33890_, _33887_);
  or _83442_ (_33893_, _33892_, _10094_);
  and _83443_ (_33894_, _14467_, _07900_);
  or _83444_ (_33895_, _33843_, _05982_);
  or _83445_ (_33896_, _33895_, _33894_);
  and _83446_ (_33897_, _33896_, _06219_);
  and _83447_ (_33898_, _33897_, _33893_);
  and _83448_ (_33899_, _07900_, _08954_);
  or _83449_ (_33900_, _33899_, _33843_);
  and _83450_ (_33901_, _33900_, _06218_);
  or _83451_ (_33903_, _33901_, _06369_);
  or _83452_ (_33904_, _33903_, _33898_);
  and _83453_ (_33905_, _14366_, _07900_);
  or _83454_ (_33906_, _33905_, _33843_);
  or _83455_ (_33907_, _33906_, _07237_);
  and _83456_ (_33908_, _33907_, _07240_);
  and _83457_ (_33909_, _33908_, _33904_);
  nor _83458_ (_33910_, _12580_, _13593_);
  or _83459_ (_33911_, _33910_, _33843_);
  nor _83460_ (_33912_, _33842_, _07240_);
  and _83461_ (_33914_, _33912_, _33911_);
  or _83462_ (_33915_, _33914_, _33909_);
  and _83463_ (_33916_, _33915_, _07242_);
  nand _83464_ (_33917_, _33900_, _06375_);
  nor _83465_ (_33918_, _33917_, _33850_);
  or _83466_ (_33919_, _33918_, _06545_);
  or _83467_ (_33920_, _33919_, _33916_);
  and _83468_ (_33921_, _33920_, _33845_);
  or _83469_ (_33922_, _33921_, _06366_);
  and _83470_ (_33923_, _14363_, _07900_);
  or _83471_ (_33925_, _33843_, _09056_);
  or _83472_ (_33926_, _33925_, _33923_);
  and _83473_ (_33927_, _33926_, _09061_);
  and _83474_ (_33928_, _33927_, _33922_);
  and _83475_ (_33929_, _33911_, _06528_);
  or _83476_ (_33930_, _33929_, _06568_);
  or _83477_ (_33931_, _33930_, _33928_);
  or _83478_ (_33932_, _33851_, _06926_);
  and _83479_ (_33933_, _33932_, _33931_);
  or _83480_ (_33934_, _33933_, _05927_);
  or _83481_ (_33936_, _33843_, _05928_);
  and _83482_ (_33937_, _33936_, _33934_);
  or _83483_ (_33938_, _33937_, _06278_);
  or _83484_ (_33939_, _33851_, _06279_);
  and _83485_ (_33940_, _33939_, _01347_);
  and _83486_ (_33941_, _33940_, _33938_);
  or _83487_ (_33942_, _33941_, _33840_);
  and _83488_ (_43304_, _33942_, _42618_);
  not _83489_ (_33943_, \oc8051_golden_model_1.IE [1]);
  nor _83490_ (_33944_, _01347_, _33943_);
  nor _83491_ (_33946_, _07900_, _33943_);
  nor _83492_ (_33947_, _11261_, _13593_);
  or _83493_ (_33948_, _33947_, _33946_);
  or _83494_ (_33949_, _33948_, _09061_);
  nand _83495_ (_33950_, _07900_, _07038_);
  or _83496_ (_33951_, _07900_, \oc8051_golden_model_1.IE [1]);
  and _83497_ (_33952_, _33951_, _06218_);
  and _83498_ (_33953_, _33952_, _33950_);
  nor _83499_ (_33954_, _13593_, _07357_);
  or _83500_ (_33955_, _33954_, _33946_);
  or _83501_ (_33957_, _33955_, _07166_);
  and _83502_ (_33958_, _14562_, _07900_);
  not _83503_ (_33959_, _33958_);
  and _83504_ (_33960_, _33959_, _33951_);
  or _83505_ (_33961_, _33960_, _07151_);
  and _83506_ (_33962_, _07900_, \oc8051_golden_model_1.ACC [1]);
  or _83507_ (_33963_, _33962_, _33946_);
  and _83508_ (_33964_, _33963_, _07141_);
  nor _83509_ (_33965_, _07141_, _33943_);
  or _83510_ (_33966_, _33965_, _06341_);
  or _83511_ (_33967_, _33966_, _33964_);
  and _83512_ (_33968_, _33967_, _06273_);
  and _83513_ (_33969_, _33968_, _33961_);
  nor _83514_ (_33970_, _08626_, _33943_);
  and _83515_ (_33971_, _14557_, _08626_);
  or _83516_ (_33972_, _33971_, _33970_);
  and _83517_ (_33973_, _33972_, _06272_);
  or _83518_ (_33974_, _33973_, _06461_);
  or _83519_ (_33975_, _33974_, _33969_);
  and _83520_ (_33976_, _33975_, _33957_);
  or _83521_ (_33978_, _33976_, _06464_);
  or _83522_ (_33979_, _33963_, _06465_);
  and _83523_ (_33980_, _33979_, _06269_);
  and _83524_ (_33981_, _33980_, _33978_);
  and _83525_ (_33982_, _14560_, _08626_);
  or _83526_ (_33983_, _33982_, _33970_);
  and _83527_ (_33984_, _33983_, _06268_);
  or _83528_ (_33985_, _33984_, _06261_);
  or _83529_ (_33986_, _33985_, _33981_);
  and _83530_ (_33987_, _33971_, _14556_);
  or _83531_ (_33989_, _33970_, _06262_);
  or _83532_ (_33990_, _33989_, _33987_);
  and _83533_ (_33991_, _33990_, _06258_);
  and _83534_ (_33992_, _33991_, _33986_);
  or _83535_ (_33993_, _33970_, _14597_);
  and _83536_ (_33994_, _33993_, _06257_);
  and _83537_ (_33995_, _33994_, _33972_);
  or _83538_ (_33996_, _33995_, _10080_);
  or _83539_ (_33997_, _33996_, _33992_);
  or _83540_ (_33998_, _33955_, _07215_);
  and _83541_ (_34000_, _33998_, _33997_);
  or _83542_ (_34001_, _34000_, _07460_);
  and _83543_ (_34002_, _09451_, _07900_);
  or _83544_ (_34003_, _33946_, _07208_);
  or _83545_ (_34004_, _34003_, _34002_);
  and _83546_ (_34005_, _34004_, _05982_);
  and _83547_ (_34006_, _34005_, _34001_);
  and _83548_ (_34007_, _14653_, _07900_);
  or _83549_ (_34008_, _34007_, _33946_);
  and _83550_ (_34009_, _34008_, _10094_);
  or _83551_ (_34011_, _34009_, _34006_);
  and _83552_ (_34012_, _34011_, _06219_);
  or _83553_ (_34013_, _34012_, _33953_);
  and _83554_ (_34014_, _34013_, _07237_);
  or _83555_ (_34015_, _14668_, _13593_);
  and _83556_ (_34016_, _33951_, _06369_);
  and _83557_ (_34017_, _34016_, _34015_);
  or _83558_ (_34018_, _34017_, _06536_);
  or _83559_ (_34019_, _34018_, _34014_);
  nand _83560_ (_34020_, _11260_, _07900_);
  and _83561_ (_34022_, _34020_, _33948_);
  or _83562_ (_34023_, _34022_, _07240_);
  and _83563_ (_34024_, _34023_, _07242_);
  and _83564_ (_34025_, _34024_, _34019_);
  or _83565_ (_34026_, _14666_, _13593_);
  and _83566_ (_34027_, _33951_, _06375_);
  and _83567_ (_34028_, _34027_, _34026_);
  or _83568_ (_34029_, _34028_, _06545_);
  or _83569_ (_34030_, _34029_, _34025_);
  nor _83570_ (_34031_, _33946_, _07234_);
  nand _83571_ (_34033_, _34031_, _34020_);
  and _83572_ (_34034_, _34033_, _09056_);
  and _83573_ (_34035_, _34034_, _34030_);
  or _83574_ (_34036_, _33950_, _08341_);
  and _83575_ (_34037_, _33951_, _06366_);
  and _83576_ (_34038_, _34037_, _34036_);
  or _83577_ (_34039_, _34038_, _06528_);
  or _83578_ (_34040_, _34039_, _34035_);
  and _83579_ (_34041_, _34040_, _33949_);
  or _83580_ (_34042_, _34041_, _06568_);
  or _83581_ (_34044_, _33960_, _06926_);
  and _83582_ (_34045_, _34044_, _05928_);
  and _83583_ (_34046_, _34045_, _34042_);
  and _83584_ (_34047_, _33983_, _05927_);
  or _83585_ (_34048_, _34047_, _06278_);
  or _83586_ (_34049_, _34048_, _34046_);
  or _83587_ (_34050_, _33946_, _06279_);
  or _83588_ (_34051_, _34050_, _33958_);
  and _83589_ (_34052_, _34051_, _01347_);
  and _83590_ (_34053_, _34052_, _34049_);
  or _83591_ (_34055_, _34053_, _33944_);
  and _83592_ (_43306_, _34055_, _42618_);
  and _83593_ (_34056_, _01351_, \oc8051_golden_model_1.IE [2]);
  and _83594_ (_34057_, _13593_, \oc8051_golden_model_1.IE [2]);
  nor _83595_ (_34058_, _13593_, _07776_);
  or _83596_ (_34059_, _34058_, _34057_);
  or _83597_ (_34060_, _34059_, _07215_);
  or _83598_ (_34061_, _34059_, _07166_);
  and _83599_ (_34062_, _14770_, _07900_);
  or _83600_ (_34063_, _34062_, _34057_);
  or _83601_ (_34065_, _34063_, _07151_);
  and _83602_ (_34066_, _07900_, \oc8051_golden_model_1.ACC [2]);
  or _83603_ (_34067_, _34066_, _34057_);
  and _83604_ (_34068_, _34067_, _07141_);
  and _83605_ (_34069_, _07142_, \oc8051_golden_model_1.IE [2]);
  or _83606_ (_34070_, _34069_, _06341_);
  or _83607_ (_34071_, _34070_, _34068_);
  and _83608_ (_34072_, _34071_, _06273_);
  and _83609_ (_34073_, _34072_, _34065_);
  and _83610_ (_34074_, _13601_, \oc8051_golden_model_1.IE [2]);
  and _83611_ (_34076_, _14774_, _08626_);
  or _83612_ (_34077_, _34076_, _34074_);
  and _83613_ (_34078_, _34077_, _06272_);
  or _83614_ (_34079_, _34078_, _06461_);
  or _83615_ (_34080_, _34079_, _34073_);
  and _83616_ (_34081_, _34080_, _34061_);
  or _83617_ (_34082_, _34081_, _06464_);
  or _83618_ (_34083_, _34067_, _06465_);
  and _83619_ (_34084_, _34083_, _06269_);
  and _83620_ (_34085_, _34084_, _34082_);
  and _83621_ (_34087_, _14756_, _08626_);
  or _83622_ (_34088_, _34087_, _34074_);
  and _83623_ (_34089_, _34088_, _06268_);
  or _83624_ (_34090_, _34089_, _06261_);
  or _83625_ (_34091_, _34090_, _34085_);
  and _83626_ (_34092_, _34076_, _14789_);
  or _83627_ (_34093_, _34074_, _06262_);
  or _83628_ (_34094_, _34093_, _34092_);
  and _83629_ (_34095_, _34094_, _06258_);
  and _83630_ (_34096_, _34095_, _34091_);
  and _83631_ (_34098_, _14804_, _08626_);
  or _83632_ (_34099_, _34098_, _34074_);
  and _83633_ (_34100_, _34099_, _06257_);
  or _83634_ (_34101_, _34100_, _10080_);
  or _83635_ (_34102_, _34101_, _34096_);
  and _83636_ (_34103_, _34102_, _34060_);
  or _83637_ (_34104_, _34103_, _07460_);
  and _83638_ (_34105_, _09450_, _07900_);
  or _83639_ (_34106_, _34057_, _07208_);
  or _83640_ (_34107_, _34106_, _34105_);
  and _83641_ (_34109_, _34107_, _05982_);
  and _83642_ (_34110_, _34109_, _34104_);
  and _83643_ (_34111_, _14859_, _07900_);
  or _83644_ (_34112_, _34111_, _34057_);
  and _83645_ (_34113_, _34112_, _10094_);
  or _83646_ (_34114_, _34113_, _06218_);
  or _83647_ (_34115_, _34114_, _34110_);
  and _83648_ (_34116_, _07900_, _08973_);
  or _83649_ (_34117_, _34116_, _34057_);
  or _83650_ (_34118_, _34117_, _06219_);
  and _83651_ (_34120_, _34118_, _34115_);
  or _83652_ (_34121_, _34120_, _06369_);
  and _83653_ (_34122_, _14751_, _07900_);
  or _83654_ (_34123_, _34122_, _34057_);
  or _83655_ (_34124_, _34123_, _07237_);
  and _83656_ (_34125_, _34124_, _07240_);
  and _83657_ (_34126_, _34125_, _34121_);
  and _83658_ (_34127_, _11259_, _07900_);
  or _83659_ (_34128_, _34127_, _34057_);
  and _83660_ (_34129_, _34128_, _06536_);
  or _83661_ (_34131_, _34129_, _34126_);
  and _83662_ (_34132_, _34131_, _07242_);
  or _83663_ (_34133_, _34057_, _08440_);
  and _83664_ (_34134_, _34117_, _06375_);
  and _83665_ (_34135_, _34134_, _34133_);
  or _83666_ (_34136_, _34135_, _34132_);
  and _83667_ (_34137_, _34136_, _07234_);
  and _83668_ (_34138_, _34067_, _06545_);
  and _83669_ (_34139_, _34138_, _34133_);
  or _83670_ (_34140_, _34139_, _06366_);
  or _83671_ (_34142_, _34140_, _34137_);
  and _83672_ (_34143_, _14748_, _07900_);
  or _83673_ (_34144_, _34057_, _09056_);
  or _83674_ (_34145_, _34144_, _34143_);
  and _83675_ (_34146_, _34145_, _09061_);
  and _83676_ (_34147_, _34146_, _34142_);
  nor _83677_ (_34148_, _11258_, _13593_);
  or _83678_ (_34149_, _34148_, _34057_);
  and _83679_ (_34150_, _34149_, _06528_);
  or _83680_ (_34151_, _34150_, _06568_);
  or _83681_ (_34153_, _34151_, _34147_);
  or _83682_ (_34154_, _34063_, _06926_);
  and _83683_ (_34155_, _34154_, _05928_);
  and _83684_ (_34156_, _34155_, _34153_);
  and _83685_ (_34157_, _34088_, _05927_);
  or _83686_ (_34158_, _34157_, _06278_);
  or _83687_ (_34159_, _34158_, _34156_);
  and _83688_ (_34160_, _14926_, _07900_);
  or _83689_ (_34161_, _34057_, _06279_);
  or _83690_ (_34162_, _34161_, _34160_);
  and _83691_ (_34164_, _34162_, _01347_);
  and _83692_ (_34165_, _34164_, _34159_);
  or _83693_ (_34166_, _34165_, _34056_);
  and _83694_ (_43307_, _34166_, _42618_);
  and _83695_ (_34167_, _01351_, \oc8051_golden_model_1.IE [3]);
  and _83696_ (_34168_, _13593_, \oc8051_golden_model_1.IE [3]);
  nor _83697_ (_34169_, _13593_, _07594_);
  or _83698_ (_34170_, _34169_, _34168_);
  or _83699_ (_34171_, _34170_, _07215_);
  and _83700_ (_34172_, _14953_, _07900_);
  or _83701_ (_34174_, _34172_, _34168_);
  or _83702_ (_34175_, _34174_, _07151_);
  and _83703_ (_34176_, _07900_, \oc8051_golden_model_1.ACC [3]);
  or _83704_ (_34177_, _34176_, _34168_);
  and _83705_ (_34178_, _34177_, _07141_);
  and _83706_ (_34179_, _07142_, \oc8051_golden_model_1.IE [3]);
  or _83707_ (_34180_, _34179_, _06341_);
  or _83708_ (_34181_, _34180_, _34178_);
  and _83709_ (_34183_, _34181_, _06273_);
  and _83710_ (_34185_, _34183_, _34175_);
  and _83711_ (_34188_, _13601_, \oc8051_golden_model_1.IE [3]);
  and _83712_ (_34190_, _14950_, _08626_);
  or _83713_ (_34192_, _34190_, _34188_);
  and _83714_ (_34194_, _34192_, _06272_);
  or _83715_ (_34196_, _34194_, _06461_);
  or _83716_ (_34198_, _34196_, _34185_);
  or _83717_ (_34200_, _34170_, _07166_);
  and _83718_ (_34202_, _34200_, _34198_);
  or _83719_ (_34203_, _34202_, _06464_);
  or _83720_ (_34204_, _34177_, _06465_);
  and _83721_ (_34206_, _34204_, _06269_);
  and _83722_ (_34207_, _34206_, _34203_);
  and _83723_ (_34208_, _14948_, _08626_);
  or _83724_ (_34209_, _34208_, _34188_);
  and _83725_ (_34210_, _34209_, _06268_);
  or _83726_ (_34211_, _34210_, _06261_);
  or _83727_ (_34212_, _34211_, _34207_);
  or _83728_ (_34213_, _34188_, _14979_);
  and _83729_ (_34214_, _34213_, _34192_);
  or _83730_ (_34215_, _34214_, _06262_);
  and _83731_ (_34217_, _34215_, _06258_);
  and _83732_ (_34218_, _34217_, _34212_);
  or _83733_ (_34219_, _34188_, _14992_);
  and _83734_ (_34220_, _34219_, _06257_);
  and _83735_ (_34221_, _34220_, _34192_);
  or _83736_ (_34222_, _34221_, _10080_);
  or _83737_ (_34223_, _34222_, _34218_);
  and _83738_ (_34224_, _34223_, _34171_);
  or _83739_ (_34225_, _34224_, _07460_);
  and _83740_ (_34226_, _09449_, _07900_);
  or _83741_ (_34228_, _34168_, _07208_);
  or _83742_ (_34229_, _34228_, _34226_);
  and _83743_ (_34230_, _34229_, _05982_);
  and _83744_ (_34231_, _34230_, _34225_);
  and _83745_ (_34232_, _15048_, _07900_);
  or _83746_ (_34233_, _34232_, _34168_);
  and _83747_ (_34234_, _34233_, _10094_);
  or _83748_ (_34235_, _34234_, _06218_);
  or _83749_ (_34236_, _34235_, _34231_);
  and _83750_ (_34237_, _07900_, _08930_);
  or _83751_ (_34239_, _34237_, _34168_);
  or _83752_ (_34240_, _34239_, _06219_);
  and _83753_ (_34241_, _34240_, _34236_);
  or _83754_ (_34242_, _34241_, _06369_);
  and _83755_ (_34243_, _14943_, _07900_);
  or _83756_ (_34244_, _34243_, _34168_);
  or _83757_ (_34245_, _34244_, _07237_);
  and _83758_ (_34246_, _34245_, _07240_);
  and _83759_ (_34247_, _34246_, _34242_);
  and _83760_ (_34248_, _12577_, _07900_);
  or _83761_ (_34250_, _34248_, _34168_);
  and _83762_ (_34251_, _34250_, _06536_);
  or _83763_ (_34252_, _34251_, _34247_);
  and _83764_ (_34253_, _34252_, _07242_);
  or _83765_ (_34254_, _34168_, _08292_);
  and _83766_ (_34255_, _34239_, _06375_);
  and _83767_ (_34256_, _34255_, _34254_);
  or _83768_ (_34257_, _34256_, _34253_);
  and _83769_ (_34258_, _34257_, _07234_);
  and _83770_ (_34259_, _34177_, _06545_);
  and _83771_ (_34261_, _34259_, _34254_);
  or _83772_ (_34262_, _34261_, _06366_);
  or _83773_ (_34263_, _34262_, _34258_);
  and _83774_ (_34264_, _14940_, _07900_);
  or _83775_ (_34265_, _34168_, _09056_);
  or _83776_ (_34266_, _34265_, _34264_);
  and _83777_ (_34267_, _34266_, _09061_);
  and _83778_ (_34268_, _34267_, _34263_);
  nor _83779_ (_34269_, _11256_, _13593_);
  or _83780_ (_34270_, _34269_, _34168_);
  and _83781_ (_34272_, _34270_, _06528_);
  or _83782_ (_34273_, _34272_, _06568_);
  or _83783_ (_34274_, _34273_, _34268_);
  or _83784_ (_34275_, _34174_, _06926_);
  and _83785_ (_34276_, _34275_, _05928_);
  and _83786_ (_34277_, _34276_, _34274_);
  and _83787_ (_34278_, _34209_, _05927_);
  or _83788_ (_34279_, _34278_, _06278_);
  or _83789_ (_34280_, _34279_, _34277_);
  and _83790_ (_34281_, _15128_, _07900_);
  or _83791_ (_34283_, _34168_, _06279_);
  or _83792_ (_34284_, _34283_, _34281_);
  and _83793_ (_34285_, _34284_, _01347_);
  and _83794_ (_34286_, _34285_, _34280_);
  or _83795_ (_34287_, _34286_, _34167_);
  and _83796_ (_43308_, _34287_, _42618_);
  and _83797_ (_34288_, _01351_, \oc8051_golden_model_1.IE [4]);
  and _83798_ (_34289_, _13593_, \oc8051_golden_model_1.IE [4]);
  nor _83799_ (_34290_, _08541_, _13593_);
  or _83800_ (_34291_, _34290_, _34289_);
  or _83801_ (_34293_, _34291_, _07215_);
  and _83802_ (_34294_, _13601_, \oc8051_golden_model_1.IE [4]);
  and _83803_ (_34295_, _15176_, _08626_);
  or _83804_ (_34296_, _34295_, _34294_);
  and _83805_ (_34297_, _34296_, _06268_);
  and _83806_ (_34298_, _15162_, _07900_);
  or _83807_ (_34299_, _34298_, _34289_);
  or _83808_ (_34300_, _34299_, _07151_);
  and _83809_ (_34301_, _07900_, \oc8051_golden_model_1.ACC [4]);
  or _83810_ (_34302_, _34301_, _34289_);
  and _83811_ (_34304_, _34302_, _07141_);
  and _83812_ (_34305_, _07142_, \oc8051_golden_model_1.IE [4]);
  or _83813_ (_34306_, _34305_, _06341_);
  or _83814_ (_34307_, _34306_, _34304_);
  and _83815_ (_34308_, _34307_, _06273_);
  and _83816_ (_34309_, _34308_, _34300_);
  and _83817_ (_34310_, _15166_, _08626_);
  or _83818_ (_34311_, _34310_, _34294_);
  and _83819_ (_34312_, _34311_, _06272_);
  or _83820_ (_34313_, _34312_, _06461_);
  or _83821_ (_34315_, _34313_, _34309_);
  or _83822_ (_34316_, _34291_, _07166_);
  and _83823_ (_34317_, _34316_, _34315_);
  or _83824_ (_34318_, _34317_, _06464_);
  or _83825_ (_34319_, _34302_, _06465_);
  and _83826_ (_34320_, _34319_, _06269_);
  and _83827_ (_34321_, _34320_, _34318_);
  or _83828_ (_34322_, _34321_, _34297_);
  and _83829_ (_34323_, _34322_, _06262_);
  and _83830_ (_34324_, _15184_, _08626_);
  or _83831_ (_34326_, _34324_, _34294_);
  and _83832_ (_34327_, _34326_, _06261_);
  or _83833_ (_34328_, _34327_, _34323_);
  and _83834_ (_34329_, _34328_, _06258_);
  and _83835_ (_34330_, _15200_, _08626_);
  or _83836_ (_34331_, _34330_, _34294_);
  and _83837_ (_34332_, _34331_, _06257_);
  or _83838_ (_34333_, _34332_, _10080_);
  or _83839_ (_34334_, _34333_, _34329_);
  and _83840_ (_34335_, _34334_, _34293_);
  or _83841_ (_34337_, _34335_, _07460_);
  and _83842_ (_34338_, _09448_, _07900_);
  or _83843_ (_34339_, _34289_, _07208_);
  or _83844_ (_34340_, _34339_, _34338_);
  and _83845_ (_34341_, _34340_, _05982_);
  and _83846_ (_34342_, _34341_, _34337_);
  and _83847_ (_34343_, _15254_, _07900_);
  or _83848_ (_34344_, _34343_, _34289_);
  and _83849_ (_34345_, _34344_, _10094_);
  or _83850_ (_34346_, _34345_, _06218_);
  or _83851_ (_34348_, _34346_, _34342_);
  and _83852_ (_34349_, _08959_, _07900_);
  or _83853_ (_34350_, _34349_, _34289_);
  or _83854_ (_34351_, _34350_, _06219_);
  and _83855_ (_34352_, _34351_, _34348_);
  or _83856_ (_34353_, _34352_, _06369_);
  and _83857_ (_34354_, _15269_, _07900_);
  or _83858_ (_34355_, _34354_, _34289_);
  or _83859_ (_34356_, _34355_, _07237_);
  and _83860_ (_34357_, _34356_, _07240_);
  and _83861_ (_34359_, _34357_, _34353_);
  and _83862_ (_34360_, _11254_, _07900_);
  or _83863_ (_34361_, _34360_, _34289_);
  and _83864_ (_34362_, _34361_, _06536_);
  or _83865_ (_34363_, _34362_, _34359_);
  and _83866_ (_34364_, _34363_, _07242_);
  or _83867_ (_34365_, _34289_, _08544_);
  and _83868_ (_34366_, _34350_, _06375_);
  and _83869_ (_34367_, _34366_, _34365_);
  or _83870_ (_34368_, _34367_, _34364_);
  and _83871_ (_34370_, _34368_, _07234_);
  and _83872_ (_34371_, _34302_, _06545_);
  and _83873_ (_34372_, _34371_, _34365_);
  or _83874_ (_34373_, _34372_, _06366_);
  or _83875_ (_34374_, _34373_, _34370_);
  and _83876_ (_34375_, _15266_, _07900_);
  or _83877_ (_34376_, _34289_, _09056_);
  or _83878_ (_34377_, _34376_, _34375_);
  and _83879_ (_34378_, _34377_, _09061_);
  and _83880_ (_34379_, _34378_, _34374_);
  nor _83881_ (_34381_, _11253_, _13593_);
  or _83882_ (_34382_, _34381_, _34289_);
  and _83883_ (_34383_, _34382_, _06528_);
  or _83884_ (_34384_, _34383_, _06568_);
  or _83885_ (_34385_, _34384_, _34379_);
  or _83886_ (_34386_, _34299_, _06926_);
  and _83887_ (_34387_, _34386_, _05928_);
  and _83888_ (_34388_, _34387_, _34385_);
  and _83889_ (_34389_, _34296_, _05927_);
  or _83890_ (_34390_, _34389_, _06278_);
  or _83891_ (_34392_, _34390_, _34388_);
  and _83892_ (_34393_, _15329_, _07900_);
  or _83893_ (_34394_, _34289_, _06279_);
  or _83894_ (_34395_, _34394_, _34393_);
  and _83895_ (_34396_, _34395_, _01347_);
  and _83896_ (_34397_, _34396_, _34392_);
  or _83897_ (_34398_, _34397_, _34288_);
  and _83898_ (_43309_, _34398_, _42618_);
  and _83899_ (_34399_, _01351_, \oc8051_golden_model_1.IE [5]);
  and _83900_ (_34400_, _13593_, \oc8051_golden_model_1.IE [5]);
  and _83901_ (_34402_, _15358_, _07900_);
  or _83902_ (_34403_, _34402_, _34400_);
  or _83903_ (_34404_, _34403_, _07151_);
  and _83904_ (_34405_, _07900_, \oc8051_golden_model_1.ACC [5]);
  or _83905_ (_34406_, _34405_, _34400_);
  and _83906_ (_34407_, _34406_, _07141_);
  and _83907_ (_34408_, _07142_, \oc8051_golden_model_1.IE [5]);
  or _83908_ (_34409_, _34408_, _06341_);
  or _83909_ (_34410_, _34409_, _34407_);
  and _83910_ (_34411_, _34410_, _06273_);
  and _83911_ (_34413_, _34411_, _34404_);
  and _83912_ (_34414_, _13601_, \oc8051_golden_model_1.IE [5]);
  and _83913_ (_34415_, _15372_, _08626_);
  or _83914_ (_34416_, _34415_, _34414_);
  and _83915_ (_34417_, _34416_, _06272_);
  or _83916_ (_34418_, _34417_, _06461_);
  or _83917_ (_34419_, _34418_, _34413_);
  nor _83918_ (_34420_, _08244_, _13593_);
  or _83919_ (_34421_, _34420_, _34400_);
  or _83920_ (_34422_, _34421_, _07166_);
  and _83921_ (_34424_, _34422_, _34419_);
  or _83922_ (_34425_, _34424_, _06464_);
  or _83923_ (_34426_, _34406_, _06465_);
  and _83924_ (_34427_, _34426_, _06269_);
  and _83925_ (_34428_, _34427_, _34425_);
  and _83926_ (_34429_, _15355_, _08626_);
  or _83927_ (_34430_, _34429_, _34414_);
  and _83928_ (_34431_, _34430_, _06268_);
  or _83929_ (_34432_, _34431_, _06261_);
  or _83930_ (_34433_, _34432_, _34428_);
  or _83931_ (_34435_, _34414_, _15387_);
  and _83932_ (_34436_, _34435_, _34416_);
  or _83933_ (_34437_, _34436_, _06262_);
  and _83934_ (_34438_, _34437_, _06258_);
  and _83935_ (_34439_, _34438_, _34433_);
  or _83936_ (_34440_, _34414_, _15403_);
  and _83937_ (_34441_, _34440_, _06257_);
  and _83938_ (_34442_, _34441_, _34416_);
  or _83939_ (_34443_, _34442_, _10080_);
  or _83940_ (_34444_, _34443_, _34439_);
  or _83941_ (_34446_, _34421_, _07215_);
  and _83942_ (_34447_, _34446_, _34444_);
  or _83943_ (_34448_, _34447_, _07460_);
  and _83944_ (_34449_, _09447_, _07900_);
  or _83945_ (_34450_, _34400_, _07208_);
  or _83946_ (_34451_, _34450_, _34449_);
  and _83947_ (_34452_, _34451_, _05982_);
  and _83948_ (_34453_, _34452_, _34448_);
  and _83949_ (_34454_, _15459_, _07900_);
  or _83950_ (_34455_, _34454_, _34400_);
  and _83951_ (_34457_, _34455_, _10094_);
  or _83952_ (_34458_, _34457_, _06218_);
  or _83953_ (_34459_, _34458_, _34453_);
  and _83954_ (_34460_, _08946_, _07900_);
  or _83955_ (_34461_, _34460_, _34400_);
  or _83956_ (_34462_, _34461_, _06219_);
  and _83957_ (_34463_, _34462_, _34459_);
  or _83958_ (_34464_, _34463_, _06369_);
  and _83959_ (_34465_, _15353_, _07900_);
  or _83960_ (_34466_, _34465_, _34400_);
  or _83961_ (_34468_, _34466_, _07237_);
  and _83962_ (_34469_, _34468_, _07240_);
  and _83963_ (_34470_, _34469_, _34464_);
  and _83964_ (_34471_, _11250_, _07900_);
  or _83965_ (_34472_, _34471_, _34400_);
  and _83966_ (_34473_, _34472_, _06536_);
  or _83967_ (_34474_, _34473_, _34470_);
  and _83968_ (_34475_, _34474_, _07242_);
  or _83969_ (_34476_, _34400_, _08247_);
  and _83970_ (_34477_, _34461_, _06375_);
  and _83971_ (_34479_, _34477_, _34476_);
  or _83972_ (_34480_, _34479_, _34475_);
  and _83973_ (_34481_, _34480_, _07234_);
  and _83974_ (_34482_, _34406_, _06545_);
  and _83975_ (_34483_, _34482_, _34476_);
  or _83976_ (_34484_, _34483_, _06366_);
  or _83977_ (_34485_, _34484_, _34481_);
  and _83978_ (_34486_, _15350_, _07900_);
  or _83979_ (_34487_, _34400_, _09056_);
  or _83980_ (_34488_, _34487_, _34486_);
  and _83981_ (_34490_, _34488_, _09061_);
  and _83982_ (_34491_, _34490_, _34485_);
  nor _83983_ (_34492_, _11249_, _13593_);
  or _83984_ (_34493_, _34492_, _34400_);
  and _83985_ (_34494_, _34493_, _06528_);
  or _83986_ (_34495_, _34494_, _06568_);
  or _83987_ (_34496_, _34495_, _34491_);
  or _83988_ (_34497_, _34403_, _06926_);
  and _83989_ (_34498_, _34497_, _05928_);
  and _83990_ (_34499_, _34498_, _34496_);
  and _83991_ (_34501_, _34430_, _05927_);
  or _83992_ (_34502_, _34501_, _06278_);
  or _83993_ (_34503_, _34502_, _34499_);
  and _83994_ (_34504_, _15532_, _07900_);
  or _83995_ (_34505_, _34400_, _06279_);
  or _83996_ (_34506_, _34505_, _34504_);
  and _83997_ (_34507_, _34506_, _01347_);
  and _83998_ (_34508_, _34507_, _34503_);
  or _83999_ (_34509_, _34508_, _34399_);
  and _84000_ (_43310_, _34509_, _42618_);
  and _84001_ (_34511_, _01351_, \oc8051_golden_model_1.IE [6]);
  and _84002_ (_34512_, _13593_, \oc8051_golden_model_1.IE [6]);
  and _84003_ (_34513_, _15554_, _07900_);
  or _84004_ (_34514_, _34513_, _34512_);
  or _84005_ (_34515_, _34514_, _07151_);
  and _84006_ (_34516_, _07900_, \oc8051_golden_model_1.ACC [6]);
  or _84007_ (_34517_, _34516_, _34512_);
  and _84008_ (_34518_, _34517_, _07141_);
  and _84009_ (_34519_, _07142_, \oc8051_golden_model_1.IE [6]);
  or _84010_ (_34520_, _34519_, _06341_);
  or _84011_ (_34522_, _34520_, _34518_);
  and _84012_ (_34523_, _34522_, _06273_);
  and _84013_ (_34524_, _34523_, _34515_);
  and _84014_ (_34525_, _13601_, \oc8051_golden_model_1.IE [6]);
  and _84015_ (_34526_, _15570_, _08626_);
  or _84016_ (_34527_, _34526_, _34525_);
  and _84017_ (_34528_, _34527_, _06272_);
  or _84018_ (_34529_, _34528_, _06461_);
  or _84019_ (_34530_, _34529_, _34524_);
  nor _84020_ (_34531_, _08142_, _13593_);
  or _84021_ (_34533_, _34531_, _34512_);
  or _84022_ (_34534_, _34533_, _07166_);
  and _84023_ (_34535_, _34534_, _34530_);
  or _84024_ (_34536_, _34535_, _06464_);
  or _84025_ (_34537_, _34517_, _06465_);
  and _84026_ (_34538_, _34537_, _06269_);
  and _84027_ (_34539_, _34538_, _34536_);
  and _84028_ (_34540_, _15551_, _08626_);
  or _84029_ (_34541_, _34540_, _34525_);
  and _84030_ (_34542_, _34541_, _06268_);
  or _84031_ (_34544_, _34542_, _06261_);
  or _84032_ (_34545_, _34544_, _34539_);
  or _84033_ (_34546_, _34525_, _15585_);
  and _84034_ (_34547_, _34546_, _34527_);
  or _84035_ (_34548_, _34547_, _06262_);
  and _84036_ (_34549_, _34548_, _06258_);
  and _84037_ (_34550_, _34549_, _34545_);
  and _84038_ (_34551_, _15602_, _08626_);
  or _84039_ (_34552_, _34551_, _34525_);
  and _84040_ (_34553_, _34552_, _06257_);
  or _84041_ (_34555_, _34553_, _10080_);
  or _84042_ (_34556_, _34555_, _34550_);
  or _84043_ (_34557_, _34533_, _07215_);
  and _84044_ (_34558_, _34557_, _34556_);
  or _84045_ (_34559_, _34558_, _07460_);
  and _84046_ (_34560_, _09446_, _07900_);
  or _84047_ (_34561_, _34512_, _07208_);
  or _84048_ (_34562_, _34561_, _34560_);
  and _84049_ (_34563_, _34562_, _05982_);
  and _84050_ (_34564_, _34563_, _34559_);
  and _84051_ (_34566_, _15657_, _07900_);
  or _84052_ (_34567_, _34566_, _34512_);
  and _84053_ (_34568_, _34567_, _10094_);
  or _84054_ (_34569_, _34568_, _06218_);
  or _84055_ (_34570_, _34569_, _34564_);
  and _84056_ (_34571_, _15664_, _07900_);
  or _84057_ (_34572_, _34571_, _34512_);
  or _84058_ (_34573_, _34572_, _06219_);
  and _84059_ (_34574_, _34573_, _34570_);
  or _84060_ (_34575_, _34574_, _06369_);
  and _84061_ (_34577_, _15549_, _07900_);
  or _84062_ (_34578_, _34577_, _34512_);
  or _84063_ (_34579_, _34578_, _07237_);
  and _84064_ (_34580_, _34579_, _07240_);
  and _84065_ (_34581_, _34580_, _34575_);
  and _84066_ (_34582_, _11247_, _07900_);
  or _84067_ (_34583_, _34582_, _34512_);
  and _84068_ (_34584_, _34583_, _06536_);
  or _84069_ (_34585_, _34584_, _34581_);
  and _84070_ (_34586_, _34585_, _07242_);
  or _84071_ (_34588_, _34512_, _08145_);
  and _84072_ (_34589_, _34572_, _06375_);
  and _84073_ (_34590_, _34589_, _34588_);
  or _84074_ (_34591_, _34590_, _34586_);
  and _84075_ (_34592_, _34591_, _07234_);
  and _84076_ (_34593_, _34517_, _06545_);
  and _84077_ (_34594_, _34593_, _34588_);
  or _84078_ (_34595_, _34594_, _06366_);
  or _84079_ (_34596_, _34595_, _34592_);
  and _84080_ (_34597_, _15546_, _07900_);
  or _84081_ (_34599_, _34512_, _09056_);
  or _84082_ (_34600_, _34599_, _34597_);
  and _84083_ (_34601_, _34600_, _09061_);
  and _84084_ (_34602_, _34601_, _34596_);
  nor _84085_ (_34603_, _11246_, _13593_);
  or _84086_ (_34604_, _34603_, _34512_);
  and _84087_ (_34605_, _34604_, _06528_);
  or _84088_ (_34606_, _34605_, _06568_);
  or _84089_ (_34607_, _34606_, _34602_);
  or _84090_ (_34608_, _34514_, _06926_);
  and _84091_ (_34610_, _34608_, _05928_);
  and _84092_ (_34611_, _34610_, _34607_);
  and _84093_ (_34612_, _34541_, _05927_);
  or _84094_ (_34613_, _34612_, _06278_);
  or _84095_ (_34614_, _34613_, _34611_);
  and _84096_ (_34615_, _15734_, _07900_);
  or _84097_ (_34616_, _34512_, _06279_);
  or _84098_ (_34617_, _34616_, _34615_);
  and _84099_ (_34618_, _34617_, _01347_);
  and _84100_ (_34619_, _34618_, _34614_);
  or _84101_ (_34621_, _34619_, _34511_);
  and _84102_ (_43311_, _34621_, _42618_);
  not _84103_ (_34622_, \oc8051_golden_model_1.SCON [0]);
  nor _84104_ (_34623_, _01347_, _34622_);
  nand _84105_ (_34624_, _11263_, _07973_);
  nor _84106_ (_34625_, _07973_, _34622_);
  nor _84107_ (_34626_, _34625_, _07234_);
  nand _84108_ (_34627_, _34626_, _34624_);
  and _84109_ (_34628_, _07973_, _07133_);
  or _84110_ (_34629_, _34628_, _34625_);
  or _84111_ (_34631_, _34629_, _07215_);
  nor _84112_ (_34632_, _08390_, _13705_);
  or _84113_ (_34633_, _34632_, _34625_);
  or _84114_ (_34634_, _34633_, _07151_);
  and _84115_ (_34635_, _07973_, \oc8051_golden_model_1.ACC [0]);
  or _84116_ (_34636_, _34635_, _34625_);
  and _84117_ (_34637_, _34636_, _07141_);
  nor _84118_ (_34638_, _07141_, _34622_);
  or _84119_ (_34639_, _34638_, _06341_);
  or _84120_ (_34640_, _34639_, _34637_);
  and _84121_ (_34642_, _34640_, _06273_);
  and _84122_ (_34643_, _34642_, _34634_);
  nor _84123_ (_34644_, _08622_, _34622_);
  and _84124_ (_34645_, _14382_, _08622_);
  or _84125_ (_34646_, _34645_, _34644_);
  and _84126_ (_34647_, _34646_, _06272_);
  or _84127_ (_34648_, _34647_, _34643_);
  and _84128_ (_34649_, _34648_, _07166_);
  and _84129_ (_34650_, _34629_, _06461_);
  or _84130_ (_34651_, _34650_, _06464_);
  or _84131_ (_34653_, _34651_, _34649_);
  or _84132_ (_34654_, _34636_, _06465_);
  and _84133_ (_34655_, _34654_, _06269_);
  and _84134_ (_34656_, _34655_, _34653_);
  and _84135_ (_34657_, _34625_, _06268_);
  or _84136_ (_34658_, _34657_, _06261_);
  or _84137_ (_34659_, _34658_, _34656_);
  or _84138_ (_34660_, _34633_, _06262_);
  and _84139_ (_34661_, _34660_, _06258_);
  and _84140_ (_34662_, _34661_, _34659_);
  and _84141_ (_34664_, _14413_, _08622_);
  or _84142_ (_34665_, _34664_, _34644_);
  and _84143_ (_34666_, _34665_, _06257_);
  or _84144_ (_34667_, _34666_, _10080_);
  or _84145_ (_34668_, _34667_, _34662_);
  and _84146_ (_34669_, _34668_, _34631_);
  or _84147_ (_34670_, _34669_, _07460_);
  and _84148_ (_34671_, _09392_, _07973_);
  or _84149_ (_34672_, _34625_, _07208_);
  or _84150_ (_34673_, _34672_, _34671_);
  and _84151_ (_34675_, _34673_, _34670_);
  or _84152_ (_34676_, _34675_, _10094_);
  and _84153_ (_34677_, _14467_, _07973_);
  or _84154_ (_34678_, _34625_, _05982_);
  or _84155_ (_34679_, _34678_, _34677_);
  and _84156_ (_34680_, _34679_, _06219_);
  and _84157_ (_34681_, _34680_, _34676_);
  and _84158_ (_34682_, _07973_, _08954_);
  or _84159_ (_34683_, _34682_, _34625_);
  and _84160_ (_34684_, _34683_, _06218_);
  or _84161_ (_34686_, _34684_, _06369_);
  or _84162_ (_34687_, _34686_, _34681_);
  and _84163_ (_34688_, _14366_, _07973_);
  or _84164_ (_34689_, _34688_, _34625_);
  or _84165_ (_34690_, _34689_, _07237_);
  and _84166_ (_34691_, _34690_, _07240_);
  and _84167_ (_34692_, _34691_, _34687_);
  nor _84168_ (_34693_, _12580_, _13705_);
  or _84169_ (_34694_, _34693_, _34625_);
  and _84170_ (_34695_, _34624_, _06536_);
  and _84171_ (_34696_, _34695_, _34694_);
  or _84172_ (_34697_, _34696_, _34692_);
  and _84173_ (_34698_, _34697_, _07242_);
  nand _84174_ (_34699_, _34683_, _06375_);
  nor _84175_ (_34700_, _34699_, _34632_);
  or _84176_ (_34701_, _34700_, _06545_);
  or _84177_ (_34702_, _34701_, _34698_);
  and _84178_ (_34703_, _34702_, _34627_);
  or _84179_ (_34704_, _34703_, _06366_);
  and _84180_ (_34705_, _14363_, _07973_);
  or _84181_ (_34707_, _34625_, _09056_);
  or _84182_ (_34708_, _34707_, _34705_);
  and _84183_ (_34709_, _34708_, _09061_);
  and _84184_ (_34710_, _34709_, _34704_);
  and _84185_ (_34711_, _34694_, _06528_);
  or _84186_ (_34712_, _34711_, _06568_);
  or _84187_ (_34713_, _34712_, _34710_);
  or _84188_ (_34714_, _34633_, _06926_);
  and _84189_ (_34715_, _34714_, _34713_);
  or _84190_ (_34716_, _34715_, _05927_);
  or _84191_ (_34718_, _34625_, _05928_);
  and _84192_ (_34719_, _34718_, _34716_);
  or _84193_ (_34720_, _34719_, _06278_);
  or _84194_ (_34721_, _34633_, _06279_);
  and _84195_ (_34722_, _34721_, _01347_);
  and _84196_ (_34723_, _34722_, _34720_);
  or _84197_ (_34724_, _34723_, _34623_);
  and _84198_ (_43313_, _34724_, _42618_);
  not _84199_ (_34725_, \oc8051_golden_model_1.SCON [1]);
  nor _84200_ (_34726_, _01347_, _34725_);
  nor _84201_ (_34728_, _07973_, _34725_);
  nor _84202_ (_34729_, _11261_, _13705_);
  or _84203_ (_34730_, _34729_, _34728_);
  or _84204_ (_34731_, _34730_, _09061_);
  nand _84205_ (_34732_, _07973_, _07038_);
  or _84206_ (_34733_, _07973_, \oc8051_golden_model_1.SCON [1]);
  and _84207_ (_34734_, _34733_, _06218_);
  and _84208_ (_34735_, _34734_, _34732_);
  nor _84209_ (_34736_, _13705_, _07357_);
  or _84210_ (_34737_, _34736_, _34728_);
  or _84211_ (_34739_, _34737_, _07166_);
  and _84212_ (_34740_, _14562_, _07973_);
  not _84213_ (_34741_, _34740_);
  and _84214_ (_34742_, _34741_, _34733_);
  or _84215_ (_34743_, _34742_, _07151_);
  and _84216_ (_34744_, _07973_, \oc8051_golden_model_1.ACC [1]);
  or _84217_ (_34745_, _34744_, _34728_);
  and _84218_ (_34746_, _34745_, _07141_);
  nor _84219_ (_34747_, _07141_, _34725_);
  or _84220_ (_34748_, _34747_, _06341_);
  or _84221_ (_34750_, _34748_, _34746_);
  and _84222_ (_34751_, _34750_, _06273_);
  and _84223_ (_34752_, _34751_, _34743_);
  nor _84224_ (_34753_, _08622_, _34725_);
  and _84225_ (_34754_, _14557_, _08622_);
  or _84226_ (_34755_, _34754_, _34753_);
  and _84227_ (_34756_, _34755_, _06272_);
  or _84228_ (_34757_, _34756_, _06461_);
  or _84229_ (_34758_, _34757_, _34752_);
  and _84230_ (_34759_, _34758_, _34739_);
  or _84231_ (_34761_, _34759_, _06464_);
  or _84232_ (_34762_, _34745_, _06465_);
  and _84233_ (_34763_, _34762_, _06269_);
  and _84234_ (_34764_, _34763_, _34761_);
  and _84235_ (_34765_, _14560_, _08622_);
  or _84236_ (_34766_, _34765_, _34753_);
  and _84237_ (_34767_, _34766_, _06268_);
  or _84238_ (_34768_, _34767_, _06261_);
  or _84239_ (_34769_, _34768_, _34764_);
  and _84240_ (_34770_, _34754_, _14556_);
  or _84241_ (_34772_, _34753_, _06262_);
  or _84242_ (_34773_, _34772_, _34770_);
  and _84243_ (_34774_, _34773_, _06258_);
  and _84244_ (_34775_, _34774_, _34769_);
  or _84245_ (_34776_, _34753_, _14597_);
  and _84246_ (_34777_, _34776_, _06257_);
  and _84247_ (_34778_, _34777_, _34755_);
  or _84248_ (_34779_, _34778_, _10080_);
  or _84249_ (_34780_, _34779_, _34775_);
  or _84250_ (_34781_, _34737_, _07215_);
  and _84251_ (_34783_, _34781_, _34780_);
  or _84252_ (_34784_, _34783_, _07460_);
  and _84253_ (_34785_, _09451_, _07973_);
  or _84254_ (_34786_, _34728_, _07208_);
  or _84255_ (_34787_, _34786_, _34785_);
  and _84256_ (_34788_, _34787_, _05982_);
  and _84257_ (_34789_, _34788_, _34784_);
  and _84258_ (_34790_, _14653_, _07973_);
  or _84259_ (_34791_, _34790_, _34728_);
  and _84260_ (_34792_, _34791_, _10094_);
  or _84261_ (_34794_, _34792_, _34789_);
  and _84262_ (_34795_, _34794_, _06219_);
  or _84263_ (_34796_, _34795_, _34735_);
  and _84264_ (_34797_, _34796_, _07237_);
  or _84265_ (_34798_, _14668_, _13705_);
  and _84266_ (_34799_, _34733_, _06369_);
  and _84267_ (_34800_, _34799_, _34798_);
  or _84268_ (_34801_, _34800_, _06536_);
  or _84269_ (_34802_, _34801_, _34797_);
  nand _84270_ (_34803_, _11260_, _07973_);
  and _84271_ (_34805_, _34803_, _34730_);
  or _84272_ (_34806_, _34805_, _07240_);
  and _84273_ (_34807_, _34806_, _07242_);
  and _84274_ (_34808_, _34807_, _34802_);
  or _84275_ (_34809_, _14666_, _13705_);
  and _84276_ (_34810_, _34733_, _06375_);
  and _84277_ (_34811_, _34810_, _34809_);
  or _84278_ (_34812_, _34811_, _06545_);
  or _84279_ (_34813_, _34812_, _34808_);
  nor _84280_ (_34814_, _34728_, _07234_);
  nand _84281_ (_34816_, _34814_, _34803_);
  and _84282_ (_34817_, _34816_, _09056_);
  and _84283_ (_34818_, _34817_, _34813_);
  or _84284_ (_34819_, _34732_, _08341_);
  and _84285_ (_34820_, _34733_, _06366_);
  and _84286_ (_34821_, _34820_, _34819_);
  or _84287_ (_34822_, _34821_, _06528_);
  or _84288_ (_34823_, _34822_, _34818_);
  and _84289_ (_34824_, _34823_, _34731_);
  or _84290_ (_34825_, _34824_, _06568_);
  or _84291_ (_34827_, _34742_, _06926_);
  and _84292_ (_34828_, _34827_, _05928_);
  and _84293_ (_34829_, _34828_, _34825_);
  and _84294_ (_34830_, _34766_, _05927_);
  or _84295_ (_34831_, _34830_, _06278_);
  or _84296_ (_34832_, _34831_, _34829_);
  or _84297_ (_34833_, _34728_, _06279_);
  or _84298_ (_34834_, _34833_, _34740_);
  and _84299_ (_34835_, _34834_, _01347_);
  and _84300_ (_34836_, _34835_, _34832_);
  or _84301_ (_34838_, _34836_, _34726_);
  and _84302_ (_43314_, _34838_, _42618_);
  and _84303_ (_34839_, _01351_, \oc8051_golden_model_1.SCON [2]);
  and _84304_ (_34840_, _13705_, \oc8051_golden_model_1.SCON [2]);
  nor _84305_ (_34841_, _13705_, _07776_);
  or _84306_ (_34842_, _34841_, _34840_);
  or _84307_ (_34843_, _34842_, _07215_);
  and _84308_ (_34844_, _34842_, _06461_);
  and _84309_ (_34845_, _13714_, \oc8051_golden_model_1.SCON [2]);
  and _84310_ (_34846_, _14774_, _08622_);
  or _84311_ (_34848_, _34846_, _34845_);
  or _84312_ (_34849_, _34848_, _06273_);
  and _84313_ (_34850_, _14770_, _07973_);
  or _84314_ (_34851_, _34850_, _34840_);
  and _84315_ (_34852_, _34851_, _06341_);
  and _84316_ (_34853_, _07142_, \oc8051_golden_model_1.SCON [2]);
  and _84317_ (_34854_, _07973_, \oc8051_golden_model_1.ACC [2]);
  or _84318_ (_34855_, _34854_, _34840_);
  and _84319_ (_34856_, _34855_, _07141_);
  or _84320_ (_34857_, _34856_, _34853_);
  and _84321_ (_34859_, _34857_, _07151_);
  or _84322_ (_34860_, _34859_, _06272_);
  or _84323_ (_34861_, _34860_, _34852_);
  and _84324_ (_34862_, _34861_, _34849_);
  and _84325_ (_34863_, _34862_, _07166_);
  or _84326_ (_34864_, _34863_, _34844_);
  or _84327_ (_34865_, _34864_, _06464_);
  or _84328_ (_34866_, _34855_, _06465_);
  and _84329_ (_34867_, _34866_, _06269_);
  and _84330_ (_34868_, _34867_, _34865_);
  and _84331_ (_34870_, _14756_, _08622_);
  or _84332_ (_34871_, _34870_, _34845_);
  and _84333_ (_34872_, _34871_, _06268_);
  or _84334_ (_34873_, _34872_, _06261_);
  or _84335_ (_34874_, _34873_, _34868_);
  or _84336_ (_34875_, _34845_, _14789_);
  and _84337_ (_34876_, _34875_, _34848_);
  or _84338_ (_34877_, _34876_, _06262_);
  and _84339_ (_34878_, _34877_, _06258_);
  and _84340_ (_34879_, _34878_, _34874_);
  and _84341_ (_34881_, _14804_, _08622_);
  or _84342_ (_34882_, _34881_, _34845_);
  and _84343_ (_34883_, _34882_, _06257_);
  or _84344_ (_34884_, _34883_, _10080_);
  or _84345_ (_34885_, _34884_, _34879_);
  and _84346_ (_34886_, _34885_, _34843_);
  or _84347_ (_34887_, _34886_, _07460_);
  and _84348_ (_34888_, _09450_, _07973_);
  or _84349_ (_34889_, _34840_, _07208_);
  or _84350_ (_34890_, _34889_, _34888_);
  and _84351_ (_34892_, _34890_, _05982_);
  and _84352_ (_34893_, _34892_, _34887_);
  and _84353_ (_34894_, _14859_, _07973_);
  or _84354_ (_34895_, _34894_, _34840_);
  and _84355_ (_34896_, _34895_, _10094_);
  or _84356_ (_34897_, _34896_, _06218_);
  or _84357_ (_34898_, _34897_, _34893_);
  and _84358_ (_34899_, _07973_, _08973_);
  or _84359_ (_34900_, _34899_, _34840_);
  or _84360_ (_34901_, _34900_, _06219_);
  and _84361_ (_34903_, _34901_, _34898_);
  or _84362_ (_34904_, _34903_, _06369_);
  and _84363_ (_34905_, _14751_, _07973_);
  or _84364_ (_34906_, _34905_, _34840_);
  or _84365_ (_34907_, _34906_, _07237_);
  and _84366_ (_34908_, _34907_, _07240_);
  and _84367_ (_34909_, _34908_, _34904_);
  and _84368_ (_34910_, _11259_, _07973_);
  or _84369_ (_34911_, _34910_, _34840_);
  and _84370_ (_34912_, _34911_, _06536_);
  or _84371_ (_34914_, _34912_, _34909_);
  and _84372_ (_34915_, _34914_, _07242_);
  or _84373_ (_34916_, _34840_, _08440_);
  and _84374_ (_34917_, _34900_, _06375_);
  and _84375_ (_34918_, _34917_, _34916_);
  or _84376_ (_34919_, _34918_, _34915_);
  and _84377_ (_34920_, _34919_, _07234_);
  and _84378_ (_34921_, _34855_, _06545_);
  and _84379_ (_34922_, _34921_, _34916_);
  or _84380_ (_34923_, _34922_, _06366_);
  or _84381_ (_34925_, _34923_, _34920_);
  and _84382_ (_34926_, _14748_, _07973_);
  or _84383_ (_34927_, _34840_, _09056_);
  or _84384_ (_34928_, _34927_, _34926_);
  and _84385_ (_34929_, _34928_, _09061_);
  and _84386_ (_34930_, _34929_, _34925_);
  nor _84387_ (_34931_, _11258_, _13705_);
  or _84388_ (_34932_, _34931_, _34840_);
  and _84389_ (_34933_, _34932_, _06528_);
  or _84390_ (_34934_, _34933_, _06568_);
  or _84391_ (_34936_, _34934_, _34930_);
  or _84392_ (_34937_, _34851_, _06926_);
  and _84393_ (_34938_, _34937_, _05928_);
  and _84394_ (_34939_, _34938_, _34936_);
  and _84395_ (_34940_, _34871_, _05927_);
  or _84396_ (_34941_, _34940_, _06278_);
  or _84397_ (_34942_, _34941_, _34939_);
  and _84398_ (_34943_, _14926_, _07973_);
  or _84399_ (_34944_, _34840_, _06279_);
  or _84400_ (_34945_, _34944_, _34943_);
  and _84401_ (_34947_, _34945_, _01347_);
  and _84402_ (_34948_, _34947_, _34942_);
  or _84403_ (_34949_, _34948_, _34839_);
  and _84404_ (_43315_, _34949_, _42618_);
  and _84405_ (_34950_, _01351_, \oc8051_golden_model_1.SCON [3]);
  and _84406_ (_34951_, _13705_, \oc8051_golden_model_1.SCON [3]);
  nor _84407_ (_34952_, _13705_, _07594_);
  or _84408_ (_34953_, _34952_, _34951_);
  or _84409_ (_34954_, _34953_, _07215_);
  and _84410_ (_34955_, _14953_, _07973_);
  or _84411_ (_34957_, _34955_, _34951_);
  or _84412_ (_34958_, _34957_, _07151_);
  and _84413_ (_34959_, _07973_, \oc8051_golden_model_1.ACC [3]);
  or _84414_ (_34960_, _34959_, _34951_);
  and _84415_ (_34961_, _34960_, _07141_);
  and _84416_ (_34962_, _07142_, \oc8051_golden_model_1.SCON [3]);
  or _84417_ (_34963_, _34962_, _06341_);
  or _84418_ (_34964_, _34963_, _34961_);
  and _84419_ (_34965_, _34964_, _06273_);
  and _84420_ (_34966_, _34965_, _34958_);
  and _84421_ (_34968_, _13714_, \oc8051_golden_model_1.SCON [3]);
  and _84422_ (_34969_, _14950_, _08622_);
  or _84423_ (_34970_, _34969_, _34968_);
  and _84424_ (_34971_, _34970_, _06272_);
  or _84425_ (_34972_, _34971_, _06461_);
  or _84426_ (_34973_, _34972_, _34966_);
  or _84427_ (_34974_, _34953_, _07166_);
  and _84428_ (_34975_, _34974_, _34973_);
  or _84429_ (_34976_, _34975_, _06464_);
  or _84430_ (_34977_, _34960_, _06465_);
  and _84431_ (_34979_, _34977_, _06269_);
  and _84432_ (_34980_, _34979_, _34976_);
  and _84433_ (_34981_, _14948_, _08622_);
  or _84434_ (_34982_, _34981_, _34968_);
  and _84435_ (_34983_, _34982_, _06268_);
  or _84436_ (_34984_, _34983_, _06261_);
  or _84437_ (_34985_, _34984_, _34980_);
  or _84438_ (_34986_, _34968_, _14979_);
  and _84439_ (_34987_, _34986_, _34970_);
  or _84440_ (_34988_, _34987_, _06262_);
  and _84441_ (_34990_, _34988_, _06258_);
  and _84442_ (_34991_, _34990_, _34985_);
  or _84443_ (_34992_, _34968_, _14992_);
  and _84444_ (_34993_, _34992_, _06257_);
  and _84445_ (_34994_, _34993_, _34970_);
  or _84446_ (_34995_, _34994_, _10080_);
  or _84447_ (_34996_, _34995_, _34991_);
  and _84448_ (_34997_, _34996_, _34954_);
  or _84449_ (_34998_, _34997_, _07460_);
  and _84450_ (_34999_, _09449_, _07973_);
  or _84451_ (_35001_, _34951_, _07208_);
  or _84452_ (_35002_, _35001_, _34999_);
  and _84453_ (_35003_, _35002_, _05982_);
  and _84454_ (_35004_, _35003_, _34998_);
  and _84455_ (_35005_, _15048_, _07973_);
  or _84456_ (_35006_, _35005_, _34951_);
  and _84457_ (_35007_, _35006_, _10094_);
  or _84458_ (_35008_, _35007_, _06218_);
  or _84459_ (_35009_, _35008_, _35004_);
  and _84460_ (_35010_, _07973_, _08930_);
  or _84461_ (_35012_, _35010_, _34951_);
  or _84462_ (_35013_, _35012_, _06219_);
  and _84463_ (_35014_, _35013_, _35009_);
  or _84464_ (_35015_, _35014_, _06369_);
  and _84465_ (_35016_, _14943_, _07973_);
  or _84466_ (_35017_, _35016_, _34951_);
  or _84467_ (_35018_, _35017_, _07237_);
  and _84468_ (_35019_, _35018_, _07240_);
  and _84469_ (_35020_, _35019_, _35015_);
  and _84470_ (_35021_, _12577_, _07973_);
  or _84471_ (_35023_, _35021_, _34951_);
  and _84472_ (_35024_, _35023_, _06536_);
  or _84473_ (_35025_, _35024_, _35020_);
  and _84474_ (_35026_, _35025_, _07242_);
  or _84475_ (_35027_, _34951_, _08292_);
  and _84476_ (_35028_, _35012_, _06375_);
  and _84477_ (_35029_, _35028_, _35027_);
  or _84478_ (_35030_, _35029_, _35026_);
  and _84479_ (_35031_, _35030_, _07234_);
  and _84480_ (_35032_, _34960_, _06545_);
  and _84481_ (_35034_, _35032_, _35027_);
  or _84482_ (_35035_, _35034_, _06366_);
  or _84483_ (_35036_, _35035_, _35031_);
  and _84484_ (_35037_, _14940_, _07973_);
  or _84485_ (_35038_, _34951_, _09056_);
  or _84486_ (_35039_, _35038_, _35037_);
  and _84487_ (_35040_, _35039_, _09061_);
  and _84488_ (_35041_, _35040_, _35036_);
  nor _84489_ (_35042_, _11256_, _13705_);
  or _84490_ (_35043_, _35042_, _34951_);
  and _84491_ (_35045_, _35043_, _06528_);
  or _84492_ (_35046_, _35045_, _06568_);
  or _84493_ (_35047_, _35046_, _35041_);
  or _84494_ (_35048_, _34957_, _06926_);
  and _84495_ (_35049_, _35048_, _05928_);
  and _84496_ (_35050_, _35049_, _35047_);
  and _84497_ (_35051_, _34982_, _05927_);
  or _84498_ (_35052_, _35051_, _06278_);
  or _84499_ (_35053_, _35052_, _35050_);
  and _84500_ (_35054_, _15128_, _07973_);
  or _84501_ (_35056_, _34951_, _06279_);
  or _84502_ (_35057_, _35056_, _35054_);
  and _84503_ (_35058_, _35057_, _01347_);
  and _84504_ (_35059_, _35058_, _35053_);
  or _84505_ (_35060_, _35059_, _34950_);
  and _84506_ (_43316_, _35060_, _42618_);
  and _84507_ (_35061_, _01351_, \oc8051_golden_model_1.SCON [4]);
  and _84508_ (_35062_, _13705_, \oc8051_golden_model_1.SCON [4]);
  nor _84509_ (_35063_, _08541_, _13705_);
  or _84510_ (_35064_, _35063_, _35062_);
  or _84511_ (_35066_, _35064_, _07215_);
  and _84512_ (_35067_, _13714_, \oc8051_golden_model_1.SCON [4]);
  and _84513_ (_35068_, _15176_, _08622_);
  or _84514_ (_35069_, _35068_, _35067_);
  and _84515_ (_35070_, _35069_, _06268_);
  and _84516_ (_35071_, _15162_, _07973_);
  or _84517_ (_35072_, _35071_, _35062_);
  or _84518_ (_35073_, _35072_, _07151_);
  and _84519_ (_35074_, _07973_, \oc8051_golden_model_1.ACC [4]);
  or _84520_ (_35075_, _35074_, _35062_);
  and _84521_ (_35077_, _35075_, _07141_);
  and _84522_ (_35078_, _07142_, \oc8051_golden_model_1.SCON [4]);
  or _84523_ (_35079_, _35078_, _06341_);
  or _84524_ (_35080_, _35079_, _35077_);
  and _84525_ (_35081_, _35080_, _06273_);
  and _84526_ (_35082_, _35081_, _35073_);
  and _84527_ (_35083_, _15166_, _08622_);
  or _84528_ (_35084_, _35083_, _35067_);
  and _84529_ (_35085_, _35084_, _06272_);
  or _84530_ (_35086_, _35085_, _06461_);
  or _84531_ (_35088_, _35086_, _35082_);
  or _84532_ (_35089_, _35064_, _07166_);
  and _84533_ (_35090_, _35089_, _35088_);
  or _84534_ (_35091_, _35090_, _06464_);
  or _84535_ (_35092_, _35075_, _06465_);
  and _84536_ (_35093_, _35092_, _06269_);
  and _84537_ (_35094_, _35093_, _35091_);
  or _84538_ (_35095_, _35094_, _35070_);
  and _84539_ (_35096_, _35095_, _06262_);
  or _84540_ (_35097_, _35067_, _15183_);
  and _84541_ (_35099_, _35097_, _06261_);
  and _84542_ (_35100_, _35099_, _35084_);
  or _84543_ (_35101_, _35100_, _35096_);
  and _84544_ (_35102_, _35101_, _06258_);
  and _84545_ (_35103_, _15200_, _08622_);
  or _84546_ (_35104_, _35103_, _35067_);
  and _84547_ (_35105_, _35104_, _06257_);
  or _84548_ (_35106_, _35105_, _10080_);
  or _84549_ (_35107_, _35106_, _35102_);
  and _84550_ (_35108_, _35107_, _35066_);
  or _84551_ (_35110_, _35108_, _07460_);
  and _84552_ (_35111_, _09448_, _07973_);
  or _84553_ (_35112_, _35062_, _07208_);
  or _84554_ (_35113_, _35112_, _35111_);
  and _84555_ (_35114_, _35113_, _05982_);
  and _84556_ (_35115_, _35114_, _35110_);
  and _84557_ (_35116_, _15254_, _07973_);
  or _84558_ (_35117_, _35116_, _35062_);
  and _84559_ (_35118_, _35117_, _10094_);
  or _84560_ (_35119_, _35118_, _06218_);
  or _84561_ (_35121_, _35119_, _35115_);
  and _84562_ (_35122_, _08959_, _07973_);
  or _84563_ (_35123_, _35122_, _35062_);
  or _84564_ (_35124_, _35123_, _06219_);
  and _84565_ (_35125_, _35124_, _35121_);
  or _84566_ (_35126_, _35125_, _06369_);
  and _84567_ (_35127_, _15269_, _07973_);
  or _84568_ (_35128_, _35127_, _35062_);
  or _84569_ (_35129_, _35128_, _07237_);
  and _84570_ (_35130_, _35129_, _07240_);
  and _84571_ (_35132_, _35130_, _35126_);
  and _84572_ (_35133_, _11254_, _07973_);
  or _84573_ (_35134_, _35133_, _35062_);
  and _84574_ (_35135_, _35134_, _06536_);
  or _84575_ (_35136_, _35135_, _35132_);
  and _84576_ (_35137_, _35136_, _07242_);
  or _84577_ (_35138_, _35062_, _08544_);
  and _84578_ (_35139_, _35123_, _06375_);
  and _84579_ (_35140_, _35139_, _35138_);
  or _84580_ (_35141_, _35140_, _35137_);
  and _84581_ (_35143_, _35141_, _07234_);
  and _84582_ (_35144_, _35075_, _06545_);
  and _84583_ (_35145_, _35144_, _35138_);
  or _84584_ (_35146_, _35145_, _06366_);
  or _84585_ (_35147_, _35146_, _35143_);
  and _84586_ (_35148_, _15266_, _07973_);
  or _84587_ (_35149_, _35062_, _09056_);
  or _84588_ (_35150_, _35149_, _35148_);
  and _84589_ (_35151_, _35150_, _09061_);
  and _84590_ (_35152_, _35151_, _35147_);
  nor _84591_ (_35154_, _11253_, _13705_);
  or _84592_ (_35155_, _35154_, _35062_);
  and _84593_ (_35156_, _35155_, _06528_);
  or _84594_ (_35157_, _35156_, _06568_);
  or _84595_ (_35158_, _35157_, _35152_);
  or _84596_ (_35159_, _35072_, _06926_);
  and _84597_ (_35160_, _35159_, _05928_);
  and _84598_ (_35161_, _35160_, _35158_);
  and _84599_ (_35162_, _35069_, _05927_);
  or _84600_ (_35163_, _35162_, _06278_);
  or _84601_ (_35165_, _35163_, _35161_);
  and _84602_ (_35166_, _15329_, _07973_);
  or _84603_ (_35167_, _35062_, _06279_);
  or _84604_ (_35168_, _35167_, _35166_);
  and _84605_ (_35169_, _35168_, _01347_);
  and _84606_ (_35170_, _35169_, _35165_);
  or _84607_ (_35171_, _35170_, _35061_);
  and _84608_ (_43317_, _35171_, _42618_);
  and _84609_ (_35172_, _01351_, \oc8051_golden_model_1.SCON [5]);
  and _84610_ (_35173_, _13705_, \oc8051_golden_model_1.SCON [5]);
  and _84611_ (_35175_, _15358_, _07973_);
  or _84612_ (_35176_, _35175_, _35173_);
  or _84613_ (_35177_, _35176_, _07151_);
  and _84614_ (_35178_, _07973_, \oc8051_golden_model_1.ACC [5]);
  or _84615_ (_35179_, _35178_, _35173_);
  and _84616_ (_35180_, _35179_, _07141_);
  and _84617_ (_35181_, _07142_, \oc8051_golden_model_1.SCON [5]);
  or _84618_ (_35182_, _35181_, _06341_);
  or _84619_ (_35183_, _35182_, _35180_);
  and _84620_ (_35184_, _35183_, _06273_);
  and _84621_ (_35186_, _35184_, _35177_);
  and _84622_ (_35187_, _13714_, \oc8051_golden_model_1.SCON [5]);
  and _84623_ (_35188_, _15372_, _08622_);
  or _84624_ (_35189_, _35188_, _35187_);
  and _84625_ (_35190_, _35189_, _06272_);
  or _84626_ (_35191_, _35190_, _06461_);
  or _84627_ (_35192_, _35191_, _35186_);
  nor _84628_ (_35193_, _08244_, _13705_);
  or _84629_ (_35194_, _35193_, _35173_);
  or _84630_ (_35195_, _35194_, _07166_);
  and _84631_ (_35197_, _35195_, _35192_);
  or _84632_ (_35198_, _35197_, _06464_);
  or _84633_ (_35199_, _35179_, _06465_);
  and _84634_ (_35200_, _35199_, _06269_);
  and _84635_ (_35201_, _35200_, _35198_);
  and _84636_ (_35202_, _15355_, _08622_);
  or _84637_ (_35203_, _35202_, _35187_);
  and _84638_ (_35204_, _35203_, _06268_);
  or _84639_ (_35205_, _35204_, _06261_);
  or _84640_ (_35206_, _35205_, _35201_);
  or _84641_ (_35208_, _35187_, _15387_);
  and _84642_ (_35209_, _35208_, _35189_);
  or _84643_ (_35210_, _35209_, _06262_);
  and _84644_ (_35211_, _35210_, _06258_);
  and _84645_ (_35212_, _35211_, _35206_);
  or _84646_ (_35213_, _35187_, _15403_);
  and _84647_ (_35214_, _35213_, _06257_);
  and _84648_ (_35215_, _35214_, _35189_);
  or _84649_ (_35216_, _35215_, _10080_);
  or _84650_ (_35217_, _35216_, _35212_);
  or _84651_ (_35219_, _35194_, _07215_);
  and _84652_ (_35220_, _35219_, _35217_);
  or _84653_ (_35221_, _35220_, _07460_);
  and _84654_ (_35222_, _09447_, _07973_);
  or _84655_ (_35223_, _35173_, _07208_);
  or _84656_ (_35224_, _35223_, _35222_);
  and _84657_ (_35225_, _35224_, _05982_);
  and _84658_ (_35226_, _35225_, _35221_);
  and _84659_ (_35227_, _15459_, _07973_);
  or _84660_ (_35228_, _35227_, _35173_);
  and _84661_ (_35230_, _35228_, _10094_);
  or _84662_ (_35231_, _35230_, _06218_);
  or _84663_ (_35232_, _35231_, _35226_);
  and _84664_ (_35233_, _08946_, _07973_);
  or _84665_ (_35234_, _35233_, _35173_);
  or _84666_ (_35235_, _35234_, _06219_);
  and _84667_ (_35236_, _35235_, _35232_);
  or _84668_ (_35237_, _35236_, _06369_);
  and _84669_ (_35238_, _15353_, _07973_);
  or _84670_ (_35239_, _35238_, _35173_);
  or _84671_ (_35241_, _35239_, _07237_);
  and _84672_ (_35242_, _35241_, _07240_);
  and _84673_ (_35243_, _35242_, _35237_);
  and _84674_ (_35244_, _11250_, _07973_);
  or _84675_ (_35245_, _35244_, _35173_);
  and _84676_ (_35246_, _35245_, _06536_);
  or _84677_ (_35247_, _35246_, _35243_);
  and _84678_ (_35248_, _35247_, _07242_);
  or _84679_ (_35249_, _35173_, _08247_);
  and _84680_ (_35250_, _35234_, _06375_);
  and _84681_ (_35252_, _35250_, _35249_);
  or _84682_ (_35253_, _35252_, _35248_);
  and _84683_ (_35254_, _35253_, _07234_);
  and _84684_ (_35255_, _35179_, _06545_);
  and _84685_ (_35256_, _35255_, _35249_);
  or _84686_ (_35257_, _35256_, _06366_);
  or _84687_ (_35258_, _35257_, _35254_);
  and _84688_ (_35259_, _15350_, _07973_);
  or _84689_ (_35260_, _35173_, _09056_);
  or _84690_ (_35261_, _35260_, _35259_);
  and _84691_ (_35263_, _35261_, _09061_);
  and _84692_ (_35264_, _35263_, _35258_);
  nor _84693_ (_35265_, _11249_, _13705_);
  or _84694_ (_35266_, _35265_, _35173_);
  and _84695_ (_35267_, _35266_, _06528_);
  or _84696_ (_35268_, _35267_, _06568_);
  or _84697_ (_35269_, _35268_, _35264_);
  or _84698_ (_35270_, _35176_, _06926_);
  and _84699_ (_35271_, _35270_, _05928_);
  and _84700_ (_35272_, _35271_, _35269_);
  and _84701_ (_35274_, _35203_, _05927_);
  or _84702_ (_35275_, _35274_, _06278_);
  or _84703_ (_35276_, _35275_, _35272_);
  and _84704_ (_35277_, _15532_, _07973_);
  or _84705_ (_35278_, _35173_, _06279_);
  or _84706_ (_35279_, _35278_, _35277_);
  and _84707_ (_35280_, _35279_, _01347_);
  and _84708_ (_35281_, _35280_, _35276_);
  or _84709_ (_35282_, _35281_, _35172_);
  and _84710_ (_43318_, _35282_, _42618_);
  and _84711_ (_35284_, _01351_, \oc8051_golden_model_1.SCON [6]);
  and _84712_ (_35285_, _13705_, \oc8051_golden_model_1.SCON [6]);
  and _84713_ (_35286_, _15554_, _07973_);
  or _84714_ (_35287_, _35286_, _35285_);
  or _84715_ (_35288_, _35287_, _07151_);
  and _84716_ (_35289_, _07973_, \oc8051_golden_model_1.ACC [6]);
  or _84717_ (_35290_, _35289_, _35285_);
  and _84718_ (_35291_, _35290_, _07141_);
  and _84719_ (_35292_, _07142_, \oc8051_golden_model_1.SCON [6]);
  or _84720_ (_35293_, _35292_, _06341_);
  or _84721_ (_35295_, _35293_, _35291_);
  and _84722_ (_35296_, _35295_, _06273_);
  and _84723_ (_35297_, _35296_, _35288_);
  and _84724_ (_35298_, _13714_, \oc8051_golden_model_1.SCON [6]);
  and _84725_ (_35299_, _15570_, _08622_);
  or _84726_ (_35300_, _35299_, _35298_);
  and _84727_ (_35301_, _35300_, _06272_);
  or _84728_ (_35302_, _35301_, _06461_);
  or _84729_ (_35303_, _35302_, _35297_);
  nor _84730_ (_35304_, _08142_, _13705_);
  or _84731_ (_35306_, _35304_, _35285_);
  or _84732_ (_35307_, _35306_, _07166_);
  and _84733_ (_35308_, _35307_, _35303_);
  or _84734_ (_35309_, _35308_, _06464_);
  or _84735_ (_35310_, _35290_, _06465_);
  and _84736_ (_35311_, _35310_, _06269_);
  and _84737_ (_35312_, _35311_, _35309_);
  and _84738_ (_35313_, _15551_, _08622_);
  or _84739_ (_35314_, _35313_, _35298_);
  and _84740_ (_35315_, _35314_, _06268_);
  or _84741_ (_35317_, _35315_, _06261_);
  or _84742_ (_35318_, _35317_, _35312_);
  or _84743_ (_35319_, _35298_, _15585_);
  and _84744_ (_35320_, _35319_, _35300_);
  or _84745_ (_35321_, _35320_, _06262_);
  and _84746_ (_35322_, _35321_, _06258_);
  and _84747_ (_35323_, _35322_, _35318_);
  and _84748_ (_35324_, _15602_, _08622_);
  or _84749_ (_35325_, _35324_, _35298_);
  and _84750_ (_35326_, _35325_, _06257_);
  or _84751_ (_35328_, _35326_, _10080_);
  or _84752_ (_35329_, _35328_, _35323_);
  or _84753_ (_35330_, _35306_, _07215_);
  and _84754_ (_35331_, _35330_, _35329_);
  or _84755_ (_35332_, _35331_, _07460_);
  and _84756_ (_35333_, _09446_, _07973_);
  or _84757_ (_35334_, _35285_, _07208_);
  or _84758_ (_35335_, _35334_, _35333_);
  and _84759_ (_35336_, _35335_, _05982_);
  and _84760_ (_35337_, _35336_, _35332_);
  and _84761_ (_35339_, _15657_, _07973_);
  or _84762_ (_35340_, _35339_, _35285_);
  and _84763_ (_35341_, _35340_, _10094_);
  or _84764_ (_35342_, _35341_, _06218_);
  or _84765_ (_35343_, _35342_, _35337_);
  and _84766_ (_35344_, _15664_, _07973_);
  or _84767_ (_35345_, _35344_, _35285_);
  or _84768_ (_35346_, _35345_, _06219_);
  and _84769_ (_35347_, _35346_, _35343_);
  or _84770_ (_35348_, _35347_, _06369_);
  and _84771_ (_35350_, _15549_, _07973_);
  or _84772_ (_35351_, _35350_, _35285_);
  or _84773_ (_35352_, _35351_, _07237_);
  and _84774_ (_35353_, _35352_, _07240_);
  and _84775_ (_35354_, _35353_, _35348_);
  and _84776_ (_35355_, _11247_, _07973_);
  or _84777_ (_35356_, _35355_, _35285_);
  and _84778_ (_35357_, _35356_, _06536_);
  or _84779_ (_35358_, _35357_, _35354_);
  and _84780_ (_35359_, _35358_, _07242_);
  or _84781_ (_35361_, _35285_, _08145_);
  and _84782_ (_35362_, _35345_, _06375_);
  and _84783_ (_35363_, _35362_, _35361_);
  or _84784_ (_35364_, _35363_, _35359_);
  and _84785_ (_35365_, _35364_, _07234_);
  and _84786_ (_35366_, _35290_, _06545_);
  and _84787_ (_35367_, _35366_, _35361_);
  or _84788_ (_35368_, _35367_, _06366_);
  or _84789_ (_35369_, _35368_, _35365_);
  and _84790_ (_35370_, _15546_, _07973_);
  or _84791_ (_35372_, _35285_, _09056_);
  or _84792_ (_35373_, _35372_, _35370_);
  and _84793_ (_35374_, _35373_, _09061_);
  and _84794_ (_35375_, _35374_, _35369_);
  nor _84795_ (_35376_, _11246_, _13705_);
  or _84796_ (_35377_, _35376_, _35285_);
  and _84797_ (_35378_, _35377_, _06528_);
  or _84798_ (_35379_, _35378_, _06568_);
  or _84799_ (_35380_, _35379_, _35375_);
  or _84800_ (_35381_, _35287_, _06926_);
  and _84801_ (_35383_, _35381_, _05928_);
  and _84802_ (_35384_, _35383_, _35380_);
  and _84803_ (_35385_, _35314_, _05927_);
  or _84804_ (_35386_, _35385_, _06278_);
  or _84805_ (_35387_, _35386_, _35384_);
  and _84806_ (_35388_, _15734_, _07973_);
  or _84807_ (_35389_, _35285_, _06279_);
  or _84808_ (_35390_, _35389_, _35388_);
  and _84809_ (_35391_, _35390_, _01347_);
  and _84810_ (_35392_, _35391_, _35387_);
  or _84811_ (_35394_, _35392_, _35284_);
  and _84812_ (_43319_, _35394_, _42618_);
  nor _84813_ (_35395_, _01347_, _06800_);
  nor _84814_ (_35396_, _07956_, _06800_);
  and _84815_ (_35397_, _07956_, \oc8051_golden_model_1.ACC [0]);
  and _84816_ (_35398_, _35397_, _08390_);
  or _84817_ (_35399_, _35398_, _35396_);
  or _84818_ (_35400_, _35399_, _07234_);
  nor _84819_ (_35401_, _08390_, _13872_);
  or _84820_ (_35402_, _35401_, _35396_);
  or _84821_ (_35404_, _35402_, _07151_);
  or _84822_ (_35405_, _35397_, _35396_);
  and _84823_ (_35406_, _35405_, _07141_);
  nor _84824_ (_35407_, _07141_, _06800_);
  or _84825_ (_35408_, _35407_, _06341_);
  or _84826_ (_35409_, _35408_, _35406_);
  and _84827_ (_35410_, _35409_, _07166_);
  nand _84828_ (_35411_, _35410_, _35404_);
  nand _84829_ (_35412_, _35411_, _06802_);
  or _84830_ (_35413_, _35405_, _06465_);
  and _84831_ (_35415_, _35413_, _07303_);
  and _84832_ (_35416_, _35415_, _35412_);
  nand _84833_ (_35417_, _07215_, _07186_);
  or _84834_ (_35418_, _35417_, _35416_);
  and _84835_ (_35419_, _08173_, _07133_);
  or _84836_ (_35420_, _35396_, _07215_);
  or _84837_ (_35421_, _35420_, _35419_);
  and _84838_ (_35422_, _35421_, _35418_);
  or _84839_ (_35423_, _35422_, _07460_);
  or _84840_ (_35424_, _35396_, _07208_);
  and _84841_ (_35426_, _09392_, _07956_);
  or _84842_ (_35427_, _35426_, _35424_);
  and _84843_ (_35428_, _35427_, _35423_);
  or _84844_ (_35429_, _35428_, _10094_);
  and _84845_ (_35430_, _14467_, _08173_);
  or _84846_ (_35431_, _35396_, _05982_);
  or _84847_ (_35432_, _35431_, _35430_);
  and _84848_ (_35433_, _35432_, _06219_);
  and _84849_ (_35434_, _35433_, _35429_);
  and _84850_ (_35435_, _07956_, _08954_);
  or _84851_ (_35437_, _35435_, _35396_);
  and _84852_ (_35438_, _35437_, _06218_);
  or _84853_ (_35439_, _35438_, _06369_);
  or _84854_ (_35440_, _35439_, _35434_);
  and _84855_ (_35441_, _14366_, _07956_);
  or _84856_ (_35442_, _35441_, _35396_);
  or _84857_ (_35443_, _35442_, _07237_);
  and _84858_ (_35444_, _35443_, _07240_);
  and _84859_ (_35445_, _35444_, _35440_);
  nor _84860_ (_35446_, _12580_, _13872_);
  or _84861_ (_35448_, _35446_, _35396_);
  nor _84862_ (_35449_, _35398_, _07240_);
  and _84863_ (_35450_, _35449_, _35448_);
  or _84864_ (_35451_, _35450_, _35445_);
  and _84865_ (_35452_, _35451_, _07242_);
  nand _84866_ (_35453_, _35437_, _06375_);
  nor _84867_ (_35454_, _35453_, _35401_);
  or _84868_ (_35455_, _35454_, _06545_);
  or _84869_ (_35456_, _35455_, _35452_);
  and _84870_ (_35457_, _35456_, _35400_);
  or _84871_ (_35459_, _35457_, _06366_);
  and _84872_ (_35460_, _14363_, _07956_);
  or _84873_ (_35461_, _35460_, _35396_);
  or _84874_ (_35462_, _35461_, _09056_);
  and _84875_ (_35463_, _35462_, _09061_);
  and _84876_ (_35464_, _35463_, _35459_);
  and _84877_ (_35465_, _35448_, _06528_);
  or _84878_ (_35466_, _35465_, _19502_);
  or _84879_ (_35467_, _35466_, _35464_);
  or _84880_ (_35468_, _35402_, _06661_);
  and _84881_ (_35470_, _35468_, _01347_);
  and _84882_ (_35471_, _35470_, _35467_);
  or _84883_ (_35472_, _35471_, _35395_);
  and _84884_ (_43321_, _35472_, _42618_);
  nand _84885_ (_35473_, _08173_, _07038_);
  or _84886_ (_35474_, _35473_, _08341_);
  or _84887_ (_35475_, _07956_, \oc8051_golden_model_1.SP [1]);
  and _84888_ (_35476_, _35475_, _06366_);
  and _84889_ (_35477_, _35476_, _35474_);
  and _84890_ (_35478_, _11260_, _08173_);
  nor _84891_ (_35479_, _07956_, _07067_);
  or _84892_ (_35480_, _35479_, _07234_);
  or _84893_ (_35481_, _35480_, _35478_);
  and _84894_ (_35482_, _14562_, _08173_);
  not _84895_ (_35483_, _35482_);
  and _84896_ (_35484_, _35483_, _35475_);
  or _84897_ (_35485_, _35484_, _07151_);
  nand _84898_ (_35486_, _06758_, \oc8051_golden_model_1.SP [1]);
  and _84899_ (_35487_, _07956_, \oc8051_golden_model_1.ACC [1]);
  or _84900_ (_35488_, _35487_, _35479_);
  and _84901_ (_35490_, _35488_, _07141_);
  nor _84902_ (_35491_, _07141_, _07067_);
  or _84903_ (_35492_, _35491_, _06758_);
  or _84904_ (_35493_, _35492_, _35490_);
  and _84905_ (_35494_, _35493_, _35486_);
  or _84906_ (_35495_, _35494_, _06341_);
  and _84907_ (_35496_, _35495_, _06010_);
  and _84908_ (_35497_, _35496_, _35485_);
  nor _84909_ (_35498_, _06010_, \oc8051_golden_model_1.SP [1]);
  or _84910_ (_35499_, _35498_, _06461_);
  or _84911_ (_35501_, _35499_, _35497_);
  nand _84912_ (_35502_, _07301_, _06461_);
  and _84913_ (_35503_, _35502_, _35501_);
  or _84914_ (_35504_, _35503_, _06464_);
  or _84915_ (_35505_, _35488_, _06465_);
  and _84916_ (_35506_, _35505_, _07303_);
  and _84917_ (_35507_, _35506_, _35504_);
  not _84918_ (_35508_, _07494_);
  or _84919_ (_35509_, _35508_, _07302_);
  or _84920_ (_35510_, _35509_, _35507_);
  or _84921_ (_35512_, _07494_, _07067_);
  and _84922_ (_35513_, _35512_, _07215_);
  and _84923_ (_35514_, _35513_, _35510_);
  nand _84924_ (_35515_, _08173_, _07357_);
  and _84925_ (_35516_, _35475_, _10080_);
  and _84926_ (_35517_, _35516_, _35515_);
  or _84927_ (_35518_, _35517_, _07460_);
  or _84928_ (_35519_, _35518_, _35514_);
  or _84929_ (_35520_, _35479_, _07208_);
  and _84930_ (_35521_, _09451_, _07956_);
  or _84931_ (_35523_, _35521_, _35520_);
  and _84932_ (_35524_, _35523_, _05982_);
  and _84933_ (_35525_, _35524_, _35519_);
  and _84934_ (_35526_, _35475_, _10094_);
  or _84935_ (_35527_, _14653_, _13872_);
  and _84936_ (_35528_, _35527_, _35526_);
  or _84937_ (_35529_, _35528_, _35525_);
  and _84938_ (_35530_, _35529_, _06219_);
  and _84939_ (_35531_, _35475_, _06218_);
  and _84940_ (_35532_, _35531_, _35473_);
  or _84941_ (_35534_, _35532_, _06217_);
  or _84942_ (_35535_, _35534_, _35530_);
  nor _84943_ (_35536_, _05952_, _07067_);
  nor _84944_ (_35537_, _35536_, _06369_);
  and _84945_ (_35538_, _35537_, _35535_);
  or _84946_ (_35539_, _14668_, _13872_);
  and _84947_ (_35540_, _35475_, _06369_);
  and _84948_ (_35541_, _35540_, _35539_);
  or _84949_ (_35542_, _35541_, _06536_);
  or _84950_ (_35543_, _35542_, _35538_);
  and _84951_ (_35545_, _11262_, _07956_);
  or _84952_ (_35546_, _35545_, _35479_);
  or _84953_ (_35547_, _35546_, _07240_);
  and _84954_ (_35548_, _35547_, _07242_);
  and _84955_ (_35549_, _35548_, _35543_);
  or _84956_ (_35550_, _14666_, _13872_);
  and _84957_ (_35551_, _35475_, _06375_);
  and _84958_ (_35552_, _35551_, _35550_);
  or _84959_ (_35553_, _35552_, _06545_);
  or _84960_ (_35554_, _35553_, _35549_);
  and _84961_ (_35556_, _35554_, _35481_);
  or _84962_ (_35557_, _35556_, _07233_);
  nor _84963_ (_35558_, _05961_, _07067_);
  nor _84964_ (_35559_, _35558_, _06366_);
  and _84965_ (_35560_, _35559_, _35557_);
  or _84966_ (_35561_, _35560_, _35477_);
  and _84967_ (_35562_, _35561_, _09061_);
  nor _84968_ (_35563_, _11261_, _13872_);
  or _84969_ (_35564_, _35563_, _35479_);
  and _84970_ (_35565_, _35564_, _06528_);
  or _84971_ (_35567_, _35565_, _06551_);
  nor _84972_ (_35568_, _35567_, _35562_);
  or _84973_ (_35569_, _35568_, _07044_);
  nor _84974_ (_35570_, _06281_, _07253_);
  nand _84975_ (_35571_, _35570_, _35569_);
  or _84976_ (_35572_, _35570_, _07067_);
  and _84977_ (_35573_, _35572_, _06926_);
  and _84978_ (_35574_, _35573_, _35571_);
  and _84979_ (_35575_, _35484_, _06568_);
  or _84980_ (_35576_, _35575_, _07695_);
  or _84981_ (_35578_, _35576_, _35574_);
  or _84982_ (_35579_, _07271_, _07067_);
  and _84983_ (_35580_, _35579_, _06279_);
  and _84984_ (_35581_, _35580_, _35578_);
  or _84985_ (_35582_, _35482_, _35479_);
  and _84986_ (_35583_, _35582_, _06278_);
  or _84987_ (_35584_, _35583_, _01351_);
  or _84988_ (_35585_, _35584_, _35581_);
  or _84989_ (_35586_, _01347_, \oc8051_golden_model_1.SP [1]);
  and _84990_ (_35587_, _35586_, _42618_);
  and _84991_ (_43322_, _35587_, _35585_);
  nor _84992_ (_35589_, _01347_, _06715_);
  or _84993_ (_35590_, _07866_, _05952_);
  nor _84994_ (_35591_, _13872_, _07776_);
  nor _84995_ (_35592_, _07956_, _06715_);
  or _84996_ (_35593_, _35592_, _07215_);
  or _84997_ (_35594_, _35593_, _35591_);
  or _84998_ (_35595_, _07866_, _06007_);
  and _84999_ (_35596_, _35595_, _05978_);
  and _85000_ (_35597_, _14770_, _08173_);
  or _85001_ (_35599_, _35597_, _35592_);
  and _85002_ (_35600_, _35599_, _06341_);
  and _85003_ (_35601_, _07956_, \oc8051_golden_model_1.ACC [2]);
  or _85004_ (_35602_, _35601_, _35592_);
  and _85005_ (_35603_, _35602_, _07141_);
  nor _85006_ (_35604_, _07141_, _06715_);
  or _85007_ (_35605_, _35604_, _06758_);
  or _85008_ (_35606_, _35605_, _35603_);
  nand _85009_ (_35607_, _16081_, _06758_);
  and _85010_ (_35608_, _35607_, _07151_);
  and _85011_ (_35610_, _35608_, _35606_);
  or _85012_ (_35611_, _35610_, _27826_);
  or _85013_ (_35612_, _35611_, _35600_);
  or _85014_ (_35613_, _07866_, _06010_);
  nand _85015_ (_35614_, _08684_, _06461_);
  and _85016_ (_35615_, _35614_, _35613_);
  and _85017_ (_35616_, _35615_, _35612_);
  or _85018_ (_35617_, _35616_, _06464_);
  or _85019_ (_35618_, _35602_, _06465_);
  and _85020_ (_35619_, _35618_, _07303_);
  and _85021_ (_35621_, _35619_, _35617_);
  or _85022_ (_35622_, _07720_, _12613_);
  or _85023_ (_35623_, _35622_, _35621_);
  and _85024_ (_35624_, _35623_, _35596_);
  or _85025_ (_35625_, _16081_, _05978_);
  nand _85026_ (_35626_, _35625_, _07215_);
  or _85027_ (_35627_, _35626_, _35624_);
  and _85028_ (_35628_, _35627_, _35594_);
  or _85029_ (_35629_, _35628_, _07460_);
  or _85030_ (_35630_, _35592_, _07208_);
  and _85031_ (_35632_, _09450_, _07956_);
  or _85032_ (_35633_, _35632_, _35630_);
  and _85033_ (_35634_, _35633_, _05982_);
  and _85034_ (_35635_, _35634_, _35629_);
  and _85035_ (_35636_, _14859_, _07956_);
  or _85036_ (_35637_, _35636_, _35592_);
  and _85037_ (_35638_, _35637_, _10094_);
  or _85038_ (_35639_, _35638_, _06218_);
  or _85039_ (_35640_, _35639_, _35635_);
  and _85040_ (_35641_, _07956_, _08973_);
  or _85041_ (_35643_, _35641_, _35592_);
  or _85042_ (_35644_, _35643_, _06219_);
  and _85043_ (_35645_, _35644_, _35640_);
  or _85044_ (_35646_, _35645_, _06217_);
  and _85045_ (_35647_, _35646_, _35590_);
  or _85046_ (_35648_, _35647_, _06369_);
  and _85047_ (_35649_, _14751_, _07956_);
  or _85048_ (_35650_, _35649_, _35592_);
  or _85049_ (_35651_, _35650_, _07237_);
  and _85050_ (_35652_, _35651_, _07240_);
  and _85051_ (_35654_, _35652_, _35648_);
  and _85052_ (_35655_, _11259_, _07956_);
  or _85053_ (_35656_, _35655_, _35592_);
  and _85054_ (_35657_, _35656_, _06536_);
  or _85055_ (_35658_, _35657_, _35654_);
  and _85056_ (_35659_, _35658_, _07242_);
  or _85057_ (_35660_, _35592_, _08440_);
  and _85058_ (_35661_, _35643_, _06375_);
  and _85059_ (_35662_, _35661_, _35660_);
  or _85060_ (_35663_, _35662_, _35659_);
  and _85061_ (_35665_, _35663_, _12772_);
  and _85062_ (_35666_, _35602_, _06545_);
  and _85063_ (_35667_, _35666_, _35660_);
  nor _85064_ (_35668_, _16081_, _05961_);
  or _85065_ (_35669_, _35668_, _06366_);
  or _85066_ (_35670_, _35669_, _35667_);
  or _85067_ (_35671_, _35670_, _35665_);
  and _85068_ (_35672_, _14748_, _07956_);
  or _85069_ (_35673_, _35672_, _35592_);
  or _85070_ (_35674_, _35673_, _09056_);
  and _85071_ (_35676_, _35674_, _35671_);
  or _85072_ (_35677_, _35676_, _06528_);
  nor _85073_ (_35678_, _11258_, _13872_);
  or _85074_ (_35679_, _35678_, _35592_);
  or _85075_ (_35680_, _35679_, _09061_);
  and _85076_ (_35681_, _35680_, _06716_);
  and _85077_ (_35682_, _35681_, _35677_);
  and _85078_ (_35683_, _16081_, _06551_);
  or _85079_ (_35684_, _35683_, _07253_);
  or _85080_ (_35685_, _35684_, _35682_);
  nor _85081_ (_35687_, _07866_, _05959_);
  nor _85082_ (_35688_, _35687_, _06281_);
  and _85083_ (_35689_, _35688_, _35685_);
  and _85084_ (_35690_, _16081_, _06281_);
  or _85085_ (_35691_, _35690_, _06568_);
  or _85086_ (_35692_, _35691_, _35689_);
  or _85087_ (_35693_, _35599_, _06926_);
  and _85088_ (_35694_, _35693_, _07271_);
  and _85089_ (_35695_, _35694_, _35692_);
  nor _85090_ (_35696_, _16081_, _07271_);
  or _85091_ (_35698_, _35696_, _06278_);
  or _85092_ (_35699_, _35698_, _35695_);
  and _85093_ (_35700_, _14926_, _08173_);
  or _85094_ (_35701_, _35592_, _06279_);
  or _85095_ (_35702_, _35701_, _35700_);
  and _85096_ (_35703_, _35702_, _01347_);
  and _85097_ (_35704_, _35703_, _35699_);
  or _85098_ (_35705_, _35704_, _35589_);
  and _85099_ (_43323_, _35705_, _42618_);
  nor _85100_ (_35706_, _01347_, _06460_);
  or _85101_ (_35708_, _07869_, _07271_);
  or _85102_ (_35709_, _07869_, _05959_);
  or _85103_ (_35710_, _07869_, _05952_);
  nor _85104_ (_35711_, _13872_, _07594_);
  nor _85105_ (_35712_, _07956_, _06460_);
  or _85106_ (_35713_, _35712_, _07460_);
  or _85107_ (_35714_, _35713_, _35711_);
  and _85108_ (_35715_, _35714_, _12659_);
  and _85109_ (_35716_, _14953_, _08173_);
  or _85110_ (_35717_, _35716_, _35712_);
  or _85111_ (_35719_, _35717_, _07151_);
  and _85112_ (_35720_, _07956_, \oc8051_golden_model_1.ACC [3]);
  or _85113_ (_35721_, _35720_, _35712_);
  or _85114_ (_35722_, _35721_, _07142_);
  or _85115_ (_35723_, _07141_, \oc8051_golden_model_1.SP [3]);
  and _85116_ (_35724_, _35723_, _07504_);
  and _85117_ (_35725_, _35724_, _35722_);
  and _85118_ (_35726_, _07869_, _06758_);
  or _85119_ (_35727_, _35726_, _06341_);
  or _85120_ (_35728_, _35727_, _35725_);
  and _85121_ (_35730_, _35728_, _06010_);
  and _85122_ (_35731_, _35730_, _35719_);
  nor _85123_ (_35732_, _15897_, _06010_);
  or _85124_ (_35733_, _35732_, _06461_);
  or _85125_ (_35734_, _35733_, _35731_);
  nand _85126_ (_35735_, _08674_, _06461_);
  and _85127_ (_35736_, _35735_, _35734_);
  or _85128_ (_35737_, _35736_, _06464_);
  or _85129_ (_35738_, _35721_, _06465_);
  and _85130_ (_35739_, _35738_, _07303_);
  and _85131_ (_35741_, _35739_, _35737_);
  or _85132_ (_35742_, _07652_, _35508_);
  or _85133_ (_35743_, _35742_, _35741_);
  or _85134_ (_35744_, _07869_, _07494_);
  and _85135_ (_35745_, _35744_, _07215_);
  and _85136_ (_35746_, _35745_, _35743_);
  or _85137_ (_35747_, _35746_, _35715_);
  or _85138_ (_35748_, _35712_, _07208_);
  and _85139_ (_35749_, _09449_, _07956_);
  or _85140_ (_35750_, _35749_, _35748_);
  and _85141_ (_35752_, _35750_, _05982_);
  and _85142_ (_35753_, _35752_, _35747_);
  and _85143_ (_35754_, _15048_, _07956_);
  or _85144_ (_35755_, _35754_, _35712_);
  and _85145_ (_35756_, _35755_, _10094_);
  or _85146_ (_35757_, _35756_, _06218_);
  or _85147_ (_35758_, _35757_, _35753_);
  and _85148_ (_35759_, _07956_, _08930_);
  or _85149_ (_35760_, _35759_, _35712_);
  or _85150_ (_35761_, _35760_, _06219_);
  and _85151_ (_35763_, _35761_, _35758_);
  or _85152_ (_35764_, _35763_, _06217_);
  and _85153_ (_35765_, _35764_, _35710_);
  or _85154_ (_35766_, _35765_, _06369_);
  and _85155_ (_35767_, _14943_, _07956_);
  or _85156_ (_35768_, _35767_, _35712_);
  or _85157_ (_35769_, _35768_, _07237_);
  and _85158_ (_35770_, _35769_, _07240_);
  and _85159_ (_35771_, _35770_, _35766_);
  and _85160_ (_35772_, _12577_, _07956_);
  or _85161_ (_35774_, _35772_, _35712_);
  and _85162_ (_35775_, _35774_, _06536_);
  or _85163_ (_35776_, _35775_, _35771_);
  and _85164_ (_35777_, _35776_, _07242_);
  or _85165_ (_35778_, _35712_, _08292_);
  and _85166_ (_35779_, _35760_, _06375_);
  and _85167_ (_35780_, _35779_, _35778_);
  or _85168_ (_35781_, _35780_, _35777_);
  and _85169_ (_35782_, _35781_, _12772_);
  and _85170_ (_35783_, _35721_, _06545_);
  and _85171_ (_35785_, _35783_, _35778_);
  nor _85172_ (_35786_, _15897_, _05961_);
  or _85173_ (_35787_, _35786_, _06366_);
  or _85174_ (_35788_, _35787_, _35785_);
  or _85175_ (_35789_, _35788_, _35782_);
  and _85176_ (_35790_, _14940_, _08173_);
  or _85177_ (_35791_, _35712_, _09056_);
  or _85178_ (_35792_, _35791_, _35790_);
  and _85179_ (_35793_, _35792_, _35789_);
  or _85180_ (_35794_, _35793_, _06528_);
  nor _85181_ (_35796_, _11256_, _13872_);
  or _85182_ (_35797_, _35796_, _35712_);
  or _85183_ (_35798_, _35797_, _09061_);
  and _85184_ (_35799_, _35798_, _06716_);
  and _85185_ (_35800_, _35799_, _35794_);
  nor _85186_ (_35801_, _08671_, _06460_);
  or _85187_ (_35802_, _35801_, _08672_);
  and _85188_ (_35803_, _35802_, _06551_);
  or _85189_ (_35804_, _35803_, _07253_);
  or _85190_ (_35805_, _35804_, _35800_);
  and _85191_ (_35807_, _35805_, _35709_);
  or _85192_ (_35808_, _35807_, _06281_);
  or _85193_ (_35809_, _35802_, _06282_);
  and _85194_ (_35810_, _35809_, _06926_);
  and _85195_ (_35811_, _35810_, _35808_);
  and _85196_ (_35812_, _35717_, _06568_);
  or _85197_ (_35813_, _35812_, _07695_);
  or _85198_ (_35814_, _35813_, _35811_);
  and _85199_ (_35815_, _35814_, _35708_);
  or _85200_ (_35816_, _35815_, _06278_);
  and _85201_ (_35818_, _15128_, _08173_);
  or _85202_ (_35819_, _35712_, _06279_);
  or _85203_ (_35820_, _35819_, _35818_);
  and _85204_ (_35821_, _35820_, _01347_);
  and _85205_ (_35822_, _35821_, _35816_);
  or _85206_ (_35823_, _35822_, _35706_);
  and _85207_ (_43325_, _35823_, _42618_);
  nor _85208_ (_35824_, _01347_, _13845_);
  nor _85209_ (_35825_, _07602_, \oc8051_golden_model_1.SP [4]);
  nor _85210_ (_35826_, _35825_, _13814_);
  or _85211_ (_35828_, _35826_, _07271_);
  nor _85212_ (_35829_, _08541_, _13872_);
  nor _85213_ (_35830_, _07956_, _13845_);
  or _85214_ (_35831_, _35830_, _07460_);
  or _85215_ (_35832_, _35831_, _35829_);
  and _85216_ (_35833_, _35832_, _12659_);
  and _85217_ (_35834_, _15162_, _08173_);
  or _85218_ (_35835_, _35834_, _35830_);
  or _85219_ (_35836_, _35835_, _07151_);
  and _85220_ (_35837_, _07956_, \oc8051_golden_model_1.ACC [4]);
  or _85221_ (_35839_, _35837_, _35830_);
  or _85222_ (_35840_, _35839_, _07142_);
  or _85223_ (_35841_, _07141_, \oc8051_golden_model_1.SP [4]);
  and _85224_ (_35842_, _35841_, _07504_);
  and _85225_ (_35843_, _35842_, _35840_);
  and _85226_ (_35844_, _35826_, _06758_);
  or _85227_ (_35845_, _35844_, _06341_);
  or _85228_ (_35846_, _35845_, _35843_);
  and _85229_ (_35847_, _35846_, _06010_);
  and _85230_ (_35848_, _35847_, _35836_);
  and _85231_ (_35850_, _35826_, _07611_);
  or _85232_ (_35851_, _35850_, _06461_);
  or _85233_ (_35852_, _35851_, _35848_);
  and _85234_ (_35853_, _13846_, _06800_);
  nor _85235_ (_35854_, _08673_, _13845_);
  nor _85236_ (_35855_, _35854_, _35853_);
  nand _85237_ (_35856_, _35855_, _06461_);
  and _85238_ (_35857_, _35856_, _35852_);
  or _85239_ (_35858_, _35857_, _06464_);
  or _85240_ (_35859_, _35839_, _06465_);
  and _85241_ (_35861_, _35859_, _07303_);
  and _85242_ (_35862_, _35861_, _35858_);
  and _85243_ (_35863_, _07603_, \oc8051_golden_model_1.SP [4]);
  nor _85244_ (_35864_, _07603_, \oc8051_golden_model_1.SP [4]);
  nor _85245_ (_35865_, _35864_, _35863_);
  nand _85246_ (_35866_, _35865_, _06267_);
  nand _85247_ (_35867_, _35866_, _07494_);
  or _85248_ (_35868_, _35867_, _35862_);
  or _85249_ (_35869_, _35826_, _07494_);
  and _85250_ (_35870_, _35869_, _07215_);
  and _85251_ (_35872_, _35870_, _35868_);
  or _85252_ (_35873_, _35872_, _35833_);
  or _85253_ (_35874_, _35830_, _07208_);
  and _85254_ (_35875_, _09448_, _07956_);
  or _85255_ (_35876_, _35875_, _35874_);
  and _85256_ (_35877_, _35876_, _05982_);
  and _85257_ (_35878_, _35877_, _35873_);
  and _85258_ (_35879_, _15254_, _07956_);
  or _85259_ (_35880_, _35879_, _35830_);
  and _85260_ (_35881_, _35880_, _10094_);
  or _85261_ (_35883_, _35881_, _06218_);
  or _85262_ (_35884_, _35883_, _35878_);
  and _85263_ (_35885_, _08959_, _07956_);
  or _85264_ (_35886_, _35885_, _35830_);
  or _85265_ (_35887_, _35886_, _06219_);
  and _85266_ (_35888_, _35887_, _35884_);
  or _85267_ (_35889_, _35888_, _06217_);
  or _85268_ (_35890_, _35826_, _05952_);
  and _85269_ (_35891_, _35890_, _35889_);
  or _85270_ (_35892_, _35891_, _06369_);
  and _85271_ (_35894_, _15269_, _07956_);
  or _85272_ (_35895_, _35894_, _35830_);
  or _85273_ (_35896_, _35895_, _07237_);
  and _85274_ (_35897_, _35896_, _07240_);
  and _85275_ (_35898_, _35897_, _35892_);
  and _85276_ (_35899_, _11254_, _07956_);
  or _85277_ (_35900_, _35899_, _35830_);
  and _85278_ (_35901_, _35900_, _06536_);
  or _85279_ (_35902_, _35901_, _35898_);
  and _85280_ (_35903_, _35902_, _07242_);
  or _85281_ (_35905_, _35830_, _08544_);
  and _85282_ (_35906_, _35886_, _06375_);
  and _85283_ (_35907_, _35906_, _35905_);
  or _85284_ (_35908_, _35907_, _35903_);
  and _85285_ (_35909_, _35908_, _12772_);
  and _85286_ (_35910_, _35839_, _06545_);
  and _85287_ (_35911_, _35910_, _35905_);
  and _85288_ (_35912_, _35826_, _07233_);
  or _85289_ (_35913_, _35912_, _06366_);
  or _85290_ (_35914_, _35913_, _35911_);
  or _85291_ (_35916_, _35914_, _35909_);
  and _85292_ (_35917_, _15266_, _07956_);
  or _85293_ (_35918_, _35917_, _35830_);
  or _85294_ (_35919_, _35918_, _09056_);
  and _85295_ (_35920_, _35919_, _35916_);
  or _85296_ (_35921_, _35920_, _06528_);
  nor _85297_ (_35922_, _11253_, _13872_);
  or _85298_ (_35923_, _35922_, _35830_);
  or _85299_ (_35924_, _35923_, _09061_);
  and _85300_ (_35925_, _35924_, _06716_);
  and _85301_ (_35927_, _35925_, _35921_);
  nor _85302_ (_35928_, _08672_, _13845_);
  or _85303_ (_35929_, _35928_, _13846_);
  and _85304_ (_35930_, _35929_, _06551_);
  or _85305_ (_35931_, _35930_, _07253_);
  or _85306_ (_35932_, _35931_, _35927_);
  or _85307_ (_35933_, _35826_, _05959_);
  and _85308_ (_35934_, _35933_, _35932_);
  or _85309_ (_35935_, _35934_, _06281_);
  or _85310_ (_35936_, _35929_, _06282_);
  and _85311_ (_35938_, _35936_, _06926_);
  and _85312_ (_35939_, _35938_, _35935_);
  and _85313_ (_35940_, _35835_, _06568_);
  or _85314_ (_35941_, _35940_, _07695_);
  or _85315_ (_35942_, _35941_, _35939_);
  and _85316_ (_35943_, _35942_, _35828_);
  or _85317_ (_35944_, _35943_, _06278_);
  and _85318_ (_35945_, _15329_, _08173_);
  or _85319_ (_35946_, _35830_, _06279_);
  or _85320_ (_35947_, _35946_, _35945_);
  and _85321_ (_35949_, _35947_, _01347_);
  and _85322_ (_35950_, _35949_, _35944_);
  or _85323_ (_35951_, _35950_, _35824_);
  and _85324_ (_43326_, _35951_, _42618_);
  nor _85325_ (_35952_, _01347_, _13844_);
  nor _85326_ (_35953_, _13814_, \oc8051_golden_model_1.SP [5]);
  nor _85327_ (_35954_, _35953_, _13815_);
  or _85328_ (_35955_, _35954_, _07271_);
  nor _85329_ (_35956_, _08244_, _13872_);
  nor _85330_ (_35957_, _07956_, _13844_);
  or _85331_ (_35959_, _35957_, _07460_);
  or _85332_ (_35960_, _35959_, _35956_);
  and _85333_ (_35961_, _35960_, _12659_);
  and _85334_ (_35962_, _15358_, _08173_);
  or _85335_ (_35963_, _35962_, _35957_);
  or _85336_ (_35964_, _35963_, _07151_);
  and _85337_ (_35965_, _07956_, \oc8051_golden_model_1.ACC [5]);
  or _85338_ (_35966_, _35965_, _35957_);
  and _85339_ (_35967_, _35966_, _07141_);
  nor _85340_ (_35968_, _07141_, _13844_);
  or _85341_ (_35970_, _35968_, _06758_);
  or _85342_ (_35971_, _35970_, _35967_);
  or _85343_ (_35972_, _35954_, _07504_);
  and _85344_ (_35973_, _35972_, _35971_);
  or _85345_ (_35974_, _35973_, _06341_);
  and _85346_ (_35975_, _35974_, _06010_);
  and _85347_ (_35976_, _35975_, _35964_);
  and _85348_ (_35977_, _35954_, _07611_);
  or _85349_ (_35978_, _35977_, _06461_);
  or _85350_ (_35979_, _35978_, _35976_);
  and _85351_ (_35981_, _13847_, _06800_);
  nor _85352_ (_35982_, _35853_, _13844_);
  nor _85353_ (_35983_, _35982_, _35981_);
  nand _85354_ (_35984_, _35983_, _06461_);
  and _85355_ (_35985_, _35984_, _35979_);
  or _85356_ (_35986_, _35985_, _06464_);
  or _85357_ (_35987_, _35966_, _06465_);
  and _85358_ (_35988_, _35987_, _07303_);
  and _85359_ (_35989_, _35988_, _35986_);
  nor _85360_ (_35990_, _35863_, \oc8051_golden_model_1.SP [5]);
  nor _85361_ (_35992_, _35990_, _13859_);
  nand _85362_ (_35993_, _35992_, _06267_);
  nand _85363_ (_35994_, _35993_, _07494_);
  or _85364_ (_35995_, _35994_, _35989_);
  or _85365_ (_35996_, _35954_, _07494_);
  and _85366_ (_35997_, _35996_, _07215_);
  and _85367_ (_35998_, _35997_, _35995_);
  or _85368_ (_35999_, _35998_, _35961_);
  or _85369_ (_36000_, _35957_, _07208_);
  and _85370_ (_36001_, _09447_, _07956_);
  or _85371_ (_36003_, _36001_, _36000_);
  and _85372_ (_36004_, _36003_, _05982_);
  and _85373_ (_36005_, _36004_, _35999_);
  and _85374_ (_36006_, _15459_, _07956_);
  or _85375_ (_36007_, _36006_, _35957_);
  and _85376_ (_36008_, _36007_, _10094_);
  or _85377_ (_36009_, _36008_, _06218_);
  or _85378_ (_36010_, _36009_, _36005_);
  and _85379_ (_36011_, _08946_, _07956_);
  or _85380_ (_36012_, _36011_, _35957_);
  or _85381_ (_36014_, _36012_, _06219_);
  and _85382_ (_36015_, _36014_, _36010_);
  or _85383_ (_36016_, _36015_, _06217_);
  or _85384_ (_36017_, _35954_, _05952_);
  and _85385_ (_36018_, _36017_, _36016_);
  or _85386_ (_36019_, _36018_, _06369_);
  and _85387_ (_36020_, _15353_, _07956_);
  or _85388_ (_36021_, _36020_, _35957_);
  or _85389_ (_36022_, _36021_, _07237_);
  and _85390_ (_36023_, _36022_, _07240_);
  and _85391_ (_36025_, _36023_, _36019_);
  and _85392_ (_36026_, _11250_, _07956_);
  or _85393_ (_36027_, _36026_, _35957_);
  and _85394_ (_36028_, _36027_, _06536_);
  or _85395_ (_36029_, _36028_, _36025_);
  and _85396_ (_36030_, _36029_, _07242_);
  or _85397_ (_36031_, _35957_, _08247_);
  and _85398_ (_36032_, _36012_, _06375_);
  and _85399_ (_36033_, _36032_, _36031_);
  or _85400_ (_36034_, _36033_, _36030_);
  and _85401_ (_36036_, _36034_, _12772_);
  and _85402_ (_36037_, _35966_, _06545_);
  and _85403_ (_36038_, _36037_, _36031_);
  and _85404_ (_36039_, _35954_, _07233_);
  or _85405_ (_36040_, _36039_, _06366_);
  or _85406_ (_36041_, _36040_, _36038_);
  or _85407_ (_36042_, _36041_, _36036_);
  and _85408_ (_36043_, _15350_, _07956_);
  or _85409_ (_36044_, _36043_, _35957_);
  or _85410_ (_36045_, _36044_, _09056_);
  and _85411_ (_36047_, _36045_, _36042_);
  or _85412_ (_36048_, _36047_, _06528_);
  nor _85413_ (_36049_, _11249_, _13872_);
  or _85414_ (_36050_, _36049_, _35957_);
  or _85415_ (_36051_, _36050_, _09061_);
  and _85416_ (_36052_, _36051_, _06716_);
  and _85417_ (_36053_, _36052_, _36048_);
  nor _85418_ (_36054_, _13846_, _13844_);
  or _85419_ (_36055_, _36054_, _13847_);
  and _85420_ (_36056_, _36055_, _06551_);
  or _85421_ (_36058_, _36056_, _07253_);
  or _85422_ (_36059_, _36058_, _36053_);
  or _85423_ (_36060_, _35954_, _05959_);
  and _85424_ (_36061_, _36060_, _36059_);
  or _85425_ (_36062_, _36061_, _06281_);
  or _85426_ (_36063_, _36055_, _06282_);
  and _85427_ (_36064_, _36063_, _06926_);
  and _85428_ (_36065_, _36064_, _36062_);
  and _85429_ (_36066_, _35963_, _06568_);
  or _85430_ (_36067_, _36066_, _07695_);
  or _85431_ (_36069_, _36067_, _36065_);
  and _85432_ (_36070_, _36069_, _35955_);
  or _85433_ (_36071_, _36070_, _06278_);
  and _85434_ (_36072_, _15532_, _08173_);
  or _85435_ (_36073_, _35957_, _06279_);
  or _85436_ (_36074_, _36073_, _36072_);
  and _85437_ (_36075_, _36074_, _01347_);
  and _85438_ (_36076_, _36075_, _36071_);
  or _85439_ (_36077_, _36076_, _35952_);
  and _85440_ (_43327_, _36077_, _42618_);
  nor _85441_ (_36079_, _01347_, _13843_);
  nor _85442_ (_36080_, _07956_, _13843_);
  and _85443_ (_36081_, _15554_, _08173_);
  or _85444_ (_36082_, _36081_, _36080_);
  or _85445_ (_36083_, _36082_, _07151_);
  and _85446_ (_36084_, _07956_, \oc8051_golden_model_1.ACC [6]);
  or _85447_ (_36085_, _36084_, _36080_);
  and _85448_ (_36086_, _36085_, _07141_);
  nor _85449_ (_36087_, _07141_, _13843_);
  or _85450_ (_36088_, _36087_, _06758_);
  or _85451_ (_36090_, _36088_, _36086_);
  nor _85452_ (_36091_, _13815_, \oc8051_golden_model_1.SP [6]);
  nor _85453_ (_36092_, _36091_, _13816_);
  or _85454_ (_36093_, _36092_, _07504_);
  and _85455_ (_36094_, _36093_, _36090_);
  or _85456_ (_36095_, _36094_, _06341_);
  and _85457_ (_36096_, _36095_, _06010_);
  and _85458_ (_36097_, _36096_, _36083_);
  and _85459_ (_36098_, _36092_, _07611_);
  or _85460_ (_36099_, _36098_, _06461_);
  or _85461_ (_36101_, _36099_, _36097_);
  nor _85462_ (_36102_, _35981_, _13843_);
  nor _85463_ (_36103_, _36102_, _13849_);
  nand _85464_ (_36104_, _36103_, _06461_);
  and _85465_ (_36105_, _36104_, _36101_);
  or _85466_ (_36106_, _36105_, _06464_);
  or _85467_ (_36107_, _36085_, _06465_);
  and _85468_ (_36108_, _36107_, _07303_);
  and _85469_ (_36109_, _36108_, _36106_);
  nor _85470_ (_36110_, _13859_, \oc8051_golden_model_1.SP [6]);
  nor _85471_ (_36112_, _36110_, _13860_);
  and _85472_ (_36113_, _36112_, _06267_);
  or _85473_ (_36114_, _36113_, _36109_);
  and _85474_ (_36115_, _36114_, _07494_);
  nand _85475_ (_36116_, _36092_, _35508_);
  nand _85476_ (_36117_, _36116_, _07215_);
  or _85477_ (_36118_, _36117_, _36115_);
  nor _85478_ (_36119_, _08142_, _13872_);
  or _85479_ (_36120_, _36080_, _07215_);
  or _85480_ (_36121_, _36120_, _36119_);
  and _85481_ (_36123_, _36121_, _36118_);
  or _85482_ (_36124_, _36123_, _07460_);
  and _85483_ (_36125_, _09446_, _07956_);
  or _85484_ (_36126_, _36080_, _07208_);
  or _85485_ (_36127_, _36126_, _36125_);
  and _85486_ (_36128_, _36127_, _05982_);
  and _85487_ (_36129_, _36128_, _36124_);
  and _85488_ (_36130_, _15657_, _08173_);
  or _85489_ (_36131_, _36130_, _36080_);
  and _85490_ (_36132_, _36131_, _10094_);
  or _85491_ (_36134_, _36132_, _06218_);
  or _85492_ (_36135_, _36134_, _36129_);
  and _85493_ (_36136_, _15664_, _07956_);
  or _85494_ (_36137_, _36136_, _36080_);
  or _85495_ (_36138_, _36137_, _06219_);
  and _85496_ (_36139_, _36138_, _36135_);
  or _85497_ (_36140_, _36139_, _06217_);
  or _85498_ (_36141_, _36092_, _05952_);
  and _85499_ (_36142_, _36141_, _36140_);
  or _85500_ (_36143_, _36142_, _06369_);
  and _85501_ (_36145_, _15549_, _07956_);
  or _85502_ (_36146_, _36145_, _36080_);
  or _85503_ (_36147_, _36146_, _07237_);
  and _85504_ (_36148_, _36147_, _07240_);
  and _85505_ (_36149_, _36148_, _36143_);
  and _85506_ (_36150_, _11247_, _07956_);
  or _85507_ (_36151_, _36150_, _36080_);
  and _85508_ (_36152_, _36151_, _06536_);
  or _85509_ (_36153_, _36152_, _36149_);
  and _85510_ (_36154_, _36153_, _07242_);
  or _85511_ (_36156_, _36080_, _08145_);
  and _85512_ (_36157_, _36137_, _06375_);
  and _85513_ (_36158_, _36157_, _36156_);
  or _85514_ (_36159_, _36158_, _36154_);
  and _85515_ (_36160_, _36159_, _12772_);
  and _85516_ (_36161_, _36085_, _06545_);
  and _85517_ (_36162_, _36161_, _36156_);
  and _85518_ (_36163_, _36092_, _07233_);
  or _85519_ (_36164_, _36163_, _06366_);
  or _85520_ (_36165_, _36164_, _36162_);
  or _85521_ (_36167_, _36165_, _36160_);
  and _85522_ (_36168_, _15546_, _07956_);
  or _85523_ (_36169_, _36168_, _36080_);
  or _85524_ (_36170_, _36169_, _09056_);
  and _85525_ (_36171_, _36170_, _36167_);
  or _85526_ (_36172_, _36171_, _06528_);
  nor _85527_ (_36173_, _11246_, _13872_);
  or _85528_ (_36174_, _36173_, _36080_);
  or _85529_ (_36175_, _36174_, _09061_);
  and _85530_ (_36176_, _36175_, _06716_);
  and _85531_ (_36178_, _36176_, _36172_);
  nor _85532_ (_36179_, _13847_, _13843_);
  or _85533_ (_36180_, _36179_, _13848_);
  and _85534_ (_36181_, _36180_, _06551_);
  or _85535_ (_36182_, _36181_, _07253_);
  or _85536_ (_36183_, _36182_, _36178_);
  nor _85537_ (_36184_, _36092_, _05959_);
  nor _85538_ (_36185_, _36184_, _06281_);
  and _85539_ (_36186_, _36185_, _36183_);
  and _85540_ (_36187_, _36180_, _06281_);
  or _85541_ (_36189_, _36187_, _06568_);
  or _85542_ (_36190_, _36189_, _36186_);
  or _85543_ (_36191_, _36082_, _06926_);
  and _85544_ (_36192_, _36191_, _07271_);
  and _85545_ (_36193_, _36192_, _36190_);
  and _85546_ (_36194_, _36092_, _07695_);
  or _85547_ (_36195_, _36194_, _06278_);
  or _85548_ (_36196_, _36195_, _36193_);
  and _85549_ (_36197_, _15734_, _08173_);
  or _85550_ (_36198_, _36080_, _06279_);
  or _85551_ (_36200_, _36198_, _36197_);
  and _85552_ (_36201_, _36200_, _01347_);
  and _85553_ (_36202_, _36201_, _36196_);
  or _85554_ (_36203_, _36202_, _36079_);
  and _85555_ (_43328_, _36203_, _42618_);
  not _85556_ (_36204_, \oc8051_golden_model_1.SBUF [0]);
  nor _85557_ (_36205_, _01347_, _36204_);
  nand _85558_ (_36206_, _11263_, _07886_);
  nor _85559_ (_36207_, _07886_, _36204_);
  nor _85560_ (_36208_, _36207_, _07234_);
  nand _85561_ (_36210_, _36208_, _36206_);
  and _85562_ (_36211_, _07886_, \oc8051_golden_model_1.ACC [0]);
  or _85563_ (_36212_, _36211_, _36207_);
  and _85564_ (_36213_, _36212_, _06464_);
  or _85565_ (_36214_, _36213_, _10080_);
  nor _85566_ (_36215_, _08390_, _13951_);
  or _85567_ (_36216_, _36215_, _36207_);
  and _85568_ (_36217_, _36216_, _06341_);
  nor _85569_ (_36218_, _07141_, _36204_);
  and _85570_ (_36219_, _36212_, _07141_);
  or _85571_ (_36220_, _36219_, _36218_);
  and _85572_ (_36221_, _36220_, _07151_);
  or _85573_ (_36222_, _36221_, _06461_);
  or _85574_ (_36223_, _36222_, _36217_);
  and _85575_ (_36224_, _36223_, _06465_);
  or _85576_ (_36225_, _36224_, _36214_);
  and _85577_ (_36226_, _07886_, _07133_);
  or _85578_ (_36227_, _36207_, _22611_);
  or _85579_ (_36228_, _36227_, _36226_);
  and _85580_ (_36229_, _36228_, _36225_);
  or _85581_ (_36231_, _36229_, _07460_);
  and _85582_ (_36232_, _09392_, _07886_);
  or _85583_ (_36233_, _36207_, _07208_);
  or _85584_ (_36234_, _36233_, _36232_);
  and _85585_ (_36235_, _36234_, _36231_);
  or _85586_ (_36236_, _36235_, _10094_);
  and _85587_ (_36237_, _14467_, _07886_);
  or _85588_ (_36238_, _36207_, _05982_);
  or _85589_ (_36239_, _36238_, _36237_);
  and _85590_ (_36240_, _36239_, _06219_);
  and _85591_ (_36242_, _36240_, _36236_);
  and _85592_ (_36243_, _07886_, _08954_);
  or _85593_ (_36244_, _36243_, _36207_);
  and _85594_ (_36245_, _36244_, _06218_);
  or _85595_ (_36246_, _36245_, _06369_);
  or _85596_ (_36247_, _36246_, _36242_);
  and _85597_ (_36248_, _14366_, _07886_);
  or _85598_ (_36249_, _36248_, _36207_);
  or _85599_ (_36250_, _36249_, _07237_);
  and _85600_ (_36251_, _36250_, _07240_);
  and _85601_ (_36253_, _36251_, _36247_);
  nor _85602_ (_36254_, _12580_, _13951_);
  or _85603_ (_36255_, _36254_, _36207_);
  and _85604_ (_36256_, _36206_, _06536_);
  and _85605_ (_36257_, _36256_, _36255_);
  or _85606_ (_36258_, _36257_, _36253_);
  and _85607_ (_36259_, _36258_, _07242_);
  nand _85608_ (_36260_, _36244_, _06375_);
  nor _85609_ (_36261_, _36260_, _36215_);
  or _85610_ (_36262_, _36261_, _06545_);
  or _85611_ (_36264_, _36262_, _36259_);
  and _85612_ (_36265_, _36264_, _36210_);
  or _85613_ (_36266_, _36265_, _06366_);
  and _85614_ (_36267_, _14363_, _07886_);
  or _85615_ (_36268_, _36207_, _09056_);
  or _85616_ (_36269_, _36268_, _36267_);
  and _85617_ (_36270_, _36269_, _09061_);
  and _85618_ (_36271_, _36270_, _36266_);
  and _85619_ (_36272_, _36255_, _06528_);
  or _85620_ (_36273_, _36272_, _19502_);
  or _85621_ (_36275_, _36273_, _36271_);
  or _85622_ (_36276_, _36216_, _06661_);
  and _85623_ (_36277_, _36276_, _01347_);
  and _85624_ (_36278_, _36277_, _36275_);
  or _85625_ (_36279_, _36278_, _36205_);
  and _85626_ (_43330_, _36279_, _42618_);
  not _85627_ (_36280_, \oc8051_golden_model_1.SBUF [1]);
  nor _85628_ (_36281_, _01347_, _36280_);
  nand _85629_ (_36282_, _07886_, _07038_);
  or _85630_ (_36283_, _07886_, \oc8051_golden_model_1.SBUF [1]);
  and _85631_ (_36285_, _36283_, _06218_);
  and _85632_ (_36286_, _36285_, _36282_);
  nor _85633_ (_36287_, _07886_, _36280_);
  nor _85634_ (_36288_, _13951_, _07357_);
  or _85635_ (_36289_, _36288_, _36287_);
  or _85636_ (_36290_, _36289_, _07215_);
  and _85637_ (_36291_, _14562_, _07886_);
  not _85638_ (_36292_, _36291_);
  and _85639_ (_36293_, _36292_, _36283_);
  or _85640_ (_36294_, _36293_, _07151_);
  and _85641_ (_36296_, _07886_, \oc8051_golden_model_1.ACC [1]);
  or _85642_ (_36297_, _36296_, _36287_);
  and _85643_ (_36298_, _36297_, _07141_);
  nor _85644_ (_36299_, _07141_, _36280_);
  or _85645_ (_36300_, _36299_, _06341_);
  or _85646_ (_36301_, _36300_, _36298_);
  and _85647_ (_36302_, _36301_, _07166_);
  and _85648_ (_36303_, _36302_, _36294_);
  and _85649_ (_36304_, _36289_, _06461_);
  or _85650_ (_36305_, _36304_, _36303_);
  and _85651_ (_36307_, _36305_, _06465_);
  and _85652_ (_36308_, _36297_, _06464_);
  or _85653_ (_36309_, _36308_, _10080_);
  or _85654_ (_36310_, _36309_, _36307_);
  and _85655_ (_36311_, _36310_, _36290_);
  or _85656_ (_36312_, _36311_, _07460_);
  and _85657_ (_36313_, _09451_, _07886_);
  or _85658_ (_36314_, _36287_, _07208_);
  or _85659_ (_36315_, _36314_, _36313_);
  and _85660_ (_36316_, _36315_, _05982_);
  and _85661_ (_36318_, _36316_, _36312_);
  or _85662_ (_36319_, _14653_, _13951_);
  and _85663_ (_36320_, _36283_, _10094_);
  and _85664_ (_36321_, _36320_, _36319_);
  or _85665_ (_36322_, _36321_, _36318_);
  and _85666_ (_36323_, _36322_, _06219_);
  or _85667_ (_36324_, _36323_, _36286_);
  and _85668_ (_36325_, _36324_, _07237_);
  or _85669_ (_36326_, _14668_, _13951_);
  and _85670_ (_36327_, _36283_, _06369_);
  and _85671_ (_36329_, _36327_, _36326_);
  or _85672_ (_36330_, _36329_, _06536_);
  or _85673_ (_36331_, _36330_, _36325_);
  nor _85674_ (_36332_, _11261_, _13951_);
  or _85675_ (_36333_, _36332_, _36287_);
  nand _85676_ (_36334_, _11260_, _07886_);
  and _85677_ (_36335_, _36334_, _36333_);
  or _85678_ (_36336_, _36335_, _07240_);
  and _85679_ (_36337_, _36336_, _07242_);
  and _85680_ (_36338_, _36337_, _36331_);
  or _85681_ (_36340_, _14666_, _13951_);
  and _85682_ (_36341_, _36283_, _06375_);
  and _85683_ (_36342_, _36341_, _36340_);
  or _85684_ (_36343_, _36342_, _06545_);
  or _85685_ (_36344_, _36343_, _36338_);
  nor _85686_ (_36345_, _36287_, _07234_);
  nand _85687_ (_36346_, _36345_, _36334_);
  and _85688_ (_36347_, _36346_, _09056_);
  and _85689_ (_36348_, _36347_, _36344_);
  or _85690_ (_36349_, _36282_, _08341_);
  and _85691_ (_36351_, _36283_, _06366_);
  and _85692_ (_36352_, _36351_, _36349_);
  or _85693_ (_36353_, _36352_, _06528_);
  or _85694_ (_36354_, _36353_, _36348_);
  or _85695_ (_36355_, _36333_, _09061_);
  and _85696_ (_36356_, _36355_, _06926_);
  and _85697_ (_36357_, _36356_, _36354_);
  and _85698_ (_36358_, _36293_, _06568_);
  or _85699_ (_36359_, _36358_, _06278_);
  or _85700_ (_36360_, _36359_, _36357_);
  or _85701_ (_36362_, _36287_, _06279_);
  or _85702_ (_36363_, _36362_, _36291_);
  and _85703_ (_36364_, _36363_, _01347_);
  and _85704_ (_36365_, _36364_, _36360_);
  or _85705_ (_36366_, _36365_, _36281_);
  and _85706_ (_43331_, _36366_, _42618_);
  and _85707_ (_36367_, _01351_, \oc8051_golden_model_1.SBUF [2]);
  and _85708_ (_36368_, _13951_, \oc8051_golden_model_1.SBUF [2]);
  and _85709_ (_36369_, _09450_, _07886_);
  or _85710_ (_36370_, _36369_, _36368_);
  and _85711_ (_36372_, _36370_, _07460_);
  and _85712_ (_36373_, _14770_, _07886_);
  or _85713_ (_36374_, _36373_, _36368_);
  or _85714_ (_36375_, _36374_, _07151_);
  and _85715_ (_36376_, _07886_, \oc8051_golden_model_1.ACC [2]);
  or _85716_ (_36377_, _36376_, _36368_);
  and _85717_ (_36378_, _36377_, _07141_);
  and _85718_ (_36379_, _07142_, \oc8051_golden_model_1.SBUF [2]);
  or _85719_ (_36380_, _36379_, _06341_);
  or _85720_ (_36381_, _36380_, _36378_);
  and _85721_ (_36383_, _36381_, _07166_);
  and _85722_ (_36384_, _36383_, _36375_);
  nor _85723_ (_36385_, _13951_, _07776_);
  or _85724_ (_36386_, _36385_, _36368_);
  and _85725_ (_36387_, _36386_, _06461_);
  or _85726_ (_36388_, _36387_, _36384_);
  and _85727_ (_36389_, _36388_, _06465_);
  and _85728_ (_36390_, _36377_, _06464_);
  or _85729_ (_36391_, _36390_, _10080_);
  or _85730_ (_36392_, _36391_, _36389_);
  or _85731_ (_36394_, _36386_, _07215_);
  and _85732_ (_36395_, _36394_, _07208_);
  and _85733_ (_36396_, _36395_, _36392_);
  or _85734_ (_36397_, _36396_, _10094_);
  or _85735_ (_36398_, _36397_, _36372_);
  and _85736_ (_36399_, _14859_, _07886_);
  or _85737_ (_36400_, _36368_, _05982_);
  or _85738_ (_36401_, _36400_, _36399_);
  and _85739_ (_36402_, _36401_, _06219_);
  and _85740_ (_36403_, _36402_, _36398_);
  and _85741_ (_36405_, _07886_, _08973_);
  or _85742_ (_36406_, _36405_, _36368_);
  and _85743_ (_36407_, _36406_, _06218_);
  or _85744_ (_36408_, _36407_, _06369_);
  or _85745_ (_36409_, _36408_, _36403_);
  and _85746_ (_36410_, _14751_, _07886_);
  or _85747_ (_36411_, _36410_, _36368_);
  or _85748_ (_36412_, _36411_, _07237_);
  and _85749_ (_36413_, _36412_, _07240_);
  and _85750_ (_36414_, _36413_, _36409_);
  and _85751_ (_36416_, _11259_, _07886_);
  or _85752_ (_36417_, _36416_, _36368_);
  and _85753_ (_36418_, _36417_, _06536_);
  or _85754_ (_36419_, _36418_, _36414_);
  and _85755_ (_36420_, _36419_, _07242_);
  or _85756_ (_36421_, _36368_, _08440_);
  and _85757_ (_36422_, _36406_, _06375_);
  and _85758_ (_36423_, _36422_, _36421_);
  or _85759_ (_36424_, _36423_, _36420_);
  and _85760_ (_36425_, _36424_, _07234_);
  and _85761_ (_36427_, _36377_, _06545_);
  and _85762_ (_36428_, _36427_, _36421_);
  or _85763_ (_36429_, _36428_, _06366_);
  or _85764_ (_36430_, _36429_, _36425_);
  and _85765_ (_36431_, _14748_, _07886_);
  or _85766_ (_36432_, _36368_, _09056_);
  or _85767_ (_36433_, _36432_, _36431_);
  and _85768_ (_36434_, _36433_, _09061_);
  and _85769_ (_36435_, _36434_, _36430_);
  nor _85770_ (_36436_, _11258_, _13951_);
  or _85771_ (_36438_, _36436_, _36368_);
  and _85772_ (_36439_, _36438_, _06528_);
  or _85773_ (_36440_, _36439_, _36435_);
  and _85774_ (_36441_, _36440_, _06926_);
  and _85775_ (_36442_, _36374_, _06568_);
  or _85776_ (_36443_, _36442_, _06278_);
  or _85777_ (_36444_, _36443_, _36441_);
  and _85778_ (_36445_, _14926_, _07886_);
  or _85779_ (_36446_, _36368_, _06279_);
  or _85780_ (_36447_, _36446_, _36445_);
  and _85781_ (_36449_, _36447_, _01347_);
  and _85782_ (_36450_, _36449_, _36444_);
  or _85783_ (_36451_, _36450_, _36367_);
  and _85784_ (_43332_, _36451_, _42618_);
  and _85785_ (_36452_, _01351_, \oc8051_golden_model_1.SBUF [3]);
  and _85786_ (_36453_, _13951_, \oc8051_golden_model_1.SBUF [3]);
  and _85787_ (_36454_, _14953_, _07886_);
  or _85788_ (_36455_, _36454_, _36453_);
  or _85789_ (_36456_, _36455_, _07151_);
  and _85790_ (_36457_, _07886_, \oc8051_golden_model_1.ACC [3]);
  or _85791_ (_36459_, _36457_, _36453_);
  and _85792_ (_36460_, _36459_, _07141_);
  and _85793_ (_36461_, _07142_, \oc8051_golden_model_1.SBUF [3]);
  or _85794_ (_36462_, _36461_, _06341_);
  or _85795_ (_36463_, _36462_, _36460_);
  and _85796_ (_36464_, _36463_, _07166_);
  and _85797_ (_36465_, _36464_, _36456_);
  nor _85798_ (_36466_, _13951_, _07594_);
  or _85799_ (_36467_, _36466_, _36453_);
  and _85800_ (_36468_, _36467_, _06461_);
  or _85801_ (_36470_, _36468_, _36465_);
  and _85802_ (_36471_, _36470_, _06465_);
  and _85803_ (_36472_, _36459_, _06464_);
  or _85804_ (_36473_, _36472_, _10080_);
  or _85805_ (_36474_, _36473_, _36471_);
  or _85806_ (_36475_, _36467_, _07215_);
  and _85807_ (_36476_, _36475_, _36474_);
  or _85808_ (_36477_, _36476_, _07460_);
  and _85809_ (_36478_, _09449_, _07886_);
  or _85810_ (_36479_, _36453_, _07208_);
  or _85811_ (_36481_, _36479_, _36478_);
  and _85812_ (_36482_, _36481_, _05982_);
  and _85813_ (_36483_, _36482_, _36477_);
  and _85814_ (_36484_, _15048_, _07886_);
  or _85815_ (_36485_, _36484_, _36453_);
  and _85816_ (_36486_, _36485_, _10094_);
  or _85817_ (_36487_, _36486_, _06218_);
  or _85818_ (_36488_, _36487_, _36483_);
  and _85819_ (_36489_, _07886_, _08930_);
  or _85820_ (_36490_, _36489_, _36453_);
  or _85821_ (_36492_, _36490_, _06219_);
  and _85822_ (_36493_, _36492_, _36488_);
  or _85823_ (_36494_, _36493_, _06369_);
  and _85824_ (_36495_, _14943_, _07886_);
  or _85825_ (_36496_, _36495_, _36453_);
  or _85826_ (_36497_, _36496_, _07237_);
  and _85827_ (_36498_, _36497_, _07240_);
  and _85828_ (_36499_, _36498_, _36494_);
  and _85829_ (_36500_, _12577_, _07886_);
  or _85830_ (_36501_, _36500_, _36453_);
  and _85831_ (_36503_, _36501_, _06536_);
  or _85832_ (_36504_, _36503_, _36499_);
  and _85833_ (_36505_, _36504_, _07242_);
  or _85834_ (_36506_, _36453_, _08292_);
  and _85835_ (_36507_, _36490_, _06375_);
  and _85836_ (_36508_, _36507_, _36506_);
  or _85837_ (_36509_, _36508_, _36505_);
  and _85838_ (_36510_, _36509_, _07234_);
  and _85839_ (_36511_, _36459_, _06545_);
  and _85840_ (_36512_, _36511_, _36506_);
  or _85841_ (_36514_, _36512_, _06366_);
  or _85842_ (_36515_, _36514_, _36510_);
  and _85843_ (_36516_, _14940_, _07886_);
  or _85844_ (_36517_, _36453_, _09056_);
  or _85845_ (_36518_, _36517_, _36516_);
  and _85846_ (_36519_, _36518_, _09061_);
  and _85847_ (_36520_, _36519_, _36515_);
  nor _85848_ (_36521_, _11256_, _13951_);
  or _85849_ (_36522_, _36521_, _36453_);
  and _85850_ (_36523_, _36522_, _06528_);
  or _85851_ (_36525_, _36523_, _36520_);
  and _85852_ (_36526_, _36525_, _06926_);
  and _85853_ (_36527_, _36455_, _06568_);
  or _85854_ (_36528_, _36527_, _06278_);
  or _85855_ (_36529_, _36528_, _36526_);
  and _85856_ (_36530_, _15128_, _07886_);
  or _85857_ (_36531_, _36453_, _06279_);
  or _85858_ (_36532_, _36531_, _36530_);
  and _85859_ (_36533_, _36532_, _01347_);
  and _85860_ (_36534_, _36533_, _36529_);
  or _85861_ (_36536_, _36534_, _36452_);
  and _85862_ (_43333_, _36536_, _42618_);
  and _85863_ (_36537_, _01351_, \oc8051_golden_model_1.SBUF [4]);
  and _85864_ (_36538_, _13951_, \oc8051_golden_model_1.SBUF [4]);
  nor _85865_ (_36539_, _08541_, _13951_);
  or _85866_ (_36540_, _36539_, _36538_);
  or _85867_ (_36541_, _36540_, _07215_);
  and _85868_ (_36542_, _15162_, _07886_);
  or _85869_ (_36543_, _36542_, _36538_);
  or _85870_ (_36544_, _36543_, _07151_);
  and _85871_ (_36546_, _07886_, \oc8051_golden_model_1.ACC [4]);
  or _85872_ (_36547_, _36546_, _36538_);
  and _85873_ (_36548_, _36547_, _07141_);
  and _85874_ (_36549_, _07142_, \oc8051_golden_model_1.SBUF [4]);
  or _85875_ (_36550_, _36549_, _06341_);
  or _85876_ (_36551_, _36550_, _36548_);
  and _85877_ (_36552_, _36551_, _07166_);
  and _85878_ (_36553_, _36552_, _36544_);
  and _85879_ (_36554_, _36540_, _06461_);
  or _85880_ (_36555_, _36554_, _36553_);
  and _85881_ (_36557_, _36555_, _06465_);
  and _85882_ (_36558_, _36547_, _06464_);
  or _85883_ (_36559_, _36558_, _10080_);
  or _85884_ (_36560_, _36559_, _36557_);
  and _85885_ (_36561_, _36560_, _07208_);
  and _85886_ (_36562_, _36561_, _36541_);
  and _85887_ (_36563_, _09448_, _07886_);
  or _85888_ (_36564_, _36563_, _36538_);
  and _85889_ (_36565_, _36564_, _07460_);
  or _85890_ (_36566_, _36565_, _10094_);
  or _85891_ (_36568_, _36566_, _36562_);
  and _85892_ (_36569_, _15254_, _07886_);
  or _85893_ (_36570_, _36538_, _05982_);
  or _85894_ (_36571_, _36570_, _36569_);
  and _85895_ (_36572_, _36571_, _06219_);
  and _85896_ (_36573_, _36572_, _36568_);
  and _85897_ (_36574_, _08959_, _07886_);
  or _85898_ (_36575_, _36574_, _36538_);
  and _85899_ (_36576_, _36575_, _06218_);
  or _85900_ (_36577_, _36576_, _06369_);
  or _85901_ (_36579_, _36577_, _36573_);
  and _85902_ (_36580_, _15269_, _07886_);
  or _85903_ (_36581_, _36580_, _36538_);
  or _85904_ (_36582_, _36581_, _07237_);
  and _85905_ (_36583_, _36582_, _07240_);
  and _85906_ (_36584_, _36583_, _36579_);
  and _85907_ (_36585_, _11254_, _07886_);
  or _85908_ (_36586_, _36585_, _36538_);
  and _85909_ (_36587_, _36586_, _06536_);
  or _85910_ (_36588_, _36587_, _36584_);
  and _85911_ (_36590_, _36588_, _07242_);
  or _85912_ (_36591_, _36538_, _08544_);
  and _85913_ (_36592_, _36575_, _06375_);
  and _85914_ (_36593_, _36592_, _36591_);
  or _85915_ (_36594_, _36593_, _36590_);
  and _85916_ (_36595_, _36594_, _07234_);
  and _85917_ (_36596_, _36547_, _06545_);
  and _85918_ (_36597_, _36596_, _36591_);
  or _85919_ (_36598_, _36597_, _06366_);
  or _85920_ (_36599_, _36598_, _36595_);
  and _85921_ (_36601_, _15266_, _07886_);
  or _85922_ (_36602_, _36538_, _09056_);
  or _85923_ (_36603_, _36602_, _36601_);
  and _85924_ (_36604_, _36603_, _09061_);
  and _85925_ (_36605_, _36604_, _36599_);
  nor _85926_ (_36606_, _11253_, _13951_);
  or _85927_ (_36607_, _36606_, _36538_);
  and _85928_ (_36608_, _36607_, _06528_);
  or _85929_ (_36609_, _36608_, _36605_);
  and _85930_ (_36610_, _36609_, _06926_);
  and _85931_ (_36612_, _36543_, _06568_);
  or _85932_ (_36613_, _36612_, _06278_);
  or _85933_ (_36614_, _36613_, _36610_);
  and _85934_ (_36615_, _15329_, _07886_);
  or _85935_ (_36616_, _36538_, _06279_);
  or _85936_ (_36617_, _36616_, _36615_);
  and _85937_ (_36618_, _36617_, _01347_);
  and _85938_ (_36619_, _36618_, _36614_);
  or _85939_ (_36620_, _36619_, _36537_);
  and _85940_ (_43334_, _36620_, _42618_);
  and _85941_ (_36622_, _01351_, \oc8051_golden_model_1.SBUF [5]);
  and _85942_ (_36623_, _13951_, \oc8051_golden_model_1.SBUF [5]);
  nor _85943_ (_36624_, _08244_, _13951_);
  or _85944_ (_36625_, _36624_, _36623_);
  or _85945_ (_36626_, _36625_, _07215_);
  and _85946_ (_36627_, _15358_, _07886_);
  or _85947_ (_36628_, _36627_, _36623_);
  or _85948_ (_36629_, _36628_, _07151_);
  and _85949_ (_36630_, _07886_, \oc8051_golden_model_1.ACC [5]);
  or _85950_ (_36631_, _36630_, _36623_);
  and _85951_ (_36633_, _36631_, _07141_);
  and _85952_ (_36634_, _07142_, \oc8051_golden_model_1.SBUF [5]);
  or _85953_ (_36635_, _36634_, _06341_);
  or _85954_ (_36636_, _36635_, _36633_);
  and _85955_ (_36637_, _36636_, _07166_);
  and _85956_ (_36638_, _36637_, _36629_);
  and _85957_ (_36639_, _36625_, _06461_);
  or _85958_ (_36640_, _36639_, _36638_);
  and _85959_ (_36641_, _36640_, _06465_);
  and _85960_ (_36642_, _36631_, _06464_);
  or _85961_ (_36644_, _36642_, _10080_);
  or _85962_ (_36645_, _36644_, _36641_);
  and _85963_ (_36646_, _36645_, _36626_);
  or _85964_ (_36647_, _36646_, _07460_);
  and _85965_ (_36648_, _09447_, _07886_);
  or _85966_ (_36649_, _36623_, _07208_);
  or _85967_ (_36650_, _36649_, _36648_);
  and _85968_ (_36651_, _36650_, _05982_);
  and _85969_ (_36652_, _36651_, _36647_);
  and _85970_ (_36653_, _15459_, _07886_);
  or _85971_ (_36655_, _36653_, _36623_);
  and _85972_ (_36656_, _36655_, _10094_);
  or _85973_ (_36657_, _36656_, _06218_);
  or _85974_ (_36658_, _36657_, _36652_);
  and _85975_ (_36659_, _08946_, _07886_);
  or _85976_ (_36660_, _36659_, _36623_);
  or _85977_ (_36661_, _36660_, _06219_);
  and _85978_ (_36662_, _36661_, _36658_);
  or _85979_ (_36663_, _36662_, _06369_);
  and _85980_ (_36664_, _15353_, _07886_);
  or _85981_ (_36666_, _36664_, _36623_);
  or _85982_ (_36667_, _36666_, _07237_);
  and _85983_ (_36668_, _36667_, _07240_);
  and _85984_ (_36669_, _36668_, _36663_);
  and _85985_ (_36670_, _11250_, _07886_);
  or _85986_ (_36671_, _36670_, _36623_);
  and _85987_ (_36672_, _36671_, _06536_);
  or _85988_ (_36673_, _36672_, _36669_);
  and _85989_ (_36674_, _36673_, _07242_);
  or _85990_ (_36675_, _36623_, _08247_);
  and _85991_ (_36677_, _36660_, _06375_);
  and _85992_ (_36678_, _36677_, _36675_);
  or _85993_ (_36679_, _36678_, _36674_);
  and _85994_ (_36680_, _36679_, _07234_);
  and _85995_ (_36681_, _36631_, _06545_);
  and _85996_ (_36682_, _36681_, _36675_);
  or _85997_ (_36683_, _36682_, _06366_);
  or _85998_ (_36684_, _36683_, _36680_);
  and _85999_ (_36685_, _15350_, _07886_);
  or _86000_ (_36686_, _36623_, _09056_);
  or _86001_ (_36688_, _36686_, _36685_);
  and _86002_ (_36689_, _36688_, _09061_);
  and _86003_ (_36690_, _36689_, _36684_);
  nor _86004_ (_36691_, _11249_, _13951_);
  or _86005_ (_36692_, _36691_, _36623_);
  and _86006_ (_36693_, _36692_, _06528_);
  or _86007_ (_36694_, _36693_, _36690_);
  and _86008_ (_36695_, _36694_, _06926_);
  and _86009_ (_36696_, _36628_, _06568_);
  or _86010_ (_36697_, _36696_, _06278_);
  or _86011_ (_36699_, _36697_, _36695_);
  and _86012_ (_36700_, _15532_, _07886_);
  or _86013_ (_36701_, _36623_, _06279_);
  or _86014_ (_36702_, _36701_, _36700_);
  and _86015_ (_36703_, _36702_, _01347_);
  and _86016_ (_36704_, _36703_, _36699_);
  or _86017_ (_36705_, _36704_, _36622_);
  and _86018_ (_43335_, _36705_, _42618_);
  and _86019_ (_36706_, _01351_, \oc8051_golden_model_1.SBUF [6]);
  and _86020_ (_36707_, _13951_, \oc8051_golden_model_1.SBUF [6]);
  and _86021_ (_36709_, _15554_, _07886_);
  or _86022_ (_36710_, _36709_, _36707_);
  or _86023_ (_36711_, _36710_, _07151_);
  and _86024_ (_36712_, _07886_, \oc8051_golden_model_1.ACC [6]);
  or _86025_ (_36713_, _36712_, _36707_);
  and _86026_ (_36714_, _36713_, _07141_);
  and _86027_ (_36715_, _07142_, \oc8051_golden_model_1.SBUF [6]);
  or _86028_ (_36716_, _36715_, _06341_);
  or _86029_ (_36717_, _36716_, _36714_);
  and _86030_ (_36718_, _36717_, _07166_);
  and _86031_ (_36720_, _36718_, _36711_);
  nor _86032_ (_36721_, _08142_, _13951_);
  or _86033_ (_36722_, _36721_, _36707_);
  and _86034_ (_36723_, _36722_, _06461_);
  or _86035_ (_36724_, _36723_, _36720_);
  and _86036_ (_36725_, _36724_, _06465_);
  and _86037_ (_36726_, _36713_, _06464_);
  or _86038_ (_36727_, _36726_, _10080_);
  or _86039_ (_36728_, _36727_, _36725_);
  or _86040_ (_36729_, _36722_, _07215_);
  and _86041_ (_36731_, _36729_, _36728_);
  or _86042_ (_36732_, _36731_, _07460_);
  and _86043_ (_36733_, _09446_, _07886_);
  or _86044_ (_36734_, _36707_, _07208_);
  or _86045_ (_36735_, _36734_, _36733_);
  and _86046_ (_36736_, _36735_, _05982_);
  and _86047_ (_36737_, _36736_, _36732_);
  and _86048_ (_36738_, _15657_, _07886_);
  or _86049_ (_36739_, _36738_, _36707_);
  and _86050_ (_36740_, _36739_, _10094_);
  or _86051_ (_36742_, _36740_, _06218_);
  or _86052_ (_36743_, _36742_, _36737_);
  and _86053_ (_36744_, _15664_, _07886_);
  or _86054_ (_36745_, _36744_, _36707_);
  or _86055_ (_36746_, _36745_, _06219_);
  and _86056_ (_36747_, _36746_, _36743_);
  or _86057_ (_36748_, _36747_, _06369_);
  and _86058_ (_36749_, _15549_, _07886_);
  or _86059_ (_36750_, _36749_, _36707_);
  or _86060_ (_36751_, _36750_, _07237_);
  and _86061_ (_36753_, _36751_, _07240_);
  and _86062_ (_36754_, _36753_, _36748_);
  and _86063_ (_36755_, _11247_, _07886_);
  or _86064_ (_36756_, _36755_, _36707_);
  and _86065_ (_36757_, _36756_, _06536_);
  or _86066_ (_36758_, _36757_, _36754_);
  and _86067_ (_36759_, _36758_, _07242_);
  or _86068_ (_36760_, _36707_, _08145_);
  and _86069_ (_36761_, _36745_, _06375_);
  and _86070_ (_36762_, _36761_, _36760_);
  or _86071_ (_36764_, _36762_, _36759_);
  and _86072_ (_36765_, _36764_, _07234_);
  and _86073_ (_36766_, _36713_, _06545_);
  and _86074_ (_36767_, _36766_, _36760_);
  or _86075_ (_36768_, _36767_, _06366_);
  or _86076_ (_36769_, _36768_, _36765_);
  and _86077_ (_36770_, _15546_, _07886_);
  or _86078_ (_36771_, _36707_, _09056_);
  or _86079_ (_36772_, _36771_, _36770_);
  and _86080_ (_36773_, _36772_, _09061_);
  and _86081_ (_36775_, _36773_, _36769_);
  nor _86082_ (_36776_, _11246_, _13951_);
  or _86083_ (_36777_, _36776_, _36707_);
  and _86084_ (_36778_, _36777_, _06528_);
  or _86085_ (_36779_, _36778_, _36775_);
  and _86086_ (_36780_, _36779_, _06926_);
  and _86087_ (_36781_, _36710_, _06568_);
  or _86088_ (_36782_, _36781_, _06278_);
  or _86089_ (_36783_, _36782_, _36780_);
  and _86090_ (_36784_, _15734_, _07886_);
  or _86091_ (_36786_, _36707_, _06279_);
  or _86092_ (_36787_, _36786_, _36784_);
  and _86093_ (_36788_, _36787_, _01347_);
  and _86094_ (_36789_, _36788_, _36783_);
  or _86095_ (_36790_, _36789_, _36706_);
  and _86096_ (_43336_, _36790_, _42618_);
  not _86097_ (_36791_, \oc8051_golden_model_1.PSW [0]);
  nor _86098_ (_36792_, _01347_, _36791_);
  nand _86099_ (_36793_, _11263_, _07935_);
  nor _86100_ (_36794_, _07935_, _36791_);
  nor _86101_ (_36796_, _36794_, _07234_);
  nand _86102_ (_36797_, _36796_, _36793_);
  and _86103_ (_36798_, _07935_, _07133_);
  or _86104_ (_36799_, _36798_, _36794_);
  or _86105_ (_36800_, _36799_, _07215_);
  nor _86106_ (_36801_, _08390_, _14045_);
  or _86107_ (_36802_, _36801_, _36794_);
  or _86108_ (_36803_, _36802_, _07151_);
  and _86109_ (_36804_, _07935_, \oc8051_golden_model_1.ACC [0]);
  or _86110_ (_36805_, _36804_, _36794_);
  and _86111_ (_36807_, _36805_, _07141_);
  nor _86112_ (_36808_, _07141_, _36791_);
  or _86113_ (_36809_, _36808_, _06341_);
  or _86114_ (_36810_, _36809_, _36807_);
  and _86115_ (_36811_, _36810_, _06273_);
  and _86116_ (_36812_, _36811_, _36803_);
  nor _86117_ (_36813_, _08630_, _36791_);
  and _86118_ (_36814_, _14382_, _08630_);
  or _86119_ (_36815_, _36814_, _36813_);
  and _86120_ (_36816_, _36815_, _06272_);
  or _86121_ (_36818_, _36816_, _36812_);
  and _86122_ (_36819_, _36818_, _07166_);
  and _86123_ (_36820_, _36799_, _06461_);
  or _86124_ (_36821_, _36820_, _06464_);
  or _86125_ (_36822_, _36821_, _36819_);
  or _86126_ (_36823_, _36805_, _06465_);
  and _86127_ (_36824_, _36823_, _06269_);
  and _86128_ (_36825_, _36824_, _36822_);
  and _86129_ (_36826_, _36794_, _06268_);
  or _86130_ (_36827_, _36826_, _06261_);
  or _86131_ (_36829_, _36827_, _36825_);
  or _86132_ (_36830_, _36802_, _06262_);
  and _86133_ (_36831_, _36830_, _06258_);
  and _86134_ (_36832_, _36831_, _36829_);
  and _86135_ (_36833_, _14413_, _08630_);
  or _86136_ (_36834_, _36833_, _36813_);
  and _86137_ (_36835_, _36834_, _06257_);
  or _86138_ (_36836_, _36835_, _10080_);
  or _86139_ (_36837_, _36836_, _36832_);
  and _86140_ (_36838_, _36837_, _36800_);
  or _86141_ (_36840_, _36838_, _07460_);
  and _86142_ (_36841_, _09392_, _07935_);
  or _86143_ (_36842_, _36794_, _07208_);
  or _86144_ (_36843_, _36842_, _36841_);
  and _86145_ (_36844_, _36843_, _36840_);
  or _86146_ (_36845_, _36844_, _10094_);
  and _86147_ (_36846_, _14467_, _07935_);
  or _86148_ (_36847_, _36794_, _05982_);
  or _86149_ (_36848_, _36847_, _36846_);
  and _86150_ (_36849_, _36848_, _06219_);
  and _86151_ (_36851_, _36849_, _36845_);
  and _86152_ (_36852_, _07935_, _08954_);
  or _86153_ (_36853_, _36852_, _36794_);
  and _86154_ (_36854_, _36853_, _06218_);
  or _86155_ (_36855_, _36854_, _06369_);
  or _86156_ (_36856_, _36855_, _36851_);
  and _86157_ (_36857_, _14366_, _07935_);
  or _86158_ (_36858_, _36857_, _36794_);
  or _86159_ (_36859_, _36858_, _07237_);
  and _86160_ (_36860_, _36859_, _07240_);
  and _86161_ (_36862_, _36860_, _36856_);
  nor _86162_ (_36863_, _12580_, _14045_);
  or _86163_ (_36864_, _36863_, _36794_);
  and _86164_ (_36865_, _36793_, _06536_);
  and _86165_ (_36866_, _36865_, _36864_);
  or _86166_ (_36867_, _36866_, _36862_);
  and _86167_ (_36868_, _36867_, _07242_);
  nand _86168_ (_36869_, _36853_, _06375_);
  nor _86169_ (_36870_, _36869_, _36801_);
  or _86170_ (_36871_, _36870_, _06545_);
  or _86171_ (_36872_, _36871_, _36868_);
  and _86172_ (_36873_, _36872_, _36797_);
  or _86173_ (_36874_, _36873_, _06366_);
  and _86174_ (_36875_, _14363_, _07935_);
  or _86175_ (_36876_, _36794_, _09056_);
  or _86176_ (_36877_, _36876_, _36875_);
  and _86177_ (_36878_, _36877_, _09061_);
  and _86178_ (_36879_, _36878_, _36874_);
  and _86179_ (_36880_, _36864_, _06528_);
  or _86180_ (_36881_, _36880_, _06568_);
  or _86181_ (_36883_, _36881_, _36879_);
  or _86182_ (_36884_, _36802_, _06926_);
  and _86183_ (_36885_, _36884_, _36883_);
  or _86184_ (_36886_, _36885_, _05927_);
  or _86185_ (_36887_, _36794_, _05928_);
  and _86186_ (_36888_, _36887_, _36886_);
  or _86187_ (_36889_, _36888_, _06278_);
  or _86188_ (_36890_, _36802_, _06279_);
  and _86189_ (_36891_, _36890_, _01347_);
  and _86190_ (_36892_, _36891_, _36889_);
  or _86191_ (_36894_, _36892_, _36792_);
  and _86192_ (_43338_, _36894_, _42618_);
  not _86193_ (_36895_, \oc8051_golden_model_1.PSW [1]);
  nor _86194_ (_36896_, _01347_, _36895_);
  nor _86195_ (_36897_, _07935_, _36895_);
  nor _86196_ (_36898_, _11261_, _14045_);
  or _86197_ (_36899_, _36898_, _36897_);
  or _86198_ (_36900_, _36899_, _09061_);
  nor _86199_ (_36901_, _14045_, _07357_);
  or _86200_ (_36902_, _36901_, _36897_);
  or _86201_ (_36904_, _36902_, _07215_);
  and _86202_ (_36905_, _36902_, _06461_);
  nor _86203_ (_36906_, _08630_, _36895_);
  and _86204_ (_36907_, _14557_, _08630_);
  or _86205_ (_36908_, _36907_, _36906_);
  or _86206_ (_36909_, _36908_, _06273_);
  or _86207_ (_36910_, _07935_, \oc8051_golden_model_1.PSW [1]);
  and _86208_ (_36911_, _14562_, _07935_);
  not _86209_ (_36912_, _36911_);
  and _86210_ (_36913_, _36912_, _36910_);
  and _86211_ (_36915_, _36913_, _06341_);
  nor _86212_ (_36916_, _07141_, _36895_);
  and _86213_ (_36917_, _07935_, \oc8051_golden_model_1.ACC [1]);
  or _86214_ (_36918_, _36917_, _36897_);
  and _86215_ (_36919_, _36918_, _07141_);
  or _86216_ (_36920_, _36919_, _36916_);
  and _86217_ (_36921_, _36920_, _07151_);
  or _86218_ (_36922_, _36921_, _06272_);
  or _86219_ (_36923_, _36922_, _36915_);
  and _86220_ (_36924_, _36923_, _36909_);
  and _86221_ (_36926_, _36924_, _07166_);
  or _86222_ (_36927_, _36926_, _36905_);
  or _86223_ (_36928_, _36927_, _06464_);
  or _86224_ (_36929_, _36918_, _06465_);
  and _86225_ (_36930_, _36929_, _06269_);
  and _86226_ (_36931_, _36930_, _36928_);
  and _86227_ (_36932_, _14560_, _08630_);
  or _86228_ (_36933_, _36932_, _36906_);
  and _86229_ (_36934_, _36933_, _06268_);
  or _86230_ (_36935_, _36934_, _06261_);
  or _86231_ (_36937_, _36935_, _36931_);
  or _86232_ (_36938_, _36906_, _14556_);
  and _86233_ (_36939_, _36938_, _36908_);
  or _86234_ (_36940_, _36939_, _06262_);
  and _86235_ (_36941_, _36940_, _06258_);
  and _86236_ (_36942_, _36941_, _36937_);
  or _86237_ (_36943_, _36906_, _14597_);
  and _86238_ (_36944_, _36943_, _06257_);
  and _86239_ (_36945_, _36944_, _36908_);
  or _86240_ (_36946_, _36945_, _10080_);
  or _86241_ (_36948_, _36946_, _36942_);
  and _86242_ (_36949_, _36948_, _36904_);
  or _86243_ (_36950_, _36949_, _07460_);
  and _86244_ (_36951_, _09451_, _07935_);
  or _86245_ (_36952_, _36897_, _07208_);
  or _86246_ (_36953_, _36952_, _36951_);
  and _86247_ (_36954_, _36953_, _05982_);
  and _86248_ (_36955_, _36954_, _36950_);
  or _86249_ (_36956_, _14653_, _14045_);
  and _86250_ (_36957_, _36910_, _10094_);
  and _86251_ (_36959_, _36957_, _36956_);
  or _86252_ (_36960_, _36959_, _36955_);
  and _86253_ (_36961_, _36960_, _06219_);
  nand _86254_ (_36962_, _07935_, _07038_);
  and _86255_ (_36963_, _36910_, _06218_);
  and _86256_ (_36964_, _36963_, _36962_);
  or _86257_ (_36965_, _36964_, _36961_);
  and _86258_ (_36966_, _36965_, _07237_);
  or _86259_ (_36967_, _14668_, _14045_);
  and _86260_ (_36968_, _36910_, _06369_);
  and _86261_ (_36970_, _36968_, _36967_);
  or _86262_ (_36971_, _36970_, _06536_);
  or _86263_ (_36972_, _36971_, _36966_);
  nand _86264_ (_36973_, _11260_, _07935_);
  and _86265_ (_36974_, _36973_, _36899_);
  or _86266_ (_36975_, _36974_, _07240_);
  and _86267_ (_36976_, _36975_, _07242_);
  and _86268_ (_36977_, _36976_, _36972_);
  or _86269_ (_36978_, _14666_, _14045_);
  and _86270_ (_36979_, _36910_, _06375_);
  and _86271_ (_36981_, _36979_, _36978_);
  or _86272_ (_36982_, _36981_, _06545_);
  or _86273_ (_36983_, _36982_, _36977_);
  nor _86274_ (_36984_, _36897_, _07234_);
  nand _86275_ (_36985_, _36984_, _36973_);
  and _86276_ (_36986_, _36985_, _09056_);
  and _86277_ (_36987_, _36986_, _36983_);
  or _86278_ (_36988_, _36962_, _08341_);
  and _86279_ (_36989_, _36910_, _06366_);
  and _86280_ (_36990_, _36989_, _36988_);
  or _86281_ (_36992_, _36990_, _06528_);
  or _86282_ (_36993_, _36992_, _36987_);
  and _86283_ (_36994_, _36993_, _36900_);
  or _86284_ (_36995_, _36994_, _06568_);
  or _86285_ (_36996_, _36913_, _06926_);
  and _86286_ (_36997_, _36996_, _05928_);
  and _86287_ (_36998_, _36997_, _36995_);
  and _86288_ (_36999_, _36933_, _05927_);
  or _86289_ (_37000_, _36999_, _06278_);
  or _86290_ (_37001_, _37000_, _36998_);
  or _86291_ (_37003_, _36897_, _06279_);
  or _86292_ (_37004_, _37003_, _36911_);
  and _86293_ (_37005_, _37004_, _01347_);
  and _86294_ (_37006_, _37005_, _37001_);
  or _86295_ (_37007_, _37006_, _36896_);
  and _86296_ (_43339_, _37007_, _42618_);
  and _86297_ (_37008_, _01351_, \oc8051_golden_model_1.PSW [2]);
  not _86298_ (_37009_, _10960_);
  and _86299_ (_37010_, _11319_, _37009_);
  or _86300_ (_37011_, _37010_, _14336_);
  nand _86301_ (_37013_, _37011_, _06926_);
  not _86302_ (_37014_, _10499_);
  nand _86303_ (_37015_, _11236_, _37014_);
  or _86304_ (_37016_, _11236_, _10498_);
  and _86305_ (_37017_, _37016_, _37015_);
  or _86306_ (_37018_, _37017_, _17800_);
  not _86307_ (_37019_, _11035_);
  nand _86308_ (_37020_, _11062_, \oc8051_golden_model_1.ACC [7]);
  nand _86309_ (_37021_, _37020_, _10666_);
  not _86310_ (_37022_, _10669_);
  and _86311_ (_37024_, _11062_, _37022_);
  nor _86312_ (_37025_, _37024_, _11064_);
  or _86313_ (_37026_, _37025_, _10666_);
  and _86314_ (_37027_, _37026_, _37021_);
  or _86315_ (_37028_, _37027_, _37019_);
  and _86316_ (_37029_, _14045_, \oc8051_golden_model_1.PSW [2]);
  nor _86317_ (_37030_, _14045_, _07776_);
  or _86318_ (_37031_, _37030_, _37029_);
  or _86319_ (_37032_, _37031_, _07215_);
  and _86320_ (_37033_, _14234_, _10522_);
  nor _86321_ (_37035_, _14234_, _10522_);
  or _86322_ (_37036_, _37035_, _37033_);
  or _86323_ (_37037_, _37036_, _10581_);
  nand _86324_ (_37038_, _37036_, _10581_);
  and _86325_ (_37039_, _37038_, _37037_);
  and _86326_ (_37040_, _37039_, _10516_);
  nor _86327_ (_37041_, _10596_, \oc8051_golden_model_1.ACC [7]);
  nor _86328_ (_37042_, _10595_, _37014_);
  nor _86329_ (_37043_, _37042_, _37041_);
  not _86330_ (_37044_, _37043_);
  or _86331_ (_37046_, _37044_, _14053_);
  nand _86332_ (_37047_, _37044_, _14053_);
  and _86333_ (_37048_, _37047_, _37046_);
  and _86334_ (_37049_, _37048_, _10654_);
  nor _86335_ (_37050_, _37048_, _10654_);
  or _86336_ (_37051_, _37050_, _37049_);
  or _86337_ (_37052_, _37051_, _10588_);
  and _86338_ (_37053_, _14209_, _10665_);
  nor _86339_ (_37054_, _14209_, _10665_);
  or _86340_ (_37055_, _37054_, _37053_);
  or _86341_ (_37057_, _37055_, _10724_);
  nand _86342_ (_37058_, _37055_, _10724_);
  and _86343_ (_37059_, _37058_, _10737_);
  and _86344_ (_37060_, _37059_, _37057_);
  or _86345_ (_37061_, _37031_, _07166_);
  and _86346_ (_37062_, _14770_, _07935_);
  or _86347_ (_37063_, _37062_, _37029_);
  or _86348_ (_37064_, _37063_, _07151_);
  and _86349_ (_37065_, _07935_, \oc8051_golden_model_1.ACC [2]);
  or _86350_ (_37066_, _37065_, _37029_);
  and _86351_ (_37068_, _37066_, _07141_);
  and _86352_ (_37069_, _07142_, \oc8051_golden_model_1.PSW [2]);
  or _86353_ (_37070_, _37069_, _06341_);
  or _86354_ (_37071_, _37070_, _37068_);
  and _86355_ (_37072_, _37071_, _06273_);
  and _86356_ (_37073_, _37072_, _37064_);
  not _86357_ (_37074_, _08630_);
  and _86358_ (_37075_, _37074_, \oc8051_golden_model_1.PSW [2]);
  and _86359_ (_37076_, _14774_, _08630_);
  or _86360_ (_37077_, _37076_, _37075_);
  and _86361_ (_37079_, _37077_, _06272_);
  or _86362_ (_37080_, _37079_, _06461_);
  or _86363_ (_37081_, _37080_, _37073_);
  and _86364_ (_37082_, _37081_, _37061_);
  or _86365_ (_37083_, _37082_, _06464_);
  or _86366_ (_37084_, _37066_, _06465_);
  and _86367_ (_37085_, _37084_, _06269_);
  and _86368_ (_37086_, _37085_, _37083_);
  and _86369_ (_37087_, _14756_, _08630_);
  or _86370_ (_37088_, _37087_, _37075_);
  and _86371_ (_37090_, _37088_, _06268_);
  or _86372_ (_37091_, _37090_, _06261_);
  or _86373_ (_37092_, _37091_, _37086_);
  and _86374_ (_37093_, _37076_, _14789_);
  or _86375_ (_37094_, _37075_, _06262_);
  or _86376_ (_37095_, _37094_, _37093_);
  and _86377_ (_37096_, _37095_, _37092_);
  or _86378_ (_37097_, _37096_, _09531_);
  or _86379_ (_37098_, _16582_, _16472_);
  or _86380_ (_37099_, _37098_, _16694_);
  or _86381_ (_37101_, _37099_, _16814_);
  or _86382_ (_37102_, _37101_, _16931_);
  or _86383_ (_37103_, _37102_, _17045_);
  or _86384_ (_37104_, _37103_, _17165_);
  or _86385_ (_37105_, _37104_, _10076_);
  and _86386_ (_37106_, _37105_, _10735_);
  and _86387_ (_37107_, _37106_, _37097_);
  or _86388_ (_37108_, _37107_, _10656_);
  or _86389_ (_37109_, _37108_, _37060_);
  and _86390_ (_37110_, _37109_, _06517_);
  and _86391_ (_37112_, _37110_, _37052_);
  nor _86392_ (_37113_, _10840_, _14329_);
  nor _86393_ (_37114_, _10841_, \oc8051_golden_model_1.ACC [7]);
  nor _86394_ (_37115_, _37114_, _37113_);
  not _86395_ (_37116_, _37115_);
  or _86396_ (_37117_, _37116_, _14223_);
  nand _86397_ (_37118_, _37116_, _14223_);
  and _86398_ (_37119_, _37118_, _37117_);
  and _86399_ (_37120_, _37119_, _10898_);
  nor _86400_ (_37121_, _37119_, _10898_);
  or _86401_ (_37123_, _37121_, _37120_);
  and _86402_ (_37124_, _37123_, _06512_);
  or _86403_ (_37125_, _37124_, _37112_);
  and _86404_ (_37126_, _37125_, _10517_);
  or _86405_ (_37127_, _37126_, _37040_);
  and _86406_ (_37128_, _37127_, _06258_);
  and _86407_ (_37129_, _14804_, _08630_);
  or _86408_ (_37130_, _37129_, _37075_);
  and _86409_ (_37131_, _37130_, _06257_);
  or _86410_ (_37132_, _37131_, _10080_);
  or _86411_ (_37134_, _37132_, _37128_);
  and _86412_ (_37135_, _37134_, _37032_);
  or _86413_ (_37136_, _37135_, _07460_);
  and _86414_ (_37137_, _09450_, _07935_);
  or _86415_ (_37138_, _37029_, _07208_);
  or _86416_ (_37139_, _37138_, _37137_);
  and _86417_ (_37140_, _37139_, _05982_);
  and _86418_ (_37141_, _37140_, _37136_);
  and _86419_ (_37142_, _14859_, _07935_);
  or _86420_ (_37143_, _37142_, _37029_);
  and _86421_ (_37145_, _37143_, _10094_);
  or _86422_ (_37146_, _37145_, _10093_);
  or _86423_ (_37147_, _37146_, _37141_);
  nand _86424_ (_37148_, _10113_, _10106_);
  nand _86425_ (_37149_, _37148_, _10093_);
  and _86426_ (_37150_, _37149_, _37147_);
  and _86427_ (_37151_, _37150_, _06219_);
  and _86428_ (_37152_, _07935_, _08973_);
  or _86429_ (_37153_, _37152_, _37029_);
  and _86430_ (_37154_, _37153_, _06218_);
  or _86431_ (_37156_, _37154_, _06369_);
  or _86432_ (_37157_, _37156_, _37151_);
  and _86433_ (_37158_, _14751_, _07935_);
  or _86434_ (_37159_, _37158_, _37029_);
  or _86435_ (_37160_, _37159_, _07237_);
  and _86436_ (_37161_, _37160_, _07240_);
  and _86437_ (_37162_, _37161_, _37157_);
  and _86438_ (_37163_, _11259_, _07935_);
  or _86439_ (_37164_, _37163_, _37029_);
  and _86440_ (_37165_, _37164_, _06536_);
  or _86441_ (_37167_, _37165_, _37162_);
  and _86442_ (_37168_, _37167_, _07242_);
  or _86443_ (_37169_, _37029_, _08440_);
  and _86444_ (_37170_, _37153_, _06375_);
  and _86445_ (_37171_, _37170_, _37169_);
  or _86446_ (_37172_, _37171_, _37168_);
  and _86447_ (_37173_, _37172_, _07234_);
  and _86448_ (_37174_, _37066_, _06545_);
  and _86449_ (_37175_, _37174_, _37169_);
  or _86450_ (_37176_, _37175_, _06366_);
  or _86451_ (_37178_, _37176_, _37173_);
  and _86452_ (_37179_, _14748_, _07935_);
  or _86453_ (_37180_, _37179_, _37029_);
  or _86454_ (_37181_, _37180_, _09056_);
  and _86455_ (_37182_, _37181_, _09061_);
  and _86456_ (_37183_, _37182_, _37178_);
  nor _86457_ (_37184_, _11258_, _14045_);
  or _86458_ (_37185_, _37184_, _37029_);
  and _86459_ (_37186_, _37185_, _06528_);
  or _86460_ (_37187_, _37186_, _11035_);
  or _86461_ (_37189_, _37187_, _37183_);
  and _86462_ (_37190_, _37189_, _37028_);
  or _86463_ (_37191_, _37190_, _11036_);
  not _86464_ (_37192_, _11036_);
  or _86465_ (_37193_, _37027_, _37192_);
  and _86466_ (_37194_, _37193_, _11069_);
  and _86467_ (_37195_, _37194_, _37191_);
  nor _86468_ (_37196_, _37044_, _14293_);
  nor _86469_ (_37197_, _37196_, _37042_);
  and _86470_ (_37198_, _37197_, _11093_);
  and _86471_ (_37200_, _37042_, _11090_);
  or _86472_ (_37201_, _37200_, _37198_);
  and _86473_ (_37202_, _37201_, _11041_);
  or _86474_ (_37203_, _37202_, _14297_);
  or _86475_ (_37204_, _37203_, _37195_);
  nor _86476_ (_37205_, _37116_, _14299_);
  nor _86477_ (_37206_, _37205_, _37113_);
  and _86478_ (_37207_, _37206_, _11121_);
  and _86479_ (_37208_, _37113_, _11118_);
  or _86480_ (_37209_, _37208_, _37207_);
  or _86481_ (_37211_, _37209_, _06541_);
  nor _86482_ (_37212_, _10521_, _37009_);
  nor _86483_ (_37213_, _10523_, \oc8051_golden_model_1.ACC [7]);
  nor _86484_ (_37214_, _37213_, _14305_);
  nor _86485_ (_37215_, _37214_, _37212_);
  and _86486_ (_37216_, _37215_, _11149_);
  and _86487_ (_37217_, _37212_, _11146_);
  or _86488_ (_37218_, _37217_, _37216_);
  or _86489_ (_37219_, _37218_, _11127_);
  and _86490_ (_37220_, _37219_, _11157_);
  and _86491_ (_37222_, _37220_, _37211_);
  and _86492_ (_37223_, _37222_, _37204_);
  or _86493_ (_37224_, _11193_, _10494_);
  nor _86494_ (_37225_, _14315_, _11192_);
  nor _86495_ (_37226_, _37225_, _11157_);
  and _86496_ (_37227_, _37226_, _37224_);
  or _86497_ (_37228_, _37227_, _11200_);
  or _86498_ (_37229_, _37228_, _37223_);
  and _86499_ (_37230_, _37229_, _37018_);
  or _86500_ (_37231_, _37230_, _11199_);
  or _86501_ (_37233_, _37017_, _18067_);
  and _86502_ (_37234_, _37233_, _13012_);
  and _86503_ (_37235_, _37234_, _37231_);
  or _86504_ (_37236_, _11277_, _08573_);
  and _86505_ (_37237_, _37236_, _14331_);
  or _86506_ (_37238_, _37237_, _37235_);
  or _86507_ (_37239_, _37238_, _37013_);
  or _86508_ (_37240_, _37063_, _06926_);
  and _86509_ (_37241_, _37240_, _05928_);
  and _86510_ (_37242_, _37241_, _37239_);
  and _86511_ (_37244_, _37088_, _05927_);
  or _86512_ (_37245_, _37244_, _06278_);
  or _86513_ (_37246_, _37245_, _37242_);
  and _86514_ (_37247_, _14926_, _07935_);
  or _86515_ (_37248_, _37029_, _06279_);
  or _86516_ (_37249_, _37248_, _37247_);
  and _86517_ (_37250_, _37249_, _01347_);
  and _86518_ (_37251_, _37250_, _37246_);
  or _86519_ (_37252_, _37251_, _37008_);
  and _86520_ (_43340_, _37252_, _42618_);
  nor _86521_ (_37254_, _01347_, _07615_);
  nor _86522_ (_37255_, _07935_, _07615_);
  nor _86523_ (_37256_, _14045_, _07594_);
  or _86524_ (_37257_, _37256_, _37255_);
  or _86525_ (_37258_, _37257_, _07215_);
  and _86526_ (_37259_, _14953_, _07935_);
  or _86527_ (_37260_, _37259_, _37255_);
  or _86528_ (_37261_, _37260_, _07151_);
  and _86529_ (_37262_, _07935_, \oc8051_golden_model_1.ACC [3]);
  or _86530_ (_37263_, _37262_, _37255_);
  and _86531_ (_37265_, _37263_, _07141_);
  nor _86532_ (_37266_, _07141_, _07615_);
  or _86533_ (_37267_, _37266_, _06341_);
  or _86534_ (_37268_, _37267_, _37265_);
  and _86535_ (_37269_, _37268_, _06273_);
  and _86536_ (_37270_, _37269_, _37261_);
  nor _86537_ (_37271_, _08630_, _07615_);
  and _86538_ (_37272_, _14950_, _08630_);
  or _86539_ (_37273_, _37272_, _37271_);
  and _86540_ (_37274_, _37273_, _06272_);
  or _86541_ (_37276_, _37274_, _06461_);
  or _86542_ (_37277_, _37276_, _37270_);
  or _86543_ (_37278_, _37257_, _07166_);
  and _86544_ (_37279_, _37278_, _37277_);
  or _86545_ (_37280_, _37279_, _06464_);
  or _86546_ (_37281_, _37263_, _06465_);
  and _86547_ (_37282_, _37281_, _06269_);
  and _86548_ (_37283_, _37282_, _37280_);
  and _86549_ (_37284_, _14948_, _08630_);
  or _86550_ (_37285_, _37284_, _37271_);
  and _86551_ (_37287_, _37285_, _06268_);
  or _86552_ (_37288_, _37287_, _06261_);
  or _86553_ (_37289_, _37288_, _37283_);
  or _86554_ (_37290_, _37271_, _14979_);
  and _86555_ (_37291_, _37290_, _37273_);
  or _86556_ (_37292_, _37291_, _06262_);
  and _86557_ (_37293_, _37292_, _06258_);
  and _86558_ (_37294_, _37293_, _37289_);
  or _86559_ (_37295_, _37271_, _14992_);
  and _86560_ (_37296_, _37295_, _06257_);
  and _86561_ (_37298_, _37296_, _37273_);
  or _86562_ (_37299_, _37298_, _10080_);
  or _86563_ (_37300_, _37299_, _37294_);
  and _86564_ (_37301_, _37300_, _37258_);
  or _86565_ (_37302_, _37301_, _07460_);
  and _86566_ (_37303_, _09449_, _07935_);
  or _86567_ (_37304_, _37255_, _07208_);
  or _86568_ (_37305_, _37304_, _37303_);
  and _86569_ (_37306_, _37305_, _05982_);
  and _86570_ (_37307_, _37306_, _37302_);
  and _86571_ (_37309_, _15048_, _07935_);
  or _86572_ (_37310_, _37309_, _37255_);
  and _86573_ (_37311_, _37310_, _10094_);
  or _86574_ (_37312_, _37311_, _06218_);
  or _86575_ (_37313_, _37312_, _37307_);
  and _86576_ (_37314_, _07935_, _08930_);
  or _86577_ (_37315_, _37314_, _37255_);
  or _86578_ (_37316_, _37315_, _06219_);
  and _86579_ (_37317_, _37316_, _37313_);
  or _86580_ (_37318_, _37317_, _06369_);
  and _86581_ (_37320_, _14943_, _07935_);
  or _86582_ (_37321_, _37320_, _37255_);
  or _86583_ (_37322_, _37321_, _07237_);
  and _86584_ (_37323_, _37322_, _07240_);
  and _86585_ (_37324_, _37323_, _37318_);
  and _86586_ (_37325_, _12577_, _07935_);
  or _86587_ (_37326_, _37325_, _37255_);
  and _86588_ (_37327_, _37326_, _06536_);
  or _86589_ (_37328_, _37327_, _37324_);
  and _86590_ (_37329_, _37328_, _07242_);
  or _86591_ (_37331_, _37255_, _08292_);
  and _86592_ (_37332_, _37315_, _06375_);
  and _86593_ (_37333_, _37332_, _37331_);
  or _86594_ (_37334_, _37333_, _37329_);
  and _86595_ (_37335_, _37334_, _07234_);
  and _86596_ (_37336_, _37263_, _06545_);
  and _86597_ (_37337_, _37336_, _37331_);
  or _86598_ (_37338_, _37337_, _06366_);
  or _86599_ (_37339_, _37338_, _37335_);
  and _86600_ (_37340_, _14940_, _07935_);
  or _86601_ (_37342_, _37255_, _09056_);
  or _86602_ (_37343_, _37342_, _37340_);
  and _86603_ (_37344_, _37343_, _09061_);
  and _86604_ (_37345_, _37344_, _37339_);
  nor _86605_ (_37346_, _11256_, _14045_);
  or _86606_ (_37347_, _37346_, _37255_);
  and _86607_ (_37348_, _37347_, _06528_);
  or _86608_ (_37349_, _37348_, _06568_);
  or _86609_ (_37350_, _37349_, _37345_);
  or _86610_ (_37351_, _37260_, _06926_);
  and _86611_ (_37353_, _37351_, _05928_);
  and _86612_ (_37354_, _37353_, _37350_);
  and _86613_ (_37355_, _37285_, _05927_);
  or _86614_ (_37356_, _37355_, _06278_);
  or _86615_ (_37357_, _37356_, _37354_);
  and _86616_ (_37358_, _15128_, _07935_);
  or _86617_ (_37359_, _37255_, _06279_);
  or _86618_ (_37360_, _37359_, _37358_);
  and _86619_ (_37361_, _37360_, _01347_);
  and _86620_ (_37362_, _37361_, _37357_);
  or _86621_ (_37364_, _37362_, _37254_);
  and _86622_ (_43341_, _37364_, _42618_);
  and _86623_ (_37365_, _01351_, \oc8051_golden_model_1.PSW [4]);
  and _86624_ (_37366_, _14045_, \oc8051_golden_model_1.PSW [4]);
  nor _86625_ (_37367_, _08541_, _14045_);
  or _86626_ (_37368_, _37367_, _37366_);
  or _86627_ (_37369_, _37368_, _07215_);
  and _86628_ (_37370_, _37074_, \oc8051_golden_model_1.PSW [4]);
  and _86629_ (_37371_, _15176_, _08630_);
  or _86630_ (_37372_, _37371_, _37370_);
  and _86631_ (_37374_, _37372_, _06268_);
  and _86632_ (_37375_, _15162_, _07935_);
  or _86633_ (_37376_, _37375_, _37366_);
  or _86634_ (_37377_, _37376_, _07151_);
  and _86635_ (_37378_, _07935_, \oc8051_golden_model_1.ACC [4]);
  or _86636_ (_37379_, _37378_, _37366_);
  and _86637_ (_37380_, _37379_, _07141_);
  and _86638_ (_37381_, _07142_, \oc8051_golden_model_1.PSW [4]);
  or _86639_ (_37382_, _37381_, _06341_);
  or _86640_ (_37383_, _37382_, _37380_);
  and _86641_ (_37385_, _37383_, _06273_);
  and _86642_ (_37386_, _37385_, _37377_);
  and _86643_ (_37387_, _15166_, _08630_);
  or _86644_ (_37388_, _37387_, _37370_);
  and _86645_ (_37389_, _37388_, _06272_);
  or _86646_ (_37390_, _37389_, _06461_);
  or _86647_ (_37391_, _37390_, _37386_);
  or _86648_ (_37392_, _37368_, _07166_);
  and _86649_ (_37393_, _37392_, _37391_);
  or _86650_ (_37394_, _37393_, _06464_);
  or _86651_ (_37396_, _37379_, _06465_);
  and _86652_ (_37397_, _37396_, _06269_);
  and _86653_ (_37398_, _37397_, _37394_);
  or _86654_ (_37399_, _37398_, _37374_);
  and _86655_ (_37400_, _37399_, _06262_);
  or _86656_ (_37401_, _37370_, _15183_);
  and _86657_ (_37402_, _37401_, _06261_);
  and _86658_ (_37403_, _37402_, _37388_);
  or _86659_ (_37404_, _37403_, _37400_);
  and _86660_ (_37405_, _37404_, _06258_);
  and _86661_ (_37407_, _15200_, _08630_);
  or _86662_ (_37408_, _37407_, _37370_);
  and _86663_ (_37409_, _37408_, _06257_);
  or _86664_ (_37410_, _37409_, _10080_);
  or _86665_ (_37411_, _37410_, _37405_);
  and _86666_ (_37412_, _37411_, _37369_);
  or _86667_ (_37413_, _37412_, _07460_);
  and _86668_ (_37414_, _09448_, _07935_);
  or _86669_ (_37415_, _37366_, _07208_);
  or _86670_ (_37416_, _37415_, _37414_);
  and _86671_ (_37418_, _37416_, _05982_);
  and _86672_ (_37419_, _37418_, _37413_);
  and _86673_ (_37420_, _15254_, _07935_);
  or _86674_ (_37421_, _37420_, _37366_);
  and _86675_ (_37422_, _37421_, _10094_);
  or _86676_ (_37423_, _37422_, _06218_);
  or _86677_ (_37424_, _37423_, _37419_);
  and _86678_ (_37425_, _08959_, _07935_);
  or _86679_ (_37426_, _37425_, _37366_);
  or _86680_ (_37427_, _37426_, _06219_);
  and _86681_ (_37429_, _37427_, _37424_);
  or _86682_ (_37430_, _37429_, _06369_);
  and _86683_ (_37431_, _15269_, _07935_);
  or _86684_ (_37432_, _37431_, _37366_);
  or _86685_ (_37433_, _37432_, _07237_);
  and _86686_ (_37434_, _37433_, _07240_);
  and _86687_ (_37435_, _37434_, _37430_);
  and _86688_ (_37436_, _11254_, _07935_);
  or _86689_ (_37437_, _37436_, _37366_);
  and _86690_ (_37438_, _37437_, _06536_);
  or _86691_ (_37440_, _37438_, _37435_);
  and _86692_ (_37441_, _37440_, _07242_);
  or _86693_ (_37442_, _37366_, _08544_);
  and _86694_ (_37443_, _37426_, _06375_);
  and _86695_ (_37444_, _37443_, _37442_);
  or _86696_ (_37445_, _37444_, _37441_);
  and _86697_ (_37446_, _37445_, _07234_);
  and _86698_ (_37447_, _37379_, _06545_);
  and _86699_ (_37448_, _37447_, _37442_);
  or _86700_ (_37449_, _37448_, _06366_);
  or _86701_ (_37451_, _37449_, _37446_);
  and _86702_ (_37452_, _15266_, _07935_);
  or _86703_ (_37453_, _37366_, _09056_);
  or _86704_ (_37454_, _37453_, _37452_);
  and _86705_ (_37455_, _37454_, _09061_);
  and _86706_ (_37456_, _37455_, _37451_);
  nor _86707_ (_37457_, _11253_, _14045_);
  or _86708_ (_37458_, _37457_, _37366_);
  and _86709_ (_37459_, _37458_, _06528_);
  or _86710_ (_37460_, _37459_, _06568_);
  or _86711_ (_37462_, _37460_, _37456_);
  or _86712_ (_37463_, _37376_, _06926_);
  and _86713_ (_37464_, _37463_, _05928_);
  and _86714_ (_37465_, _37464_, _37462_);
  and _86715_ (_37466_, _37372_, _05927_);
  or _86716_ (_37467_, _37466_, _06278_);
  or _86717_ (_37468_, _37467_, _37465_);
  and _86718_ (_37469_, _15329_, _07935_);
  or _86719_ (_37470_, _37366_, _06279_);
  or _86720_ (_37471_, _37470_, _37469_);
  and _86721_ (_37473_, _37471_, _01347_);
  and _86722_ (_37474_, _37473_, _37468_);
  or _86723_ (_37475_, _37474_, _37365_);
  and _86724_ (_43342_, _37475_, _42618_);
  and _86725_ (_37476_, _01351_, \oc8051_golden_model_1.PSW [5]);
  and _86726_ (_37477_, _14045_, \oc8051_golden_model_1.PSW [5]);
  and _86727_ (_37478_, _15358_, _07935_);
  or _86728_ (_37479_, _37478_, _37477_);
  or _86729_ (_37480_, _37479_, _07151_);
  and _86730_ (_37481_, _07935_, \oc8051_golden_model_1.ACC [5]);
  or _86731_ (_37483_, _37481_, _37477_);
  and _86732_ (_37484_, _37483_, _07141_);
  and _86733_ (_37485_, _07142_, \oc8051_golden_model_1.PSW [5]);
  or _86734_ (_37486_, _37485_, _06341_);
  or _86735_ (_37487_, _37486_, _37484_);
  and _86736_ (_37488_, _37487_, _06273_);
  and _86737_ (_37489_, _37488_, _37480_);
  and _86738_ (_37490_, _37074_, \oc8051_golden_model_1.PSW [5]);
  and _86739_ (_37491_, _15372_, _08630_);
  or _86740_ (_37492_, _37491_, _37490_);
  and _86741_ (_37494_, _37492_, _06272_);
  or _86742_ (_37495_, _37494_, _06461_);
  or _86743_ (_37496_, _37495_, _37489_);
  nor _86744_ (_37497_, _08244_, _14045_);
  or _86745_ (_37498_, _37497_, _37477_);
  or _86746_ (_37499_, _37498_, _07166_);
  and _86747_ (_37500_, _37499_, _37496_);
  or _86748_ (_37501_, _37500_, _06464_);
  or _86749_ (_37502_, _37483_, _06465_);
  and _86750_ (_37503_, _37502_, _06269_);
  and _86751_ (_37505_, _37503_, _37501_);
  and _86752_ (_37506_, _15355_, _08630_);
  or _86753_ (_37507_, _37506_, _37490_);
  and _86754_ (_37508_, _37507_, _06268_);
  or _86755_ (_37509_, _37508_, _06261_);
  or _86756_ (_37510_, _37509_, _37505_);
  or _86757_ (_37511_, _37490_, _15387_);
  and _86758_ (_37512_, _37511_, _37492_);
  or _86759_ (_37513_, _37512_, _06262_);
  and _86760_ (_37514_, _37513_, _06258_);
  and _86761_ (_37516_, _37514_, _37510_);
  or _86762_ (_37517_, _37490_, _15403_);
  and _86763_ (_37518_, _37517_, _06257_);
  and _86764_ (_37519_, _37518_, _37492_);
  or _86765_ (_37520_, _37519_, _10080_);
  or _86766_ (_37521_, _37520_, _37516_);
  or _86767_ (_37522_, _37498_, _07215_);
  and _86768_ (_37523_, _37522_, _07208_);
  and _86769_ (_37524_, _37523_, _37521_);
  and _86770_ (_37525_, _09447_, _07935_);
  or _86771_ (_37527_, _37525_, _37477_);
  and _86772_ (_37528_, _37527_, _07460_);
  or _86773_ (_37529_, _37528_, _10094_);
  or _86774_ (_37530_, _37529_, _37524_);
  and _86775_ (_37531_, _15459_, _07935_);
  or _86776_ (_37532_, _37477_, _05982_);
  or _86777_ (_37533_, _37532_, _37531_);
  and _86778_ (_37534_, _37533_, _06219_);
  and _86779_ (_37535_, _37534_, _37530_);
  and _86780_ (_37536_, _08946_, _07935_);
  or _86781_ (_37538_, _37536_, _37477_);
  and _86782_ (_37539_, _37538_, _06218_);
  or _86783_ (_37540_, _37539_, _06369_);
  or _86784_ (_37541_, _37540_, _37535_);
  and _86785_ (_37542_, _15353_, _07935_);
  or _86786_ (_37543_, _37542_, _37477_);
  or _86787_ (_37544_, _37543_, _07237_);
  and _86788_ (_37545_, _37544_, _07240_);
  and _86789_ (_37546_, _37545_, _37541_);
  and _86790_ (_37547_, _11250_, _07935_);
  or _86791_ (_37549_, _37547_, _37477_);
  and _86792_ (_37550_, _37549_, _06536_);
  or _86793_ (_37551_, _37550_, _37546_);
  and _86794_ (_37552_, _37551_, _07242_);
  or _86795_ (_37553_, _37477_, _08247_);
  and _86796_ (_37554_, _37538_, _06375_);
  and _86797_ (_37555_, _37554_, _37553_);
  or _86798_ (_37556_, _37555_, _37552_);
  and _86799_ (_37557_, _37556_, _07234_);
  and _86800_ (_37558_, _37483_, _06545_);
  and _86801_ (_37560_, _37558_, _37553_);
  or _86802_ (_37561_, _37560_, _06366_);
  or _86803_ (_37562_, _37561_, _37557_);
  and _86804_ (_37563_, _15350_, _07935_);
  or _86805_ (_37564_, _37477_, _09056_);
  or _86806_ (_37565_, _37564_, _37563_);
  and _86807_ (_37566_, _37565_, _09061_);
  and _86808_ (_37567_, _37566_, _37562_);
  nor _86809_ (_37568_, _11249_, _14045_);
  or _86810_ (_37569_, _37568_, _37477_);
  and _86811_ (_37571_, _37569_, _06528_);
  or _86812_ (_37572_, _37571_, _06568_);
  or _86813_ (_37573_, _37572_, _37567_);
  or _86814_ (_37574_, _37479_, _06926_);
  and _86815_ (_37575_, _37574_, _05928_);
  and _86816_ (_37576_, _37575_, _37573_);
  and _86817_ (_37577_, _37507_, _05927_);
  or _86818_ (_37578_, _37577_, _06278_);
  or _86819_ (_37579_, _37578_, _37576_);
  and _86820_ (_37580_, _15532_, _07935_);
  or _86821_ (_37582_, _37477_, _06279_);
  or _86822_ (_37583_, _37582_, _37580_);
  and _86823_ (_37584_, _37583_, _01347_);
  and _86824_ (_37585_, _37584_, _37579_);
  or _86825_ (_37586_, _37585_, _37476_);
  and _86826_ (_43344_, _37586_, _42618_);
  nor _86827_ (_37587_, _01347_, _18157_);
  or _86828_ (_37588_, _11140_, _10519_);
  and _86829_ (_37589_, _37588_, _11097_);
  or _86830_ (_37590_, _11069_, _10592_);
  or _86831_ (_37592_, _37590_, _11084_);
  not _86832_ (_37593_, _11033_);
  or _86833_ (_37594_, _11056_, _10661_);
  or _86834_ (_37595_, _37594_, _37593_);
  nor _86835_ (_37596_, _07935_, _18157_);
  nor _86836_ (_37597_, _08142_, _14045_);
  or _86837_ (_37598_, _37597_, _37596_);
  or _86838_ (_37599_, _37598_, _07215_);
  nor _86839_ (_37600_, _08630_, _18157_);
  and _86840_ (_37601_, _15570_, _08630_);
  or _86841_ (_37603_, _37601_, _37600_);
  or _86842_ (_37604_, _37600_, _15585_);
  and _86843_ (_37605_, _37604_, _37603_);
  or _86844_ (_37606_, _37605_, _06262_);
  and _86845_ (_37607_, _15554_, _07935_);
  or _86846_ (_37608_, _37607_, _37596_);
  or _86847_ (_37609_, _37608_, _07151_);
  and _86848_ (_37610_, _07935_, \oc8051_golden_model_1.ACC [6]);
  or _86849_ (_37611_, _37610_, _37596_);
  and _86850_ (_37612_, _37611_, _07141_);
  nor _86851_ (_37614_, _07141_, _18157_);
  or _86852_ (_37615_, _37614_, _06341_);
  or _86853_ (_37616_, _37615_, _37612_);
  and _86854_ (_37617_, _37616_, _06273_);
  and _86855_ (_37618_, _37617_, _37609_);
  and _86856_ (_37619_, _37603_, _06272_);
  or _86857_ (_37620_, _37619_, _06461_);
  or _86858_ (_37621_, _37620_, _37618_);
  or _86859_ (_37622_, _37598_, _07166_);
  and _86860_ (_37623_, _37622_, _37621_);
  or _86861_ (_37625_, _37623_, _06464_);
  or _86862_ (_37626_, _37611_, _06465_);
  and _86863_ (_37627_, _37626_, _06269_);
  and _86864_ (_37628_, _37627_, _37625_);
  and _86865_ (_37629_, _15551_, _08630_);
  or _86866_ (_37630_, _37629_, _37600_);
  and _86867_ (_37631_, _37630_, _06268_);
  or _86868_ (_37632_, _37631_, _06261_);
  or _86869_ (_37633_, _37632_, _37628_);
  and _86870_ (_37634_, _37633_, _37606_);
  and _86871_ (_37636_, _37634_, _10735_);
  or _86872_ (_37637_, _10661_, _10656_);
  or _86873_ (_37638_, _37637_, _10717_);
  and _86874_ (_37639_, _37638_, _26197_);
  or _86875_ (_37640_, _37639_, _37636_);
  or _86876_ (_37641_, _10592_, _10588_);
  or _86877_ (_37642_, _37641_, _10641_);
  and _86878_ (_37643_, _37642_, _37640_);
  or _86879_ (_37644_, _37643_, _12644_);
  or _86880_ (_37645_, _10837_, _06517_);
  or _86881_ (_37647_, _37645_, _10888_);
  or _86882_ (_37648_, _10519_, _10517_);
  or _86883_ (_37649_, _37648_, _10574_);
  and _86884_ (_37650_, _37649_, _06258_);
  and _86885_ (_37651_, _37650_, _37647_);
  and _86886_ (_37652_, _37651_, _37644_);
  and _86887_ (_37653_, _15602_, _08630_);
  or _86888_ (_37654_, _37653_, _37600_);
  and _86889_ (_37655_, _37654_, _06257_);
  or _86890_ (_37656_, _37655_, _10080_);
  or _86891_ (_37658_, _37656_, _37652_);
  and _86892_ (_37659_, _37658_, _37599_);
  or _86893_ (_37660_, _37659_, _07460_);
  and _86894_ (_37661_, _09446_, _07935_);
  or _86895_ (_37662_, _37596_, _07208_);
  or _86896_ (_37663_, _37662_, _37661_);
  and _86897_ (_37664_, _37663_, _05982_);
  and _86898_ (_37665_, _37664_, _37660_);
  and _86899_ (_37666_, _15657_, _07935_);
  or _86900_ (_37667_, _37666_, _37596_);
  and _86901_ (_37669_, _37667_, _10094_);
  or _86902_ (_37670_, _37669_, _06218_);
  or _86903_ (_37671_, _37670_, _37665_);
  and _86904_ (_37672_, _15664_, _07935_);
  or _86905_ (_37673_, _37672_, _37596_);
  or _86906_ (_37674_, _37673_, _06219_);
  and _86907_ (_37675_, _37674_, _37671_);
  or _86908_ (_37676_, _37675_, _06369_);
  and _86909_ (_37677_, _15549_, _07935_);
  or _86910_ (_37678_, _37677_, _37596_);
  or _86911_ (_37680_, _37678_, _07237_);
  and _86912_ (_37681_, _37680_, _07240_);
  and _86913_ (_37682_, _37681_, _37676_);
  and _86914_ (_37683_, _11247_, _07935_);
  or _86915_ (_37684_, _37683_, _37596_);
  and _86916_ (_37685_, _37684_, _06536_);
  or _86917_ (_37686_, _37685_, _37682_);
  and _86918_ (_37687_, _37686_, _07242_);
  or _86919_ (_37688_, _37596_, _08145_);
  and _86920_ (_37689_, _37673_, _06375_);
  and _86921_ (_37691_, _37689_, _37688_);
  or _86922_ (_37692_, _37691_, _37687_);
  and _86923_ (_37693_, _37692_, _07234_);
  and _86924_ (_37694_, _37611_, _06545_);
  and _86925_ (_37695_, _37694_, _37688_);
  or _86926_ (_37696_, _37695_, _06366_);
  or _86927_ (_37697_, _37696_, _37693_);
  and _86928_ (_37698_, _15546_, _07935_);
  or _86929_ (_37699_, _37698_, _37596_);
  or _86930_ (_37700_, _37699_, _09056_);
  and _86931_ (_37702_, _37700_, _37697_);
  or _86932_ (_37703_, _37702_, _06528_);
  nor _86933_ (_37704_, _11246_, _14045_);
  or _86934_ (_37705_, _37704_, _37596_);
  nor _86935_ (_37706_, _37705_, _09061_);
  nor _86936_ (_37707_, _37706_, _11034_);
  and _86937_ (_37708_, _37707_, _37703_);
  and _86938_ (_37709_, _37594_, _11034_);
  or _86939_ (_37710_, _37709_, _11033_);
  or _86940_ (_37711_, _37710_, _37708_);
  and _86941_ (_37713_, _37711_, _37595_);
  or _86942_ (_37714_, _37713_, _17504_);
  not _86943_ (_37715_, _17504_);
  or _86944_ (_37716_, _37594_, _37715_);
  and _86945_ (_37717_, _37716_, _17724_);
  and _86946_ (_37718_, _37717_, _37714_);
  and _86947_ (_37719_, _37594_, _17723_);
  or _86948_ (_37720_, _37719_, _11041_);
  or _86949_ (_37721_, _37720_, _37718_);
  and _86950_ (_37722_, _37721_, _37592_);
  or _86951_ (_37724_, _37722_, _06540_);
  or _86952_ (_37725_, _10837_, _06541_);
  or _86953_ (_37726_, _37725_, _11112_);
  and _86954_ (_37727_, _37726_, _11127_);
  and _86955_ (_37728_, _37727_, _37724_);
  or _86956_ (_37729_, _37728_, _37589_);
  and _86957_ (_37730_, _37729_, _11157_);
  and _86958_ (_37731_, _11186_, _18059_);
  or _86959_ (_37732_, _37731_, _11201_);
  or _86960_ (_37733_, _37732_, _37730_);
  or _86961_ (_37735_, _11230_, _11203_);
  and _86962_ (_37736_, _37735_, _06285_);
  and _86963_ (_37737_, _37736_, _37733_);
  and _86964_ (_37738_, _11270_, _06283_);
  or _86965_ (_37739_, _37738_, _11243_);
  or _86966_ (_37740_, _37739_, _37737_);
  or _86967_ (_37741_, _11313_, _11321_);
  and _86968_ (_37742_, _37741_, _37740_);
  or _86969_ (_37743_, _37742_, _06568_);
  or _86970_ (_37744_, _37608_, _06926_);
  and _86971_ (_37746_, _37744_, _05928_);
  and _86972_ (_37747_, _37746_, _37743_);
  and _86973_ (_37748_, _37630_, _05927_);
  or _86974_ (_37749_, _37748_, _06278_);
  or _86975_ (_37750_, _37749_, _37747_);
  and _86976_ (_37751_, _15734_, _07935_);
  or _86977_ (_37752_, _37596_, _06279_);
  or _86978_ (_37753_, _37752_, _37751_);
  and _86979_ (_37754_, _37753_, _01347_);
  and _86980_ (_37755_, _37754_, _37750_);
  or _86981_ (_37757_, _37755_, _37587_);
  and _86982_ (_43345_, _37757_, _42618_);
  and _86983_ (_37758_, _05938_, op0_cnst);
  or _86984_ (_00000_, _37758_, rst);
  and _86985_ (_37759_, _37758_, _01347_);
  and _86986_ (_37760_, _25696_, _01960_);
  nor _86987_ (_37761_, _25696_, _01960_);
  or _86988_ (_37762_, _37761_, _37760_);
  and _86989_ (_37763_, _26055_, _01964_);
  nor _86990_ (_37764_, _26055_, _01964_);
  nand _86991_ (_37766_, _26747_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _86992_ (_37767_, _26747_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _86993_ (_37768_, _37767_, _37766_);
  nor _86994_ (_37769_, _27450_, _01979_);
  and _86995_ (_37770_, _27450_, _01979_);
  or _86996_ (_37771_, _37770_, _37769_);
  nor _86997_ (_37772_, _27099_, _01975_);
  nor _86998_ (_37773_, _26404_, _01968_);
  and _86999_ (_37774_, _27099_, _01975_);
  or _87000_ (_37775_, _37774_, _37773_);
  or _87001_ (_37777_, _37775_, _37772_);
  nor _87002_ (_37778_, _27805_, _01983_);
  and _87003_ (_37779_, _28456_, _38291_);
  nor _87004_ (_37780_, _28456_, _38291_);
  nor _87005_ (_37781_, _28133_, _38285_);
  and _87006_ (_37782_, _28133_, _38285_);
  and _87007_ (_37783_, _29063_, _38281_);
  nor _87008_ (_37784_, _29063_, _38281_);
  nor _87009_ (_37785_, _29667_, _38307_);
  or _87010_ (_37786_, _37785_, _37784_);
  or _87011_ (_37788_, _37786_, _37783_);
  nor _87012_ (_37789_, _13073_, _38317_);
  and _87013_ (_37790_, _13073_, _38317_);
  and _87014_ (_37791_, _29667_, _38307_);
  and _87015_ (_37792_, _28759_, _38296_);
  and _87016_ (_37793_, _25306_, _01956_);
  nor _87017_ (_37794_, _25306_, _01956_);
  or _87018_ (_37795_, _37794_, _37793_);
  nor _87019_ (_37796_, _28759_, _38296_);
  or _87020_ (_37797_, _37796_, _37795_);
  or _87021_ (_37799_, _37797_, _37792_);
  and _87022_ (_37800_, _29366_, _38302_);
  nor _87023_ (_37801_, _29366_, _38302_);
  or _87024_ (_37802_, _37801_, _37800_);
  and _87025_ (_37803_, _29970_, _38312_);
  nor _87026_ (_37804_, _29970_, _38312_);
  or _87027_ (_37805_, _37804_, _37803_);
  or _87028_ (_37806_, _37805_, _37802_);
  or _87029_ (_37807_, _37806_, _37799_);
  or _87030_ (_37808_, _37807_, _37791_);
  or _87031_ (_37810_, _37808_, _37790_);
  or _87032_ (_37811_, _37810_, _37789_);
  or _87033_ (_37812_, _37811_, _37788_);
  or _87034_ (_37813_, _37812_, _37782_);
  or _87035_ (_37814_, _37813_, _37781_);
  or _87036_ (_37815_, _37814_, _37780_);
  or _87037_ (_37816_, _37815_, _37779_);
  or _87038_ (_37817_, _37816_, _37778_);
  and _87039_ (_37818_, _26404_, _01968_);
  and _87040_ (_37819_, _27805_, _01983_);
  or _87041_ (_37821_, _37819_, _37818_);
  or _87042_ (_37822_, _37821_, _37817_);
  or _87043_ (_37823_, _37822_, _37777_);
  or _87044_ (_37824_, _37823_, _37771_);
  or _87045_ (_37825_, _37824_, _37768_);
  or _87046_ (_37826_, _37825_, _37764_);
  or _87047_ (_37827_, _37826_, _37763_);
  or _87048_ (_37828_, _37827_, _37762_);
  and _87049_ (property_invalid_pc, _37828_, _37759_);
  buf _87050_ (_00543_, _42621_);
  buf _87051_ (_05076_, _42618_);
  buf _87052_ (_05127_, _42618_);
  buf _87053_ (_05179_, _42618_);
  buf _87054_ (_05230_, _42618_);
  buf _87055_ (_05282_, _42618_);
  buf _87056_ (_05334_, _42618_);
  buf _87057_ (_05385_, _42618_);
  buf _87058_ (_05437_, _42618_);
  buf _87059_ (_05488_, _42618_);
  buf _87060_ (_05540_, _42618_);
  buf _87061_ (_05591_, _42618_);
  buf _87062_ (_05644_, _42618_);
  buf _87063_ (_05697_, _42618_);
  buf _87064_ (_05750_, _42618_);
  buf _87065_ (_05803_, _42618_);
  buf _87066_ (_05856_, _42618_);
  buf _87067_ (_38745_, _38644_);
  buf _87068_ (_38747_, _38646_);
  buf _87069_ (_38760_, _38644_);
  buf _87070_ (_38761_, _38646_);
  buf _87071_ (_39074_, _38664_);
  buf _87072_ (_39075_, _38665_);
  buf _87073_ (_39076_, _38667_);
  buf _87074_ (_39077_, _38668_);
  buf _87075_ (_39078_, _38669_);
  buf _87076_ (_39079_, _38670_);
  buf _87077_ (_39080_, _38671_);
  buf _87078_ (_39081_, _38673_);
  buf _87079_ (_39082_, _38674_);
  buf _87080_ (_39084_, _38675_);
  buf _87081_ (_39085_, _38676_);
  buf _87082_ (_39086_, _38677_);
  buf _87083_ (_39087_, _38679_);
  buf _87084_ (_39088_, _38680_);
  buf _87085_ (_39140_, _38664_);
  buf _87086_ (_39141_, _38665_);
  buf _87087_ (_39142_, _38667_);
  buf _87088_ (_39143_, _38668_);
  buf _87089_ (_39144_, _38669_);
  buf _87090_ (_39145_, _38670_);
  buf _87091_ (_39146_, _38671_);
  buf _87092_ (_39147_, _38673_);
  buf _87093_ (_39148_, _38674_);
  buf _87094_ (_39150_, _38675_);
  buf _87095_ (_39151_, _38676_);
  buf _87096_ (_39152_, _38677_);
  buf _87097_ (_39153_, _38679_);
  buf _87098_ (_39154_, _38680_);
  buf _87099_ (_39685_, _39457_);
  buf _87100_ (_39845_, _39457_);
  dff _87101_ (op0_cnst, _00000_, clk);
  dff _87102_ (\oc8051_gm_cxrom_1.cell0.data [0], _05080_, clk);
  dff _87103_ (\oc8051_gm_cxrom_1.cell0.data [1], _05083_, clk);
  dff _87104_ (\oc8051_gm_cxrom_1.cell0.data [2], _05087_, clk);
  dff _87105_ (\oc8051_gm_cxrom_1.cell0.data [3], _05091_, clk);
  dff _87106_ (\oc8051_gm_cxrom_1.cell0.data [4], _05095_, clk);
  dff _87107_ (\oc8051_gm_cxrom_1.cell0.data [5], _05099_, clk);
  dff _87108_ (\oc8051_gm_cxrom_1.cell0.data [6], _05103_, clk);
  dff _87109_ (\oc8051_gm_cxrom_1.cell0.data [7], _05073_, clk);
  dff _87110_ (\oc8051_gm_cxrom_1.cell0.valid , _05076_, clk);
  dff _87111_ (\oc8051_gm_cxrom_1.cell1.data [0], _05131_, clk);
  dff _87112_ (\oc8051_gm_cxrom_1.cell1.data [1], _05135_, clk);
  dff _87113_ (\oc8051_gm_cxrom_1.cell1.data [2], _05139_, clk);
  dff _87114_ (\oc8051_gm_cxrom_1.cell1.data [3], _05143_, clk);
  dff _87115_ (\oc8051_gm_cxrom_1.cell1.data [4], _05147_, clk);
  dff _87116_ (\oc8051_gm_cxrom_1.cell1.data [5], _05151_, clk);
  dff _87117_ (\oc8051_gm_cxrom_1.cell1.data [6], _05155_, clk);
  dff _87118_ (\oc8051_gm_cxrom_1.cell1.data [7], _05124_, clk);
  dff _87119_ (\oc8051_gm_cxrom_1.cell1.valid , _05127_, clk);
  dff _87120_ (\oc8051_gm_cxrom_1.cell10.data [0], _05595_, clk);
  dff _87121_ (\oc8051_gm_cxrom_1.cell10.data [1], _05599_, clk);
  dff _87122_ (\oc8051_gm_cxrom_1.cell10.data [2], _05603_, clk);
  dff _87123_ (\oc8051_gm_cxrom_1.cell10.data [3], _05607_, clk);
  dff _87124_ (\oc8051_gm_cxrom_1.cell10.data [4], _05611_, clk);
  dff _87125_ (\oc8051_gm_cxrom_1.cell10.data [5], _05615_, clk);
  dff _87126_ (\oc8051_gm_cxrom_1.cell10.data [6], _05619_, clk);
  dff _87127_ (\oc8051_gm_cxrom_1.cell10.data [7], _05589_, clk);
  dff _87128_ (\oc8051_gm_cxrom_1.cell10.valid , _05591_, clk);
  dff _87129_ (\oc8051_gm_cxrom_1.cell11.data [0], _05648_, clk);
  dff _87130_ (\oc8051_gm_cxrom_1.cell11.data [1], _05652_, clk);
  dff _87131_ (\oc8051_gm_cxrom_1.cell11.data [2], _05656_, clk);
  dff _87132_ (\oc8051_gm_cxrom_1.cell11.data [3], _05660_, clk);
  dff _87133_ (\oc8051_gm_cxrom_1.cell11.data [4], _05664_, clk);
  dff _87134_ (\oc8051_gm_cxrom_1.cell11.data [5], _05668_, clk);
  dff _87135_ (\oc8051_gm_cxrom_1.cell11.data [6], _05672_, clk);
  dff _87136_ (\oc8051_gm_cxrom_1.cell11.data [7], _05641_, clk);
  dff _87137_ (\oc8051_gm_cxrom_1.cell11.valid , _05644_, clk);
  dff _87138_ (\oc8051_gm_cxrom_1.cell12.data [0], _05701_, clk);
  dff _87139_ (\oc8051_gm_cxrom_1.cell12.data [1], _05705_, clk);
  dff _87140_ (\oc8051_gm_cxrom_1.cell12.data [2], _05709_, clk);
  dff _87141_ (\oc8051_gm_cxrom_1.cell12.data [3], _05713_, clk);
  dff _87142_ (\oc8051_gm_cxrom_1.cell12.data [4], _05717_, clk);
  dff _87143_ (\oc8051_gm_cxrom_1.cell12.data [5], _05721_, clk);
  dff _87144_ (\oc8051_gm_cxrom_1.cell12.data [6], _05725_, clk);
  dff _87145_ (\oc8051_gm_cxrom_1.cell12.data [7], _05694_, clk);
  dff _87146_ (\oc8051_gm_cxrom_1.cell12.valid , _05697_, clk);
  dff _87147_ (\oc8051_gm_cxrom_1.cell13.data [0], _05754_, clk);
  dff _87148_ (\oc8051_gm_cxrom_1.cell13.data [1], _05758_, clk);
  dff _87149_ (\oc8051_gm_cxrom_1.cell13.data [2], _05762_, clk);
  dff _87150_ (\oc8051_gm_cxrom_1.cell13.data [3], _05766_, clk);
  dff _87151_ (\oc8051_gm_cxrom_1.cell13.data [4], _05770_, clk);
  dff _87152_ (\oc8051_gm_cxrom_1.cell13.data [5], _05774_, clk);
  dff _87153_ (\oc8051_gm_cxrom_1.cell13.data [6], _05778_, clk);
  dff _87154_ (\oc8051_gm_cxrom_1.cell13.data [7], _05747_, clk);
  dff _87155_ (\oc8051_gm_cxrom_1.cell13.valid , _05750_, clk);
  dff _87156_ (\oc8051_gm_cxrom_1.cell14.data [0], _05807_, clk);
  dff _87157_ (\oc8051_gm_cxrom_1.cell14.data [1], _05811_, clk);
  dff _87158_ (\oc8051_gm_cxrom_1.cell14.data [2], _05815_, clk);
  dff _87159_ (\oc8051_gm_cxrom_1.cell14.data [3], _05819_, clk);
  dff _87160_ (\oc8051_gm_cxrom_1.cell14.data [4], _05823_, clk);
  dff _87161_ (\oc8051_gm_cxrom_1.cell14.data [5], _05827_, clk);
  dff _87162_ (\oc8051_gm_cxrom_1.cell14.data [6], _05831_, clk);
  dff _87163_ (\oc8051_gm_cxrom_1.cell14.data [7], _05800_, clk);
  dff _87164_ (\oc8051_gm_cxrom_1.cell14.valid , _05803_, clk);
  dff _87165_ (\oc8051_gm_cxrom_1.cell15.data [0], _05860_, clk);
  dff _87166_ (\oc8051_gm_cxrom_1.cell15.data [1], _05864_, clk);
  dff _87167_ (\oc8051_gm_cxrom_1.cell15.data [2], _05868_, clk);
  dff _87168_ (\oc8051_gm_cxrom_1.cell15.data [3], _05872_, clk);
  dff _87169_ (\oc8051_gm_cxrom_1.cell15.data [4], _05876_, clk);
  dff _87170_ (\oc8051_gm_cxrom_1.cell15.data [5], _05880_, clk);
  dff _87171_ (\oc8051_gm_cxrom_1.cell15.data [6], _05884_, clk);
  dff _87172_ (\oc8051_gm_cxrom_1.cell15.data [7], _05853_, clk);
  dff _87173_ (\oc8051_gm_cxrom_1.cell15.valid , _05856_, clk);
  dff _87174_ (\oc8051_gm_cxrom_1.cell2.data [0], _05183_, clk);
  dff _87175_ (\oc8051_gm_cxrom_1.cell2.data [1], _05187_, clk);
  dff _87176_ (\oc8051_gm_cxrom_1.cell2.data [2], _05191_, clk);
  dff _87177_ (\oc8051_gm_cxrom_1.cell2.data [3], _05194_, clk);
  dff _87178_ (\oc8051_gm_cxrom_1.cell2.data [4], _05198_, clk);
  dff _87179_ (\oc8051_gm_cxrom_1.cell2.data [5], _05202_, clk);
  dff _87180_ (\oc8051_gm_cxrom_1.cell2.data [6], _05206_, clk);
  dff _87181_ (\oc8051_gm_cxrom_1.cell2.data [7], _05176_, clk);
  dff _87182_ (\oc8051_gm_cxrom_1.cell2.valid , _05179_, clk);
  dff _87183_ (\oc8051_gm_cxrom_1.cell3.data [0], _05234_, clk);
  dff _87184_ (\oc8051_gm_cxrom_1.cell3.data [1], _05238_, clk);
  dff _87185_ (\oc8051_gm_cxrom_1.cell3.data [2], _05242_, clk);
  dff _87186_ (\oc8051_gm_cxrom_1.cell3.data [3], _05246_, clk);
  dff _87187_ (\oc8051_gm_cxrom_1.cell3.data [4], _05250_, clk);
  dff _87188_ (\oc8051_gm_cxrom_1.cell3.data [5], _05254_, clk);
  dff _87189_ (\oc8051_gm_cxrom_1.cell3.data [6], _05258_, clk);
  dff _87190_ (\oc8051_gm_cxrom_1.cell3.data [7], _05227_, clk);
  dff _87191_ (\oc8051_gm_cxrom_1.cell3.valid , _05230_, clk);
  dff _87192_ (\oc8051_gm_cxrom_1.cell4.data [0], _05286_, clk);
  dff _87193_ (\oc8051_gm_cxrom_1.cell4.data [1], _05290_, clk);
  dff _87194_ (\oc8051_gm_cxrom_1.cell4.data [2], _05294_, clk);
  dff _87195_ (\oc8051_gm_cxrom_1.cell4.data [3], _05298_, clk);
  dff _87196_ (\oc8051_gm_cxrom_1.cell4.data [4], _05301_, clk);
  dff _87197_ (\oc8051_gm_cxrom_1.cell4.data [5], _05305_, clk);
  dff _87198_ (\oc8051_gm_cxrom_1.cell4.data [6], _05309_, clk);
  dff _87199_ (\oc8051_gm_cxrom_1.cell4.data [7], _05279_, clk);
  dff _87200_ (\oc8051_gm_cxrom_1.cell4.valid , _05282_, clk);
  dff _87201_ (\oc8051_gm_cxrom_1.cell5.data [0], _05337_, clk);
  dff _87202_ (\oc8051_gm_cxrom_1.cell5.data [1], _05341_, clk);
  dff _87203_ (\oc8051_gm_cxrom_1.cell5.data [2], _05345_, clk);
  dff _87204_ (\oc8051_gm_cxrom_1.cell5.data [3], _05349_, clk);
  dff _87205_ (\oc8051_gm_cxrom_1.cell5.data [4], _05353_, clk);
  dff _87206_ (\oc8051_gm_cxrom_1.cell5.data [5], _05357_, clk);
  dff _87207_ (\oc8051_gm_cxrom_1.cell5.data [6], _05361_, clk);
  dff _87208_ (\oc8051_gm_cxrom_1.cell5.data [7], _05331_, clk);
  dff _87209_ (\oc8051_gm_cxrom_1.cell5.valid , _05334_, clk);
  dff _87210_ (\oc8051_gm_cxrom_1.cell6.data [0], _05389_, clk);
  dff _87211_ (\oc8051_gm_cxrom_1.cell6.data [1], _05393_, clk);
  dff _87212_ (\oc8051_gm_cxrom_1.cell6.data [2], _05397_, clk);
  dff _87213_ (\oc8051_gm_cxrom_1.cell6.data [3], _05401_, clk);
  dff _87214_ (\oc8051_gm_cxrom_1.cell6.data [4], _05405_, clk);
  dff _87215_ (\oc8051_gm_cxrom_1.cell6.data [5], _05409_, clk);
  dff _87216_ (\oc8051_gm_cxrom_1.cell6.data [6], _05412_, clk);
  dff _87217_ (\oc8051_gm_cxrom_1.cell6.data [7], _05382_, clk);
  dff _87218_ (\oc8051_gm_cxrom_1.cell6.valid , _05385_, clk);
  dff _87219_ (\oc8051_gm_cxrom_1.cell7.data [0], _05441_, clk);
  dff _87220_ (\oc8051_gm_cxrom_1.cell7.data [1], _05445_, clk);
  dff _87221_ (\oc8051_gm_cxrom_1.cell7.data [2], _05448_, clk);
  dff _87222_ (\oc8051_gm_cxrom_1.cell7.data [3], _05452_, clk);
  dff _87223_ (\oc8051_gm_cxrom_1.cell7.data [4], _05456_, clk);
  dff _87224_ (\oc8051_gm_cxrom_1.cell7.data [5], _05460_, clk);
  dff _87225_ (\oc8051_gm_cxrom_1.cell7.data [6], _05464_, clk);
  dff _87226_ (\oc8051_gm_cxrom_1.cell7.data [7], _05434_, clk);
  dff _87227_ (\oc8051_gm_cxrom_1.cell7.valid , _05437_, clk);
  dff _87228_ (\oc8051_gm_cxrom_1.cell8.data [0], _05492_, clk);
  dff _87229_ (\oc8051_gm_cxrom_1.cell8.data [1], _05496_, clk);
  dff _87230_ (\oc8051_gm_cxrom_1.cell8.data [2], _05500_, clk);
  dff _87231_ (\oc8051_gm_cxrom_1.cell8.data [3], _05504_, clk);
  dff _87232_ (\oc8051_gm_cxrom_1.cell8.data [4], _05508_, clk);
  dff _87233_ (\oc8051_gm_cxrom_1.cell8.data [5], _05512_, clk);
  dff _87234_ (\oc8051_gm_cxrom_1.cell8.data [6], _05516_, clk);
  dff _87235_ (\oc8051_gm_cxrom_1.cell8.data [7], _05485_, clk);
  dff _87236_ (\oc8051_gm_cxrom_1.cell8.valid , _05488_, clk);
  dff _87237_ (\oc8051_gm_cxrom_1.cell9.data [0], _05544_, clk);
  dff _87238_ (\oc8051_gm_cxrom_1.cell9.data [1], _05548_, clk);
  dff _87239_ (\oc8051_gm_cxrom_1.cell9.data [2], _05552_, clk);
  dff _87240_ (\oc8051_gm_cxrom_1.cell9.data [3], _05555_, clk);
  dff _87241_ (\oc8051_gm_cxrom_1.cell9.data [4], _05559_, clk);
  dff _87242_ (\oc8051_gm_cxrom_1.cell9.data [5], _05563_, clk);
  dff _87243_ (\oc8051_gm_cxrom_1.cell9.data [6], _05567_, clk);
  dff _87244_ (\oc8051_gm_cxrom_1.cell9.data [7], _05537_, clk);
  dff _87245_ (\oc8051_gm_cxrom_1.cell9.valid , _05540_, clk);
  dff _87246_ (\oc8051_golden_model_1.IRAM[15] [0], _40795_, clk);
  dff _87247_ (\oc8051_golden_model_1.IRAM[15] [1], _40796_, clk);
  dff _87248_ (\oc8051_golden_model_1.IRAM[15] [2], _40797_, clk);
  dff _87249_ (\oc8051_golden_model_1.IRAM[15] [3], _40799_, clk);
  dff _87250_ (\oc8051_golden_model_1.IRAM[15] [4], _40800_, clk);
  dff _87251_ (\oc8051_golden_model_1.IRAM[15] [5], _40801_, clk);
  dff _87252_ (\oc8051_golden_model_1.IRAM[15] [6], _40802_, clk);
  dff _87253_ (\oc8051_golden_model_1.IRAM[15] [7], _40572_, clk);
  dff _87254_ (\oc8051_golden_model_1.IRAM[14] [0], _40783_, clk);
  dff _87255_ (\oc8051_golden_model_1.IRAM[14] [1], _40784_, clk);
  dff _87256_ (\oc8051_golden_model_1.IRAM[14] [2], _40785_, clk);
  dff _87257_ (\oc8051_golden_model_1.IRAM[14] [3], _40787_, clk);
  dff _87258_ (\oc8051_golden_model_1.IRAM[14] [4], _40788_, clk);
  dff _87259_ (\oc8051_golden_model_1.IRAM[14] [5], _40789_, clk);
  dff _87260_ (\oc8051_golden_model_1.IRAM[14] [6], _40790_, clk);
  dff _87261_ (\oc8051_golden_model_1.IRAM[14] [7], _40791_, clk);
  dff _87262_ (\oc8051_golden_model_1.IRAM[13] [0], _40771_, clk);
  dff _87263_ (\oc8051_golden_model_1.IRAM[13] [1], _40772_, clk);
  dff _87264_ (\oc8051_golden_model_1.IRAM[13] [2], _40773_, clk);
  dff _87265_ (\oc8051_golden_model_1.IRAM[13] [3], _40774_, clk);
  dff _87266_ (\oc8051_golden_model_1.IRAM[13] [4], _40776_, clk);
  dff _87267_ (\oc8051_golden_model_1.IRAM[13] [5], _40777_, clk);
  dff _87268_ (\oc8051_golden_model_1.IRAM[13] [6], _40778_, clk);
  dff _87269_ (\oc8051_golden_model_1.IRAM[13] [7], _40779_, clk);
  dff _87270_ (\oc8051_golden_model_1.IRAM[12] [0], _40759_, clk);
  dff _87271_ (\oc8051_golden_model_1.IRAM[12] [1], _40760_, clk);
  dff _87272_ (\oc8051_golden_model_1.IRAM[12] [2], _40761_, clk);
  dff _87273_ (\oc8051_golden_model_1.IRAM[12] [3], _40762_, clk);
  dff _87274_ (\oc8051_golden_model_1.IRAM[12] [4], _40764_, clk);
  dff _87275_ (\oc8051_golden_model_1.IRAM[12] [5], _40765_, clk);
  dff _87276_ (\oc8051_golden_model_1.IRAM[12] [6], _40766_, clk);
  dff _87277_ (\oc8051_golden_model_1.IRAM[12] [7], _40767_, clk);
  dff _87278_ (\oc8051_golden_model_1.IRAM[11] [0], _40746_, clk);
  dff _87279_ (\oc8051_golden_model_1.IRAM[11] [1], _40748_, clk);
  dff _87280_ (\oc8051_golden_model_1.IRAM[11] [2], _40749_, clk);
  dff _87281_ (\oc8051_golden_model_1.IRAM[11] [3], _40750_, clk);
  dff _87282_ (\oc8051_golden_model_1.IRAM[11] [4], _40751_, clk);
  dff _87283_ (\oc8051_golden_model_1.IRAM[11] [5], _40752_, clk);
  dff _87284_ (\oc8051_golden_model_1.IRAM[11] [6], _40754_, clk);
  dff _87285_ (\oc8051_golden_model_1.IRAM[11] [7], _40755_, clk);
  dff _87286_ (\oc8051_golden_model_1.IRAM[10] [0], _40734_, clk);
  dff _87287_ (\oc8051_golden_model_1.IRAM[10] [1], _40736_, clk);
  dff _87288_ (\oc8051_golden_model_1.IRAM[10] [2], _40737_, clk);
  dff _87289_ (\oc8051_golden_model_1.IRAM[10] [3], _40738_, clk);
  dff _87290_ (\oc8051_golden_model_1.IRAM[10] [4], _40739_, clk);
  dff _87291_ (\oc8051_golden_model_1.IRAM[10] [5], _40740_, clk);
  dff _87292_ (\oc8051_golden_model_1.IRAM[10] [6], _40742_, clk);
  dff _87293_ (\oc8051_golden_model_1.IRAM[10] [7], _40743_, clk);
  dff _87294_ (\oc8051_golden_model_1.IRAM[9] [0], _40723_, clk);
  dff _87295_ (\oc8051_golden_model_1.IRAM[9] [1], _40724_, clk);
  dff _87296_ (\oc8051_golden_model_1.IRAM[9] [2], _40726_, clk);
  dff _87297_ (\oc8051_golden_model_1.IRAM[9] [3], _40727_, clk);
  dff _87298_ (\oc8051_golden_model_1.IRAM[9] [4], _40728_, clk);
  dff _87299_ (\oc8051_golden_model_1.IRAM[9] [5], _40729_, clk);
  dff _87300_ (\oc8051_golden_model_1.IRAM[9] [6], _40730_, clk);
  dff _87301_ (\oc8051_golden_model_1.IRAM[9] [7], _40732_, clk);
  dff _87302_ (\oc8051_golden_model_1.IRAM[8] [0], _40711_, clk);
  dff _87303_ (\oc8051_golden_model_1.IRAM[8] [1], _40712_, clk);
  dff _87304_ (\oc8051_golden_model_1.IRAM[8] [2], _40714_, clk);
  dff _87305_ (\oc8051_golden_model_1.IRAM[8] [3], _40715_, clk);
  dff _87306_ (\oc8051_golden_model_1.IRAM[8] [4], _40716_, clk);
  dff _87307_ (\oc8051_golden_model_1.IRAM[8] [5], _40717_, clk);
  dff _87308_ (\oc8051_golden_model_1.IRAM[8] [6], _40718_, clk);
  dff _87309_ (\oc8051_golden_model_1.IRAM[8] [7], _40720_, clk);
  dff _87310_ (\oc8051_golden_model_1.IRAM[7] [0], _40698_, clk);
  dff _87311_ (\oc8051_golden_model_1.IRAM[7] [1], _40700_, clk);
  dff _87312_ (\oc8051_golden_model_1.IRAM[7] [2], _40701_, clk);
  dff _87313_ (\oc8051_golden_model_1.IRAM[7] [3], _40702_, clk);
  dff _87314_ (\oc8051_golden_model_1.IRAM[7] [4], _40703_, clk);
  dff _87315_ (\oc8051_golden_model_1.IRAM[7] [5], _40704_, clk);
  dff _87316_ (\oc8051_golden_model_1.IRAM[7] [6], _40706_, clk);
  dff _87317_ (\oc8051_golden_model_1.IRAM[7] [7], _40707_, clk);
  dff _87318_ (\oc8051_golden_model_1.IRAM[6] [0], _40685_, clk);
  dff _87319_ (\oc8051_golden_model_1.IRAM[6] [1], _40688_, clk);
  dff _87320_ (\oc8051_golden_model_1.IRAM[6] [2], _40689_, clk);
  dff _87321_ (\oc8051_golden_model_1.IRAM[6] [3], _40690_, clk);
  dff _87322_ (\oc8051_golden_model_1.IRAM[6] [4], _40691_, clk);
  dff _87323_ (\oc8051_golden_model_1.IRAM[6] [5], _40692_, clk);
  dff _87324_ (\oc8051_golden_model_1.IRAM[6] [6], _40694_, clk);
  dff _87325_ (\oc8051_golden_model_1.IRAM[6] [7], _40695_, clk);
  dff _87326_ (\oc8051_golden_model_1.IRAM[5] [0], _40673_, clk);
  dff _87327_ (\oc8051_golden_model_1.IRAM[5] [1], _40674_, clk);
  dff _87328_ (\oc8051_golden_model_1.IRAM[5] [2], _40677_, clk);
  dff _87329_ (\oc8051_golden_model_1.IRAM[5] [3], _40678_, clk);
  dff _87330_ (\oc8051_golden_model_1.IRAM[5] [4], _40679_, clk);
  dff _87331_ (\oc8051_golden_model_1.IRAM[5] [5], _40680_, clk);
  dff _87332_ (\oc8051_golden_model_1.IRAM[5] [6], _40681_, clk);
  dff _87333_ (\oc8051_golden_model_1.IRAM[5] [7], _40683_, clk);
  dff _87334_ (\oc8051_golden_model_1.IRAM[4] [0], _40662_, clk);
  dff _87335_ (\oc8051_golden_model_1.IRAM[4] [1], _40663_, clk);
  dff _87336_ (\oc8051_golden_model_1.IRAM[4] [2], _40665_, clk);
  dff _87337_ (\oc8051_golden_model_1.IRAM[4] [3], _40666_, clk);
  dff _87338_ (\oc8051_golden_model_1.IRAM[4] [4], _40667_, clk);
  dff _87339_ (\oc8051_golden_model_1.IRAM[4] [5], _40668_, clk);
  dff _87340_ (\oc8051_golden_model_1.IRAM[4] [6], _40669_, clk);
  dff _87341_ (\oc8051_golden_model_1.IRAM[4] [7], _40671_, clk);
  dff _87342_ (\oc8051_golden_model_1.IRAM[3] [0], _40649_, clk);
  dff _87343_ (\oc8051_golden_model_1.IRAM[3] [1], _40651_, clk);
  dff _87344_ (\oc8051_golden_model_1.IRAM[3] [2], _40652_, clk);
  dff _87345_ (\oc8051_golden_model_1.IRAM[3] [3], _40653_, clk);
  dff _87346_ (\oc8051_golden_model_1.IRAM[3] [4], _40654_, clk);
  dff _87347_ (\oc8051_golden_model_1.IRAM[3] [5], _40655_, clk);
  dff _87348_ (\oc8051_golden_model_1.IRAM[3] [6], _40657_, clk);
  dff _87349_ (\oc8051_golden_model_1.IRAM[3] [7], _40658_, clk);
  dff _87350_ (\oc8051_golden_model_1.IRAM[2] [0], _40637_, clk);
  dff _87351_ (\oc8051_golden_model_1.IRAM[2] [1], _40638_, clk);
  dff _87352_ (\oc8051_golden_model_1.IRAM[2] [2], _40640_, clk);
  dff _87353_ (\oc8051_golden_model_1.IRAM[2] [3], _40641_, clk);
  dff _87354_ (\oc8051_golden_model_1.IRAM[2] [4], _40642_, clk);
  dff _87355_ (\oc8051_golden_model_1.IRAM[2] [5], _40643_, clk);
  dff _87356_ (\oc8051_golden_model_1.IRAM[2] [6], _40644_, clk);
  dff _87357_ (\oc8051_golden_model_1.IRAM[2] [7], _40646_, clk);
  dff _87358_ (\oc8051_golden_model_1.IRAM[1] [0], _40623_, clk);
  dff _87359_ (\oc8051_golden_model_1.IRAM[1] [1], _40626_, clk);
  dff _87360_ (\oc8051_golden_model_1.IRAM[1] [2], _40627_, clk);
  dff _87361_ (\oc8051_golden_model_1.IRAM[1] [3], _40628_, clk);
  dff _87362_ (\oc8051_golden_model_1.IRAM[1] [4], _40629_, clk);
  dff _87363_ (\oc8051_golden_model_1.IRAM[1] [5], _40630_, clk);
  dff _87364_ (\oc8051_golden_model_1.IRAM[1] [6], _40632_, clk);
  dff _87365_ (\oc8051_golden_model_1.IRAM[1] [7], _40633_, clk);
  dff _87366_ (\oc8051_golden_model_1.B [0], _43153_, clk);
  dff _87367_ (\oc8051_golden_model_1.B [1], _43154_, clk);
  dff _87368_ (\oc8051_golden_model_1.B [2], _43155_, clk);
  dff _87369_ (\oc8051_golden_model_1.B [3], _43156_, clk);
  dff _87370_ (\oc8051_golden_model_1.B [4], _43157_, clk);
  dff _87371_ (\oc8051_golden_model_1.B [5], _43159_, clk);
  dff _87372_ (\oc8051_golden_model_1.B [6], _43160_, clk);
  dff _87373_ (\oc8051_golden_model_1.B [7], _40573_, clk);
  dff _87374_ (\oc8051_golden_model_1.ACC [0], _43161_, clk);
  dff _87375_ (\oc8051_golden_model_1.ACC [1], _43163_, clk);
  dff _87376_ (\oc8051_golden_model_1.ACC [2], _43164_, clk);
  dff _87377_ (\oc8051_golden_model_1.ACC [3], _43165_, clk);
  dff _87378_ (\oc8051_golden_model_1.ACC [4], _43166_, clk);
  dff _87379_ (\oc8051_golden_model_1.ACC [5], _43167_, clk);
  dff _87380_ (\oc8051_golden_model_1.ACC [6], _43168_, clk);
  dff _87381_ (\oc8051_golden_model_1.ACC [7], _40574_, clk);
  dff _87382_ (\oc8051_golden_model_1.PCON [0], _43170_, clk);
  dff _87383_ (\oc8051_golden_model_1.PCON [1], _43171_, clk);
  dff _87384_ (\oc8051_golden_model_1.PCON [2], _43172_, clk);
  dff _87385_ (\oc8051_golden_model_1.PCON [3], _43173_, clk);
  dff _87386_ (\oc8051_golden_model_1.PCON [4], _43174_, clk);
  dff _87387_ (\oc8051_golden_model_1.PCON [5], _43175_, clk);
  dff _87388_ (\oc8051_golden_model_1.PCON [6], _43176_, clk);
  dff _87389_ (\oc8051_golden_model_1.PCON [7], _40575_, clk);
  dff _87390_ (\oc8051_golden_model_1.TMOD [0], _43178_, clk);
  dff _87391_ (\oc8051_golden_model_1.TMOD [1], _43179_, clk);
  dff _87392_ (\oc8051_golden_model_1.TMOD [2], _43180_, clk);
  dff _87393_ (\oc8051_golden_model_1.TMOD [3], _43182_, clk);
  dff _87394_ (\oc8051_golden_model_1.TMOD [4], _43183_, clk);
  dff _87395_ (\oc8051_golden_model_1.TMOD [5], _43184_, clk);
  dff _87396_ (\oc8051_golden_model_1.TMOD [6], _43185_, clk);
  dff _87397_ (\oc8051_golden_model_1.TMOD [7], _40576_, clk);
  dff _87398_ (\oc8051_golden_model_1.DPL [0], _43187_, clk);
  dff _87399_ (\oc8051_golden_model_1.DPL [1], _43188_, clk);
  dff _87400_ (\oc8051_golden_model_1.DPL [2], _43189_, clk);
  dff _87401_ (\oc8051_golden_model_1.DPL [3], _43190_, clk);
  dff _87402_ (\oc8051_golden_model_1.DPL [4], _43191_, clk);
  dff _87403_ (\oc8051_golden_model_1.DPL [5], _43192_, clk);
  dff _87404_ (\oc8051_golden_model_1.DPL [6], _43193_, clk);
  dff _87405_ (\oc8051_golden_model_1.DPL [7], _40577_, clk);
  dff _87406_ (\oc8051_golden_model_1.DPH [0], _43195_, clk);
  dff _87407_ (\oc8051_golden_model_1.DPH [1], _43196_, clk);
  dff _87408_ (\oc8051_golden_model_1.DPH [2], _43197_, clk);
  dff _87409_ (\oc8051_golden_model_1.DPH [3], _43198_, clk);
  dff _87410_ (\oc8051_golden_model_1.DPH [4], _43199_, clk);
  dff _87411_ (\oc8051_golden_model_1.DPH [5], _43200_, clk);
  dff _87412_ (\oc8051_golden_model_1.DPH [6], _43201_, clk);
  dff _87413_ (\oc8051_golden_model_1.DPH [7], _40580_, clk);
  dff _87414_ (\oc8051_golden_model_1.TL1 [0], _43202_, clk);
  dff _87415_ (\oc8051_golden_model_1.TL1 [1], _43204_, clk);
  dff _87416_ (\oc8051_golden_model_1.TL1 [2], _43205_, clk);
  dff _87417_ (\oc8051_golden_model_1.TL1 [3], _43206_, clk);
  dff _87418_ (\oc8051_golden_model_1.TL1 [4], _43207_, clk);
  dff _87419_ (\oc8051_golden_model_1.TL1 [5], _43208_, clk);
  dff _87420_ (\oc8051_golden_model_1.TL1 [6], _43209_, clk);
  dff _87421_ (\oc8051_golden_model_1.TL1 [7], _40581_, clk);
  dff _87422_ (\oc8051_golden_model_1.TL0 [0], _43211_, clk);
  dff _87423_ (\oc8051_golden_model_1.TL0 [1], _43212_, clk);
  dff _87424_ (\oc8051_golden_model_1.TL0 [2], _43213_, clk);
  dff _87425_ (\oc8051_golden_model_1.TL0 [3], _43214_, clk);
  dff _87426_ (\oc8051_golden_model_1.TL0 [4], _43215_, clk);
  dff _87427_ (\oc8051_golden_model_1.TL0 [5], _43216_, clk);
  dff _87428_ (\oc8051_golden_model_1.TL0 [6], _43217_, clk);
  dff _87429_ (\oc8051_golden_model_1.TL0 [7], _40582_, clk);
  dff _87430_ (\oc8051_golden_model_1.TCON [0], _43219_, clk);
  dff _87431_ (\oc8051_golden_model_1.TCON [1], _43220_, clk);
  dff _87432_ (\oc8051_golden_model_1.TCON [2], _43221_, clk);
  dff _87433_ (\oc8051_golden_model_1.TCON [3], _43223_, clk);
  dff _87434_ (\oc8051_golden_model_1.TCON [4], _43224_, clk);
  dff _87435_ (\oc8051_golden_model_1.TCON [5], _43225_, clk);
  dff _87436_ (\oc8051_golden_model_1.TCON [6], _43226_, clk);
  dff _87437_ (\oc8051_golden_model_1.TCON [7], _40583_, clk);
  dff _87438_ (\oc8051_golden_model_1.TH1 [0], _43228_, clk);
  dff _87439_ (\oc8051_golden_model_1.TH1 [1], _43229_, clk);
  dff _87440_ (\oc8051_golden_model_1.TH1 [2], _43230_, clk);
  dff _87441_ (\oc8051_golden_model_1.TH1 [3], _43231_, clk);
  dff _87442_ (\oc8051_golden_model_1.TH1 [4], _43232_, clk);
  dff _87443_ (\oc8051_golden_model_1.TH1 [5], _43233_, clk);
  dff _87444_ (\oc8051_golden_model_1.TH1 [6], _43234_, clk);
  dff _87445_ (\oc8051_golden_model_1.TH1 [7], _40584_, clk);
  dff _87446_ (\oc8051_golden_model_1.TH0 [0], _43236_, clk);
  dff _87447_ (\oc8051_golden_model_1.TH0 [1], _43237_, clk);
  dff _87448_ (\oc8051_golden_model_1.TH0 [2], _43238_, clk);
  dff _87449_ (\oc8051_golden_model_1.TH0 [3], _43239_, clk);
  dff _87450_ (\oc8051_golden_model_1.TH0 [4], _43240_, clk);
  dff _87451_ (\oc8051_golden_model_1.TH0 [5], _43242_, clk);
  dff _87452_ (\oc8051_golden_model_1.TH0 [6], _43243_, clk);
  dff _87453_ (\oc8051_golden_model_1.TH0 [7], _40585_, clk);
  dff _87454_ (\oc8051_golden_model_1.PC [0], _43245_, clk);
  dff _87455_ (\oc8051_golden_model_1.PC [1], _43246_, clk);
  dff _87456_ (\oc8051_golden_model_1.PC [2], _43247_, clk);
  dff _87457_ (\oc8051_golden_model_1.PC [3], _43249_, clk);
  dff _87458_ (\oc8051_golden_model_1.PC [4], _43250_, clk);
  dff _87459_ (\oc8051_golden_model_1.PC [5], _43251_, clk);
  dff _87460_ (\oc8051_golden_model_1.PC [6], _43252_, clk);
  dff _87461_ (\oc8051_golden_model_1.PC [7], _43253_, clk);
  dff _87462_ (\oc8051_golden_model_1.PC [8], _43254_, clk);
  dff _87463_ (\oc8051_golden_model_1.PC [9], _43255_, clk);
  dff _87464_ (\oc8051_golden_model_1.PC [10], _43256_, clk);
  dff _87465_ (\oc8051_golden_model_1.PC [11], _43257_, clk);
  dff _87466_ (\oc8051_golden_model_1.PC [12], _43258_, clk);
  dff _87467_ (\oc8051_golden_model_1.PC [13], _43260_, clk);
  dff _87468_ (\oc8051_golden_model_1.PC [14], _43261_, clk);
  dff _87469_ (\oc8051_golden_model_1.PC [15], _40586_, clk);
  dff _87470_ (\oc8051_golden_model_1.P2 [0], _43262_, clk);
  dff _87471_ (\oc8051_golden_model_1.P2 [1], _43264_, clk);
  dff _87472_ (\oc8051_golden_model_1.P2 [2], _43265_, clk);
  dff _87473_ (\oc8051_golden_model_1.P2 [3], _43266_, clk);
  dff _87474_ (\oc8051_golden_model_1.P2 [4], _43267_, clk);
  dff _87475_ (\oc8051_golden_model_1.P2 [5], _43268_, clk);
  dff _87476_ (\oc8051_golden_model_1.P2 [6], _43269_, clk);
  dff _87477_ (\oc8051_golden_model_1.P2 [7], _40587_, clk);
  dff _87478_ (\oc8051_golden_model_1.P3 [0], _43271_, clk);
  dff _87479_ (\oc8051_golden_model_1.P3 [1], _43272_, clk);
  dff _87480_ (\oc8051_golden_model_1.P3 [2], _43273_, clk);
  dff _87481_ (\oc8051_golden_model_1.P3 [3], _43274_, clk);
  dff _87482_ (\oc8051_golden_model_1.P3 [4], _43275_, clk);
  dff _87483_ (\oc8051_golden_model_1.P3 [5], _43276_, clk);
  dff _87484_ (\oc8051_golden_model_1.P3 [6], _43277_, clk);
  dff _87485_ (\oc8051_golden_model_1.P3 [7], _40588_, clk);
  dff _87486_ (\oc8051_golden_model_1.P0 [0], _43279_, clk);
  dff _87487_ (\oc8051_golden_model_1.P0 [1], _43280_, clk);
  dff _87488_ (\oc8051_golden_model_1.P0 [2], _43281_, clk);
  dff _87489_ (\oc8051_golden_model_1.P0 [3], _43283_, clk);
  dff _87490_ (\oc8051_golden_model_1.P0 [4], _43284_, clk);
  dff _87491_ (\oc8051_golden_model_1.P0 [5], _43285_, clk);
  dff _87492_ (\oc8051_golden_model_1.P0 [6], _43286_, clk);
  dff _87493_ (\oc8051_golden_model_1.P0 [7], _40589_, clk);
  dff _87494_ (\oc8051_golden_model_1.P1 [0], _43288_, clk);
  dff _87495_ (\oc8051_golden_model_1.P1 [1], _43289_, clk);
  dff _87496_ (\oc8051_golden_model_1.P1 [2], _43290_, clk);
  dff _87497_ (\oc8051_golden_model_1.P1 [3], _43291_, clk);
  dff _87498_ (\oc8051_golden_model_1.P1 [4], _43292_, clk);
  dff _87499_ (\oc8051_golden_model_1.P1 [5], _43293_, clk);
  dff _87500_ (\oc8051_golden_model_1.P1 [6], _43294_, clk);
  dff _87501_ (\oc8051_golden_model_1.P1 [7], _40591_, clk);
  dff _87502_ (\oc8051_golden_model_1.IP [0], _43296_, clk);
  dff _87503_ (\oc8051_golden_model_1.IP [1], _43297_, clk);
  dff _87504_ (\oc8051_golden_model_1.IP [2], _43298_, clk);
  dff _87505_ (\oc8051_golden_model_1.IP [3], _43299_, clk);
  dff _87506_ (\oc8051_golden_model_1.IP [4], _43300_, clk);
  dff _87507_ (\oc8051_golden_model_1.IP [5], _43302_, clk);
  dff _87508_ (\oc8051_golden_model_1.IP [6], _43303_, clk);
  dff _87509_ (\oc8051_golden_model_1.IP [7], _40592_, clk);
  dff _87510_ (\oc8051_golden_model_1.IE [0], _43304_, clk);
  dff _87511_ (\oc8051_golden_model_1.IE [1], _43306_, clk);
  dff _87512_ (\oc8051_golden_model_1.IE [2], _43307_, clk);
  dff _87513_ (\oc8051_golden_model_1.IE [3], _43308_, clk);
  dff _87514_ (\oc8051_golden_model_1.IE [4], _43309_, clk);
  dff _87515_ (\oc8051_golden_model_1.IE [5], _43310_, clk);
  dff _87516_ (\oc8051_golden_model_1.IE [6], _43311_, clk);
  dff _87517_ (\oc8051_golden_model_1.IE [7], _40593_, clk);
  dff _87518_ (\oc8051_golden_model_1.SCON [0], _43313_, clk);
  dff _87519_ (\oc8051_golden_model_1.SCON [1], _43314_, clk);
  dff _87520_ (\oc8051_golden_model_1.SCON [2], _43315_, clk);
  dff _87521_ (\oc8051_golden_model_1.SCON [3], _43316_, clk);
  dff _87522_ (\oc8051_golden_model_1.SCON [4], _43317_, clk);
  dff _87523_ (\oc8051_golden_model_1.SCON [5], _43318_, clk);
  dff _87524_ (\oc8051_golden_model_1.SCON [6], _43319_, clk);
  dff _87525_ (\oc8051_golden_model_1.SCON [7], _40594_, clk);
  dff _87526_ (\oc8051_golden_model_1.SP [0], _43321_, clk);
  dff _87527_ (\oc8051_golden_model_1.SP [1], _43322_, clk);
  dff _87528_ (\oc8051_golden_model_1.SP [2], _43323_, clk);
  dff _87529_ (\oc8051_golden_model_1.SP [3], _43325_, clk);
  dff _87530_ (\oc8051_golden_model_1.SP [4], _43326_, clk);
  dff _87531_ (\oc8051_golden_model_1.SP [5], _43327_, clk);
  dff _87532_ (\oc8051_golden_model_1.SP [6], _43328_, clk);
  dff _87533_ (\oc8051_golden_model_1.SP [7], _40595_, clk);
  dff _87534_ (\oc8051_golden_model_1.SBUF [0], _43330_, clk);
  dff _87535_ (\oc8051_golden_model_1.SBUF [1], _43331_, clk);
  dff _87536_ (\oc8051_golden_model_1.SBUF [2], _43332_, clk);
  dff _87537_ (\oc8051_golden_model_1.SBUF [3], _43333_, clk);
  dff _87538_ (\oc8051_golden_model_1.SBUF [4], _43334_, clk);
  dff _87539_ (\oc8051_golden_model_1.SBUF [5], _43335_, clk);
  dff _87540_ (\oc8051_golden_model_1.SBUF [6], _43336_, clk);
  dff _87541_ (\oc8051_golden_model_1.SBUF [7], _40597_, clk);
  dff _87542_ (\oc8051_golden_model_1.PSW [0], _43338_, clk);
  dff _87543_ (\oc8051_golden_model_1.PSW [1], _43339_, clk);
  dff _87544_ (\oc8051_golden_model_1.PSW [2], _43340_, clk);
  dff _87545_ (\oc8051_golden_model_1.PSW [3], _43341_, clk);
  dff _87546_ (\oc8051_golden_model_1.PSW [4], _43342_, clk);
  dff _87547_ (\oc8051_golden_model_1.PSW [5], _43344_, clk);
  dff _87548_ (\oc8051_golden_model_1.PSW [6], _43345_, clk);
  dff _87549_ (\oc8051_golden_model_1.PSW [7], _40598_, clk);
  dff _87550_ (\oc8051_golden_model_1.IRAM[0] [0], _40612_, clk);
  dff _87551_ (\oc8051_golden_model_1.IRAM[0] [1], _40613_, clk);
  dff _87552_ (\oc8051_golden_model_1.IRAM[0] [2], _40614_, clk);
  dff _87553_ (\oc8051_golden_model_1.IRAM[0] [3], _40615_, clk);
  dff _87554_ (\oc8051_golden_model_1.IRAM[0] [4], _40616_, clk);
  dff _87555_ (\oc8051_golden_model_1.IRAM[0] [5], _40618_, clk);
  dff _87556_ (\oc8051_golden_model_1.IRAM[0] [6], _40619_, clk);
  dff _87557_ (\oc8051_golden_model_1.IRAM[0] [7], _40620_, clk);
  dff _87558_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02836_, clk);
  dff _87559_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02848_, clk);
  dff _87560_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02870_, clk);
  dff _87561_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02894_, clk);
  dff _87562_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02916_, clk);
  dff _87563_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00951_, clk);
  dff _87564_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02927_, clk);
  dff _87565_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00925_, clk);
  dff _87566_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02940_, clk);
  dff _87567_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02954_, clk);
  dff _87568_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02967_, clk);
  dff _87569_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02981_, clk);
  dff _87570_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _02995_, clk);
  dff _87571_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03008_, clk);
  dff _87572_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03022_, clk);
  dff _87573_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00971_, clk);
  dff _87574_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02354_, clk);
  dff _87575_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22124_, clk);
  dff _87576_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02542_, clk);
  dff _87577_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02700_, clk);
  dff _87578_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02882_, clk);
  dff _87579_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03125_, clk);
  dff _87580_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03328_, clk);
  dff _87581_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03527_, clk);
  dff _87582_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03728_, clk);
  dff _87583_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03927_, clk);
  dff _87584_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04023_, clk);
  dff _87585_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04123_, clk);
  dff _87586_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04222_, clk);
  dff _87587_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04321_, clk);
  dff _87588_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04414_, clk);
  dff _87589_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04512_, clk);
  dff _87590_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04611_, clk);
  dff _87591_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24283_, clk);
  dff _87592_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38656_, clk);
  dff _87593_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38658_, clk);
  dff _87594_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38659_, clk);
  dff _87595_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38660_, clk);
  dff _87596_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38661_, clk);
  dff _87597_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38662_, clk);
  dff _87598_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38663_, clk);
  dff _87599_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38643_, clk);
  dff _87600_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38664_, clk);
  dff _87601_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38665_, clk);
  dff _87602_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38667_, clk);
  dff _87603_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38668_, clk);
  dff _87604_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38669_, clk);
  dff _87605_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38670_, clk);
  dff _87606_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38671_, clk);
  dff _87607_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38644_, clk);
  dff _87608_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38673_, clk);
  dff _87609_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38674_, clk);
  dff _87610_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38675_, clk);
  dff _87611_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38676_, clk);
  dff _87612_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38677_, clk);
  dff _87613_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38679_, clk);
  dff _87614_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38680_, clk);
  dff _87615_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38646_, clk);
  dff _87616_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34184_, clk);
  dff _87617_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34187_, clk);
  dff _87618_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09680_, clk);
  dff _87619_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34189_, clk);
  dff _87620_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34191_, clk);
  dff _87621_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09683_, clk);
  dff _87622_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34193_, clk);
  dff _87623_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09686_, clk);
  dff _87624_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34195_, clk);
  dff _87625_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34197_, clk);
  dff _87626_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34199_, clk);
  dff _87627_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09689_, clk);
  dff _87628_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34201_, clk);
  dff _87629_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09692_, clk);
  dff _87630_ (\oc8051_top_1.oc8051_decoder1.wr , _09695_, clk);
  dff _87631_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09754_, clk);
  dff _87632_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09756_, clk);
  dff _87633_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09659_, clk);
  dff _87634_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09759_, clk);
  dff _87635_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09762_, clk);
  dff _87636_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09662_, clk);
  dff _87637_ (\oc8051_top_1.oc8051_decoder1.state [0], _09765_, clk);
  dff _87638_ (\oc8051_top_1.oc8051_decoder1.state [1], _09665_, clk);
  dff _87639_ (\oc8051_top_1.oc8051_decoder1.op [0], _09768_, clk);
  dff _87640_ (\oc8051_top_1.oc8051_decoder1.op [1], _09771_, clk);
  dff _87641_ (\oc8051_top_1.oc8051_decoder1.op [2], _09774_, clk);
  dff _87642_ (\oc8051_top_1.oc8051_decoder1.op [3], _09777_, clk);
  dff _87643_ (\oc8051_top_1.oc8051_decoder1.op [4], _09780_, clk);
  dff _87644_ (\oc8051_top_1.oc8051_decoder1.op [5], _09783_, clk);
  dff _87645_ (\oc8051_top_1.oc8051_decoder1.op [6], _09786_, clk);
  dff _87646_ (\oc8051_top_1.oc8051_decoder1.op [7], _09668_, clk);
  dff _87647_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09671_, clk);
  dff _87648_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34182_, clk);
  dff _87649_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09677_, clk);
  dff _87650_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09789_, clk);
  dff _87651_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09674_, clk);
  dff _87652_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39457_, clk);
  dff _87653_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _39555_, clk);
  dff _87654_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _39556_, clk);
  dff _87655_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _39557_, clk);
  dff _87656_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _39558_, clk);
  dff _87657_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _39559_, clk);
  dff _87658_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _39560_, clk);
  dff _87659_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _39561_, clk);
  dff _87660_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39458_, clk);
  dff _87661_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _39562_, clk);
  dff _87662_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _39563_, clk);
  dff _87663_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _39564_, clk);
  dff _87664_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _39566_, clk);
  dff _87665_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _39567_, clk);
  dff _87666_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _39568_, clk);
  dff _87667_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _39569_, clk);
  dff _87668_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39459_, clk);
  dff _87669_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _39570_, clk);
  dff _87670_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _39571_, clk);
  dff _87671_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _39572_, clk);
  dff _87672_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _39573_, clk);
  dff _87673_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _39574_, clk);
  dff _87674_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _39575_, clk);
  dff _87675_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _39577_, clk);
  dff _87676_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39460_, clk);
  dff _87677_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _39578_, clk);
  dff _87678_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _39579_, clk);
  dff _87679_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _39580_, clk);
  dff _87680_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _39581_, clk);
  dff _87681_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _39582_, clk);
  dff _87682_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _39583_, clk);
  dff _87683_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _39584_, clk);
  dff _87684_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39462_, clk);
  dff _87685_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _39585_, clk);
  dff _87686_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _39586_, clk);
  dff _87687_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _39588_, clk);
  dff _87688_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _39589_, clk);
  dff _87689_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _39590_, clk);
  dff _87690_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _39591_, clk);
  dff _87691_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _39592_, clk);
  dff _87692_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _39463_, clk);
  dff _87693_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _39593_, clk);
  dff _87694_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _39594_, clk);
  dff _87695_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _39595_, clk);
  dff _87696_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _39596_, clk);
  dff _87697_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _39597_, clk);
  dff _87698_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _39599_, clk);
  dff _87699_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _39600_, clk);
  dff _87700_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _39464_, clk);
  dff _87701_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _39601_, clk);
  dff _87702_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _39602_, clk);
  dff _87703_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _39603_, clk);
  dff _87704_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _39604_, clk);
  dff _87705_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _39605_, clk);
  dff _87706_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _39606_, clk);
  dff _87707_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _39607_, clk);
  dff _87708_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _39465_, clk);
  dff _87709_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _39608_, clk);
  dff _87710_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _39610_, clk);
  dff _87711_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _39611_, clk);
  dff _87712_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _39612_, clk);
  dff _87713_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _39613_, clk);
  dff _87714_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _39614_, clk);
  dff _87715_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _39615_, clk);
  dff _87716_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _39466_, clk);
  dff _87717_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39027_, clk);
  dff _87718_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39028_, clk);
  dff _87719_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39029_, clk);
  dff _87720_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39030_, clk);
  dff _87721_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38743_, clk);
  dff _87722_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38816_, clk);
  dff _87723_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38817_, clk);
  dff _87724_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38818_, clk);
  dff _87725_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38819_, clk);
  dff _87726_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38820_, clk);
  dff _87727_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38822_, clk);
  dff _87728_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38823_, clk);
  dff _87729_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38824_, clk);
  dff _87730_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38825_, clk);
  dff _87731_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38826_, clk);
  dff _87732_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38827_, clk);
  dff _87733_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38828_, clk);
  dff _87734_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38829_, clk);
  dff _87735_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _38830_, clk);
  dff _87736_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _38831_, clk);
  dff _87737_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38705_, clk);
  dff _87738_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _38836_, clk);
  dff _87739_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _38837_, clk);
  dff _87740_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _38838_, clk);
  dff _87741_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _38839_, clk);
  dff _87742_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _38840_, clk);
  dff _87743_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _38841_, clk);
  dff _87744_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _38842_, clk);
  dff _87745_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _38843_, clk);
  dff _87746_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _38844_, clk);
  dff _87747_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _38845_, clk);
  dff _87748_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _38847_, clk);
  dff _87749_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _38848_, clk);
  dff _87750_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _38849_, clk);
  dff _87751_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _38850_, clk);
  dff _87752_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _38851_, clk);
  dff _87753_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38706_, clk);
  dff _87754_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39031_, clk);
  dff _87755_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39032_, clk);
  dff _87756_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39033_, clk);
  dff _87757_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39034_, clk);
  dff _87758_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39036_, clk);
  dff _87759_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39037_, clk);
  dff _87760_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39038_, clk);
  dff _87761_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39039_, clk);
  dff _87762_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39040_, clk);
  dff _87763_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39041_, clk);
  dff _87764_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39042_, clk);
  dff _87765_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39043_, clk);
  dff _87766_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39044_, clk);
  dff _87767_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39045_, clk);
  dff _87768_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39047_, clk);
  dff _87769_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39048_, clk);
  dff _87770_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39049_, clk);
  dff _87771_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39050_, clk);
  dff _87772_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39051_, clk);
  dff _87773_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39052_, clk);
  dff _87774_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39053_, clk);
  dff _87775_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39054_, clk);
  dff _87776_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39055_, clk);
  dff _87777_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39056_, clk);
  dff _87778_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39058_, clk);
  dff _87779_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39059_, clk);
  dff _87780_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39060_, clk);
  dff _87781_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39061_, clk);
  dff _87782_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39062_, clk);
  dff _87783_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39063_, clk);
  dff _87784_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39064_, clk);
  dff _87785_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38768_, clk);
  dff _87786_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38741_, clk);
  dff _87787_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _87788_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39065_, clk);
  dff _87789_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39067_, clk);
  dff _87790_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39068_, clk);
  dff _87791_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39069_, clk);
  dff _87792_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39070_, clk);
  dff _87793_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39071_, clk);
  dff _87794_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39073_, clk);
  dff _87795_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38744_, clk);
  dff _87796_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39074_, clk);
  dff _87797_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39075_, clk);
  dff _87798_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39076_, clk);
  dff _87799_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39077_, clk);
  dff _87800_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39078_, clk);
  dff _87801_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39079_, clk);
  dff _87802_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39080_, clk);
  dff _87803_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38745_, clk);
  dff _87804_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39081_, clk);
  dff _87805_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39082_, clk);
  dff _87806_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39084_, clk);
  dff _87807_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39085_, clk);
  dff _87808_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39086_, clk);
  dff _87809_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39087_, clk);
  dff _87810_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39088_, clk);
  dff _87811_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38747_, clk);
  dff _87812_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38748_, clk);
  dff _87813_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38749_, clk);
  dff _87814_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39089_, clk);
  dff _87815_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39090_, clk);
  dff _87816_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39091_, clk);
  dff _87817_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39092_, clk);
  dff _87818_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39093_, clk);
  dff _87819_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39095_, clk);
  dff _87820_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39096_, clk);
  dff _87821_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38750_, clk);
  dff _87822_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39097_, clk);
  dff _87823_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39098_, clk);
  dff _87824_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39099_, clk);
  dff _87825_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39100_, clk);
  dff _87826_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39101_, clk);
  dff _87827_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39102_, clk);
  dff _87828_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39103_, clk);
  dff _87829_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39104_, clk);
  dff _87830_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39106_, clk);
  dff _87831_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39107_, clk);
  dff _87832_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39108_, clk);
  dff _87833_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39109_, clk);
  dff _87834_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39110_, clk);
  dff _87835_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39111_, clk);
  dff _87836_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39112_, clk);
  dff _87837_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38751_, clk);
  dff _87838_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39113_, clk);
  dff _87839_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39114_, clk);
  dff _87840_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39115_, clk);
  dff _87841_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39117_, clk);
  dff _87842_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39118_, clk);
  dff _87843_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39119_, clk);
  dff _87844_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39120_, clk);
  dff _87845_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39121_, clk);
  dff _87846_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39122_, clk);
  dff _87847_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39123_, clk);
  dff _87848_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39124_, clk);
  dff _87849_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39125_, clk);
  dff _87850_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39126_, clk);
  dff _87851_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39128_, clk);
  dff _87852_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39129_, clk);
  dff _87853_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38753_, clk);
  dff _87854_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38754_, clk);
  dff _87855_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38756_, clk);
  dff _87856_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38755_, clk);
  dff _87857_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39130_, clk);
  dff _87858_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39131_, clk);
  dff _87859_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39132_, clk);
  dff _87860_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39133_, clk);
  dff _87861_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39134_, clk);
  dff _87862_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39135_, clk);
  dff _87863_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39136_, clk);
  dff _87864_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38758_, clk);
  dff _87865_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39137_, clk);
  dff _87866_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39139_, clk);
  dff _87867_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38759_, clk);
  dff _87868_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39140_, clk);
  dff _87869_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39141_, clk);
  dff _87870_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39142_, clk);
  dff _87871_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39143_, clk);
  dff _87872_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39144_, clk);
  dff _87873_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39145_, clk);
  dff _87874_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39146_, clk);
  dff _87875_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38760_, clk);
  dff _87876_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39147_, clk);
  dff _87877_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39148_, clk);
  dff _87878_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39150_, clk);
  dff _87879_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39151_, clk);
  dff _87880_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39152_, clk);
  dff _87881_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39153_, clk);
  dff _87882_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39154_, clk);
  dff _87883_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38761_, clk);
  dff _87884_ (\oc8051_top_1.oc8051_memory_interface1.reti , _38762_, clk);
  dff _87885_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39155_, clk);
  dff _87886_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39156_, clk);
  dff _87887_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39157_, clk);
  dff _87888_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39158_, clk);
  dff _87889_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39159_, clk);
  dff _87890_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39161_, clk);
  dff _87891_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39162_, clk);
  dff _87892_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38763_, clk);
  dff _87893_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _38765_, clk);
  dff _87894_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38766_, clk);
  dff _87895_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39163_, clk);
  dff _87896_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39164_, clk);
  dff _87897_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39165_, clk);
  dff _87898_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38767_, clk);
  dff _87899_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39166_, clk);
  dff _87900_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39167_, clk);
  dff _87901_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39168_, clk);
  dff _87902_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39169_, clk);
  dff _87903_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39170_, clk);
  dff _87904_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39171_, clk);
  dff _87905_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39172_, clk);
  dff _87906_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39173_, clk);
  dff _87907_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39174_, clk);
  dff _87908_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39175_, clk);
  dff _87909_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39176_, clk);
  dff _87910_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39177_, clk);
  dff _87911_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39178_, clk);
  dff _87912_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39179_, clk);
  dff _87913_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39180_, clk);
  dff _87914_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39182_, clk);
  dff _87915_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39183_, clk);
  dff _87916_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39184_, clk);
  dff _87917_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39185_, clk);
  dff _87918_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39186_, clk);
  dff _87919_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39187_, clk);
  dff _87920_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39188_, clk);
  dff _87921_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39189_, clk);
  dff _87922_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39190_, clk);
  dff _87923_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39191_, clk);
  dff _87924_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39193_, clk);
  dff _87925_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39194_, clk);
  dff _87926_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39195_, clk);
  dff _87927_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39196_, clk);
  dff _87928_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39197_, clk);
  dff _87929_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39198_, clk);
  dff _87930_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38769_, clk);
  dff _87931_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39199_, clk);
  dff _87932_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39200_, clk);
  dff _87933_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39201_, clk);
  dff _87934_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39202_, clk);
  dff _87935_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39204_, clk);
  dff _87936_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39205_, clk);
  dff _87937_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39206_, clk);
  dff _87938_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38770_, clk);
  dff _87939_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38771_, clk);
  dff _87940_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38773_, clk);
  dff _87941_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39207_, clk);
  dff _87942_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39208_, clk);
  dff _87943_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39209_, clk);
  dff _87944_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39210_, clk);
  dff _87945_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39211_, clk);
  dff _87946_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39212_, clk);
  dff _87947_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39213_, clk);
  dff _87948_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39215_, clk);
  dff _87949_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39216_, clk);
  dff _87950_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39217_, clk);
  dff _87951_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39218_, clk);
  dff _87952_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39219_, clk);
  dff _87953_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39220_, clk);
  dff _87954_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39221_, clk);
  dff _87955_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39222_, clk);
  dff _87956_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38774_, clk);
  dff _87957_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38775_, clk);
  dff _87958_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38776_, clk);
  dff _87959_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38777_, clk);
  dff _87960_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39223_, clk);
  dff _87961_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39224_, clk);
  dff _87962_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39226_, clk);
  dff _87963_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39227_, clk);
  dff _87964_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39228_, clk);
  dff _87965_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39229_, clk);
  dff _87966_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39230_, clk);
  dff _87967_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39231_, clk);
  dff _87968_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39232_, clk);
  dff _87969_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39233_, clk);
  dff _87970_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39234_, clk);
  dff _87971_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39235_, clk);
  dff _87972_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39237_, clk);
  dff _87973_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39238_, clk);
  dff _87974_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39239_, clk);
  dff _87975_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38778_, clk);
  dff _87976_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38779_, clk);
  dff _87977_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39843_, clk);
  dff _87978_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39864_, clk);
  dff _87979_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39865_, clk);
  dff _87980_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39866_, clk);
  dff _87981_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39867_, clk);
  dff _87982_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39868_, clk);
  dff _87983_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39869_, clk);
  dff _87984_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39870_, clk);
  dff _87985_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39844_, clk);
  dff _87986_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39845_, clk);
  dff _87987_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39871_, clk);
  dff _87988_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39872_, clk);
  dff _87989_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39846_, clk);
  dff _87990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02798_, clk);
  dff _87991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02803_, clk);
  dff _87992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02809_, clk);
  dff _87993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02814_, clk);
  dff _87994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02819_, clk);
  dff _87995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02824_, clk);
  dff _87996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02829_, clk);
  dff _87997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02831_, clk);
  dff _87998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02839_, clk);
  dff _87999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02842_, clk);
  dff _88000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02846_, clk);
  dff _88001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02850_, clk);
  dff _88002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02853_, clk);
  dff _88003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02856_, clk);
  dff _88004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02860_, clk);
  dff _88005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02862_, clk);
  dff _88006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02868_, clk);
  dff _88007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02873_, clk);
  dff _88008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02876_, clk);
  dff _88009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02879_, clk);
  dff _88010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02884_, clk);
  dff _88011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02887_, clk);
  dff _88012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02890_, clk);
  dff _88013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02893_, clk);
  dff _88014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02929_, clk);
  dff _88015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02933_, clk);
  dff _88016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02937_, clk);
  dff _88017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02941_, clk);
  dff _88018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02945_, clk);
  dff _88019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02948_, clk);
  dff _88020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02952_, clk);
  dff _88021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02956_, clk);
  dff _88022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02898_, clk);
  dff _88023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02902_, clk);
  dff _88024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02905_, clk);
  dff _88025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02908_, clk);
  dff _88026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02911_, clk);
  dff _88027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02915_, clk);
  dff _88028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02918_, clk);
  dff _88029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02921_, clk);
  dff _88030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03140_, clk);
  dff _88031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03143_, clk);
  dff _88032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03146_, clk);
  dff _88033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03149_, clk);
  dff _88034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03153_, clk);
  dff _88035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03156_, clk);
  dff _88036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03159_, clk);
  dff _88037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03162_, clk);
  dff _88038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03112_, clk);
  dff _88039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03115_, clk);
  dff _88040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03119_, clk);
  dff _88041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03122_, clk);
  dff _88042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03126_, clk);
  dff _88043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03130_, clk);
  dff _88044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03133_, clk);
  dff _88045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03136_, clk);
  dff _88046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03083_, clk);
  dff _88047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03087_, clk);
  dff _88048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03090_, clk);
  dff _88049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03094_, clk);
  dff _88050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03097_, clk);
  dff _88051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03101_, clk);
  dff _88052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03104_, clk);
  dff _88053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03107_, clk);
  dff _88054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03055_, clk);
  dff _88055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03058_, clk);
  dff _88056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03062_, clk);
  dff _88057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03065_, clk);
  dff _88058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03069_, clk);
  dff _88059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03072_, clk);
  dff _88060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03076_, clk);
  dff _88061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03079_, clk);
  dff _88062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03026_, clk);
  dff _88063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03030_, clk);
  dff _88064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03033_, clk);
  dff _88065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03037_, clk);
  dff _88066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03040_, clk);
  dff _88067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03043_, clk);
  dff _88068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03046_, clk);
  dff _88069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03049_, clk);
  dff _88070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02993_, clk);
  dff _88071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _02998_, clk);
  dff _88072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03002_, clk);
  dff _88073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03005_, clk);
  dff _88074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03010_, clk);
  dff _88075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03014_, clk);
  dff _88076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03017_, clk);
  dff _88077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03020_, clk);
  dff _88078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02960_, clk);
  dff _88079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02964_, clk);
  dff _88080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02969_, clk);
  dff _88081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02973_, clk);
  dff _88082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02977_, clk);
  dff _88083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02982_, clk);
  dff _88084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02986_, clk);
  dff _88085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02988_, clk);
  dff _88086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03248_, clk);
  dff _88087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03251_, clk);
  dff _88088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03255_, clk);
  dff _88089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03258_, clk);
  dff _88090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03261_, clk);
  dff _88091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03264_, clk);
  dff _88092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03268_, clk);
  dff _88093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02574_, clk);
  dff _88094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03221_, clk);
  dff _88095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03225_, clk);
  dff _88096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03228_, clk);
  dff _88097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03232_, clk);
  dff _88098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03235_, clk);
  dff _88099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03238_, clk);
  dff _88100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03242_, clk);
  dff _88101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03244_, clk);
  dff _88102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03193_, clk);
  dff _88103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03196_, clk);
  dff _88104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03200_, clk);
  dff _88105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03204_, clk);
  dff _88106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03207_, clk);
  dff _88107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03211_, clk);
  dff _88108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03214_, clk);
  dff _88109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03217_, clk);
  dff _88110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03166_, clk);
  dff _88111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03170_, clk);
  dff _88112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03173_, clk);
  dff _88113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03176_, clk);
  dff _88114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03179_, clk);
  dff _88115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03183_, clk);
  dff _88116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03186_, clk);
  dff _88117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03188_, clk);
  dff _88118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05053_, clk);
  dff _88119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05055_, clk);
  dff _88120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05057_, clk);
  dff _88121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05059_, clk);
  dff _88122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05061_, clk);
  dff _88123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05063_, clk);
  dff _88124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05065_, clk);
  dff _88125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02564_, clk);
  dff _88126_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0], clk);
  dff _88127_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1], clk);
  dff _88128_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2], clk);
  dff _88129_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3], clk);
  dff _88130_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4], clk);
  dff _88131_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5], clk);
  dff _88132_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6], clk);
  dff _88133_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7], clk);
  dff _88134_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8], clk);
  dff _88135_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9], clk);
  dff _88136_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10], clk);
  dff _88137_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11], clk);
  dff _88138_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12], clk);
  dff _88139_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13], clk);
  dff _88140_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14], clk);
  dff _88141_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15], clk);
  dff _88142_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16], clk);
  dff _88143_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17], clk);
  dff _88144_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18], clk);
  dff _88145_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19], clk);
  dff _88146_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20], clk);
  dff _88147_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21], clk);
  dff _88148_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22], clk);
  dff _88149_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23], clk);
  dff _88150_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24], clk);
  dff _88151_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25], clk);
  dff _88152_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26], clk);
  dff _88153_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27], clk);
  dff _88154_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28], clk);
  dff _88155_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29], clk);
  dff _88156_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30], clk);
  dff _88157_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31], clk);
  dff _88158_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _88159_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _39679_, clk);
  dff _88160_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _39764_, clk);
  dff _88161_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _39765_, clk);
  dff _88162_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _39766_, clk);
  dff _88163_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _39681_, clk);
  dff _88164_ (\oc8051_top_1.oc8051_sfr1.bit_out , _39682_, clk);
  dff _88165_ (\oc8051_top_1.oc8051_sfr1.wait_data , _39683_, clk);
  dff _88166_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39768_, clk);
  dff _88167_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39769_, clk);
  dff _88168_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39770_, clk);
  dff _88169_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39771_, clk);
  dff _88170_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39772_, clk);
  dff _88171_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39773_, clk);
  dff _88172_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39774_, clk);
  dff _88173_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39684_, clk);
  dff _88174_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39685_, clk);
  dff _88175_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19757_, clk);
  dff _88176_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19769_, clk);
  dff _88177_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19780_, clk);
  dff _88178_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19792_, clk);
  dff _88179_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19804_, clk);
  dff _88180_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19816_, clk);
  dff _88181_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19828_, clk);
  dff _88182_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17963_, clk);
  dff _88183_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08867_, clk);
  dff _88184_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08878_, clk);
  dff _88185_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08889_, clk);
  dff _88186_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08900_, clk);
  dff _88187_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08911_, clk);
  dff _88188_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08922_, clk);
  dff _88189_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08933_, clk);
  dff _88190_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06626_, clk);
  dff _88191_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13613_, clk);
  dff _88192_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13624_, clk);
  dff _88193_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13635_, clk);
  dff _88194_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13646_, clk);
  dff _88195_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13657_, clk);
  dff _88196_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13668_, clk);
  dff _88197_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13679_, clk);
  dff _88198_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12677_, clk);
  dff _88199_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13690_, clk);
  dff _88200_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13701_, clk);
  dff _88201_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13711_, clk);
  dff _88202_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13722_, clk);
  dff _88203_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13733_, clk);
  dff _88204_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13744_, clk);
  dff _88205_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13755_, clk);
  dff _88206_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12698_, clk);
  dff _88207_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _42623_, clk);
  dff _88208_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _42621_, clk);
  dff _88209_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _88210_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _42618_, clk);
  dff _88211_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00130_, clk);
  dff _88212_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00132_, clk);
  dff _88213_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00134_, clk);
  dff _88214_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00136_, clk);
  dff _88215_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00138_, clk);
  dff _88216_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00139_, clk);
  dff _88217_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00141_, clk);
  dff _88218_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42616_, clk);
  dff _88219_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00143_, clk);
  dff _88220_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _42615_, clk);
  dff _88221_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _42613_, clk);
  dff _88222_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00145_, clk);
  dff _88223_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00147_, clk);
  dff _88224_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _42611_, clk);
  dff _88225_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00149_, clk);
  dff _88226_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00150_, clk);
  dff _88227_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _42609_, clk);
  dff _88228_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00152_, clk);
  dff _88229_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42607_, clk);
  dff _88230_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00154_, clk);
  dff _88231_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42605_, clk);
  dff _88232_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _42570_, clk);
  dff _88233_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _42568_, clk);
  dff _88234_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _42566_, clk);
  dff _88235_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _42564_, clk);
  dff _88236_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00156_, clk);
  dff _88237_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00158_, clk);
  dff _88238_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00160_, clk);
  dff _88239_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _42561_, clk);
  dff _88240_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00161_, clk);
  dff _88241_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00163_, clk);
  dff _88242_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00165_, clk);
  dff _88243_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00167_, clk);
  dff _88244_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00169_, clk);
  dff _88245_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00171_, clk);
  dff _88246_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00173_, clk);
  dff _88247_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _42559_, clk);
  dff _88248_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00174_, clk);
  dff _88249_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00176_, clk);
  dff _88250_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00178_, clk);
  dff _88251_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00180_, clk);
  dff _88252_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00182_, clk);
  dff _88253_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00184_, clk);
  dff _88254_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00185_, clk);
  dff _88255_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _42556_, clk);
  dff _88256_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40308_, clk);
  dff _88257_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40310_, clk);
  dff _88258_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40312_, clk);
  dff _88259_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40314_, clk);
  dff _88260_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40316_, clk);
  dff _88261_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40318_, clk);
  dff _88262_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40320_, clk);
  dff _88263_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31034_, clk);
  dff _88264_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40322_, clk);
  dff _88265_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40324_, clk);
  dff _88266_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40326_, clk);
  dff _88267_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40327_, clk);
  dff _88268_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40329_, clk);
  dff _88269_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40331_, clk);
  dff _88270_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40333_, clk);
  dff _88271_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31057_, clk);
  dff _88272_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40335_, clk);
  dff _88273_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40337_, clk);
  dff _88274_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40339_, clk);
  dff _88275_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40341_, clk);
  dff _88276_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40343_, clk);
  dff _88277_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40345_, clk);
  dff _88278_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40347_, clk);
  dff _88279_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31079_, clk);
  dff _88280_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40349_, clk);
  dff _88281_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40351_, clk);
  dff _88282_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40353_, clk);
  dff _88283_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40355_, clk);
  dff _88284_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40356_, clk);
  dff _88285_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40358_, clk);
  dff _88286_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40360_, clk);
  dff _88287_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31102_, clk);
  dff _88288_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17339_, clk);
  dff _88289_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17350_, clk);
  dff _88290_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17361_, clk);
  dff _88291_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17372_, clk);
  dff _88292_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17383_, clk);
  dff _88293_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17394_, clk);
  dff _88294_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15158_, clk);
  dff _88295_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09484_, clk);
  dff _88296_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10660_, clk);
  dff _88297_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10671_, clk);
  dff _88298_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10682_, clk);
  dff _88299_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10693_, clk);
  dff _88300_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10704_, clk);
  dff _88301_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10715_, clk);
  dff _88302_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10726_, clk);
  dff _88303_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09504_, clk);
  dff _88304_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _40810_, clk);
  dff _88305_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _40813_, clk);
  dff _88306_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41323_, clk);
  dff _88307_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41325_, clk);
  dff _88308_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41327_, clk);
  dff _88309_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41328_, clk);
  dff _88310_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41330_, clk);
  dff _88311_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41332_, clk);
  dff _88312_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41334_, clk);
  dff _88313_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _40816_, clk);
  dff _88314_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41336_, clk);
  dff _88315_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41338_, clk);
  dff _88316_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41340_, clk);
  dff _88317_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41342_, clk);
  dff _88318_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41344_, clk);
  dff _88319_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41345_, clk);
  dff _88320_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41347_, clk);
  dff _88321_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _40819_, clk);
  dff _88322_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _40822_, clk);
  dff _88323_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _40825_, clk);
  dff _88324_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41349_, clk);
  dff _88325_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41351_, clk);
  dff _88326_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41353_, clk);
  dff _88327_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41355_, clk);
  dff _88328_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41357_, clk);
  dff _88329_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41359_, clk);
  dff _88330_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41361_, clk);
  dff _88331_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _40828_, clk);
  dff _88332_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41362_, clk);
  dff _88333_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41364_, clk);
  dff _88334_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41366_, clk);
  dff _88335_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41368_, clk);
  dff _88336_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41370_, clk);
  dff _88337_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41372_, clk);
  dff _88338_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41374_, clk);
  dff _88339_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _40831_, clk);
  dff _88340_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _40834_, clk);
  dff _88341_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41376_, clk);
  dff _88342_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41378_, clk);
  dff _88343_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41379_, clk);
  dff _88344_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41381_, clk);
  dff _88345_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41383_, clk);
  dff _88346_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41385_, clk);
  dff _88347_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41387_, clk);
  dff _88348_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _40837_, clk);
  dff _88349_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01626_, clk);
  dff _88350_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01628_, clk);
  dff _88351_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01631_, clk);
  dff _88352_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01634_, clk);
  dff _88353_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02111_, clk);
  dff _88354_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02113_, clk);
  dff _88355_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02115_, clk);
  dff _88356_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02117_, clk);
  dff _88357_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02118_, clk);
  dff _88358_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02120_, clk);
  dff _88359_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02122_, clk);
  dff _88360_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01637_, clk);
  dff _88361_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02124_, clk);
  dff _88362_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02125_, clk);
  dff _88363_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02127_, clk);
  dff _88364_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02129_, clk);
  dff _88365_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02131_, clk);
  dff _88366_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02132_, clk);
  dff _88367_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02134_, clk);
  dff _88368_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01640_, clk);
  dff _88369_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01643_, clk);
  dff _88370_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02136_, clk);
  dff _88371_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02138_, clk);
  dff _88372_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02139_, clk);
  dff _88373_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02141_, clk);
  dff _88374_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02143_, clk);
  dff _88375_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02145_, clk);
  dff _88376_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02146_, clk);
  dff _88377_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01646_, clk);
  dff _88378_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02148_, clk);
  dff _88379_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02150_, clk);
  dff _88380_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02152_, clk);
  dff _88381_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02153_, clk);
  dff _88382_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02155_, clk);
  dff _88383_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02157_, clk);
  dff _88384_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02159_, clk);
  dff _88385_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01649_, clk);
  dff _88386_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01652_, clk);
  dff _88387_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02160_, clk);
  dff _88388_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02162_, clk);
  dff _88389_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02164_, clk);
  dff _88390_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02166_, clk);
  dff _88391_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02167_, clk);
  dff _88392_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02169_, clk);
  dff _88393_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02171_, clk);
  dff _88394_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01655_, clk);
  dff _88395_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01206_, clk);
  dff _88396_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01208_, clk);
  dff _88397_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01210_, clk);
  dff _88398_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01212_, clk);
  dff _88399_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01214_, clk);
  dff _88400_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01216_, clk);
  dff _88401_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01218_, clk);
  dff _88402_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01220_, clk);
  dff _88403_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01221_, clk);
  dff _88404_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01223_, clk);
  dff _88405_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01225_, clk);
  dff _88406_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00567_, clk);
  dff _88407_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00543_, clk);
  dff _88408_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00545_, clk);
  dff _88409_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00548_, clk);
  dff _88410_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00551_, clk);
  dff _88411_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00554_, clk);
  dff _88412_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00556_, clk);
  dff _88413_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01227_, clk);
  dff _88414_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00559_, clk);
  dff _88415_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01229_, clk);
  dff _88416_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01231_, clk);
  dff _88417_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01233_, clk);
  dff _88418_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00562_, clk);
  dff _88419_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01235_, clk);
  dff _88420_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01237_, clk);
  dff _88421_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01239_, clk);
  dff _88422_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01241_, clk);
  dff _88423_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01243_, clk);
  dff _88424_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01245_, clk);
  dff _88425_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01247_, clk);
  dff _88426_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00564_, clk);
  dff _88427_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00570_, clk);
  dff _88428_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00572_, clk);
  dff _88429_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00575_, clk);
  dff _88430_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00578_, clk);
  dff _88431_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00580_, clk);
  dff _88432_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01249_, clk);
  dff _88433_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01251_, clk);
  dff _88434_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01253_, clk);
  dff _88435_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00583_, clk);
  dff _88436_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01255_, clk);
  dff _88437_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01256_, clk);
  dff _88438_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01258_, clk);
  dff _88439_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01260_, clk);
  dff _88440_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01262_, clk);
  dff _88441_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01264_, clk);
  dff _88442_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01266_, clk);
  dff _88443_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01268_, clk);
  dff _88444_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01270_, clk);
  dff _88445_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01272_, clk);
  dff _88446_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00586_, clk);
  dff _88447_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01274_, clk);
  dff _88448_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01276_, clk);
  dff _88449_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01278_, clk);
  dff _88450_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01280_, clk);
  dff _88451_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01282_, clk);
  dff _88452_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01284_, clk);
  dff _88453_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01286_, clk);
  dff _88454_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00588_, clk);
  dff _88455_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01288_, clk);
  dff _88456_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01290_, clk);
  dff _88457_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01291_, clk);
  dff _88458_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01293_, clk);
  dff _88459_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01295_, clk);
  dff _88460_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01297_, clk);
  dff _88461_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01299_, clk);
  dff _88462_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00591_, clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1071 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1071 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1071 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1071 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1073 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1075 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1075 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1076 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1076 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1077 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1077 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1078 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1078 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1079 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1079 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1080 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1080 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1081 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1118 , \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.n1146 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1147 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1147 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1147 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1147 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1147 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1147 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1148 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1148 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1148 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1148 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1148 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1148 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1149 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1149 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1149 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1149 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1149 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1149 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1149 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1149 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1150 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1151 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1152 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1152 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1152 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1153 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1154 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1154 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1155 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1155 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1155 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1155 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1155 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1155 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1181 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1181 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1181 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1181 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1181 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1181 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1181 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1181 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1181 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1181 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1181 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1181 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1181 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1183 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1183 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1183 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1183 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1183 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1183 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1185 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1185 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1185 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1185 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1185 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1185 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1185 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1189 [8], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1190 , \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1191 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1191 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1191 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1191 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1192 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1192 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1192 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1196 [4], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1197 , \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1198 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1198 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1198 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1198 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1198 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1198 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1198 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1198 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1198 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1206 , \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.n1207 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1207 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1207 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1207 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1207 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1212 , \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1217 [4], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1218 , \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1226 , \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.n1227 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1227 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1227 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1227 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1227 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1229 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1229 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1229 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1229 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1229 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1229 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1229 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1229 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1229 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1231 [8], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1232 , \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1233 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1233 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1233 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1233 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1234 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1234 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1234 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1236 [4], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1237 , \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1238 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1238 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1238 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1238 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1238 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1238 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1238 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1238 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1238 [8], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1249 [8], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1257 , \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.n1258 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1258 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1258 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1258 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1258 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1260 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1262 [8], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1276 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1278 [4], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1279 , \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1280 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1280 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1280 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1280 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1280 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1280 [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1282 [8], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1290 , \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1291 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1291 [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1291 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1291 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1291 [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1292 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1292 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1292 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1292 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1292 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1295 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1295 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1295 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1295 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1295 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1295 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1295 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1295 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1295 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1296 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1296 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1296 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1296 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1296 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1296 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1297 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1297 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1297 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1297 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1297 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1297 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1297 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1297 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1298 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1299 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1299 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1299 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1299 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1299 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1299 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1299 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1299 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1300 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1300 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1303 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1305 [8], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1306 , \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1307 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1307 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1309 [4], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1310 , \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1317 , \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.n1318 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1318 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1318 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1318 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1318 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1322 [8], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1323 , \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.n1334 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1334 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1334 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1334 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1334 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1338 [8], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1339 , \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1350 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1350 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1354 [8], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1357 [4], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1358 , \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1365 , \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1520 , \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1521 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1521 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1521 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1521 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1521 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1521 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1521 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1553 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1553 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1553 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1553 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.n1555 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1555 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1555 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1555 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1555 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1555 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1555 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1680 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1683 , \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.n1685 , \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.n1691 , \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.n1692 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1692 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1692 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1692 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1692 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1696 , \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.n1698 , \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1709 , \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.n1711 , \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.n1717 , \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.n1718 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1718 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1718 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1718 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1718 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1722 , \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.n1724 , \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.n1730 , \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.n1731 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1731 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1731 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1731 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1731 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1733 , \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.n1734 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1734 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1734 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1734 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1734 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1734 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1734 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1739 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1739 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1739 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1739 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1739 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1739 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1739 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1739 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1739 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1745 , \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.n1746 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1746 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1746 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1746 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1746 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1746 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1746 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1749 , \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.n1750 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1750 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1750 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1750 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1750 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1750 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1750 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1765 , \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.n1766 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1766 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1766 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1766 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1766 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1766 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1766 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1771 , \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.n1772 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1772 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1772 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1772 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1772 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1772 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1772 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.n1778 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1778 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1778 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1778 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1778 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1778 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1778 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1783 , \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.n1784 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1784 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1784 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1784 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1784 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1784 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1784 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1789 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1791 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1791 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1791 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1791 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1791 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1791 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1792 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1792 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1792 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1792 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1793 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1793 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1793 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1793 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1793 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1793 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1828 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1828 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1828 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1828 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1828 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1828 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1828 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1828 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1847 , \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.n1848 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1848 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1848 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1848 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1848 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1848 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1848 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1852 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1854 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1854 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1854 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1854 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
